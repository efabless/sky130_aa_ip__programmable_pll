magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect -1962 760 -1621 796
rect -162 761 111 796
rect -2082 692 -1609 760
rect -215 693 258 761
rect 656 760 3392 797
rect -1962 332 -1621 692
rect -162 343 111 693
rect 584 692 3392 760
rect 656 343 3392 692
rect -163 -651 678 -645
rect -163 -1000 3379 -651
rect -205 -1068 3379 -1000
rect -163 -1104 3379 -1068
rect 643 -1105 3379 -1104
<< locali >>
rect -2082 692 -1609 760
rect -215 693 258 761
rect 584 692 1057 760
rect 2476 695 3580 763
rect 737 464 985 509
rect 737 330 782 464
rect 3324 333 3449 335
rect -1900 322 -1840 326
rect -1987 319 -1764 322
rect -2610 -131 -2571 300
rect -1987 285 -1887 319
rect -1853 285 -1764 319
rect -1987 280 -1764 285
rect -1900 241 -1840 280
rect -225 271 63 328
rect 654 295 782 330
rect 654 285 730 295
rect -1900 207 -1887 241
rect -1853 207 -1840 241
rect -1900 194 -1840 207
rect 717 261 730 285
rect 764 285 782 295
rect 832 326 892 327
rect 832 320 975 326
rect 832 286 845 320
rect 879 286 975 320
rect 764 261 777 285
rect 717 217 777 261
rect 717 183 730 217
rect 764 183 777 217
rect 832 268 975 286
rect 2442 278 2814 331
rect 3324 296 3450 333
rect 832 242 892 268
rect 832 208 845 242
rect 879 208 892 242
rect 832 195 892 208
rect -2251 52 -2114 65
rect -2251 18 -2244 52
rect -2210 18 -2166 52
rect -2132 18 -2114 52
rect -2251 5 -2114 18
rect -2015 2 -1518 70
rect -250 43 -204 175
rect 717 170 777 183
rect 376 51 513 64
rect 376 17 383 51
rect 417 17 461 51
rect 495 17 513 51
rect 376 4 513 17
rect 613 2 1133 70
rect 2980 55 3112 68
rect 2980 21 2987 55
rect 3021 21 3065 55
rect 3099 21 3112 55
rect 2980 8 3112 21
rect -1941 -45 -1809 -34
rect 2582 -45 2714 -32
rect -1941 -47 2589 -45
rect -1941 -81 -1934 -47
rect -1900 -81 -1856 -47
rect -1822 -79 2589 -47
rect 2623 -79 2667 -45
rect 2701 -79 3120 -45
rect 3402 -62 3450 296
rect -1822 -81 3120 -79
rect -1941 -84 3120 -81
rect 3391 -69 3451 -62
rect -1941 -94 -1809 -84
rect 2582 -92 2714 -84
rect 3391 -103 3404 -69
rect 3438 -103 3451 -69
rect -137 -131 -5 -120
rect 804 -131 941 -121
rect -2610 -133 3120 -131
rect -2610 -167 -130 -133
rect -96 -167 -52 -133
rect -18 -134 3120 -133
rect -18 -167 811 -134
rect -2610 -168 811 -167
rect 845 -168 889 -134
rect 923 -168 3120 -134
rect -2610 -170 3120 -168
rect 3391 -147 3451 -103
rect -137 -180 -5 -170
rect 804 -181 941 -170
rect 3391 -181 3404 -147
rect 3438 -181 3451 -147
rect 3391 -199 3451 -181
rect -2264 -217 -2132 -204
rect -2264 -223 -2257 -217
rect -2265 -251 -2257 -223
rect -2223 -251 -2179 -217
rect -2145 -223 -2132 -217
rect 369 -217 506 -204
rect 369 -223 376 -217
rect -2145 -251 376 -223
rect 410 -251 454 -217
rect 488 -223 506 -217
rect 2966 -223 3103 -210
rect 488 -251 2973 -223
rect -2265 -257 2973 -251
rect 3007 -257 3051 -223
rect 3085 -257 3120 -223
rect -2265 -262 3120 -257
rect -2264 -264 -2132 -262
rect -506 -357 -395 -262
rect 369 -264 506 -262
rect -220 -376 300 -308
rect 372 -351 483 -264
rect 2170 -355 2281 -262
rect 2966 -270 3103 -262
rect 2491 -378 2845 -310
rect 2981 -356 3092 -270
rect -94 -419 -34 -412
rect -94 -453 -81 -419
rect -47 -453 -34 -419
rect -94 -497 -34 -453
rect -94 -531 -81 -497
rect -47 -531 -34 -497
rect -1715 -568 -1583 -555
rect -1715 -602 -1708 -568
rect -1674 -602 -1630 -568
rect -1596 -602 -1583 -568
rect -1715 -615 -1583 -602
rect -94 -634 -34 -531
rect 2618 -434 2678 -427
rect 2618 -468 2631 -434
rect 2665 -468 2678 -434
rect 2618 -512 2678 -468
rect 2618 -546 2631 -512
rect 2665 -546 2678 -512
rect 969 -570 1106 -557
rect 3 -652 141 -582
rect 633 -591 765 -578
rect 633 -625 640 -591
rect 674 -625 718 -591
rect 752 -625 765 -591
rect 969 -604 976 -570
rect 1010 -604 1054 -570
rect 1088 -604 1106 -570
rect 2618 -571 2678 -546
rect 2606 -576 2678 -571
rect 969 -617 1106 -604
rect 633 -638 765 -625
rect 2618 -633 2678 -576
rect 2714 -652 2841 -582
rect 3402 -615 3450 -199
rect 3 -781 65 -652
rect -123 -843 65 -781
rect 2714 -782 2760 -652
rect 2582 -831 2760 -782
rect 3491 -1000 3580 695
rect -205 -1068 268 -1000
rect 636 -1068 1109 -1000
rect 2478 -1068 3580 -1000
<< viali >>
rect -1887 285 -1853 319
rect -1887 207 -1853 241
rect 730 261 764 295
rect 845 286 879 320
rect 730 183 764 217
rect 845 208 879 242
rect -2244 18 -2210 52
rect -2166 18 -2132 52
rect 383 17 417 51
rect 461 17 495 51
rect 2987 21 3021 55
rect 3065 21 3099 55
rect -1934 -81 -1900 -47
rect -1856 -81 -1822 -47
rect 2589 -79 2623 -45
rect 2667 -79 2701 -45
rect 3404 -103 3438 -69
rect -130 -167 -96 -133
rect -52 -167 -18 -133
rect 811 -168 845 -134
rect 889 -168 923 -134
rect 3404 -181 3438 -147
rect -2257 -251 -2223 -217
rect -2179 -251 -2145 -217
rect 376 -251 410 -217
rect 454 -251 488 -217
rect 2973 -257 3007 -223
rect 3051 -257 3085 -223
rect -81 -453 -47 -419
rect -81 -531 -47 -497
rect -1708 -602 -1674 -568
rect -1630 -602 -1596 -568
rect 2631 -468 2665 -434
rect 2631 -546 2665 -512
rect 640 -625 674 -591
rect 718 -625 752 -591
rect 976 -604 1010 -570
rect 1054 -604 1088 -570
<< metal1 >>
rect -1900 319 -1840 326
rect -1900 285 -1887 319
rect -1853 285 -1840 319
rect -1900 241 -1840 285
rect -1900 207 -1887 241
rect -1853 207 -1840 241
rect -1900 194 -1840 207
rect -2251 52 -2114 65
rect -2251 18 -2244 52
rect -2210 18 -2166 52
rect -2132 18 -2114 52
rect -2251 5 -2114 18
rect -2244 -204 -2149 5
rect -1900 -34 -1842 194
rect -1941 -47 -1809 -34
rect -1941 -81 -1934 -47
rect -1900 -81 -1856 -47
rect -1822 -81 -1809 -47
rect -1941 -94 -1809 -81
rect -1759 -142 -1702 423
rect 832 320 892 327
rect 717 295 777 302
rect 717 261 730 295
rect 764 261 777 295
rect 717 217 777 261
rect 717 215 730 217
rect 716 183 730 215
rect 764 183 777 217
rect -832 -22 -790 90
rect -636 -22 -594 93
rect -441 -22 -399 89
rect -250 -22 -204 175
rect 716 170 777 183
rect 832 286 845 320
rect 879 286 892 320
rect 832 242 892 286
rect 832 208 845 242
rect 879 208 892 242
rect 376 51 513 64
rect 376 17 383 51
rect 417 17 461 51
rect 495 17 513 51
rect 376 4 513 17
rect -1968 -199 -1702 -142
rect -964 -68 -204 -22
rect -2264 -217 -2132 -204
rect -2264 -251 -2257 -217
rect -2223 -251 -2179 -217
rect -2145 -251 -2132 -217
rect -2264 -264 -2132 -251
rect -1968 -320 -1911 -199
rect -964 -234 -918 -68
rect -137 -133 -5 -120
rect -137 -167 -130 -133
rect -96 -167 -52 -133
rect -18 -167 -5 -133
rect -137 -180 -5 -167
rect -1729 -235 -918 -234
rect -2652 -377 -1911 -320
rect -1737 -280 -918 -235
rect -1737 -555 -1691 -280
rect -94 -419 -34 -180
rect 400 -204 495 4
rect 369 -217 506 -204
rect 369 -251 376 -217
rect 410 -251 454 -217
rect 488 -251 506 -217
rect 369 -264 506 -251
rect -94 -453 -81 -419
rect -47 -453 -34 -419
rect -94 -497 -34 -453
rect -94 -531 -81 -497
rect -47 -531 -34 -497
rect -94 -544 -34 -531
rect -1737 -568 -1583 -555
rect -1737 -602 -1708 -568
rect -1674 -602 -1630 -568
rect -1596 -602 -1583 -568
rect 716 -578 776 170
rect 832 -121 892 208
rect 1861 -24 1922 94
rect 2052 -24 2113 96
rect 2248 -24 2309 94
rect 2453 -24 2501 130
rect 2980 55 3112 68
rect 2980 21 2987 55
rect 3021 21 3065 55
rect 3099 21 3112 55
rect 2980 8 3112 21
rect 970 -72 2501 -24
rect 2582 -45 2714 -32
rect 804 -134 941 -121
rect 804 -168 811 -134
rect 845 -168 889 -134
rect 923 -168 941 -134
rect 804 -181 941 -168
rect 970 -557 1011 -72
rect 2582 -79 2589 -45
rect 2623 -79 2667 -45
rect 2701 -79 2714 -45
rect 2582 -92 2714 -79
rect 2618 -434 2678 -92
rect 2993 -210 3088 8
rect 3391 -69 3451 -62
rect 3391 -103 3404 -69
rect 3438 -88 3451 -69
rect 3438 -103 3660 -88
rect 3391 -147 3660 -103
rect 3391 -181 3404 -147
rect 3438 -152 3660 -147
rect 3438 -181 3451 -152
rect 3391 -199 3451 -181
rect 2966 -223 3103 -210
rect 2966 -257 2973 -223
rect 3007 -257 3051 -223
rect 3085 -257 3103 -223
rect 2966 -270 3103 -257
rect 2618 -468 2631 -434
rect 2665 -468 2678 -434
rect 2618 -512 2678 -468
rect 2618 -546 2631 -512
rect 2665 -546 2678 -512
rect -1737 -615 -1583 -602
rect 633 -591 776 -578
rect 633 -625 640 -591
rect 674 -625 718 -591
rect 752 -625 776 -591
rect 969 -570 1106 -557
rect 2618 -559 2678 -546
rect 969 -604 976 -570
rect 1010 -604 1054 -570
rect 1088 -604 1106 -570
rect 969 -617 1106 -604
rect 970 -618 1011 -617
rect 633 -638 776 -625
rect 716 -644 776 -638
use inverter  inverter_0
timestamp 1726359333
transform 1 0 -225 0 1 429
box 220 -453 904 367
use inverter  inverter_1
timestamp 1726359333
transform 1 0 -2850 0 1 429
box 220 -453 904 367
use inverter  inverter_2
timestamp 1726359333
transform -1 0 963 0 -1 -737
box 220 -453 904 367
use inverter  inverter_3
timestamp 1726359333
transform 1 0 2475 0 1 429
box 220 -453 904 367
use inverter  inverter_4
timestamp 1726359333
transform -1 0 3663 0 -1 -737
box 220 -453 904 367
use TG_MAGIC  TG_MAGIC_0
timestamp 1726359333
transform 1 0 -1727 0 1 -3
box -56 -27 1568 799
use TG_MAGIC  TG_MAGIC_1
timestamp 1726359333
transform -1 0 -115 0 -1 -305
box -56 -27 1568 799
use TG_MAGIC  TG_MAGIC_2
timestamp 1726359333
transform 1 0 973 0 1 -3
box -56 -27 1568 799
use TG_MAGIC  TG_MAGIC_3
timestamp 1726359333
transform -1 0 2585 0 -1 -305
box -56 -27 1568 799
<< labels >>
flabel locali s -40 730 -40 730 0 FreeSans 2443 0 0 0 VDD
flabel metal1 s 3621 -119 3621 -119 0 FreeSans 2443 0 0 0 Q
flabel metal1 s -2612 -356 -2612 -356 0 FreeSans 2443 0 0 0 D
flabel locali s -2587 -114 -2587 -114 0 FreeSans 2443 0 0 0 CLK
flabel locali s -1815 -241 -1815 -241 0 FreeSans 2443 0 0 0 VSS
<< end >>
