magic
tech sky130A
magscale 1 2
timestamp 1717685973
<< nwell >>
rect -223 -162 223 162
<< pmos >>
rect -129 -100 -29 100
rect 29 -100 129 100
<< pdiff >>
rect -187 85 -129 100
rect -187 51 -175 85
rect -141 51 -129 85
rect -187 17 -129 51
rect -187 -17 -175 17
rect -141 -17 -129 17
rect -187 -51 -129 -17
rect -187 -85 -175 -51
rect -141 -85 -129 -51
rect -187 -100 -129 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 129 85 187 100
rect 129 51 141 85
rect 175 51 187 85
rect 129 17 187 51
rect 129 -17 141 17
rect 175 -17 187 17
rect 129 -51 187 -17
rect 129 -85 141 -51
rect 175 -85 187 -51
rect 129 -100 187 -85
<< pdiffc >>
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
<< poly >>
rect -129 100 -29 126
rect 29 100 129 126
rect -129 -126 -29 -100
rect 29 -126 129 -100
<< locali >>
rect -175 85 -141 104
rect -175 17 -141 19
rect -175 -19 -141 -17
rect -175 -104 -141 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 141 85 175 104
rect 141 17 175 19
rect 141 -19 175 -17
rect 141 -104 175 -85
<< viali >>
rect -175 51 -141 53
rect -175 19 -141 51
rect -175 -51 -141 -19
rect -175 -53 -141 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 141 51 175 53
rect 141 19 175 51
rect 141 -51 175 -19
rect 141 -53 175 -51
<< metal1 >>
rect -181 53 -135 100
rect -181 19 -175 53
rect -141 19 -135 53
rect -181 -19 -135 19
rect -181 -53 -175 -19
rect -141 -53 -135 -19
rect -181 -100 -135 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 135 53 181 100
rect 135 19 141 53
rect 175 19 181 53
rect 135 -19 181 19
rect 135 -53 141 -19
rect 175 -53 181 -19
rect 135 -100 181 -53
<< properties >>
string GDS_END 39760
string GDS_FILE /home/shahid/Sky130Projects/top_layout/VCO.gds
string GDS_START 38092
<< end >>
