magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< pwell >>
rect -104 -176 104 176
<< nmos >>
rect -20 -150 20 150
<< ndiff >>
rect -78 119 -20 150
rect -78 85 -66 119
rect -32 85 -20 119
rect -78 51 -20 85
rect -78 17 -66 51
rect -32 17 -20 51
rect -78 -17 -20 17
rect -78 -51 -66 -17
rect -32 -51 -20 -17
rect -78 -85 -20 -51
rect -78 -119 -66 -85
rect -32 -119 -20 -85
rect -78 -150 -20 -119
rect 20 119 78 150
rect 20 85 32 119
rect 66 85 78 119
rect 20 51 78 85
rect 20 17 32 51
rect 66 17 78 51
rect 20 -17 78 17
rect 20 -51 32 -17
rect 66 -51 78 -17
rect 20 -85 78 -51
rect 20 -119 32 -85
rect 66 -119 78 -85
rect 20 -150 78 -119
<< ndiffc >>
rect -66 85 -32 119
rect -66 17 -32 51
rect -66 -51 -32 -17
rect -66 -119 -32 -85
rect 32 85 66 119
rect 32 17 66 51
rect 32 -51 66 -17
rect 32 -119 66 -85
<< poly >>
rect -20 150 20 176
rect -20 -176 20 -150
<< locali >>
rect -66 125 -32 154
rect -66 53 -32 85
rect -66 -17 -32 17
rect -66 -85 -32 -53
rect -66 -154 -32 -125
rect 32 125 66 154
rect 32 53 66 85
rect 32 -17 66 17
rect 32 -85 66 -53
rect 32 -154 66 -125
<< viali >>
rect -66 119 -32 125
rect -66 91 -32 119
rect -66 51 -32 53
rect -66 19 -32 51
rect -66 -51 -32 -19
rect -66 -53 -32 -51
rect -66 -119 -32 -91
rect -66 -125 -32 -119
rect 32 119 66 125
rect 32 91 66 119
rect 32 51 66 53
rect 32 19 66 51
rect 32 -51 66 -19
rect 32 -53 66 -51
rect 32 -119 66 -91
rect 32 -125 66 -119
<< metal1 >>
rect -72 125 -26 150
rect -72 91 -66 125
rect -32 91 -26 125
rect -72 53 -26 91
rect -72 19 -66 53
rect -32 19 -26 53
rect -72 -19 -26 19
rect -72 -53 -66 -19
rect -32 -53 -26 -19
rect -72 -91 -26 -53
rect -72 -125 -66 -91
rect -32 -125 -26 -91
rect -72 -150 -26 -125
rect 26 125 72 150
rect 26 91 32 125
rect 66 91 72 125
rect 26 53 72 91
rect 26 19 32 53
rect 66 19 72 53
rect 26 -19 72 19
rect 26 -53 32 -19
rect 66 -53 72 -19
rect 26 -91 72 -53
rect 26 -125 32 -91
rect 66 -125 72 -91
rect 26 -150 72 -125
<< end >>
