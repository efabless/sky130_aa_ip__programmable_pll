magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< pwell >>
rect -1771 -426 1771 426
<< nmos >>
rect -1687 -400 -887 400
rect -829 -400 -29 400
rect 29 -400 829 400
rect 887 -400 1687 400
<< ndiff >>
rect -1745 357 -1687 400
rect -1745 323 -1733 357
rect -1699 323 -1687 357
rect -1745 289 -1687 323
rect -1745 255 -1733 289
rect -1699 255 -1687 289
rect -1745 221 -1687 255
rect -1745 187 -1733 221
rect -1699 187 -1687 221
rect -1745 153 -1687 187
rect -1745 119 -1733 153
rect -1699 119 -1687 153
rect -1745 85 -1687 119
rect -1745 51 -1733 85
rect -1699 51 -1687 85
rect -1745 17 -1687 51
rect -1745 -17 -1733 17
rect -1699 -17 -1687 17
rect -1745 -51 -1687 -17
rect -1745 -85 -1733 -51
rect -1699 -85 -1687 -51
rect -1745 -119 -1687 -85
rect -1745 -153 -1733 -119
rect -1699 -153 -1687 -119
rect -1745 -187 -1687 -153
rect -1745 -221 -1733 -187
rect -1699 -221 -1687 -187
rect -1745 -255 -1687 -221
rect -1745 -289 -1733 -255
rect -1699 -289 -1687 -255
rect -1745 -323 -1687 -289
rect -1745 -357 -1733 -323
rect -1699 -357 -1687 -323
rect -1745 -400 -1687 -357
rect -887 357 -829 400
rect -887 323 -875 357
rect -841 323 -829 357
rect -887 289 -829 323
rect -887 255 -875 289
rect -841 255 -829 289
rect -887 221 -829 255
rect -887 187 -875 221
rect -841 187 -829 221
rect -887 153 -829 187
rect -887 119 -875 153
rect -841 119 -829 153
rect -887 85 -829 119
rect -887 51 -875 85
rect -841 51 -829 85
rect -887 17 -829 51
rect -887 -17 -875 17
rect -841 -17 -829 17
rect -887 -51 -829 -17
rect -887 -85 -875 -51
rect -841 -85 -829 -51
rect -887 -119 -829 -85
rect -887 -153 -875 -119
rect -841 -153 -829 -119
rect -887 -187 -829 -153
rect -887 -221 -875 -187
rect -841 -221 -829 -187
rect -887 -255 -829 -221
rect -887 -289 -875 -255
rect -841 -289 -829 -255
rect -887 -323 -829 -289
rect -887 -357 -875 -323
rect -841 -357 -829 -323
rect -887 -400 -829 -357
rect -29 357 29 400
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -400 29 -357
rect 829 357 887 400
rect 829 323 841 357
rect 875 323 887 357
rect 829 289 887 323
rect 829 255 841 289
rect 875 255 887 289
rect 829 221 887 255
rect 829 187 841 221
rect 875 187 887 221
rect 829 153 887 187
rect 829 119 841 153
rect 875 119 887 153
rect 829 85 887 119
rect 829 51 841 85
rect 875 51 887 85
rect 829 17 887 51
rect 829 -17 841 17
rect 875 -17 887 17
rect 829 -51 887 -17
rect 829 -85 841 -51
rect 875 -85 887 -51
rect 829 -119 887 -85
rect 829 -153 841 -119
rect 875 -153 887 -119
rect 829 -187 887 -153
rect 829 -221 841 -187
rect 875 -221 887 -187
rect 829 -255 887 -221
rect 829 -289 841 -255
rect 875 -289 887 -255
rect 829 -323 887 -289
rect 829 -357 841 -323
rect 875 -357 887 -323
rect 829 -400 887 -357
rect 1687 357 1745 400
rect 1687 323 1699 357
rect 1733 323 1745 357
rect 1687 289 1745 323
rect 1687 255 1699 289
rect 1733 255 1745 289
rect 1687 221 1745 255
rect 1687 187 1699 221
rect 1733 187 1745 221
rect 1687 153 1745 187
rect 1687 119 1699 153
rect 1733 119 1745 153
rect 1687 85 1745 119
rect 1687 51 1699 85
rect 1733 51 1745 85
rect 1687 17 1745 51
rect 1687 -17 1699 17
rect 1733 -17 1745 17
rect 1687 -51 1745 -17
rect 1687 -85 1699 -51
rect 1733 -85 1745 -51
rect 1687 -119 1745 -85
rect 1687 -153 1699 -119
rect 1733 -153 1745 -119
rect 1687 -187 1745 -153
rect 1687 -221 1699 -187
rect 1733 -221 1745 -187
rect 1687 -255 1745 -221
rect 1687 -289 1699 -255
rect 1733 -289 1745 -255
rect 1687 -323 1745 -289
rect 1687 -357 1699 -323
rect 1733 -357 1745 -323
rect 1687 -400 1745 -357
<< ndiffc >>
rect -1733 323 -1699 357
rect -1733 255 -1699 289
rect -1733 187 -1699 221
rect -1733 119 -1699 153
rect -1733 51 -1699 85
rect -1733 -17 -1699 17
rect -1733 -85 -1699 -51
rect -1733 -153 -1699 -119
rect -1733 -221 -1699 -187
rect -1733 -289 -1699 -255
rect -1733 -357 -1699 -323
rect -875 323 -841 357
rect -875 255 -841 289
rect -875 187 -841 221
rect -875 119 -841 153
rect -875 51 -841 85
rect -875 -17 -841 17
rect -875 -85 -841 -51
rect -875 -153 -841 -119
rect -875 -221 -841 -187
rect -875 -289 -841 -255
rect -875 -357 -841 -323
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect 841 323 875 357
rect 841 255 875 289
rect 841 187 875 221
rect 841 119 875 153
rect 841 51 875 85
rect 841 -17 875 17
rect 841 -85 875 -51
rect 841 -153 875 -119
rect 841 -221 875 -187
rect 841 -289 875 -255
rect 841 -357 875 -323
rect 1699 323 1733 357
rect 1699 255 1733 289
rect 1699 187 1733 221
rect 1699 119 1733 153
rect 1699 51 1733 85
rect 1699 -17 1733 17
rect 1699 -85 1733 -51
rect 1699 -153 1733 -119
rect 1699 -221 1733 -187
rect 1699 -289 1733 -255
rect 1699 -357 1733 -323
<< poly >>
rect -1687 400 -887 426
rect -829 400 -29 426
rect 29 400 829 426
rect 887 400 1687 426
rect -1687 -426 -887 -400
rect -829 -426 -29 -400
rect 29 -426 829 -400
rect 887 -426 1687 -400
<< locali >>
rect -1733 377 -1699 404
rect -1733 305 -1699 323
rect -1733 233 -1699 255
rect -1733 161 -1699 187
rect -1733 89 -1699 119
rect -1733 17 -1699 51
rect -1733 -51 -1699 -17
rect -1733 -119 -1699 -89
rect -1733 -187 -1699 -161
rect -1733 -255 -1699 -233
rect -1733 -323 -1699 -305
rect -1733 -404 -1699 -377
rect -875 377 -841 404
rect -875 305 -841 323
rect -875 233 -841 255
rect -875 161 -841 187
rect -875 89 -841 119
rect -875 17 -841 51
rect -875 -51 -841 -17
rect -875 -119 -841 -89
rect -875 -187 -841 -161
rect -875 -255 -841 -233
rect -875 -323 -841 -305
rect -875 -404 -841 -377
rect -17 377 17 404
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -404 17 -377
rect 841 377 875 404
rect 841 305 875 323
rect 841 233 875 255
rect 841 161 875 187
rect 841 89 875 119
rect 841 17 875 51
rect 841 -51 875 -17
rect 841 -119 875 -89
rect 841 -187 875 -161
rect 841 -255 875 -233
rect 841 -323 875 -305
rect 841 -404 875 -377
rect 1699 377 1733 404
rect 1699 305 1733 323
rect 1699 233 1733 255
rect 1699 161 1733 187
rect 1699 89 1733 119
rect 1699 17 1733 51
rect 1699 -51 1733 -17
rect 1699 -119 1733 -89
rect 1699 -187 1733 -161
rect 1699 -255 1733 -233
rect 1699 -323 1733 -305
rect 1699 -404 1733 -377
<< viali >>
rect -1733 357 -1699 377
rect -1733 343 -1699 357
rect -1733 289 -1699 305
rect -1733 271 -1699 289
rect -1733 221 -1699 233
rect -1733 199 -1699 221
rect -1733 153 -1699 161
rect -1733 127 -1699 153
rect -1733 85 -1699 89
rect -1733 55 -1699 85
rect -1733 -17 -1699 17
rect -1733 -85 -1699 -55
rect -1733 -89 -1699 -85
rect -1733 -153 -1699 -127
rect -1733 -161 -1699 -153
rect -1733 -221 -1699 -199
rect -1733 -233 -1699 -221
rect -1733 -289 -1699 -271
rect -1733 -305 -1699 -289
rect -1733 -357 -1699 -343
rect -1733 -377 -1699 -357
rect -875 357 -841 377
rect -875 343 -841 357
rect -875 289 -841 305
rect -875 271 -841 289
rect -875 221 -841 233
rect -875 199 -841 221
rect -875 153 -841 161
rect -875 127 -841 153
rect -875 85 -841 89
rect -875 55 -841 85
rect -875 -17 -841 17
rect -875 -85 -841 -55
rect -875 -89 -841 -85
rect -875 -153 -841 -127
rect -875 -161 -841 -153
rect -875 -221 -841 -199
rect -875 -233 -841 -221
rect -875 -289 -841 -271
rect -875 -305 -841 -289
rect -875 -357 -841 -343
rect -875 -377 -841 -357
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect 841 357 875 377
rect 841 343 875 357
rect 841 289 875 305
rect 841 271 875 289
rect 841 221 875 233
rect 841 199 875 221
rect 841 153 875 161
rect 841 127 875 153
rect 841 85 875 89
rect 841 55 875 85
rect 841 -17 875 17
rect 841 -85 875 -55
rect 841 -89 875 -85
rect 841 -153 875 -127
rect 841 -161 875 -153
rect 841 -221 875 -199
rect 841 -233 875 -221
rect 841 -289 875 -271
rect 841 -305 875 -289
rect 841 -357 875 -343
rect 841 -377 875 -357
rect 1699 357 1733 377
rect 1699 343 1733 357
rect 1699 289 1733 305
rect 1699 271 1733 289
rect 1699 221 1733 233
rect 1699 199 1733 221
rect 1699 153 1733 161
rect 1699 127 1733 153
rect 1699 85 1733 89
rect 1699 55 1733 85
rect 1699 -17 1733 17
rect 1699 -85 1733 -55
rect 1699 -89 1733 -85
rect 1699 -153 1733 -127
rect 1699 -161 1733 -153
rect 1699 -221 1733 -199
rect 1699 -233 1733 -221
rect 1699 -289 1733 -271
rect 1699 -305 1733 -289
rect 1699 -357 1733 -343
rect 1699 -377 1733 -357
<< metal1 >>
rect -1739 377 -1693 400
rect -1739 343 -1733 377
rect -1699 343 -1693 377
rect -1739 305 -1693 343
rect -1739 271 -1733 305
rect -1699 271 -1693 305
rect -1739 233 -1693 271
rect -1739 199 -1733 233
rect -1699 199 -1693 233
rect -1739 161 -1693 199
rect -1739 127 -1733 161
rect -1699 127 -1693 161
rect -1739 89 -1693 127
rect -1739 55 -1733 89
rect -1699 55 -1693 89
rect -1739 17 -1693 55
rect -1739 -17 -1733 17
rect -1699 -17 -1693 17
rect -1739 -55 -1693 -17
rect -1739 -89 -1733 -55
rect -1699 -89 -1693 -55
rect -1739 -127 -1693 -89
rect -1739 -161 -1733 -127
rect -1699 -161 -1693 -127
rect -1739 -199 -1693 -161
rect -1739 -233 -1733 -199
rect -1699 -233 -1693 -199
rect -1739 -271 -1693 -233
rect -1739 -305 -1733 -271
rect -1699 -305 -1693 -271
rect -1739 -343 -1693 -305
rect -1739 -377 -1733 -343
rect -1699 -377 -1693 -343
rect -1739 -400 -1693 -377
rect -881 377 -835 400
rect -881 343 -875 377
rect -841 343 -835 377
rect -881 305 -835 343
rect -881 271 -875 305
rect -841 271 -835 305
rect -881 233 -835 271
rect -881 199 -875 233
rect -841 199 -835 233
rect -881 161 -835 199
rect -881 127 -875 161
rect -841 127 -835 161
rect -881 89 -835 127
rect -881 55 -875 89
rect -841 55 -835 89
rect -881 17 -835 55
rect -881 -17 -875 17
rect -841 -17 -835 17
rect -881 -55 -835 -17
rect -881 -89 -875 -55
rect -841 -89 -835 -55
rect -881 -127 -835 -89
rect -881 -161 -875 -127
rect -841 -161 -835 -127
rect -881 -199 -835 -161
rect -881 -233 -875 -199
rect -841 -233 -835 -199
rect -881 -271 -835 -233
rect -881 -305 -875 -271
rect -841 -305 -835 -271
rect -881 -343 -835 -305
rect -881 -377 -875 -343
rect -841 -377 -835 -343
rect -881 -400 -835 -377
rect -23 377 23 400
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -400 23 -377
rect 835 377 881 400
rect 835 343 841 377
rect 875 343 881 377
rect 835 305 881 343
rect 835 271 841 305
rect 875 271 881 305
rect 835 233 881 271
rect 835 199 841 233
rect 875 199 881 233
rect 835 161 881 199
rect 835 127 841 161
rect 875 127 881 161
rect 835 89 881 127
rect 835 55 841 89
rect 875 55 881 89
rect 835 17 881 55
rect 835 -17 841 17
rect 875 -17 881 17
rect 835 -55 881 -17
rect 835 -89 841 -55
rect 875 -89 881 -55
rect 835 -127 881 -89
rect 835 -161 841 -127
rect 875 -161 881 -127
rect 835 -199 881 -161
rect 835 -233 841 -199
rect 875 -233 881 -199
rect 835 -271 881 -233
rect 835 -305 841 -271
rect 875 -305 881 -271
rect 835 -343 881 -305
rect 835 -377 841 -343
rect 875 -377 881 -343
rect 835 -400 881 -377
rect 1693 377 1739 400
rect 1693 343 1699 377
rect 1733 343 1739 377
rect 1693 305 1739 343
rect 1693 271 1699 305
rect 1733 271 1739 305
rect 1693 233 1739 271
rect 1693 199 1699 233
rect 1733 199 1739 233
rect 1693 161 1739 199
rect 1693 127 1699 161
rect 1733 127 1739 161
rect 1693 89 1739 127
rect 1693 55 1699 89
rect 1733 55 1739 89
rect 1693 17 1739 55
rect 1693 -17 1699 17
rect 1733 -17 1739 17
rect 1693 -55 1739 -17
rect 1693 -89 1699 -55
rect 1733 -89 1739 -55
rect 1693 -127 1739 -89
rect 1693 -161 1699 -127
rect 1733 -161 1739 -127
rect 1693 -199 1739 -161
rect 1693 -233 1699 -199
rect 1733 -233 1739 -199
rect 1693 -271 1739 -233
rect 1693 -305 1699 -271
rect 1733 -305 1739 -271
rect 1693 -343 1739 -305
rect 1693 -377 1699 -343
rect 1733 -377 1739 -343
rect 1693 -400 1739 -377
<< end >>
