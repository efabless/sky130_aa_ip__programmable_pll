magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect 0 458 1425 459
rect 0 324 1456 458
rect 0 302 1425 324
rect 259 0 1425 302
<< pwell >>
rect 22 -929 1348 -812
<< psubdiff >>
rect 48 -854 1322 -838
rect 48 -888 106 -854
rect 140 -888 174 -854
rect 208 -888 306 -854
rect 340 -888 374 -854
rect 408 -888 506 -854
rect 540 -888 574 -854
rect 608 -888 706 -854
rect 740 -888 774 -854
rect 808 -888 906 -854
rect 940 -888 974 -854
rect 1008 -888 1106 -854
rect 1140 -888 1174 -854
rect 1208 -888 1322 -854
rect 48 -903 1322 -888
<< nsubdiff >>
rect 53 405 669 423
rect 53 371 104 405
rect 138 371 172 405
rect 206 371 240 405
rect 274 371 308 405
rect 342 371 376 405
rect 410 371 444 405
rect 478 371 512 405
rect 546 371 580 405
rect 614 371 669 405
rect 53 354 669 371
rect 1173 403 1418 417
rect 1173 369 1237 403
rect 1271 369 1305 403
rect 1339 369 1418 403
rect 1173 350 1418 369
<< psubdiffcont >>
rect 106 -888 140 -854
rect 174 -888 208 -854
rect 306 -888 340 -854
rect 374 -888 408 -854
rect 506 -888 540 -854
rect 574 -888 608 -854
rect 706 -888 740 -854
rect 774 -888 808 -854
rect 906 -888 940 -854
rect 974 -888 1008 -854
rect 1106 -888 1140 -854
rect 1174 -888 1208 -854
<< nsubdiffcont >>
rect 104 371 138 405
rect 172 371 206 405
rect 240 371 274 405
rect 308 371 342 405
rect 376 371 410 405
rect 444 371 478 405
rect 512 371 546 405
rect 580 371 614 405
rect 1237 369 1271 403
rect 1305 369 1339 403
<< poly >>
rect 94 19 134 41
rect -29 9 134 19
rect -29 -25 -13 9
rect 21 -25 56 9
rect 90 -25 134 9
rect -29 -35 134 -25
rect 94 -259 134 -35
rect 192 -259 232 41
rect 290 -18 330 36
rect 388 -18 428 36
rect 486 -3 624 36
rect 290 -49 444 -18
rect 307 -73 444 -49
rect 307 -107 323 -73
rect 357 -107 392 -73
rect 426 -107 444 -73
rect 307 -117 444 -107
rect 94 -299 232 -259
rect 94 -321 134 -299
rect 192 -321 232 -299
rect 404 -289 444 -117
rect 583 -141 624 -3
rect 1224 -8 1362 37
rect 495 -151 630 -141
rect 1224 -143 1264 -8
rect 495 -185 511 -151
rect 545 -185 580 -151
rect 614 -185 630 -151
rect 495 -186 630 -185
rect 1106 -153 1264 -143
rect 495 -195 753 -186
rect 583 -226 753 -195
rect 1106 -187 1122 -153
rect 1156 -187 1191 -153
rect 1225 -187 1264 -153
rect 1106 -197 1264 -187
rect 713 -281 753 -226
rect 404 -320 542 -289
rect 713 -320 851 -281
rect 404 -329 444 -320
rect 713 -324 753 -320
rect 1224 -427 1264 -197
<< polycont >>
rect -13 -25 21 9
rect 56 -25 90 9
rect 323 -107 357 -73
rect 392 -107 426 -73
rect 511 -185 545 -151
rect 580 -185 614 -151
rect 1122 -187 1156 -153
rect 1191 -187 1225 -153
<< locali >>
rect 48 405 669 423
rect 48 371 104 405
rect 138 371 172 405
rect 206 371 240 405
rect 274 371 308 405
rect 342 371 376 405
rect 410 371 444 405
rect 478 371 512 405
rect 546 371 580 405
rect 614 383 669 405
rect 1173 403 1418 417
rect 614 371 670 383
rect 48 354 670 371
rect 48 266 82 354
rect 244 266 278 354
rect 440 266 474 354
rect 636 266 670 354
rect 1173 369 1237 403
rect 1271 369 1305 403
rect 1339 369 1418 403
rect 1173 350 1418 369
rect 1178 266 1212 350
rect 1374 266 1408 350
rect 146 22 180 58
rect 342 22 376 60
rect 538 22 572 58
rect -29 11 106 19
rect -48 9 106 11
rect -48 -25 -13 9
rect 21 -25 56 9
rect 90 -25 106 9
rect 146 -15 701 22
rect -48 -26 106 -25
rect -29 -35 106 -26
rect 307 -72 442 -63
rect -48 -73 442 -72
rect -48 -107 323 -73
rect 357 -107 392 -73
rect 426 -107 442 -73
rect -48 -110 442 -107
rect 307 -117 442 -110
rect 495 -151 630 -141
rect 495 -154 511 -151
rect -46 -185 511 -154
rect 545 -185 580 -151
rect 614 -185 630 -151
rect -46 -188 630 -185
rect 495 -195 630 -188
rect 664 -153 701 -15
rect 1106 -153 1241 -143
rect 664 -187 1122 -153
rect 1156 -187 1191 -153
rect 1225 -187 1241 -153
rect 664 -190 1241 -187
rect 664 -244 701 -190
rect 1106 -197 1241 -190
rect 48 -278 491 -244
rect 664 -278 897 -244
rect 48 -341 82 -278
rect 244 -279 491 -278
rect 244 -341 278 -279
rect 456 -342 491 -279
rect 667 -342 701 -278
rect 863 -342 897 -278
rect 1276 -458 1310 62
rect 146 -838 180 -647
rect 358 -745 393 -641
rect 554 -745 589 -639
rect 358 -748 589 -745
rect 765 -748 799 -646
rect 358 -782 799 -748
rect 1178 -838 1212 -637
rect 48 -854 1322 -838
rect 48 -888 106 -854
rect 140 -888 174 -854
rect 208 -888 306 -854
rect 340 -888 374 -854
rect 408 -888 506 -854
rect 540 -888 574 -854
rect 608 -888 706 -854
rect 740 -888 774 -854
rect 808 -888 906 -854
rect 940 -888 974 -854
rect 1008 -888 1106 -854
rect 1140 -888 1174 -854
rect 1208 -888 1322 -854
rect 48 -903 1322 -888
use sky130_fd_pr__nfet_01v8_FQGQPX  sky130_fd_pr__nfet_01v8_FQGQPX_0
timestamp 1717691374
transform 1 0 212 0 1 -495
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPX  sky130_fd_pr__nfet_01v8_FQGQPX_1
timestamp 1717691374
transform 1 0 114 0 1 -495
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPX  sky130_fd_pr__nfet_01v8_FQGQPX_2
timestamp 1717691374
transform 1 0 424 0 1 -496
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPX  sky130_fd_pr__nfet_01v8_FQGQPX_3
timestamp 1717691374
transform 1 0 522 0 1 -496
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPX  sky130_fd_pr__nfet_01v8_FQGQPX_4
timestamp 1717691374
transform 1 0 733 0 1 -496
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPX  sky130_fd_pr__nfet_01v8_FQGQPX_6
timestamp 1717691374
transform 1 0 831 0 1 -496
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_NUEGCF  sky130_fd_pr__nfet_01v8_NUEGCF_0
timestamp 1717691374
transform 1 0 1244 0 1 -546
box -104 -126 104 126
use sky130_fd_pr__pfet_01v8_ES6JQB  sky130_fd_pr__pfet_01v8_ES6JQB_0
timestamp 1717691374
transform 1 0 1342 0 1 162
box -114 -162 114 162
use sky130_fd_pr__pfet_01v8_ES6JQB  sky130_fd_pr__pfet_01v8_ES6JQB_1
timestamp 1717691374
transform 1 0 114 0 1 162
box -114 -162 114 162
use sky130_fd_pr__pfet_01v8_ES6JQB  sky130_fd_pr__pfet_01v8_ES6JQB_2
timestamp 1717691374
transform 1 0 212 0 1 162
box -114 -162 114 162
use sky130_fd_pr__pfet_01v8_ES6JQB  sky130_fd_pr__pfet_01v8_ES6JQB_3
timestamp 1717691374
transform 1 0 310 0 1 162
box -114 -162 114 162
use sky130_fd_pr__pfet_01v8_ES6JQB  sky130_fd_pr__pfet_01v8_ES6JQB_5
timestamp 1717691374
transform 1 0 506 0 1 162
box -114 -162 114 162
use sky130_fd_pr__pfet_01v8_ES6JQB  sky130_fd_pr__pfet_01v8_ES6JQB_6
timestamp 1717691374
transform 1 0 604 0 1 162
box -114 -162 114 162
use sky130_fd_pr__pfet_01v8_ES6JQB  sky130_fd_pr__pfet_01v8_ES6JQB_7
timestamp 1717691374
transform 1 0 1244 0 1 162
box -114 -162 114 162
use sky130_fd_pr__pfet_01v8_ES6JQB  sky130_fd_pr__pfet_01v8_ES6JQB_8
timestamp 1717691374
transform 1 0 408 0 1 162
box -114 -162 114 162
<< labels >>
flabel locali s 317 406 317 406 0 FreeSans 1250 0 0 0 VDD
flabel locali s 259 -893 259 -893 0 FreeSans 1250 0 0 0 VSS
flabel locali s -42 -7 -42 -7 0 FreeSans 750 0 0 0 C
flabel locali s -44 -91 -44 -91 0 FreeSans 750 0 0 0 B
flabel locali s -38 -170 -38 -170 0 FreeSans 750 0 0 0 A
flabel locali s 1305 -178 1305 -178 0 FreeSans 750 0 0 0 VOUT
<< end >>
