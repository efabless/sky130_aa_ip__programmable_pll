magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect -336 464 1539 500
rect 1757 464 1848 500
rect -336 371 1712 464
rect -336 369 1576 371
rect 1720 370 1886 464
rect -336 294 1539 369
rect -336 83 0 294
rect 136 236 170 294
rect 182 291 477 294
rect 204 276 476 291
rect 211 269 476 276
rect 212 258 476 269
rect 312 236 346 258
rect 488 221 554 294
rect 488 220 522 221
rect -336 48 -231 83
rect -119 48 0 83
rect 595 81 657 86
rect 859 80 880 294
rect 1041 269 1539 294
rect 1107 146 1539 269
rect 1041 109 1101 146
rect 1106 109 1539 146
rect 969 86 1029 87
rect 765 79 888 80
rect 946 79 1029 86
rect 765 76 1029 79
rect 804 75 1029 76
rect 804 74 1008 75
rect 1025 74 1029 75
rect 1101 74 1106 87
rect 741 59 789 68
rect 804 62 1029 74
rect 1107 67 1539 109
rect 1107 62 1655 67
rect 804 48 1655 62
rect 1757 48 1848 370
rect 804 4 1008 48
<< pwell >>
rect -348 -315 -95 -294
rect 1516 -315 2078 -215
rect -374 -329 240 -315
rect 622 -329 2078 -315
rect -374 -462 2078 -329
<< psubdiff >>
rect -322 -341 -121 -320
rect 1542 -341 2052 -241
rect -348 -355 214 -341
rect 648 -355 2052 -341
rect -348 -372 2052 -355
rect -348 -406 -313 -372
rect -279 -406 -221 -372
rect -187 -406 -129 -372
rect -95 -406 -37 -372
rect -3 -406 55 -372
rect 89 -406 147 -372
rect 181 -406 239 -372
rect 273 -406 331 -372
rect 365 -406 423 -372
rect 457 -406 515 -372
rect 549 -406 607 -372
rect 641 -406 699 -372
rect 733 -406 791 -372
rect 825 -406 883 -372
rect 917 -406 975 -372
rect 1009 -406 1067 -372
rect 1101 -406 1157 -372
rect 1191 -406 1295 -372
rect 1329 -406 1422 -372
rect 1456 -406 1571 -372
rect 1605 -406 1663 -372
rect 1697 -406 1755 -372
rect 1789 -406 1847 -372
rect 1881 -406 1939 -372
rect 1973 -406 2052 -372
rect -348 -436 2052 -406
<< nsubdiff >>
rect -155 435 47 464
rect -155 401 -109 435
rect -75 401 -17 435
rect 17 401 47 435
rect -155 374 47 401
rect 597 441 1712 464
rect 1720 441 1886 464
rect 597 436 1886 441
rect 597 435 1193 436
rect 597 401 627 435
rect 661 401 719 435
rect 753 401 811 435
rect 845 401 903 435
rect 937 401 995 435
rect 1029 401 1087 435
rect 1121 402 1193 435
rect 1227 402 1261 436
rect 1295 402 1329 436
rect 1363 402 1397 436
rect 1431 435 1886 436
rect 1431 402 1499 435
rect 1121 401 1499 402
rect 1533 401 1707 435
rect 1741 401 1799 435
rect 1833 401 1886 435
rect 597 395 1886 401
rect 597 374 1712 395
rect -155 370 -119 374
rect 1539 371 1712 374
rect 1539 370 1576 371
rect 1720 370 1886 395
<< psubdiffcont >>
rect -313 -406 -279 -372
rect -221 -406 -187 -372
rect -129 -406 -95 -372
rect -37 -406 -3 -372
rect 55 -406 89 -372
rect 147 -406 181 -372
rect 239 -406 273 -372
rect 331 -406 365 -372
rect 423 -406 457 -372
rect 515 -406 549 -372
rect 607 -406 641 -372
rect 699 -406 733 -372
rect 791 -406 825 -372
rect 883 -406 917 -372
rect 975 -406 1009 -372
rect 1067 -406 1101 -372
rect 1157 -406 1191 -372
rect 1295 -406 1329 -372
rect 1422 -406 1456 -372
rect 1571 -406 1605 -372
rect 1663 -406 1697 -372
rect 1755 -406 1789 -372
rect 1847 -406 1881 -372
rect 1939 -406 1973 -372
<< nsubdiffcont >>
rect -109 401 -75 435
rect -17 401 17 435
rect 627 401 661 435
rect 719 401 753 435
rect 811 401 845 435
rect 903 401 937 435
rect 995 401 1029 435
rect 1087 401 1121 435
rect 1193 402 1227 436
rect 1261 402 1295 436
rect 1329 402 1363 436
rect 1397 402 1431 436
rect 1499 401 1533 435
rect 1707 401 1741 435
rect 1799 401 1833 435
<< poly >>
rect 182 333 476 367
rect 182 332 398 333
rect 182 298 221 332
rect 255 299 398 332
rect 432 299 476 333
rect 255 298 476 299
rect 182 258 476 298
rect 182 257 212 258
rect 657 86 677 96
rect 94 43 124 86
rect 94 10 300 43
rect 240 -33 300 10
rect 358 -33 388 86
rect 518 59 678 86
rect 735 78 765 87
rect 518 57 622 59
rect 518 23 540 57
rect 574 25 622 57
rect 656 25 678 59
rect 574 23 678 25
rect 518 7 678 23
rect 648 -39 678 7
rect 722 76 765 78
rect 969 77 1106 87
rect 722 56 804 76
rect 722 22 748 56
rect 782 22 804 56
rect 722 6 804 22
rect 941 59 1106 77
rect 941 25 968 59
rect 1002 25 1048 59
rect 1082 25 1106 59
rect 941 9 1106 25
rect -18 -235 64 -203
rect 446 -205 476 -204
rect -18 -269 5 -235
rect 39 -269 64 -235
rect -18 -291 64 -269
rect 112 -235 191 -205
rect 112 -269 135 -235
rect 169 -269 191 -235
rect 112 -290 191 -269
rect 240 -249 300 -205
rect 446 -238 531 -205
rect 446 -249 475 -238
rect 240 -272 475 -249
rect 509 -272 531 -238
rect 648 -242 766 -200
rect 240 -291 531 -272
rect 683 -246 766 -242
rect 683 -280 709 -246
rect 743 -280 766 -246
rect 683 -302 766 -280
rect 938 -248 1376 -217
rect 938 -282 981 -248
rect 1015 -249 1376 -248
rect 1015 -282 1088 -249
rect 938 -283 1088 -282
rect 1122 -250 1376 -249
rect 1122 -283 1210 -250
rect 938 -284 1210 -283
rect 1244 -284 1376 -250
rect 938 -307 1376 -284
<< polycont >>
rect 221 298 255 332
rect 398 299 432 333
rect 540 23 574 57
rect 622 25 656 59
rect 748 22 782 56
rect 968 25 1002 59
rect 1048 25 1082 59
rect 5 -269 39 -235
rect 135 -269 169 -235
rect 475 -272 509 -238
rect 709 -280 743 -246
rect 981 -282 1015 -248
rect 1088 -283 1122 -249
rect 1210 -284 1244 -250
<< locali >>
rect -118 488 1539 500
rect 1757 488 1848 500
rect -118 464 2047 488
rect -155 436 2047 464
rect -155 435 1193 436
rect -155 401 -109 435
rect -75 401 -17 435
rect 17 401 627 435
rect 661 401 719 435
rect 753 401 811 435
rect 845 401 903 435
rect 937 401 995 435
rect 1029 401 1087 435
rect 1121 402 1193 435
rect 1227 402 1261 436
rect 1295 402 1329 436
rect 1363 402 1397 436
rect 1431 435 2047 436
rect 1431 402 1499 435
rect 1121 401 1499 402
rect 1533 401 1707 435
rect 1741 401 1799 435
rect 1833 401 2047 435
rect -155 392 2047 401
rect -155 370 170 392
rect -118 355 170 370
rect 136 236 170 355
rect 204 337 276 357
rect 204 332 222 337
rect 204 298 221 332
rect 256 303 276 337
rect 255 298 276 303
rect 204 276 276 298
rect 312 236 346 392
rect 381 338 453 358
rect 381 333 399 338
rect 381 299 398 333
rect 433 304 453 338
rect 432 299 453 304
rect 381 277 453 299
rect 488 355 2047 392
rect 488 221 522 355
rect 777 296 811 355
rect 923 296 957 355
rect 1757 340 1848 355
rect 1041 269 1186 306
rect 1152 146 1186 269
rect 224 47 258 109
rect 400 47 434 110
rect 601 74 635 120
rect 1041 109 1186 146
rect 518 59 678 74
rect 518 57 622 59
rect 518 47 540 57
rect -448 8 -334 47
rect -177 23 540 47
rect 574 25 622 57
rect 656 25 678 59
rect 574 23 678 25
rect -444 -497 -405 8
rect -177 -1 678 23
rect 722 57 804 74
rect 722 22 748 57
rect 782 22 804 57
rect 945 59 1106 74
rect 945 42 968 59
rect 722 8 804 22
rect 846 25 968 42
rect 1002 25 1048 59
rect 1082 25 1106 59
rect 846 7 1106 25
rect 488 -56 522 -1
rect -18 -235 62 -217
rect -18 -238 5 -235
rect -18 -272 4 -238
rect 39 -269 62 -235
rect 38 -272 62 -269
rect -18 -291 62 -272
rect 113 -233 191 -217
rect 113 -235 136 -233
rect 113 -269 135 -235
rect 170 -267 191 -233
rect 169 -269 191 -267
rect 113 -290 191 -269
rect -322 -341 -121 -320
rect 312 -341 346 -183
rect 453 -238 531 -217
rect 453 -276 475 -238
rect 509 -276 531 -238
rect 453 -291 531 -276
rect 602 -341 636 -183
rect 687 -242 766 -223
rect 846 -242 881 7
rect 945 -26 1106 7
rect 1152 40 1186 109
rect 1152 6 1525 40
rect 2080 8 2335 47
rect 1152 -67 1186 6
rect 1388 -67 1422 6
rect 1708 -1 1810 8
rect 687 -246 881 -242
rect 687 -280 709 -246
rect 743 -280 881 -246
rect 687 -284 881 -280
rect 939 -248 1372 -229
rect 1587 -241 1621 -152
rect 1896 -241 1930 -160
rect 939 -250 981 -248
rect 1015 -249 1372 -248
rect 939 -284 962 -250
rect 1015 -282 1088 -249
rect 1122 -250 1372 -249
rect 1122 -252 1210 -250
rect 996 -283 1088 -282
rect 996 -284 1091 -283
rect 687 -303 766 -284
rect 939 -286 1091 -284
rect 1125 -284 1210 -252
rect 1244 -253 1372 -250
rect 1125 -286 1213 -284
rect 939 -287 1213 -286
rect 1247 -287 1372 -253
rect 939 -307 1372 -287
rect 1542 -341 2052 -241
rect -348 -372 2052 -341
rect -348 -406 -313 -372
rect -279 -406 -221 -372
rect -187 -406 -129 -372
rect -95 -406 -37 -372
rect -3 -406 55 -372
rect 89 -406 147 -372
rect 181 -406 239 -372
rect 273 -406 331 -372
rect 365 -406 423 -372
rect 457 -406 515 -372
rect 549 -406 607 -372
rect 641 -406 699 -372
rect 733 -406 791 -372
rect 825 -406 883 -372
rect 917 -406 975 -372
rect 1009 -406 1067 -372
rect 1101 -406 1157 -372
rect 1191 -406 1295 -372
rect 1329 -406 1422 -372
rect 1456 -406 1571 -372
rect 1605 -406 1663 -372
rect 1697 -406 1755 -372
rect 1789 -406 1847 -372
rect 1881 -406 1939 -372
rect 1973 -406 2052 -372
rect -348 -436 2052 -406
rect -175 -497 62 -470
rect -444 -531 -124 -497
rect -90 -531 -13 -497
rect 21 -531 62 -497
rect -444 -536 62 -531
rect -175 -566 62 -536
rect 121 -503 1099 -474
rect 121 -505 1040 -503
rect 121 -507 941 -505
rect 121 -541 142 -507
rect 176 -541 245 -507
rect 279 -539 941 -507
rect 975 -537 1040 -505
rect 1074 -537 1099 -503
rect 975 -539 1099 -537
rect 279 -541 1099 -539
rect 121 -570 1099 -541
<< viali >>
rect 222 332 256 337
rect 222 303 255 332
rect 255 303 256 332
rect 399 333 433 338
rect 399 304 432 333
rect 432 304 433 333
rect 748 56 782 57
rect 748 23 782 56
rect 4 -269 5 -238
rect 5 -269 38 -238
rect 4 -272 38 -269
rect 136 -235 170 -233
rect 136 -267 169 -235
rect 169 -267 170 -235
rect 475 -272 509 -242
rect 475 -276 509 -272
rect 962 -282 981 -250
rect 981 -282 996 -250
rect 962 -284 996 -282
rect 1091 -283 1122 -252
rect 1122 -283 1125 -252
rect 1091 -286 1125 -283
rect 1213 -284 1244 -253
rect 1244 -284 1247 -253
rect 1213 -287 1247 -284
rect -124 -531 -90 -497
rect -13 -531 21 -497
rect 142 -541 176 -507
rect 245 -541 279 -507
rect 941 -539 975 -505
rect 1040 -537 1074 -503
<< metal1 >>
rect 207 357 273 360
rect 384 358 450 361
rect 204 352 276 357
rect 381 352 453 358
rect 42 338 453 352
rect 42 337 399 338
rect 42 306 222 337
rect 42 231 88 306
rect 204 303 222 306
rect 256 306 399 337
rect 256 303 276 306
rect 204 276 276 303
rect 381 304 399 306
rect 433 304 453 338
rect 381 277 453 304
rect 42 62 88 113
rect -48 16 88 62
rect 725 57 820 74
rect 1035 72 1081 113
rect 725 23 748 57
rect 782 23 820 57
rect -48 -67 -2 16
rect 725 6 820 23
rect 910 26 1081 72
rect 910 -71 956 26
rect 1028 -39 1936 -3
rect 1028 -72 1074 -39
rect 1264 -71 1310 -39
rect 805 -103 919 -79
rect 805 -150 924 -103
rect -43 -238 62 -208
rect -43 -272 4 -238
rect 38 -272 62 -238
rect -43 -470 62 -272
rect -175 -497 62 -470
rect -175 -531 -124 -497
rect -90 -531 -13 -497
rect 21 -531 62 -497
rect -175 -566 62 -531
rect 108 -233 199 -214
rect 108 -267 136 -233
rect 170 -267 199 -233
rect 108 -474 199 -267
rect 438 -242 544 -208
rect 438 -276 475 -242
rect 509 -276 544 -242
rect 108 -507 344 -474
rect 108 -541 142 -507
rect 176 -541 245 -507
rect 279 -541 344 -507
rect 108 -570 344 -541
rect 438 -610 544 -276
rect 939 -250 1372 -229
rect 939 -284 962 -250
rect 996 -252 1372 -250
rect 996 -284 1091 -252
rect 939 -286 1091 -284
rect 1125 -253 1372 -252
rect 1125 -286 1213 -253
rect 939 -287 1213 -286
rect 1247 -287 1372 -253
rect 939 -307 1372 -287
rect 1008 -474 1099 -307
rect 1478 -425 1514 -39
rect 1890 -70 1936 -39
rect 1478 -461 1929 -425
rect 910 -503 1099 -474
rect 910 -505 1040 -503
rect 910 -539 941 -505
rect 975 -537 1040 -505
rect 1074 -537 1099 -503
rect 975 -539 1099 -537
rect 910 -570 1099 -539
use PFD_INV  PFD_INV_0
timestamp 1717691374
transform -1 0 -118 0 1 48
box -65 -394 271 452
use PFD_INV  PFD_INV_1
timestamp 1717691374
transform 1 0 1848 0 1 48
box -65 -394 271 452
use PFD_INV  PFD_INV_2
timestamp 1717691374
transform 1 0 1539 0 1 48
box -65 -394 271 452
use sky130_fd_pr__nfet_01v8_FB3UY2  sky130_fd_pr__nfet_01v8_FB3UY2_0
timestamp 1717691374
transform 1 0 461 0 1 -119
box -99 -86 99 86
use sky130_fd_pr__nfet_01v8_FB3UY2  sky130_fd_pr__nfet_01v8_FB3UY2_1
timestamp 1717691374
transform 1 0 373 0 1 -119
box -99 -86 99 86
use sky130_fd_pr__nfet_01v8_FB3UY2  sky130_fd_pr__nfet_01v8_FB3UY2_2
timestamp 1717691374
transform 1 0 751 0 1 -124
box -99 -86 99 86
use sky130_fd_pr__nfet_01v8_FB3UY2  sky130_fd_pr__nfet_01v8_FB3UY2_3
timestamp 1717691374
transform 1 0 663 0 1 -124
box -99 -86 99 86
use sky130_fd_pr__nfet_01v8_R2UA5N  sky130_fd_pr__nfet_01v8_R2UA5N_0
timestamp 1717691374
transform 1 0 270 0 1 -119
box -114 -86 114 86
use sky130_fd_pr__nfet_01v8_R2UA5N  sky130_fd_pr__nfet_01v8_R2UA5N_1
timestamp 1717691374
transform 1 0 34 0 1 -119
box -114 -86 114 86
use sky130_fd_pr__nfet_01v8_R2UA5N  sky130_fd_pr__nfet_01v8_R2UA5N_2
timestamp 1717691374
transform 1 0 152 0 1 -119
box -114 -86 114 86
use sky130_fd_pr__nfet_01v8_R2UA5N  sky130_fd_pr__nfet_01v8_R2UA5N_3
timestamp 1717691374
transform 1 0 1110 0 1 -131
box -114 -86 114 86
use sky130_fd_pr__nfet_01v8_R2UA5N  sky130_fd_pr__nfet_01v8_R2UA5N_4
timestamp 1717691374
transform 1 0 992 0 1 -131
box -114 -86 114 86
use sky130_fd_pr__nfet_01v8_R2UA5N  sky130_fd_pr__nfet_01v8_R2UA5N_5
timestamp 1717691374
transform 1 0 1228 0 1 -131
box -114 -86 114 86
use sky130_fd_pr__nfet_01v8_R2UA5N  sky130_fd_pr__nfet_01v8_R2UA5N_6
timestamp 1717691374
transform 1 0 1346 0 1 -131
box -114 -86 114 86
use sky130_fd_pr__pfet_01v8_5AY9XA  sky130_fd_pr__pfet_01v8_5AY9XA_1
timestamp 1717691374
transform 1 0 662 0 1 202
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AY9XA  sky130_fd_pr__pfet_01v8_5AY9XA_2
timestamp 1717691374
transform 1 0 750 0 1 202
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_58P8XA  sky130_fd_pr__pfet_01v8_58P8XA_1
timestamp 1717691374
transform 1 0 109 0 1 172
box -109 -122 109 122
use sky130_fd_pr__pfet_01v8_58P8XA  sky130_fd_pr__pfet_01v8_58P8XA_2
timestamp 1717691374
transform 1 0 197 0 1 172
box -109 -122 109 122
use sky130_fd_pr__pfet_01v8_58P8XA  sky130_fd_pr__pfet_01v8_58P8XA_3
timestamp 1717691374
transform 1 0 285 0 1 172
box -109 -122 109 122
use sky130_fd_pr__pfet_01v8_58P8XA  sky130_fd_pr__pfet_01v8_58P8XA_4
timestamp 1717691374
transform 1 0 373 0 1 172
box -109 -122 109 122
use sky130_fd_pr__pfet_01v8_58P8XA  sky130_fd_pr__pfet_01v8_58P8XA_5
timestamp 1717691374
transform 1 0 461 0 1 172
box -109 -122 109 122
use sky130_fd_pr__pfet_01v8_EP25JC  sky130_fd_pr__pfet_01v8_EP25JC_0
timestamp 1717691374
transform 1 0 999 0 1 202
box -124 -152 124 152
<< end >>
