magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< pwell >>
rect -8109 4481 13970 4728
rect -8109 -228 -7862 4481
rect 13723 -228 13970 4481
rect -8109 -475 13970 -228
<< psubdiff >>
rect -8083 4649 13944 4702
rect -8083 4547 -7779 4649
rect 13675 4547 13944 4649
rect -8083 4507 13944 4547
rect -8083 4426 -7888 4507
rect -8083 -164 -8031 4426
rect -7929 -164 -7888 4426
rect -8083 -254 -7888 -164
rect 13749 4414 13944 4507
rect 13749 -176 13798 4414
rect 13900 -176 13944 4414
rect 13749 -254 13944 -176
rect -8083 -303 13944 -254
rect -8083 -405 -7783 -303
rect 13603 -405 13944 -303
rect -8083 -449 13944 -405
<< psubdiffcont >>
rect -7779 4547 13675 4649
rect -8031 -164 -7929 4426
rect 13798 -176 13900 4414
rect -7783 -405 13603 -303
<< locali >>
rect -8117 4753 -7298 4754
rect -8117 4649 13984 4753
rect -8117 4547 -7779 4649
rect 13675 4547 13984 4649
rect -8117 4459 13984 4547
rect -8117 4426 -7822 4459
rect -7401 4458 13984 4459
rect -8117 -164 -8031 4426
rect -7929 -164 -7822 4426
rect -5865 3275 -5676 3833
rect -391 3664 15 4458
rect 13689 4414 13984 4458
rect -2082 3615 1395 3664
rect -2082 3539 1396 3615
rect 2639 3523 3127 3616
rect 4360 3523 5248 3619
rect 5184 3382 5248 3523
rect 5090 3364 5282 3382
rect 5090 3330 5109 3364
rect 5143 3330 5228 3364
rect 5262 3330 5282 3364
rect 5090 3276 5282 3330
rect -6652 3206 -6102 3248
rect 5090 3242 5108 3276
rect 5142 3242 5227 3276
rect 5261 3242 5282 3276
rect -6652 3172 -6371 3206
rect -6337 3172 -6162 3206
rect -6128 3172 -6102 3206
rect -6652 3120 -6102 3172
rect -5899 3192 -5738 3215
rect -5899 3158 -5889 3192
rect -5855 3191 -5738 3192
rect -5855 3158 -5798 3191
rect -5899 3157 -5798 3158
rect -5764 3184 -5738 3191
rect -1043 3185 -878 3208
rect -5764 3157 -5684 3184
rect -5899 3154 -5684 3157
rect -5899 3136 -5643 3154
rect -5777 3115 -5643 3136
rect -1043 3151 -1033 3185
rect -999 3184 -878 3185
rect -999 3151 -942 3184
rect -1043 3150 -942 3151
rect -908 3150 -878 3184
rect -1043 3147 -878 3150
rect 5090 3183 5282 3242
rect 5090 3149 5112 3183
rect 5146 3149 5231 3183
rect 5265 3149 5282 3183
rect -1043 3128 -788 3147
rect -948 3108 -788 3128
rect 5090 3124 5282 3149
rect -4048 2897 -3541 2979
rect 844 2919 1189 3001
rect 4739 2970 4931 2988
rect 4739 2936 4758 2970
rect 4792 2936 4877 2970
rect 4911 2936 4931 2970
rect -4048 2734 -3966 2897
rect -2073 2869 -1699 2903
rect -7412 2051 -7220 2069
rect -7412 2017 -7393 2051
rect -7359 2017 -7274 2051
rect -7240 2017 -7220 2051
rect -7412 1963 -7220 2017
rect -7412 1929 -7394 1963
rect -7360 1929 -7275 1963
rect -7241 1929 -6558 1963
rect -7412 1898 -6558 1929
rect -1760 1915 -1699 2869
rect 844 2737 926 2919
rect 2688 2891 2938 2925
rect 4739 2917 4931 2936
rect 5463 2917 5555 3162
rect 4739 2882 5555 2917
rect 4409 2848 4757 2882
rect 4791 2848 4876 2882
rect 4910 2848 5555 2882
rect 4739 2825 5555 2848
rect 4739 2789 4931 2825
rect 4739 2755 4761 2789
rect 4795 2755 4880 2789
rect 4914 2755 4931 2789
rect 4739 2730 4931 2755
rect 12925 2743 13130 2813
rect 1375 1945 1409 2306
rect 1691 1949 1725 2301
rect 2007 1926 2041 2337
rect 2323 1908 2357 2335
rect 2658 2310 3115 2338
rect 2639 2274 3115 2310
rect 2639 1986 2673 2274
rect 4359 2217 6408 2301
rect 13002 2204 13174 2270
rect 2639 1923 3111 1986
rect 2654 1922 3111 1923
rect -7412 1870 -7220 1898
rect -7412 1836 -7390 1870
rect -7356 1836 -7271 1870
rect -7237 1836 -7220 1870
rect -7412 1811 -7220 1836
rect -7449 1503 -7257 1521
rect -7449 1469 -7430 1503
rect -7396 1469 -7311 1503
rect -7277 1469 -7257 1503
rect -7449 1415 -7257 1469
rect -4284 1468 -3893 1550
rect 4761 1522 4953 1540
rect -7449 1381 -7431 1415
rect -7397 1381 -7312 1415
rect -7278 1381 -7257 1415
rect -7449 1342 -7257 1381
rect -7449 1322 -6560 1342
rect -7449 1288 -7427 1322
rect -7393 1288 -7308 1322
rect -7274 1301 -6560 1322
rect -3975 1333 -3893 1468
rect 579 1440 926 1522
rect -2035 1335 -1973 1361
rect 844 1356 926 1440
rect 4761 1488 4780 1522
rect 4814 1488 4899 1522
rect 4933 1488 4953 1522
rect 4761 1458 4953 1488
rect 4761 1434 4967 1458
rect 4761 1427 4779 1434
rect 4396 1400 4779 1427
rect 4813 1400 4898 1434
rect 4932 1400 4967 1434
rect 4396 1393 4967 1400
rect -7274 1288 -7257 1301
rect -7449 1263 -7257 1288
rect -3975 1251 -3515 1333
rect -2035 1294 -1653 1335
rect -1531 1294 -1522 1335
rect 844 1274 1227 1356
rect 2688 1350 2952 1384
rect 4761 1355 4967 1393
rect 4761 1341 4953 1355
rect 4761 1307 4783 1341
rect 4817 1307 4902 1341
rect 4936 1307 4953 1341
rect 4761 1282 4953 1307
rect -6702 906 -6386 937
rect -6805 883 -6386 906
rect -6805 849 -6672 883
rect -6638 849 -6463 883
rect -6429 849 -6386 883
rect -6805 826 -6386 849
rect -6085 883 -5923 906
rect -6085 849 -6075 883
rect -6041 882 -5923 883
rect -6041 849 -5984 882
rect -6085 848 -5984 849
rect -5950 848 -5923 882
rect -6085 826 -5923 848
rect -1229 880 -1067 903
rect -1229 846 -1219 880
rect -1185 879 -1067 880
rect -1185 846 -1128 879
rect -1229 845 -1128 846
rect -1094 845 -1067 879
rect -6702 809 -6386 826
rect -1229 823 -1067 845
rect -8117 -180 -7822 -164
rect -6153 -180 -5964 764
rect -4107 742 -3341 793
rect -4107 684 -3332 742
rect -2093 702 -1191 758
rect -2096 668 -1191 702
rect 730 715 812 777
rect 730 681 1409 715
rect 2639 710 3127 765
rect 13689 -176 13798 4414
rect 13900 -176 13984 4414
rect 13689 -180 13984 -176
rect -8117 -303 13984 -180
rect -8117 -405 -7783 -303
rect 13603 -405 13984 -303
rect -8117 -475 13984 -405
<< viali >>
rect 5109 3330 5143 3364
rect 5228 3330 5262 3364
rect 5108 3242 5142 3276
rect 5227 3242 5261 3276
rect -6371 3172 -6337 3206
rect -6162 3172 -6128 3206
rect -5889 3158 -5855 3192
rect -5798 3157 -5764 3191
rect -1033 3151 -999 3185
rect -942 3150 -908 3184
rect 5112 3149 5146 3183
rect 5231 3149 5265 3183
rect 4758 2936 4792 2970
rect 4877 2936 4911 2970
rect -7393 2017 -7359 2051
rect -7274 2017 -7240 2051
rect -7394 1929 -7360 1963
rect -7275 1929 -7241 1963
rect 4757 2848 4791 2882
rect 4876 2848 4910 2882
rect 4761 2755 4795 2789
rect 4880 2755 4914 2789
rect -7390 1836 -7356 1870
rect -7271 1836 -7237 1870
rect -7430 1469 -7396 1503
rect -7311 1469 -7277 1503
rect -7431 1381 -7397 1415
rect -7312 1381 -7278 1415
rect -7427 1288 -7393 1322
rect -7308 1288 -7274 1322
rect 4780 1488 4814 1522
rect 4899 1488 4933 1522
rect 4779 1400 4813 1434
rect 4898 1400 4932 1434
rect 4783 1307 4817 1341
rect 4902 1307 4936 1341
rect -6672 849 -6638 883
rect -6463 849 -6429 883
rect -6075 849 -6041 883
rect -5984 848 -5950 882
rect -1219 846 -1185 880
rect -1128 845 -1094 879
<< metal1 >>
rect -7366 3992 4900 4128
rect -7366 2069 -7230 3992
rect -6089 3546 -1579 3627
rect -6089 3253 -6008 3546
rect -6418 3206 -6008 3253
rect -6418 3172 -6371 3206
rect -6337 3172 -6162 3206
rect -6128 3201 -6008 3206
rect -5899 3201 -5738 3215
rect -6128 3192 -5738 3201
rect -6128 3172 -5889 3192
rect -6418 3158 -5889 3172
rect -5855 3191 -5738 3192
rect -5855 3158 -5798 3191
rect -6418 3157 -5798 3158
rect -5764 3157 -5738 3191
rect -6418 3146 -5738 3157
rect -6418 3120 -6038 3146
rect -5899 3136 -5738 3146
rect -1660 3208 -1579 3546
rect -1660 3185 -881 3208
rect -1660 3151 -1033 3185
rect -999 3184 -881 3185
rect -999 3151 -942 3184
rect -1660 3150 -942 3151
rect -908 3150 -881 3184
rect -1660 3128 -881 3150
rect -1660 3127 -1010 3128
rect 4764 2988 4900 3992
rect 5115 3382 5251 3383
rect 5090 3364 5282 3382
rect 5090 3330 5109 3364
rect 5143 3330 5228 3364
rect 5262 3330 5282 3364
rect 5090 3276 5282 3330
rect 5090 3242 5108 3276
rect 5142 3242 5227 3276
rect 5261 3263 5282 3276
rect 5261 3242 5865 3263
rect 5090 3183 5865 3242
rect 5090 3149 5112 3183
rect 5146 3149 5231 3183
rect 5265 3168 5865 3183
rect 5265 3149 5282 3168
rect 11610 3153 11611 3217
rect 5090 3124 5282 3149
rect 4739 2970 4931 2988
rect 4739 2936 4758 2970
rect 4792 2936 4877 2970
rect 4911 2936 4931 2970
rect 4739 2882 4931 2936
rect 4739 2848 4757 2882
rect 4791 2848 4876 2882
rect 4910 2848 4931 2882
rect 860 2768 906 2816
rect -4221 2692 -3561 2738
rect 665 2722 906 2768
rect 4739 2789 4931 2848
rect 4739 2755 4761 2789
rect 4795 2755 4880 2789
rect 4914 2755 4931 2789
rect 4739 2730 4931 2755
rect -4221 2656 -4175 2692
rect -3607 2386 -3561 2692
rect -3366 2386 -3320 2431
rect -3607 2340 -3320 2386
rect -2102 2392 -2056 2433
rect -1120 2392 -1074 2440
rect -2102 2346 -1074 2392
rect -7412 2051 -7220 2069
rect -7412 2017 -7393 2051
rect -7359 2017 -7274 2051
rect -7240 2017 -7220 2051
rect -7412 1963 -7220 2017
rect -7412 1929 -7394 1963
rect -7360 1929 -7275 1963
rect -7241 1929 -7220 1963
rect -7412 1870 -7220 1929
rect 860 1945 906 2722
rect 860 1899 1415 1945
rect -7412 1836 -7390 1870
rect -7356 1836 -7271 1870
rect -7237 1836 -7220 1870
rect 1369 1838 1415 1899
rect -7412 1811 -7220 1836
rect 4761 1522 4953 1540
rect -7449 1503 -7257 1521
rect -7449 1469 -7430 1503
rect -7396 1469 -7311 1503
rect -7277 1469 -7257 1503
rect -7449 1415 -7257 1469
rect -7449 1381 -7431 1415
rect -7397 1381 -7312 1415
rect -7278 1381 -7257 1415
rect -7449 1322 -7257 1381
rect -7449 1288 -7427 1322
rect -7393 1288 -7308 1322
rect -7274 1288 -7257 1322
rect -7449 1263 -7257 1288
rect 4761 1488 4780 1522
rect 4814 1488 4899 1522
rect 4933 1488 4953 1522
rect 4761 1434 4953 1488
rect 4761 1400 4779 1434
rect 4813 1400 4898 1434
rect 4932 1400 4953 1434
rect 4761 1341 4953 1400
rect 4761 1307 4783 1341
rect 4817 1307 4902 1341
rect 4936 1307 4953 1341
rect 4761 1282 4953 1307
rect -7411 355 -7275 1263
rect -6702 906 -6386 937
rect -6702 883 -5923 906
rect -6702 849 -6672 883
rect -6638 849 -6463 883
rect -6429 849 -6075 883
rect -6041 882 -5923 883
rect -6041 849 -5984 882
rect -6702 848 -5984 849
rect -5950 848 -5923 882
rect -6702 826 -5923 848
rect -1824 880 -1067 903
rect -1824 846 -1219 880
rect -1185 879 -1067 880
rect -1185 846 -1128 879
rect -1824 845 -1128 846
rect -1094 845 -1067 879
rect -6702 809 -6386 826
rect -6300 669 -6220 826
rect -1824 823 -1067 845
rect -1824 669 -1744 823
rect -6300 589 -1744 669
rect 4791 355 4927 1282
rect -7411 219 4927 355
use DelayCell_1  DelayCell_1_0
timestamp 1726359333
transform 1 0 -774 0 1 2763
box -994 -2079 1786 587
use DelayCell_1  DelayCell_1_1
timestamp 1726359333
transform 1 0 -5629 0 1 2770
box -994 -2079 1786 587
use Divide_By_2_magic  Divide_By_2_magic_0
timestamp 1726359333
transform 1 0 8014 0 1 3305
box -2665 -1159 5054 829
use INV_1_mag  INV_1_mag_0
timestamp 1726359333
transform 1 0 1327 0 1 1376
box -142 -903 1395 763
use INV_1_mag  INV_1_mag_1
timestamp 1726359333
transform 1 0 3048 0 1 1419
box -142 -903 1395 763
use INV_1_mag  INV_1_mag_2
timestamp 1726359333
transform 1 0 -3408 0 -1 2877
box -142 -903 1395 763
use INV_1_mag  INV_1_mag_3
timestamp 1726359333
transform 1 0 -3408 0 1 1353
box -142 -903 1395 763
use INV_1_mag  INV_1_mag_4
timestamp 1726359333
transform 1 0 3048 0 -1 2856
box -142 -903 1395 763
use INV_1_mag  INV_1_mag_5
timestamp 1726359333
transform 1 0 1327 0 -1 2899
box -142 -903 1395 763
<< labels >>
flabel locali s -6585 3183 -6585 3183 0 FreeSans 1250 0 0 0 VCTRL
flabel locali s -6763 859 -6763 859 0 FreeSans 1250 0 0 0 VCTRL2
flabel locali s -5786 3775 -5786 3775 0 FreeSans 1250 0 0 0 VDD
flabel locali s -6062 415 -6062 415 0 FreeSans 1250 0 0 0 VSS
flabel locali s 13144 2239 13144 2239 0 FreeSans 1250 0 0 0 OUT
flabel locali s 13087 2777 13087 2777 0 FreeSans 1250 0 0 0 OUTB
<< end >>
