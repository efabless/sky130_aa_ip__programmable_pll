magic
tech sky130A
magscale 1 2
timestamp 1717685973
<< nwell >>
rect 0 521 1394 763
rect 364 466 398 521
rect 680 463 714 521
rect 996 464 1030 521
rect 1312 464 1346 521
rect 838 36 872 61
rect 1154 36 1188 62
rect 94 0 1300 36
<< pwell >>
rect -3 -903 1385 -726
<< psubdiff >>
rect 23 -798 1359 -752
rect 23 -832 56 -798
rect 90 -832 124 -798
rect 158 -832 192 -798
rect 226 -832 260 -798
rect 294 -832 328 -798
rect 362 -832 396 -798
rect 430 -832 464 -798
rect 498 -832 532 -798
rect 566 -832 600 -798
rect 634 -832 668 -798
rect 702 -832 736 -798
rect 770 -832 804 -798
rect 838 -832 872 -798
rect 906 -832 940 -798
rect 974 -832 1008 -798
rect 1042 -832 1076 -798
rect 1110 -832 1144 -798
rect 1178 -832 1212 -798
rect 1246 -832 1280 -798
rect 1314 -832 1359 -798
rect 23 -877 1359 -832
<< nsubdiff >>
rect 39 686 1346 723
rect 39 652 84 686
rect 118 652 152 686
rect 186 652 220 686
rect 254 652 288 686
rect 322 652 356 686
rect 390 652 424 686
rect 458 652 492 686
rect 526 652 560 686
rect 594 652 628 686
rect 662 652 696 686
rect 730 652 764 686
rect 798 652 832 686
rect 866 652 900 686
rect 934 652 968 686
rect 1002 652 1036 686
rect 1070 652 1104 686
rect 1138 652 1172 686
rect 1206 652 1240 686
rect 1274 652 1346 686
rect 39 616 1346 652
<< psubdiffcont >>
rect 56 -832 90 -798
rect 124 -832 158 -798
rect 192 -832 226 -798
rect 260 -832 294 -798
rect 328 -832 362 -798
rect 396 -832 430 -798
rect 464 -832 498 -798
rect 532 -832 566 -798
rect 600 -832 634 -798
rect 668 -832 702 -798
rect 736 -832 770 -798
rect 804 -832 838 -798
rect 872 -832 906 -798
rect 940 -832 974 -798
rect 1008 -832 1042 -798
rect 1076 -832 1110 -798
rect 1144 -832 1178 -798
rect 1212 -832 1246 -798
rect 1280 -832 1314 -798
<< nsubdiffcont >>
rect 84 652 118 686
rect 152 652 186 686
rect 220 652 254 686
rect 288 652 322 686
rect 356 652 390 686
rect 424 652 458 686
rect 492 652 526 686
rect 560 652 594 686
rect 628 652 662 686
rect 696 652 730 686
rect 764 652 798 686
rect 832 652 866 686
rect 900 652 934 686
rect 968 652 1002 686
rect 1036 652 1070 686
rect 1104 652 1138 686
rect 1172 652 1206 686
rect 1240 652 1274 686
<< poly >>
rect 94 61 120 62
rect 94 36 194 61
rect 252 36 352 64
rect 410 36 510 65
rect 568 36 668 65
rect 94 0 1300 36
rect 94 -20 194 0
rect -93 -46 194 -20
rect -93 -48 85 -46
rect -93 -82 -65 -48
rect -31 -80 85 -48
rect 119 -80 194 -46
rect -31 -82 194 -80
rect -93 -102 194 -82
rect 94 -173 194 -102
rect 252 -170 352 0
rect 410 -169 510 0
rect 568 -169 668 0
rect 887 -109 1290 -85
rect 887 -111 1229 -109
rect 887 -113 1065 -111
rect 887 -138 915 -113
rect 726 -147 915 -138
rect 949 -145 1065 -113
rect 1099 -143 1229 -111
rect 1263 -138 1290 -109
rect 1263 -143 1300 -138
rect 1099 -145 1300 -143
rect 949 -147 1300 -145
rect 726 -168 1300 -147
rect 94 -183 120 -173
<< polycont >>
rect -65 -82 -31 -48
rect 85 -80 119 -46
rect 915 -147 949 -113
rect 1065 -145 1099 -111
rect 1229 -143 1263 -109
<< locali >>
rect 39 686 1346 723
rect 39 652 84 686
rect 118 652 152 686
rect 186 652 220 686
rect 254 652 288 686
rect 322 652 356 686
rect 390 652 424 686
rect 458 652 492 686
rect 526 652 560 686
rect 594 652 628 686
rect 662 652 696 686
rect 730 652 764 686
rect 798 652 832 686
rect 866 652 900 686
rect 934 652 968 686
rect 1002 652 1036 686
rect 1070 652 1104 686
rect 1138 652 1172 686
rect 1206 652 1240 686
rect 1274 652 1346 686
rect 39 616 1346 652
rect 48 465 82 616
rect 364 466 398 616
rect 680 463 714 616
rect 996 464 1030 616
rect 1312 464 1346 616
rect -142 -46 155 -20
rect -142 -48 85 -46
rect -142 -82 -65 -48
rect -31 -80 85 -48
rect 119 -80 155 -46
rect -31 -82 155 -80
rect -142 -102 155 -82
rect 206 -80 240 71
rect 522 8 556 64
rect 838 8 872 61
rect 1154 8 1188 62
rect 522 -26 1395 8
rect 522 -80 556 -26
rect 206 -114 556 -80
rect 206 -202 240 -114
rect 522 -198 556 -114
rect 887 -109 1290 -85
rect 887 -111 1229 -109
rect 887 -113 1065 -111
rect 887 -138 915 -113
rect 838 -147 915 -138
rect 949 -145 1065 -113
rect 1099 -143 1229 -111
rect 1263 -138 1290 -109
rect 1263 -143 1346 -138
rect 1099 -145 1346 -143
rect 949 -147 1346 -145
rect 838 -172 1346 -147
rect 838 -200 872 -172
rect 996 -191 1030 -172
rect 1154 -206 1188 -172
rect 1312 -208 1346 -172
rect 48 -752 82 -597
rect 364 -752 398 -597
rect 680 -752 714 -597
rect 996 -752 1030 -597
rect 1312 -752 1346 -597
rect 23 -798 1359 -752
rect 23 -832 56 -798
rect 90 -832 124 -798
rect 158 -832 192 -798
rect 226 -832 260 -798
rect 294 -832 328 -798
rect 362 -832 396 -798
rect 430 -832 464 -798
rect 498 -832 532 -798
rect 566 -832 600 -798
rect 634 -832 668 -798
rect 702 -832 736 -798
rect 770 -832 804 -798
rect 838 -832 872 -798
rect 906 -832 940 -798
rect 974 -832 1008 -798
rect 1042 -832 1076 -798
rect 1110 -832 1144 -798
rect 1178 -832 1212 -798
rect 1246 -832 1280 -798
rect 1314 -832 1359 -798
rect 23 -877 1359 -832
use sky130_fd_pr__nfet_01v8_TMD3M2  sky130_fd_pr__nfet_01v8_TMD3M2_0
timestamp 1717685973
transform -1 0 1013 0 1 -394
box -371 -226 371 226
use sky130_fd_pr__nfet_01v8_TMD3M2  sky130_fd_pr__nfet_01v8_TMD3M2_1
timestamp 1717685973
transform 1 0 381 0 1 -394
box -371 -226 371 226
use sky130_fd_pr__pfet_01v8_2P97UG  sky130_fd_pr__pfet_01v8_2P97UG_0
timestamp 1717685973
transform -1 0 697 0 1 262
box -697 -262 697 262
<< labels >>
flabel locali s -123 -66 -123 -66 0 FreeSans 1250 0 0 0 IN
flabel locali s 1381 -11 1381 -11 0 FreeSans 1250 0 0 0 OUT
flabel locali s 696 708 696 708 0 FreeSans 1250 0 0 0 VDD
flabel locali s 679 -853 679 -853 0 FreeSans 1250 0 0 0 VSS
<< properties >>
string GDS_END 88274
string GDS_FILE /home/shahid/Sky130Projects/top_layout/VCO.gds
string GDS_START 81158
<< end >>
