magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< pwell >>
rect -484 -426 484 426
<< nmos >>
rect -400 -400 400 400
<< ndiff >>
rect -458 357 -400 400
rect -458 323 -446 357
rect -412 323 -400 357
rect -458 289 -400 323
rect -458 255 -446 289
rect -412 255 -400 289
rect -458 221 -400 255
rect -458 187 -446 221
rect -412 187 -400 221
rect -458 153 -400 187
rect -458 119 -446 153
rect -412 119 -400 153
rect -458 85 -400 119
rect -458 51 -446 85
rect -412 51 -400 85
rect -458 17 -400 51
rect -458 -17 -446 17
rect -412 -17 -400 17
rect -458 -51 -400 -17
rect -458 -85 -446 -51
rect -412 -85 -400 -51
rect -458 -119 -400 -85
rect -458 -153 -446 -119
rect -412 -153 -400 -119
rect -458 -187 -400 -153
rect -458 -221 -446 -187
rect -412 -221 -400 -187
rect -458 -255 -400 -221
rect -458 -289 -446 -255
rect -412 -289 -400 -255
rect -458 -323 -400 -289
rect -458 -357 -446 -323
rect -412 -357 -400 -323
rect -458 -400 -400 -357
rect 400 357 458 400
rect 400 323 412 357
rect 446 323 458 357
rect 400 289 458 323
rect 400 255 412 289
rect 446 255 458 289
rect 400 221 458 255
rect 400 187 412 221
rect 446 187 458 221
rect 400 153 458 187
rect 400 119 412 153
rect 446 119 458 153
rect 400 85 458 119
rect 400 51 412 85
rect 446 51 458 85
rect 400 17 458 51
rect 400 -17 412 17
rect 446 -17 458 17
rect 400 -51 458 -17
rect 400 -85 412 -51
rect 446 -85 458 -51
rect 400 -119 458 -85
rect 400 -153 412 -119
rect 446 -153 458 -119
rect 400 -187 458 -153
rect 400 -221 412 -187
rect 446 -221 458 -187
rect 400 -255 458 -221
rect 400 -289 412 -255
rect 446 -289 458 -255
rect 400 -323 458 -289
rect 400 -357 412 -323
rect 446 -357 458 -323
rect 400 -400 458 -357
<< ndiffc >>
rect -446 323 -412 357
rect -446 255 -412 289
rect -446 187 -412 221
rect -446 119 -412 153
rect -446 51 -412 85
rect -446 -17 -412 17
rect -446 -85 -412 -51
rect -446 -153 -412 -119
rect -446 -221 -412 -187
rect -446 -289 -412 -255
rect -446 -357 -412 -323
rect 412 323 446 357
rect 412 255 446 289
rect 412 187 446 221
rect 412 119 446 153
rect 412 51 446 85
rect 412 -17 446 17
rect 412 -85 446 -51
rect 412 -153 446 -119
rect 412 -221 446 -187
rect 412 -289 446 -255
rect 412 -357 446 -323
<< poly >>
rect -400 400 400 426
rect -400 -426 400 -400
<< locali >>
rect -446 377 -412 404
rect -446 305 -412 323
rect -446 233 -412 255
rect -446 161 -412 187
rect -446 89 -412 119
rect -446 17 -412 51
rect -446 -51 -412 -17
rect -446 -119 -412 -89
rect -446 -187 -412 -161
rect -446 -255 -412 -233
rect -446 -323 -412 -305
rect -446 -404 -412 -377
rect 412 377 446 404
rect 412 305 446 323
rect 412 233 446 255
rect 412 161 446 187
rect 412 89 446 119
rect 412 17 446 51
rect 412 -51 446 -17
rect 412 -119 446 -89
rect 412 -187 446 -161
rect 412 -255 446 -233
rect 412 -323 446 -305
rect 412 -404 446 -377
<< viali >>
rect -446 357 -412 377
rect -446 343 -412 357
rect -446 289 -412 305
rect -446 271 -412 289
rect -446 221 -412 233
rect -446 199 -412 221
rect -446 153 -412 161
rect -446 127 -412 153
rect -446 85 -412 89
rect -446 55 -412 85
rect -446 -17 -412 17
rect -446 -85 -412 -55
rect -446 -89 -412 -85
rect -446 -153 -412 -127
rect -446 -161 -412 -153
rect -446 -221 -412 -199
rect -446 -233 -412 -221
rect -446 -289 -412 -271
rect -446 -305 -412 -289
rect -446 -357 -412 -343
rect -446 -377 -412 -357
rect 412 357 446 377
rect 412 343 446 357
rect 412 289 446 305
rect 412 271 446 289
rect 412 221 446 233
rect 412 199 446 221
rect 412 153 446 161
rect 412 127 446 153
rect 412 85 446 89
rect 412 55 446 85
rect 412 -17 446 17
rect 412 -85 446 -55
rect 412 -89 446 -85
rect 412 -153 446 -127
rect 412 -161 446 -153
rect 412 -221 446 -199
rect 412 -233 446 -221
rect 412 -289 446 -271
rect 412 -305 446 -289
rect 412 -357 446 -343
rect 412 -377 446 -357
<< metal1 >>
rect -452 377 -406 400
rect -452 343 -446 377
rect -412 343 -406 377
rect -452 305 -406 343
rect -452 271 -446 305
rect -412 271 -406 305
rect -452 233 -406 271
rect -452 199 -446 233
rect -412 199 -406 233
rect -452 161 -406 199
rect -452 127 -446 161
rect -412 127 -406 161
rect -452 89 -406 127
rect -452 55 -446 89
rect -412 55 -406 89
rect -452 17 -406 55
rect -452 -17 -446 17
rect -412 -17 -406 17
rect -452 -55 -406 -17
rect -452 -89 -446 -55
rect -412 -89 -406 -55
rect -452 -127 -406 -89
rect -452 -161 -446 -127
rect -412 -161 -406 -127
rect -452 -199 -406 -161
rect -452 -233 -446 -199
rect -412 -233 -406 -199
rect -452 -271 -406 -233
rect -452 -305 -446 -271
rect -412 -305 -406 -271
rect -452 -343 -406 -305
rect -452 -377 -446 -343
rect -412 -377 -406 -343
rect -452 -400 -406 -377
rect 406 377 452 400
rect 406 343 412 377
rect 446 343 452 377
rect 406 305 452 343
rect 406 271 412 305
rect 446 271 452 305
rect 406 233 452 271
rect 406 199 412 233
rect 446 199 452 233
rect 406 161 452 199
rect 406 127 412 161
rect 446 127 452 161
rect 406 89 452 127
rect 406 55 412 89
rect 446 55 452 89
rect 406 17 452 55
rect 406 -17 412 17
rect 446 -17 452 17
rect 406 -55 452 -17
rect 406 -89 412 -55
rect 446 -89 452 -55
rect 406 -127 452 -89
rect 406 -161 412 -127
rect 446 -161 452 -127
rect 406 -199 452 -161
rect 406 -233 412 -199
rect 446 -233 452 -199
rect 406 -271 452 -233
rect 406 -305 412 -271
rect 446 -305 452 -271
rect 406 -343 452 -305
rect 406 -377 412 -343
rect 446 -377 452 -343
rect 406 -400 452 -377
<< end >>
