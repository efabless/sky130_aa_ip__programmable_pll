magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect -32616 3266 -31841 3358
<< locali >>
rect -3644 13816 16487 14578
rect -17873 12651 -17182 12662
rect -20204 12562 -17182 12651
rect -3644 12613 -2882 13816
rect -2298 13246 8970 13579
rect -2298 12868 -2037 13246
rect -2298 12762 -2256 12868
rect -2078 12762 -2037 12868
rect -17875 12469 -17182 12562
rect -34192 11775 -25170 11988
rect -34192 11765 -32133 11775
rect -34192 10024 -33920 11765
rect -30632 11658 -29305 11775
rect -17839 11764 -17707 11800
rect -17839 11730 -17825 11764
rect -17791 11730 -17753 11764
rect -17719 11730 -17707 11764
rect -17839 11729 -17707 11730
rect -18047 11693 -17707 11729
rect -33425 11595 -33364 11625
rect -33425 11561 -33412 11595
rect -33378 11561 -33364 11595
rect -19082 11573 -18712 11616
rect -17953 11588 -17547 11622
rect -33534 11509 -33473 11539
rect -33534 11475 -33521 11509
rect -33487 11475 -33473 11509
rect -33725 11430 -33664 11460
rect -33725 11396 -33712 11430
rect -33678 11396 -33664 11430
rect -33725 11358 -33664 11396
rect -33725 11324 -33712 11358
rect -33678 11324 -33664 11358
rect -33725 11286 -33664 11324
rect -33534 11437 -33473 11475
rect -33534 11403 -33521 11437
rect -33487 11403 -33473 11437
rect -33534 11365 -33473 11403
rect -33425 11523 -33364 11561
rect -33425 11489 -33412 11523
rect -33378 11489 -33364 11523
rect -33425 11451 -33364 11489
rect -33425 11417 -33412 11451
rect -33378 11422 -33364 11451
rect -33378 11417 -32640 11422
rect -33425 11387 -32640 11417
rect -33534 11331 -33521 11365
rect -33487 11339 -33473 11365
rect -29273 11383 -29077 11384
rect -29273 11371 -29013 11383
rect -33487 11331 -32619 11339
rect -33534 11301 -32619 11331
rect -29273 11337 -29135 11371
rect -29101 11337 -29063 11371
rect -29029 11337 -29013 11371
rect -29273 11325 -29013 11337
rect -29273 11314 -29077 11325
rect -33725 11252 -33712 11286
rect -33678 11257 -33664 11286
rect -33678 11252 -32634 11257
rect -33725 11223 -32634 11252
rect -33725 11222 -33664 11223
rect -30895 11201 -30758 11213
rect -30895 11167 -30880 11201
rect -30846 11167 -30808 11201
rect -30774 11167 -30758 11201
rect -30895 11155 -30758 11167
rect -29440 11164 -28282 11225
rect -30800 11094 -30663 11106
rect -30800 11060 -30785 11094
rect -30751 11060 -30713 11094
rect -30679 11060 -30663 11094
rect -29440 11081 -29379 11164
rect -18965 11106 -18687 11130
rect -30800 11048 -30663 11060
rect -26078 11034 -25727 11077
rect -18965 11072 -18933 11106
rect -18899 11072 -18687 11106
rect -18965 11047 -18687 11072
rect -33213 10508 -33152 10527
rect -31634 10510 -29678 10662
rect -33213 10474 -33200 10508
rect -33166 10474 -33152 10508
rect -33326 10430 -33266 10459
rect -33326 10396 -33313 10430
rect -33279 10396 -33266 10430
rect -33326 10383 -33266 10396
rect -33213 10436 -33152 10474
rect -33213 10402 -33200 10436
rect -33166 10402 -33152 10436
rect -33326 10358 -33258 10383
rect -33326 10324 -33313 10358
rect -33279 10343 -33258 10358
rect -33213 10364 -33152 10402
rect -33279 10324 -33266 10343
rect -33873 10261 -33772 10301
rect -33873 10227 -33841 10261
rect -33807 10227 -33772 10261
rect -33873 10189 -33772 10227
rect -33326 10286 -33266 10324
rect -33213 10330 -33200 10364
rect -33166 10349 -33152 10364
rect -30925 10434 -30872 10445
rect -30925 10400 -30918 10434
rect -30884 10400 -30872 10434
rect -30925 10362 -30872 10400
rect -30925 10349 -30918 10362
rect -33166 10330 -30918 10349
rect -33213 10328 -30918 10330
rect -30884 10328 -30872 10362
rect -33213 10313 -30872 10328
rect -33213 10311 -33152 10313
rect -33326 10252 -33313 10286
rect -33279 10266 -33266 10286
rect -30909 10268 -30777 10275
rect -30909 10266 -30894 10268
rect -33279 10252 -30894 10266
rect -33326 10234 -30894 10252
rect -30860 10234 -30822 10268
rect -30788 10234 -30777 10268
rect -33326 10226 -30777 10234
rect -33326 10222 -33266 10226
rect -30909 10222 -30777 10226
rect -33873 10155 -33841 10189
rect -33807 10155 -33772 10189
rect -33873 10128 -33772 10155
rect -29363 10128 -29306 10680
rect -33873 10117 -29306 10128
rect -33873 10083 -33841 10117
rect -33807 10083 -29306 10117
rect -33873 10065 -29306 10083
rect -33873 10058 -33772 10065
rect -34192 9911 -28709 10024
rect -34192 9891 -29379 9911
rect -34192 9792 -29420 9891
rect -32954 9457 -32894 9486
rect -32954 9423 -32941 9457
rect -32907 9423 -32894 9457
rect -31186 9451 -30809 9486
rect -32954 9385 -32894 9423
rect -30941 9403 -30883 9411
rect -32954 9351 -32941 9385
rect -32907 9351 -32894 9385
rect -30967 9395 -30776 9403
rect -30967 9365 -30929 9395
rect -32954 9313 -32894 9351
rect -32954 9279 -32941 9313
rect -32907 9287 -32894 9313
rect -30941 9361 -30929 9365
rect -30895 9365 -30776 9395
rect -30895 9361 -30883 9365
rect -30941 9323 -30883 9361
rect -30941 9289 -30929 9323
rect -30895 9289 -30883 9323
rect -32907 9279 -32784 9287
rect -32954 9251 -32784 9279
rect -31038 9264 -30980 9280
rect -30941 9274 -30883 9289
rect -32954 9249 -32894 9251
rect -31038 9230 -31026 9264
rect -30992 9230 -30980 9264
rect -33080 9153 -32684 9193
rect -31038 9192 -30980 9230
rect -31252 9167 -31194 9183
rect -33080 9048 -33040 9153
rect -31252 9133 -31240 9167
rect -31206 9133 -31194 9167
rect -31038 9158 -31026 9192
rect -30992 9180 -30980 9192
rect -30843 9180 -30809 9321
rect -29521 9226 -29043 9260
rect -30992 9158 -30809 9180
rect -31038 9146 -30809 9158
rect -31038 9143 -30980 9146
rect -31252 9095 -31194 9133
rect -31252 9061 -31240 9095
rect -31206 9061 -31194 9095
rect -33097 9019 -33037 9048
rect -31252 9046 -31194 9061
rect -33097 8985 -33084 9019
rect -33050 8985 -33037 9019
rect -33097 8947 -33037 8985
rect -33097 8913 -33084 8947
rect -33050 8913 -33037 8947
rect -33097 8875 -33037 8913
rect -33097 8841 -33084 8875
rect -33050 8841 -33037 8875
rect -33097 8811 -33037 8841
rect -28072 8787 -27986 8811
rect -31932 8713 -30931 8767
rect -32101 8652 -30931 8713
rect -28072 8664 -27862 8787
rect -31046 8634 -30931 8652
rect -31046 8624 -30586 8634
rect -29820 8624 -27862 8664
rect -31046 8509 -27862 8624
rect -26940 8675 -26672 8725
rect -25910 8675 -25727 11034
rect -26940 8672 -25727 8675
rect -26940 8494 -26850 8672
rect -26744 8494 -25727 8672
rect -26940 8492 -25727 8494
rect -24767 9088 -24614 10850
rect -21150 10058 -18798 10101
rect -18974 10056 -18798 10058
rect -18974 10022 -18937 10056
rect -18903 10022 -18865 10056
rect -18831 10022 -18798 10056
rect -18974 9979 -18798 10022
rect -24500 9734 -24314 9761
rect -24500 9628 -24459 9734
rect -24353 9628 -24314 9734
rect -24500 9607 -24314 9628
rect -17581 9329 -17547 11588
rect -2298 11124 -2037 12762
rect -1813 12244 -1613 12278
rect -1813 12215 5950 12244
rect -1813 11965 -1770 12215
rect -1664 12072 5950 12215
rect -1664 11965 -1613 12072
rect -1813 11907 -1613 11965
rect 5373 11346 5665 11347
rect -1601 11297 5665 11346
rect -1601 11295 -1031 11297
rect -1601 11261 -1555 11295
rect -1521 11261 -1483 11295
rect -1449 11261 -1411 11295
rect -1377 11261 -1339 11295
rect -1305 11263 -1031 11295
rect -997 11263 -959 11297
rect -925 11263 -887 11297
rect -853 11263 -815 11297
rect -781 11293 5665 11297
rect -781 11263 5429 11293
rect -1305 11261 5429 11263
rect -1601 11259 5429 11261
rect 5463 11259 5501 11293
rect 5535 11259 5573 11293
rect 5607 11259 5665 11293
rect -1601 11207 5665 11259
rect 6109 11295 6209 11326
rect 6109 11261 6142 11295
rect 6176 11261 6209 11295
rect 6109 11231 6209 11261
rect 8425 11163 8970 13246
rect 15384 12307 16487 13816
rect 18 10702 556 10743
rect 18 10524 79 10702
rect 257 10524 556 10702
rect 18 10496 556 10524
rect 389 10302 551 10307
rect 389 10124 417 10302
rect 523 10124 551 10302
rect 389 10120 551 10124
rect -1573 9733 -1355 9741
rect 5603 9733 5756 9772
rect -1573 9712 5756 9733
rect -1573 9709 5659 9712
rect -1573 9675 -1554 9709
rect -1520 9675 -1482 9709
rect -1448 9675 -1410 9709
rect -1376 9678 5659 9709
rect 5693 9678 5756 9712
rect -1376 9675 5756 9678
rect -1573 9658 5756 9675
rect -1573 9652 -1355 9658
rect 5603 9621 5756 9658
rect 6333 9749 6430 9772
rect 6333 9715 6361 9749
rect 6395 9715 6430 9749
rect 6333 9677 6430 9715
rect 6333 9643 6361 9677
rect 6395 9643 6430 9677
rect 6333 9621 6430 9643
rect -591 9512 -541 9518
rect 4921 9512 5019 9526
rect -600 9505 5019 9512
rect -600 9471 -585 9505
rect -551 9497 5019 9505
rect -551 9471 4954 9497
rect -600 9463 4954 9471
rect 4988 9463 5019 9497
rect -600 9431 5019 9463
rect -600 9397 -584 9431
rect -550 9425 5019 9431
rect -550 9397 4954 9425
rect -600 9391 4954 9397
rect 4988 9391 5019 9425
rect -600 9389 5019 9391
rect -591 9385 -541 9389
rect 4921 9362 5019 9389
rect -17581 9313 -17397 9329
rect -17581 9279 -17533 9313
rect -17499 9279 -17461 9313
rect -17427 9279 -17397 9313
rect -17581 9266 -17397 9279
rect -17560 9265 -17397 9266
rect -24767 8935 -23812 9088
rect -26940 8460 -26672 8492
rect -29326 8275 -25788 8324
rect -29326 8268 -25946 8275
rect -29326 8162 -29272 8268
rect -29166 8169 -25946 8268
rect -25840 8169 -25788 8275
rect -29166 8162 -25788 8169
rect -29326 8118 -25788 8162
rect -25996 8116 -25788 8118
rect -26935 7858 -26667 7905
rect -34338 7853 -26667 7858
rect -34338 7675 -26858 7853
rect -26752 7675 -26667 7853
rect -34338 7672 -26667 7675
rect -26935 7640 -26667 7672
rect -24767 7641 -24614 8935
rect -17355 7710 -17266 8433
rect -21151 7625 -17266 7710
rect -17355 7510 -17266 7625
rect -17355 7421 -17265 7510
rect -17355 7264 -17266 7421
rect -17067 7370 -16798 8390
rect -16398 8387 -16330 8391
rect -16521 7367 -16252 8387
rect -15644 7379 -15375 8399
rect -14782 7373 -14513 8393
rect -13879 7375 -13610 8395
rect -12848 7379 -12579 8399
rect -16398 7353 -16330 7367
rect -11896 7067 -11598 8414
rect -10287 7195 -10026 8472
rect -9450 7195 -9189 8461
rect -8410 7195 -8149 8480
rect -6952 7195 -6691 8495
rect -5738 7195 -5477 8468
rect -3792 7195 -3531 8507
rect -2298 7131 -2037 8600
rect -753 7258 -689 7281
rect 4612 7258 4695 7495
rect -753 7237 4695 7258
rect -753 7203 -739 7237
rect -705 7203 4695 7237
rect -753 7175 4695 7203
rect -753 7163 -689 7175
rect -32776 6966 -25139 6995
rect -32776 6860 -29375 6966
rect -29269 6860 -25139 6966
rect -1074 6954 -1015 6961
rect -1074 6930 2902 6954
rect -1074 6896 -1062 6930
rect -1028 6896 2902 6930
rect -1074 6871 2902 6896
rect -1074 6866 -1015 6871
rect -32776 6828 -25139 6860
rect -32406 6595 -31624 6828
rect -31248 6657 -30730 6828
rect -30359 6660 -29806 6828
rect -17839 6820 -17707 6847
rect -17839 6795 -17788 6820
rect -18015 6786 -17788 6795
rect -17754 6786 -17707 6820
rect -18015 6759 -17707 6786
rect -17564 6689 -17422 6705
rect -17564 6688 -17543 6689
rect -19068 6639 -18688 6682
rect -17930 6655 -17543 6688
rect -17509 6655 -17471 6689
rect -17437 6655 -17422 6689
rect -17930 6654 -17422 6655
rect -17564 6641 -17422 6654
rect -2297 6507 -1143 6768
rect 2819 6648 2902 6871
rect -1706 6309 -1561 6355
rect -1706 6275 -1651 6309
rect -1617 6275 -1561 6309
rect -29476 6164 -28210 6225
rect -1706 6220 -1561 6275
rect -17565 6195 -17460 6201
rect -17980 6171 -17460 6195
rect -31431 6078 -31373 6094
rect -31431 6044 -31419 6078
rect -31385 6044 -31373 6078
rect -31431 6006 -31373 6044
rect -31431 5972 -31419 6006
rect -31385 5999 -31373 6006
rect -30515 6077 -30457 6093
rect -30515 6043 -30503 6077
rect -30469 6043 -30457 6077
rect -30515 6005 -30457 6043
rect -31385 5972 -31256 5999
rect -31431 5963 -31256 5972
rect -30515 5971 -30503 6005
rect -30469 5998 -30457 6005
rect -30469 5971 -30366 5998
rect -31431 5957 -31373 5963
rect -30515 5962 -30366 5971
rect -30515 5956 -30457 5962
rect -33725 5889 -33665 5918
rect -33725 5855 -33712 5889
rect -33678 5855 -33665 5889
rect -33725 5817 -33665 5855
rect -33725 5783 -33712 5817
rect -33678 5783 -33665 5817
rect -31356 5907 -31298 5923
rect -31356 5873 -31344 5907
rect -31310 5873 -31298 5907
rect -31356 5835 -31298 5873
rect -30740 5917 -30603 5929
rect -30740 5883 -30725 5917
rect -30691 5883 -30653 5917
rect -30619 5883 -30603 5917
rect -30740 5871 -30603 5883
rect -30438 5905 -30380 5921
rect -30438 5871 -30426 5905
rect -30392 5871 -30380 5905
rect -31356 5801 -31344 5835
rect -31310 5801 -31298 5835
rect -31356 5786 -31298 5801
rect -30438 5833 -30380 5871
rect -29809 5916 -29672 5928
rect -29809 5882 -29794 5916
rect -29760 5882 -29722 5916
rect -29688 5882 -29672 5916
rect -29809 5870 -29672 5882
rect -30438 5799 -30426 5833
rect -30392 5799 -30380 5833
rect -29476 5806 -29415 6164
rect -25975 6115 -25838 6147
rect -25975 6077 -25957 6115
rect -26104 6034 -25957 6077
rect -25975 6009 -25957 6034
rect -25851 6009 -25838 6115
rect -17980 6137 -17529 6171
rect -17495 6137 -17460 6171
rect -17980 6113 -17460 6137
rect -17565 6106 -17460 6113
rect -25975 5981 -25838 6009
rect -30438 5784 -30380 5799
rect -33725 5745 -33665 5783
rect -33725 5711 -33712 5745
rect -33678 5737 -33665 5745
rect -29863 5745 -29415 5806
rect -33678 5711 -32523 5737
rect -33725 5696 -32523 5711
rect -33725 5681 -33665 5696
rect -33534 5648 -33474 5661
rect -33534 5632 -32496 5648
rect -33534 5598 -33521 5632
rect -33487 5607 -32496 5632
rect -33487 5598 -33474 5607
rect -33534 5560 -33474 5598
rect -33534 5526 -33521 5560
rect -33487 5526 -33474 5560
rect -31627 5568 -31490 5580
rect -33534 5488 -33474 5526
rect -33534 5454 -33521 5488
rect -33487 5454 -33474 5488
rect -33534 5424 -33474 5454
rect -33424 5556 -33364 5558
rect -33424 5529 -32540 5556
rect -33424 5495 -33411 5529
rect -33377 5515 -32540 5529
rect -31627 5534 -31612 5568
rect -31578 5534 -31540 5568
rect -31506 5534 -31490 5568
rect -31627 5522 -31490 5534
rect -33377 5495 -33364 5515
rect -33424 5457 -33364 5495
rect -33424 5423 -33411 5457
rect -33377 5423 -33364 5457
rect -33424 5385 -33364 5423
rect -33424 5351 -33411 5385
rect -33377 5351 -33364 5385
rect -33424 5321 -33364 5351
rect -31841 5369 -30000 5485
rect -29863 5467 -29802 5745
rect -29548 5680 -29431 5695
rect -29548 5650 -29306 5680
rect -29548 5616 -29507 5650
rect -29473 5644 -29306 5650
rect -29473 5616 -29431 5644
rect -29548 5572 -29431 5616
rect -31841 5188 -31725 5369
rect -1989 5205 -1866 5206
rect -1990 5201 -1866 5205
rect -32499 5165 -31695 5188
rect -32499 5059 -32449 5165
rect -31767 5059 -31695 5165
rect -1990 5167 -1982 5201
rect -1948 5167 -1908 5201
rect -1874 5167 -1866 5201
rect -1990 5162 -1866 5167
rect -33326 5032 -33268 5048
rect -32499 5038 -31695 5059
rect -33326 4998 -33314 5032
rect -33280 4998 -33268 5032
rect -33326 4960 -33268 4998
rect -33326 4926 -33314 4960
rect -33280 4952 -33268 4960
rect -31451 5032 -31393 5048
rect -31451 4998 -31439 5032
rect -31405 4998 -31393 5032
rect -31451 4960 -31393 4998
rect -30188 5030 -28612 5064
rect -31451 4952 -31439 4960
rect -33280 4926 -31439 4952
rect -31405 4926 -31393 4960
rect -33326 4911 -31393 4926
rect -31358 4953 -31300 4969
rect -31358 4919 -31346 4953
rect -31312 4919 -31300 4953
rect -31358 4881 -31300 4919
rect -30188 4924 -29341 5030
rect -29235 4924 -28612 5030
rect -30188 4892 -28612 4924
rect -33213 4873 -33155 4876
rect -31358 4873 -31346 4881
rect -33213 4860 -31346 4873
rect -33213 4826 -33201 4860
rect -33167 4847 -31346 4860
rect -31312 4847 -31300 4881
rect -33167 4832 -31300 4847
rect -30537 4874 -30479 4890
rect -30537 4840 -30525 4874
rect -30491 4840 -30479 4874
rect -33167 4826 -33155 4832
rect -33213 4788 -33155 4826
rect -30537 4802 -30479 4840
rect -33213 4754 -33201 4788
rect -33167 4754 -33155 4788
rect -33213 4739 -33155 4754
rect -33099 4794 -33041 4795
rect -30537 4794 -30525 4802
rect -33099 4779 -30525 4794
rect -33099 4745 -33087 4779
rect -33053 4768 -30525 4779
rect -30491 4768 -30479 4802
rect -33053 4753 -30479 4768
rect -30444 4797 -30386 4813
rect -30444 4763 -30432 4797
rect -30398 4763 -30386 4797
rect -33053 4745 -33041 4753
rect -33099 4707 -33041 4745
rect -30444 4725 -30386 4763
rect -30444 4717 -30432 4725
rect -33099 4673 -33087 4707
rect -33053 4673 -33041 4707
rect -33099 4658 -33041 4673
rect -32954 4691 -30432 4717
rect -30398 4691 -30386 4725
rect -32954 4676 -30386 4691
rect -32954 4651 -32896 4676
rect -32954 4617 -32942 4651
rect -32908 4617 -32896 4651
rect -32954 4580 -32896 4617
rect -32712 4581 -31729 4626
rect -32712 4547 -32675 4581
rect -32641 4547 -32603 4581
rect -32569 4547 -32531 4581
rect -32497 4547 -32459 4581
rect -32425 4547 -32387 4581
rect -32353 4547 -32315 4581
rect -32281 4547 -32243 4581
rect -32209 4547 -32171 4581
rect -32137 4547 -32099 4581
rect -32065 4547 -32027 4581
rect -31993 4547 -31955 4581
rect -31921 4547 -31883 4581
rect -31849 4547 -31811 4581
rect -31777 4547 -31729 4581
rect -32712 4511 -31729 4547
rect -31387 3967 -31329 3983
rect -31387 3933 -31375 3967
rect -31341 3933 -31329 3967
rect -31387 3895 -31329 3933
rect -31387 3861 -31375 3895
rect -31341 3861 -31329 3895
rect -31387 3846 -31329 3861
rect -30657 3885 -30599 3901
rect -30188 3897 -30016 4892
rect -1990 4354 -1932 5162
rect -1846 4643 -1723 4648
rect -1846 4609 -1839 4643
rect -1805 4609 -1765 4643
rect -1731 4609 -1723 4643
rect -1846 4604 -1723 4609
rect -29647 4303 -29589 4304
rect -29647 4288 -29056 4303
rect -29647 4254 -29635 4288
rect -29601 4254 -29056 4288
rect -29647 4235 -29056 4254
rect -29647 4216 -29589 4235
rect -29647 4182 -29635 4216
rect -29601 4182 -29589 4216
rect -29647 4167 -29589 4182
rect -30657 3851 -30645 3885
rect -30611 3851 -30599 3885
rect -30657 3813 -30599 3851
rect -30657 3802 -30645 3813
rect -31419 3779 -30645 3802
rect -30611 3779 -30599 3813
rect -30190 3869 -30014 3897
rect -30190 3835 -30154 3869
rect -30120 3835 -30082 3869
rect -30048 3835 -30014 3869
rect -30190 3810 -30014 3835
rect -31419 3764 -30599 3779
rect -29732 3799 -29674 3815
rect -29732 3765 -29720 3799
rect -29686 3765 -29674 3799
rect -29732 3727 -29674 3765
rect -29732 3718 -29720 3727
rect -31373 3693 -29720 3718
rect -29686 3693 -29674 3727
rect -31373 3683 -29674 3693
rect -29732 3678 -29674 3683
rect -18987 3562 -18787 3586
rect -29368 3552 -18787 3562
rect -29368 3511 -18935 3552
rect -29368 3477 -29349 3511
rect -29315 3477 -29277 3511
rect -29243 3477 -18935 3511
rect -29368 3446 -18935 3477
rect -18829 3446 -18787 3552
rect -29368 3426 -18787 3446
rect -18987 3415 -18787 3426
rect -32616 3328 -30014 3358
rect -32616 3294 -30156 3328
rect -30122 3294 -30084 3328
rect -30050 3294 -30014 3328
rect -17850 3308 -17687 3328
rect -32616 3266 -30014 3294
rect -29545 3293 -17687 3308
rect -29545 3291 -17822 3293
rect -29545 3185 -29531 3291
rect -29425 3187 -17822 3291
rect -17716 3187 -17687 3293
rect -29425 3185 -17687 3187
rect -29545 3172 -17687 3185
rect -29545 3171 -29407 3172
rect -32751 3126 -32593 3159
rect -17850 3153 -17687 3172
rect -29683 3126 -29546 3131
rect -32751 3119 -29546 3126
rect -32751 3113 -29668 3119
rect -32751 3079 -32729 3113
rect -32695 3079 -32657 3113
rect -32623 3085 -29668 3113
rect -29634 3085 -29596 3119
rect -29562 3085 -29546 3119
rect -32623 3079 -29546 3085
rect -32751 3074 -29546 3079
rect -32751 3043 -32593 3074
rect -29683 3073 -29546 3074
rect -1989 2944 -1933 4354
rect -1890 4096 -1825 4113
rect -1890 4062 -1882 4096
rect -1848 4062 -1825 4096
rect -1890 4022 -1825 4062
rect -1890 3988 -1882 4022
rect -1848 3988 -1825 4022
rect -1890 3976 -1825 3988
rect -1887 3332 -1833 3976
rect -1887 3298 -1881 3332
rect -1847 3298 -1833 3332
rect -1887 3258 -1833 3298
rect -1887 3224 -1881 3258
rect -1847 3224 -1833 3258
rect -1887 3216 -1833 3224
rect -1782 3334 -1728 4604
rect -1782 3300 -1772 3334
rect -1738 3300 -1728 3334
rect -1782 3260 -1728 3300
rect -1782 3226 -1772 3260
rect -1738 3226 -1728 3260
rect -1782 3216 -1728 3226
rect -1683 3117 -1627 6220
rect -1404 5713 -1143 6507
rect -921 6151 -852 6169
rect 4292 6151 4403 6400
rect -921 6116 4403 6151
rect -921 6082 -904 6116
rect -870 6082 4403 6116
rect -921 6040 4403 6082
rect -921 6030 -852 6040
rect 6703 5826 8225 5895
rect -1404 5452 -434 5713
rect -1412 5339 -1221 5345
rect -1412 5307 -849 5339
rect -1412 5273 -1370 5307
rect -1336 5273 -1298 5307
rect -1264 5273 -849 5307
rect -1412 5256 -849 5273
rect -1412 5238 -1221 5256
rect -1256 5051 -1108 5057
rect -1256 5017 -1241 5051
rect -1207 5017 -1167 5051
rect -1133 5017 -1108 5051
rect -1256 5009 -1108 5017
rect -1412 4913 -1289 4918
rect -1412 4879 -1404 4913
rect -1370 4879 -1330 4913
rect -1296 4879 -1289 4913
rect -1412 4874 -1289 4879
rect -1571 4782 -1414 4787
rect -1571 4748 -1529 4782
rect -1495 4748 -1455 4782
rect -1421 4748 -1414 4782
rect -1571 4747 -1414 4748
rect -1571 3334 -1517 4747
rect -1357 4443 -1303 4874
rect -1571 3300 -1561 3334
rect -1527 3300 -1517 3334
rect -1571 3260 -1517 3300
rect -1571 3226 -1561 3260
rect -1527 3226 -1517 3260
rect -1571 3216 -1517 3226
rect -1456 4389 -1303 4443
rect -1456 3334 -1402 4389
rect -1456 3300 -1446 3334
rect -1412 3300 -1402 3334
rect -1456 3260 -1402 3300
rect -1456 3226 -1446 3260
rect -1412 3226 -1402 3260
rect -1456 3216 -1402 3226
rect -1312 3307 -1298 3341
rect -1264 3311 -1258 3341
rect -1214 3311 -1160 5009
rect -932 3391 -849 5256
rect -695 3672 -434 5452
rect 6703 5326 6829 5826
rect 18 4509 313 4559
rect 18 4403 38 4509
rect 288 4461 313 4509
rect 288 4422 700 4461
rect 288 4403 313 4422
rect 18 4356 313 4403
rect 1089 3672 1350 4352
rect -695 3411 1350 3672
rect -1264 3307 -1160 3311
rect -1312 3267 -1160 3307
rect -1312 3233 -1298 3267
rect -1264 3257 -1160 3267
rect -956 3354 -828 3391
rect -956 3320 -909 3354
rect -875 3320 -828 3354
rect -956 3282 -828 3320
rect -1264 3233 -1258 3257
rect -1312 3216 -1258 3233
rect -956 3248 -909 3282
rect -875 3248 -828 3282
rect -956 3212 -828 3248
rect -1683 3083 -1672 3117
rect -1638 3083 -1627 3117
rect -1683 3043 -1627 3083
rect -1683 3009 -1672 3043
rect -1638 3009 -1627 3043
rect -1683 2999 -1627 3009
rect -34598 2928 983 2944
rect -34598 2889 -25647 2928
rect -34598 2855 -33733 2889
rect -33699 2855 -25647 2889
rect -34598 2822 -25647 2855
rect -25541 2822 983 2928
rect -34598 2808 983 2822
rect -34598 2695 1180 2745
rect -34598 2690 -1903 2695
rect -34598 2656 -33542 2690
rect -33508 2661 -1903 2690
rect -1869 2661 1180 2695
rect -33508 2656 1180 2661
rect -34598 2609 1180 2656
rect -34598 2462 1218 2512
rect -34598 2457 -1797 2462
rect -34598 2423 -33436 2457
rect -33402 2428 -1797 2457
rect -1763 2428 1218 2462
rect -33402 2423 1218 2428
rect -34598 2376 1218 2423
rect -34598 2205 965 2257
rect -34598 2200 -1704 2205
rect -34598 2166 -33343 2200
rect -33309 2171 -1704 2200
rect -1670 2171 965 2205
rect -33309 2166 965 2171
rect -34598 2121 965 2166
rect -1552 1971 -1416 1973
rect -34598 1925 1034 1971
rect -34598 1920 -1597 1925
rect -34598 1886 -33236 1920
rect -33202 1891 -1597 1920
rect -1563 1891 1034 1925
rect -33202 1886 1034 1891
rect -34598 1835 1034 1886
rect -34598 1830 -32782 1835
rect -34598 1620 1011 1672
rect -34598 1615 -1438 1620
rect -34598 1581 -33077 1615
rect -33043 1586 -1438 1615
rect -1404 1586 1011 1620
rect -33043 1581 1011 1586
rect -34598 1536 1011 1581
rect -34598 1253 1042 1302
rect -34598 1248 -1287 1253
rect -34598 1214 -32926 1248
rect -32892 1219 -1287 1248
rect -1253 1219 1042 1253
rect -32892 1214 1042 1219
rect -34598 1166 1042 1214
rect -34042 1058 -33829 1090
rect -34598 1043 313 1058
rect -34598 937 -33995 1043
rect -33889 1042 313 1043
rect -33889 937 42 1042
rect -34598 936 42 937
rect 292 936 313 1042
rect -34598 922 313 936
rect -34042 912 -33829 922
rect -17848 783 7096 798
rect -17848 677 -17826 783
rect -17720 782 7096 783
rect -17720 677 6977 782
rect -17848 676 6977 677
rect 7083 676 7096 782
rect -17848 662 7096 676
rect -34598 546 570 560
rect -34598 440 421 546
rect 527 440 570 546
rect -34598 425 570 440
<< viali >>
rect -2256 12762 -2078 12868
rect -17825 11730 -17791 11764
rect -17753 11730 -17719 11764
rect -33412 11561 -33378 11595
rect -33521 11475 -33487 11509
rect -33712 11396 -33678 11430
rect -33712 11324 -33678 11358
rect -33521 11403 -33487 11437
rect -33412 11489 -33378 11523
rect -33412 11417 -33378 11451
rect -33521 11331 -33487 11365
rect -29135 11337 -29101 11371
rect -29063 11337 -29029 11371
rect -33712 11252 -33678 11286
rect -30880 11167 -30846 11201
rect -30808 11167 -30774 11201
rect -30785 11060 -30751 11094
rect -30713 11060 -30679 11094
rect -18933 11072 -18899 11106
rect -33200 10474 -33166 10508
rect -33313 10396 -33279 10430
rect -33200 10402 -33166 10436
rect -33313 10324 -33279 10358
rect -33841 10227 -33807 10261
rect -33200 10330 -33166 10364
rect -30918 10400 -30884 10434
rect -30918 10328 -30884 10362
rect -33313 10252 -33279 10286
rect -30894 10234 -30860 10268
rect -30822 10234 -30788 10268
rect -33841 10155 -33807 10189
rect -33841 10083 -33807 10117
rect -32941 9423 -32907 9457
rect -32941 9351 -32907 9385
rect -32941 9279 -32907 9313
rect -30929 9361 -30895 9395
rect -30929 9289 -30895 9323
rect -31026 9230 -30992 9264
rect -31240 9133 -31206 9167
rect -31026 9158 -30992 9192
rect -31240 9061 -31206 9095
rect -33084 8985 -33050 9019
rect -33084 8913 -33050 8947
rect -33084 8841 -33050 8875
rect -26850 8494 -26744 8672
rect -18937 10022 -18903 10056
rect -18865 10022 -18831 10056
rect -24459 9628 -24353 9734
rect -1770 11965 -1664 12215
rect -1555 11261 -1521 11295
rect -1483 11261 -1449 11295
rect -1411 11261 -1377 11295
rect -1339 11261 -1305 11295
rect -1031 11263 -997 11297
rect -959 11263 -925 11297
rect -887 11263 -853 11297
rect -815 11263 -781 11297
rect 5429 11259 5463 11293
rect 5501 11259 5535 11293
rect 5573 11259 5607 11293
rect 6142 11261 6176 11295
rect 79 10524 257 10702
rect 417 10124 523 10302
rect -1554 9675 -1520 9709
rect -1482 9675 -1448 9709
rect -1410 9675 -1376 9709
rect 5659 9678 5693 9712
rect 6361 9715 6395 9749
rect 6361 9643 6395 9677
rect -585 9471 -551 9505
rect 4954 9463 4988 9497
rect -584 9397 -550 9431
rect 4954 9391 4988 9425
rect -17533 9279 -17499 9313
rect -17461 9279 -17427 9313
rect -29272 8162 -29166 8268
rect -25946 8169 -25840 8275
rect -26858 7675 -26752 7853
rect -739 7203 -705 7237
rect -29375 6860 -29269 6966
rect -1062 6896 -1028 6930
rect -17788 6786 -17754 6820
rect -17543 6655 -17509 6689
rect -17471 6655 -17437 6689
rect -1651 6275 -1617 6309
rect -31419 6044 -31385 6078
rect -31419 5972 -31385 6006
rect -30503 6043 -30469 6077
rect -30503 5971 -30469 6005
rect -33712 5855 -33678 5889
rect -33712 5783 -33678 5817
rect -31344 5873 -31310 5907
rect -30725 5883 -30691 5917
rect -30653 5883 -30619 5917
rect -30426 5871 -30392 5905
rect -31344 5801 -31310 5835
rect -29794 5882 -29760 5916
rect -29722 5882 -29688 5916
rect -30426 5799 -30392 5833
rect -25957 6009 -25851 6115
rect -17529 6137 -17495 6171
rect -33712 5711 -33678 5745
rect -33521 5598 -33487 5632
rect -33521 5526 -33487 5560
rect -33521 5454 -33487 5488
rect -33411 5495 -33377 5529
rect -31612 5534 -31578 5568
rect -31540 5534 -31506 5568
rect -33411 5423 -33377 5457
rect -33411 5351 -33377 5385
rect -29507 5616 -29473 5650
rect -32449 5059 -31767 5165
rect -1982 5167 -1948 5201
rect -1908 5167 -1874 5201
rect -33314 4998 -33280 5032
rect -33314 4926 -33280 4960
rect -31439 4998 -31405 5032
rect -31439 4926 -31405 4960
rect -31346 4919 -31312 4953
rect -29341 4924 -29235 5030
rect -33201 4826 -33167 4860
rect -31346 4847 -31312 4881
rect -30525 4840 -30491 4874
rect -33201 4754 -33167 4788
rect -33087 4745 -33053 4779
rect -30525 4768 -30491 4802
rect -30432 4763 -30398 4797
rect -33087 4673 -33053 4707
rect -30432 4691 -30398 4725
rect -32942 4617 -32908 4651
rect -32675 4547 -32641 4581
rect -32603 4547 -32569 4581
rect -32531 4547 -32497 4581
rect -32459 4547 -32425 4581
rect -32387 4547 -32353 4581
rect -32315 4547 -32281 4581
rect -32243 4547 -32209 4581
rect -32171 4547 -32137 4581
rect -32099 4547 -32065 4581
rect -32027 4547 -31993 4581
rect -31955 4547 -31921 4581
rect -31883 4547 -31849 4581
rect -31811 4547 -31777 4581
rect -31375 3933 -31341 3967
rect -31375 3861 -31341 3895
rect -1839 4609 -1805 4643
rect -1765 4609 -1731 4643
rect -29635 4254 -29601 4288
rect -29635 4182 -29601 4216
rect -30645 3851 -30611 3885
rect -30645 3779 -30611 3813
rect -30154 3835 -30120 3869
rect -30082 3835 -30048 3869
rect -29720 3765 -29686 3799
rect -29720 3693 -29686 3727
rect -29349 3477 -29315 3511
rect -29277 3477 -29243 3511
rect -18935 3446 -18829 3552
rect -30156 3294 -30122 3328
rect -30084 3294 -30050 3328
rect -29531 3185 -29425 3291
rect -17822 3187 -17716 3293
rect -32729 3079 -32695 3113
rect -32657 3079 -32623 3113
rect -29668 3085 -29634 3119
rect -29596 3085 -29562 3119
rect -1882 4062 -1848 4096
rect -1882 3988 -1848 4022
rect -1881 3298 -1847 3332
rect -1881 3224 -1847 3258
rect -1772 3300 -1738 3334
rect -1772 3226 -1738 3260
rect -904 6082 -870 6116
rect -1370 5273 -1336 5307
rect -1298 5273 -1264 5307
rect -1241 5017 -1207 5051
rect -1167 5017 -1133 5051
rect -1404 4879 -1370 4913
rect -1330 4879 -1296 4913
rect -1529 4748 -1495 4782
rect -1455 4748 -1421 4782
rect -1561 3300 -1527 3334
rect -1561 3226 -1527 3260
rect -1446 3300 -1412 3334
rect -1446 3226 -1412 3260
rect -1298 3307 -1264 3341
rect 38 4403 288 4509
rect -1298 3233 -1264 3267
rect -909 3320 -875 3354
rect -909 3248 -875 3282
rect -1672 3083 -1638 3117
rect -1672 3009 -1638 3043
rect -33733 2855 -33699 2889
rect -25647 2822 -25541 2928
rect -33542 2656 -33508 2690
rect -1903 2661 -1869 2695
rect -33436 2423 -33402 2457
rect -1797 2428 -1763 2462
rect -33343 2166 -33309 2200
rect -1704 2171 -1670 2205
rect -33236 1886 -33202 1920
rect -1597 1891 -1563 1925
rect -33077 1581 -33043 1615
rect -1438 1586 -1404 1620
rect -32926 1214 -32892 1248
rect -1287 1219 -1253 1253
rect -33995 937 -33889 1043
rect 42 936 292 1042
rect -17826 677 -17720 783
rect 6977 676 7083 782
rect 421 440 527 546
<< metal1 >>
rect 18196 15412 22119 15696
rect 17053 14479 20405 14790
rect 17328 14029 19301 14206
rect 11547 13470 13403 13691
rect 12074 12913 14120 13139
rect -26445 12868 -2037 12912
rect -26445 12762 -2256 12868
rect -2078 12762 -2037 12868
rect -26445 12722 -2037 12762
rect -33425 11595 -33364 11625
rect -33425 11561 -33412 11595
rect -33378 11561 -33364 11595
rect -33534 11509 -33473 11539
rect -33534 11475 -33521 11509
rect -33487 11475 -33473 11509
rect -33725 11430 -33664 11460
rect -33725 11396 -33712 11430
rect -33678 11396 -33664 11430
rect -33725 11358 -33664 11396
rect -33725 11324 -33712 11358
rect -33678 11324 -33664 11358
rect -33725 11286 -33664 11324
rect -33725 11252 -33712 11286
rect -33678 11252 -33664 11286
rect -33873 10261 -33772 10301
rect -33873 10246 -33841 10261
rect -34025 10227 -33841 10246
rect -33807 10227 -33772 10261
rect -34025 10189 -33772 10227
rect -34025 10155 -33841 10189
rect -33807 10155 -33772 10189
rect -34025 10117 -33772 10155
rect -34025 10083 -33841 10117
rect -33807 10083 -33772 10117
rect -34025 10058 -33772 10083
rect -34025 10015 -33785 10058
rect -34025 1090 -33889 10015
rect -33725 5889 -33664 11252
rect -33725 5855 -33712 5889
rect -33678 5855 -33664 5889
rect -33725 5817 -33664 5855
rect -33725 5783 -33712 5817
rect -33678 5783 -33664 5817
rect -33725 5745 -33664 5783
rect -33725 5711 -33712 5745
rect -33678 5711 -33664 5745
rect -33725 2933 -33664 5711
rect -33534 11437 -33473 11475
rect -33534 11403 -33521 11437
rect -33487 11403 -33473 11437
rect -33534 11365 -33473 11403
rect -33534 11331 -33521 11365
rect -33487 11331 -33473 11365
rect -33534 5632 -33473 11331
rect -33534 5598 -33521 5632
rect -33487 5598 -33473 5632
rect -33534 5560 -33473 5598
rect -33534 5526 -33521 5560
rect -33487 5526 -33473 5560
rect -33534 5488 -33473 5526
rect -33534 5454 -33521 5488
rect -33487 5454 -33473 5488
rect -33778 2889 -33655 2933
rect -33778 2855 -33733 2889
rect -33699 2855 -33655 2889
rect -33778 2810 -33655 2855
rect -33534 2734 -33473 5454
rect -33425 11523 -33364 11561
rect -26445 11555 -26255 12722
rect -25362 11635 -25245 11699
rect -18965 11686 -18870 12722
rect 12331 12433 14070 12698
rect -1813 12215 -1613 12278
rect -1813 11965 -1770 12215
rect -1664 11965 -1613 12215
rect 17522 12027 20097 12276
rect -1813 11926 -1613 11965
rect -2221 11898 -244 11926
rect -33425 11489 -33412 11523
rect -33378 11489 -33364 11523
rect -33425 11451 -33364 11489
rect -33425 11417 -33412 11451
rect -33378 11417 -33364 11451
rect -33425 11387 -33364 11417
rect -33425 5558 -33365 11387
rect -29159 11371 -29013 11383
rect -29159 11337 -29135 11371
rect -29101 11337 -29063 11371
rect -29029 11337 -29013 11371
rect -29159 11325 -29013 11337
rect -29159 11299 -29078 11325
rect -29471 11264 -29078 11299
rect -30895 11201 -30758 11213
rect -30895 11196 -30880 11201
rect -30923 11167 -30880 11196
rect -30846 11167 -30808 11201
rect -30774 11167 -30758 11201
rect -30923 11155 -30758 11167
rect -31342 10814 -30998 10849
rect -33213 10508 -33152 10527
rect -33213 10474 -33200 10508
rect -33166 10474 -33152 10508
rect -33326 10430 -33265 10460
rect -33326 10396 -33313 10430
rect -33279 10396 -33265 10430
rect -33326 10358 -33265 10396
rect -33326 10324 -33313 10358
rect -33279 10324 -33265 10358
rect -33326 10286 -33265 10324
rect -33326 10252 -33313 10286
rect -33279 10252 -33265 10286
rect -33425 5529 -33364 5558
rect -33425 5495 -33411 5529
rect -33377 5495 -33364 5529
rect -33425 5457 -33364 5495
rect -33425 5423 -33411 5457
rect -33377 5423 -33364 5457
rect -33425 5385 -33364 5423
rect -33425 5351 -33411 5385
rect -33377 5351 -33364 5385
rect -33425 5321 -33364 5351
rect -33587 2690 -33464 2734
rect -33587 2656 -33542 2690
rect -33508 2656 -33464 2690
rect -33587 2611 -33464 2656
rect -33425 2501 -33365 5321
rect -33326 5032 -33265 10252
rect -33326 4998 -33314 5032
rect -33280 4998 -33265 5032
rect -33326 4960 -33265 4998
rect -33326 4926 -33314 4960
rect -33280 4926 -33265 4960
rect -33481 2457 -33358 2501
rect -33481 2423 -33436 2457
rect -33402 2423 -33358 2457
rect -33481 2378 -33358 2423
rect -33326 2244 -33265 4926
rect -33213 10436 -33152 10474
rect -33213 10402 -33200 10436
rect -33166 10402 -33152 10436
rect -33213 10364 -33152 10402
rect -33213 10330 -33200 10364
rect -33166 10330 -33152 10364
rect -33213 4860 -33152 10330
rect -32954 9457 -32894 9486
rect -32954 9423 -32941 9457
rect -32907 9423 -32894 9457
rect -32954 9385 -32894 9423
rect -32954 9351 -32941 9385
rect -32907 9351 -32894 9385
rect -32954 9313 -32894 9351
rect -32954 9279 -32941 9313
rect -32907 9279 -32894 9313
rect -31033 9280 -30998 10814
rect -30923 10445 -30887 11155
rect -30800 11094 -30663 11106
rect -30800 11060 -30785 11094
rect -30751 11060 -30713 11094
rect -30679 11060 -30663 11094
rect -30800 11048 -30663 11060
rect -30925 10434 -30872 10445
rect -30925 10400 -30918 10434
rect -30884 10400 -30872 10434
rect -30925 10362 -30872 10400
rect -30925 10328 -30918 10362
rect -30884 10328 -30872 10362
rect -30925 10313 -30872 10328
rect -30793 10275 -30753 11048
rect -30909 10268 -30753 10275
rect -30909 10266 -30894 10268
rect -30956 10234 -30894 10266
rect -30860 10234 -30822 10268
rect -30788 10234 -30753 10268
rect -30956 10226 -30753 10234
rect -30909 10222 -30777 10226
rect -29471 10194 -29436 11264
rect -30967 10159 -29436 10194
rect -30967 9411 -30932 10159
rect -25362 9719 -25298 11635
rect -19499 11591 -18870 11686
rect -18965 11106 -18870 11591
rect -18965 11072 -18933 11106
rect -18899 11072 -18870 11106
rect -18965 10657 -18870 11072
rect -17839 11764 -17707 11800
rect -17839 11730 -17825 11764
rect -17791 11730 -17753 11764
rect -17719 11730 -17707 11764
rect -2200 11761 -318 11789
rect -21391 10544 -18869 10657
rect -24500 9734 -24314 9761
rect -24500 9719 -24459 9734
rect -25362 9655 -24459 9719
rect -24500 9628 -24459 9655
rect -24353 9628 -24314 9734
rect -24500 9607 -24314 9628
rect -30967 9395 -30883 9411
rect -30967 9365 -30929 9395
rect -30941 9361 -30929 9365
rect -30895 9361 -30883 9395
rect -30941 9323 -30883 9361
rect -30941 9289 -30929 9323
rect -30895 9289 -30883 9323
rect -33213 4826 -33201 4860
rect -33167 4826 -33152 4860
rect -33213 4788 -33152 4826
rect -33213 4754 -33201 4788
rect -33167 4754 -33152 4788
rect -33388 2200 -33264 2244
rect -33388 2166 -33343 2200
rect -33309 2166 -33264 2200
rect -33388 2121 -33264 2166
rect -33213 1960 -33152 4754
rect -33282 1959 -33152 1960
rect -33099 9019 -33035 9055
rect -33099 8985 -33084 9019
rect -33050 8985 -33035 9019
rect -33099 8947 -33035 8985
rect -33099 8913 -33084 8947
rect -33050 8913 -33035 8947
rect -33099 8875 -33035 8913
rect -33099 8841 -33084 8875
rect -33050 8841 -33035 8875
rect -33099 4779 -33035 8841
rect -33099 4745 -33087 4779
rect -33053 4745 -33035 4779
rect -33099 4707 -33035 4745
rect -33099 4673 -33087 4707
rect -33053 4673 -33035 4707
rect -33282 1926 -33151 1959
rect -33281 1920 -33151 1926
rect -33281 1886 -33236 1920
rect -33202 1886 -33151 1920
rect -33281 1841 -33151 1886
rect -33099 1832 -33035 4673
rect -33101 1660 -33035 1832
rect -33122 1659 -33035 1660
rect -32954 4651 -32894 9279
rect -31038 9264 -30980 9280
rect -30941 9274 -30883 9289
rect -31038 9230 -31026 9264
rect -30992 9230 -30980 9264
rect -31038 9192 -30980 9230
rect -31252 9167 -31194 9183
rect -31252 9133 -31240 9167
rect -31206 9133 -31194 9167
rect -31038 9158 -31026 9192
rect -30992 9158 -30980 9192
rect -31038 9143 -30980 9158
rect -31252 9095 -31194 9133
rect -31252 9061 -31240 9095
rect -31206 9061 -31194 9095
rect -31252 9046 -31194 9061
rect -29326 8268 -29086 8886
rect -26940 8672 -26672 8725
rect -26940 8494 -26850 8672
rect -26744 8494 -26672 8672
rect -26940 8460 -26672 8494
rect -29326 8162 -29272 8268
rect -29166 8162 -29086 8268
rect -29326 8118 -29086 8162
rect -26891 7905 -26703 8460
rect -26935 7853 -26667 7905
rect -26935 7675 -26858 7853
rect -26752 7675 -26667 7853
rect -26935 7640 -26667 7675
rect -29411 6966 -29232 6995
rect -29411 6860 -29375 6966
rect -29269 6860 -29232 6966
rect -29411 6828 -29232 6860
rect -31431 6078 -31373 6094
rect -31431 6044 -31419 6078
rect -31385 6044 -31373 6078
rect -31431 6006 -31373 6044
rect -31431 5972 -31419 6006
rect -31385 5972 -31373 6006
rect -31431 5957 -31373 5972
rect -30515 6077 -30457 6093
rect -30515 6043 -30503 6077
rect -30469 6043 -30457 6077
rect -30515 6005 -30457 6043
rect -30515 5971 -30503 6005
rect -30469 5971 -30457 6005
rect -31627 5568 -31490 5580
rect -31627 5534 -31612 5568
rect -31578 5534 -31540 5568
rect -31506 5534 -31490 5568
rect -31627 5522 -31490 5534
rect -32499 5165 -31695 5188
rect -32499 5059 -32449 5165
rect -31767 5059 -31695 5165
rect -32499 5038 -31695 5059
rect -32954 4617 -32942 4651
rect -32908 4617 -32894 4651
rect -32487 4626 -32400 5038
rect -32307 4626 -32220 5038
rect -32134 4626 -32047 5038
rect -31950 4626 -31863 5038
rect -31825 4626 -31738 5038
rect -33122 1615 -32999 1659
rect -33122 1581 -33077 1615
rect -33043 1581 -32999 1615
rect -33122 1536 -32999 1581
rect -32954 1292 -32894 4617
rect -32712 4581 -31729 4626
rect -32712 4547 -32675 4581
rect -32641 4547 -32603 4581
rect -32569 4547 -32531 4581
rect -32497 4547 -32459 4581
rect -32425 4547 -32387 4581
rect -32353 4547 -32315 4581
rect -32281 4547 -32243 4581
rect -32209 4547 -32171 4581
rect -32137 4547 -32099 4581
rect -32065 4547 -32027 4581
rect -31993 4547 -31955 4581
rect -31921 4547 -31883 4581
rect -31849 4547 -31811 4581
rect -31777 4547 -31729 4581
rect -32712 4511 -31729 4547
rect -31615 4524 -31525 5522
rect -31431 5048 -31396 5957
rect -30515 5956 -30457 5971
rect -31356 5919 -31298 5923
rect -31357 5907 -31298 5919
rect -31357 5873 -31344 5907
rect -31310 5873 -31298 5907
rect -31357 5835 -31298 5873
rect -30740 5917 -30603 5929
rect -30740 5883 -30725 5917
rect -30691 5883 -30653 5917
rect -30619 5883 -30603 5917
rect -30740 5871 -30603 5883
rect -31357 5801 -31344 5835
rect -31310 5801 -31298 5835
rect -31357 5786 -31298 5801
rect -31451 5032 -31393 5048
rect -31451 4998 -31439 5032
rect -31405 4998 -31393 5032
rect -31451 4960 -31393 4998
rect -31357 4969 -31314 5786
rect -31451 4926 -31439 4960
rect -31405 4926 -31393 4960
rect -31451 4911 -31393 4926
rect -31358 4953 -31300 4969
rect -31358 4919 -31346 4953
rect -31312 4919 -31300 4953
rect -31358 4881 -31300 4919
rect -31358 4847 -31346 4881
rect -31312 4847 -31300 4881
rect -31358 4832 -31300 4847
rect -31615 4434 -31298 4524
rect -31388 3967 -31298 4434
rect -31388 3933 -31375 3967
rect -31341 3933 -31298 3967
rect -31388 3895 -31298 3933
rect -30649 3901 -30614 5871
rect -30515 4890 -30480 5956
rect -30438 5905 -30380 5921
rect -30438 5871 -30426 5905
rect -30392 5871 -30380 5905
rect -30438 5833 -30380 5871
rect -29809 5916 -29672 5928
rect -29809 5882 -29794 5916
rect -29760 5882 -29722 5916
rect -29688 5882 -29672 5916
rect -29809 5870 -29672 5882
rect -30438 5799 -30426 5833
rect -30392 5799 -30380 5833
rect -30438 5784 -30380 5799
rect -30537 4874 -30479 4890
rect -30537 4840 -30525 4874
rect -30491 4840 -30479 4874
rect -30537 4802 -30479 4840
rect -30438 4813 -30403 5784
rect -30537 4768 -30525 4802
rect -30491 4768 -30479 4802
rect -30537 4753 -30479 4768
rect -30444 4797 -30386 4813
rect -30444 4763 -30432 4797
rect -30398 4763 -30386 4797
rect -30444 4725 -30386 4763
rect -30444 4691 -30432 4725
rect -30398 4691 -30386 4725
rect -30444 4676 -30386 4691
rect -31388 3861 -31375 3895
rect -31341 3861 -31298 3895
rect -31388 3846 -31298 3861
rect -30657 3885 -30599 3901
rect -30657 3851 -30645 3885
rect -30611 3851 -30599 3885
rect -30657 3813 -30599 3851
rect -30657 3779 -30645 3813
rect -30611 3779 -30599 3813
rect -30657 3764 -30599 3779
rect -30190 3869 -30014 3897
rect -30190 3835 -30154 3869
rect -30120 3835 -30082 3869
rect -30048 3835 -30014 3869
rect -32701 3159 -32658 3506
rect -30190 3328 -30014 3835
rect -29724 3815 -29689 5870
rect -29548 5650 -29431 5695
rect -29548 5616 -29507 5650
rect -29473 5616 -29431 5650
rect -29548 5572 -29431 5616
rect -29647 4288 -29589 4304
rect -29647 4254 -29635 4288
rect -29601 4254 -29589 4288
rect -29647 4216 -29589 4254
rect -29647 4182 -29635 4216
rect -29601 4182 -29589 4216
rect -29647 4167 -29589 4182
rect -29732 3799 -29674 3815
rect -29732 3765 -29720 3799
rect -29686 3765 -29674 3799
rect -29732 3727 -29674 3765
rect -29732 3693 -29720 3727
rect -29686 3693 -29674 3727
rect -29732 3678 -29674 3693
rect -30190 3294 -30156 3328
rect -30122 3294 -30084 3328
rect -30050 3294 -30014 3328
rect -30190 3266 -30014 3294
rect -32751 3113 -32593 3159
rect -29646 3131 -29607 4167
rect -29545 3308 -29453 5572
rect -29384 5064 -29258 6828
rect -26262 6353 -26149 9406
rect -25684 8547 -24047 8723
rect -25996 8275 -25788 8324
rect -25996 8169 -25946 8275
rect -25840 8169 -25788 8275
rect -25996 6115 -25788 8169
rect -25996 6009 -25957 6115
rect -25851 6009 -25788 6115
rect -25996 5928 -25788 6009
rect -29385 5030 -29193 5064
rect -29385 4924 -29341 5030
rect -29235 4924 -29193 5030
rect -29385 4892 -29193 4924
rect -29338 3562 -29284 3886
rect -29368 3511 -29224 3562
rect -29368 3477 -29349 3511
rect -29315 3477 -29277 3511
rect -29243 3477 -29224 3511
rect -29368 3426 -29224 3477
rect -29545 3291 -29407 3308
rect -29545 3185 -29531 3291
rect -29425 3185 -29407 3291
rect -29545 3171 -29407 3185
rect -32751 3079 -32729 3113
rect -32695 3079 -32657 3113
rect -32623 3079 -32593 3113
rect -32751 3043 -32593 3079
rect -29683 3119 -29546 3131
rect -29683 3085 -29668 3119
rect -29634 3085 -29596 3119
rect -29562 3085 -29546 3119
rect -29683 3073 -29546 3085
rect -25684 2928 -25508 8547
rect -25420 7856 -24202 7910
rect -25420 6772 -25366 7856
rect -25420 6708 -25239 6772
rect -19500 6669 -19405 10544
rect -18974 10056 -18798 10101
rect -18974 10022 -18937 10056
rect -18903 10022 -18865 10056
rect -18831 10022 -18798 10056
rect -18974 3586 -18798 10022
rect -17839 6820 -17707 11730
rect -1601 11297 -409 11340
rect -1601 11295 -1031 11297
rect -1601 11261 -1555 11295
rect -1521 11261 -1483 11295
rect -1449 11261 -1411 11295
rect -1377 11261 -1339 11295
rect -1305 11263 -1031 11295
rect -997 11263 -959 11297
rect -925 11263 -887 11297
rect -853 11263 -815 11297
rect -781 11263 -409 11297
rect -1305 11261 -409 11263
rect -1601 11223 -409 11261
rect -1601 11207 -400 11223
rect -1524 11195 -400 11207
rect -1545 11135 -469 11163
rect -1492 11052 -553 11090
rect -1540 10988 -628 11016
rect -1488 10925 -705 10953
rect -1474 10868 -790 10896
rect -1548 10789 -864 10840
rect -1544 10721 -949 10757
rect -1590 10639 -1020 10690
rect -1608 10560 -1116 10611
rect -1501 10303 -1241 10354
rect -1573 9709 -1355 9741
rect -1573 9675 -1554 9709
rect -1520 9675 -1482 9709
rect -1448 9675 -1410 9709
rect -1376 9675 -1355 9709
rect -1573 9652 -1355 9675
rect -1487 9495 -1436 9546
rect -17581 9313 -17397 9329
rect -17581 9279 -17533 9313
rect -17499 9279 -17461 9313
rect -17427 9279 -17397 9313
rect -17581 9266 -17397 9279
rect -17560 9265 -17397 9266
rect -17839 6786 -17788 6820
rect -17754 6786 -17707 6820
rect -18987 3552 -18787 3586
rect -18987 3446 -18935 3552
rect -18829 3446 -18787 3552
rect -18987 3415 -18787 3446
rect -17839 3328 -17707 6786
rect -17572 6689 -17397 6724
rect -17572 6655 -17543 6689
rect -17509 6655 -17471 6689
rect -17437 6655 -17397 6689
rect -17572 6410 -17397 6655
rect -16863 6375 -16768 6516
rect -17350 6280 -16768 6375
rect -1706 6309 -1561 6355
rect -17350 6201 -17255 6280
rect -1706 6275 -1651 6309
rect -1617 6275 -1561 6309
rect -1706 6220 -1561 6275
rect -1474 6232 -1446 9495
rect -17565 6171 -17255 6201
rect -17565 6137 -17529 6171
rect -17495 6137 -17255 6171
rect -17565 6106 -17255 6137
rect -1406 6116 -1378 9652
rect -1507 6088 -1378 6116
rect -1292 5467 -1241 10303
rect -1554 5416 -1241 5467
rect -1292 5345 -1241 5416
rect -1412 5307 -1221 5345
rect -1412 5273 -1370 5307
rect -1336 5273 -1298 5307
rect -1264 5273 -1221 5307
rect -1412 5238 -1221 5273
rect -1167 5210 -1116 10560
rect -1071 6961 -1020 10639
rect -1074 6930 -1015 6961
rect -1074 6896 -1062 6930
rect -1028 6896 -1015 6930
rect -1074 6866 -1015 6896
rect -1989 5201 -1866 5206
rect -1989 5167 -1982 5201
rect -1948 5167 -1908 5201
rect -1874 5167 -1866 5201
rect -1989 5162 -1866 5167
rect -1519 5159 -1116 5210
rect -1071 5131 -1020 6866
rect -1507 5085 -1020 5131
rect -1256 5051 -1108 5057
rect -1256 5049 -1241 5051
rect -1482 5017 -1241 5049
rect -1207 5017 -1167 5051
rect -1133 5049 -1108 5051
rect -985 5049 -949 10721
rect -915 6169 -864 10789
rect -921 6116 -852 6169
rect -921 6082 -904 6116
rect -870 6082 -852 6116
rect -921 6030 -852 6082
rect -1133 5017 -949 5049
rect -1482 5013 -949 5017
rect -1256 5009 -1108 5013
rect -915 4981 -864 6030
rect -1505 4950 -864 4981
rect -1251 4943 -864 4950
rect -1416 4913 -1273 4920
rect -1416 4902 -1404 4913
rect -1494 4879 -1404 4902
rect -1370 4879 -1330 4913
rect -1296 4902 -1273 4913
rect -818 4902 -790 10868
rect -733 7281 -705 10925
rect -753 7237 -689 7281
rect -753 7203 -739 7237
rect -705 7203 -689 7237
rect -753 7163 -689 7203
rect -1296 4879 -790 4902
rect -1494 4874 -790 4879
rect -1416 4873 -1273 4874
rect -733 4845 -705 7163
rect -1494 4817 -705 4845
rect -1542 4782 -1398 4789
rect -656 4782 -628 10988
rect -1542 4748 -1529 4782
rect -1495 4748 -1455 4782
rect -1421 4754 -628 4782
rect -591 9518 -553 11052
rect -591 9505 -541 9518
rect -591 9471 -585 9505
rect -551 9471 -541 9505
rect -591 9431 -541 9471
rect -591 9397 -584 9431
rect -550 9397 -541 9431
rect -591 9385 -541 9397
rect -1421 4748 -1398 4754
rect -1542 4742 -1398 4748
rect -591 4718 -553 9385
rect -1356 4708 -553 4718
rect -1505 4680 -553 4708
rect -1855 4643 -1716 4650
rect -1855 4609 -1839 4643
rect -1805 4609 -1765 4643
rect -1731 4609 -1716 4643
rect -497 4635 -469 11135
rect -1855 4603 -1716 4609
rect -1508 4607 -469 4635
rect -428 4575 -400 11195
rect -1485 4547 -400 4575
rect -1890 4096 -1825 4113
rect -1890 4062 -1882 4096
rect -1848 4062 -1825 4096
rect -1890 4022 -1825 4062
rect -1890 4009 -1882 4022
rect -2292 3988 -1882 4009
rect -1848 4009 -1825 4022
rect -346 4009 -318 11761
rect -1848 3988 -318 4009
rect -2292 3981 -318 3988
rect -1890 3976 -1825 3981
rect -272 3872 -244 11898
rect 5658 11347 6223 11348
rect 5373 11295 6223 11347
rect 5373 11293 6142 11295
rect 5373 11259 5429 11293
rect 5463 11259 5501 11293
rect 5535 11259 5573 11293
rect 5607 11261 6142 11293
rect 6176 11261 6223 11295
rect 5607 11259 6223 11261
rect 5373 11207 6223 11259
rect -2303 3844 -244 3872
rect 18 10702 313 10743
rect 18 10524 79 10702
rect 257 10524 313 10702
rect 18 4509 313 10524
rect 18 4403 38 4509
rect 288 4403 313 4509
rect 18 3453 313 4403
rect -1895 3332 -1834 3343
rect -1777 3339 -1733 3342
rect -17850 3293 -17687 3328
rect -17850 3187 -17822 3293
rect -17716 3187 -17687 3293
rect -17850 3153 -17687 3187
rect -1895 3298 -1881 3332
rect -1847 3298 -1834 3332
rect -1895 3258 -1834 3298
rect -1895 3224 -1881 3258
rect -1847 3224 -1834 3258
rect -25684 2822 -25647 2928
rect -25541 2822 -25508 2928
rect -25684 2808 -25508 2822
rect -32971 1248 -32848 1292
rect -32971 1214 -32926 1248
rect -32892 1214 -32848 1248
rect -32971 1169 -32848 1214
rect -34042 1043 -33829 1090
rect -34042 937 -33995 1043
rect -33889 937 -33829 1043
rect -34042 912 -33829 937
rect -17839 798 -17707 3153
rect -1895 2739 -1834 3224
rect -1786 3334 -1726 3339
rect -1786 3300 -1772 3334
rect -1738 3300 -1726 3334
rect -1786 3260 -1726 3300
rect -1786 3226 -1772 3260
rect -1738 3226 -1726 3260
rect -1948 2695 -1825 2739
rect -1948 2661 -1903 2695
rect -1869 2661 -1825 2695
rect -1948 2616 -1825 2661
rect -1786 2506 -1726 3226
rect -1574 3334 -1513 3342
rect -1574 3300 -1561 3334
rect -1527 3300 -1513 3334
rect -1574 3260 -1513 3300
rect -1574 3226 -1561 3260
rect -1527 3226 -1513 3260
rect -1687 3117 -1626 3196
rect -1687 3083 -1672 3117
rect -1638 3083 -1626 3117
rect -1687 3043 -1626 3083
rect -1687 3009 -1672 3043
rect -1638 3009 -1626 3043
rect -1842 2462 -1719 2506
rect -1842 2428 -1797 2462
rect -1763 2428 -1719 2462
rect -1842 2383 -1719 2428
rect -1687 2249 -1626 3009
rect -1749 2205 -1625 2249
rect -1749 2171 -1704 2205
rect -1670 2171 -1625 2205
rect -1749 2126 -1625 2171
rect -1574 1965 -1513 3226
rect -1643 1964 -1513 1965
rect -1460 3334 -1396 3346
rect -1460 3300 -1446 3334
rect -1412 3300 -1396 3334
rect -1460 3260 -1396 3300
rect -1460 3226 -1446 3260
rect -1412 3226 -1396 3260
rect -1643 1931 -1512 1964
rect -1642 1925 -1512 1931
rect -1642 1891 -1597 1925
rect -1563 1891 -1512 1925
rect -1642 1846 -1512 1891
rect -1460 1837 -1396 3226
rect -1462 1665 -1396 1837
rect -1483 1664 -1396 1665
rect -1315 3341 -1255 3382
rect -1315 3307 -1298 3341
rect -1264 3307 -1255 3341
rect -1315 3267 -1255 3307
rect -1315 3233 -1298 3267
rect -1264 3233 -1255 3267
rect -1483 1620 -1360 1664
rect -1483 1586 -1438 1620
rect -1404 1586 -1360 1620
rect -1483 1541 -1360 1586
rect -1315 1297 -1255 3233
rect -1034 3354 313 3453
rect -1034 3320 -909 3354
rect -875 3320 313 3354
rect -1034 3282 313 3320
rect -1034 3248 -909 3282
rect -875 3248 313 3282
rect -1034 3184 313 3248
rect -1332 1253 -1209 1297
rect -1332 1219 -1287 1253
rect -1253 1219 -1209 1253
rect -1332 1174 -1209 1219
rect 18 1042 313 3184
rect 18 936 42 1042
rect 292 936 313 1042
rect 18 922 313 936
rect 370 10302 570 10328
rect 370 10124 417 10302
rect 523 10124 570 10302
rect 370 4272 570 10124
rect 5603 9749 6430 9772
rect 5603 9715 6361 9749
rect 6395 9715 6430 9749
rect 5603 9712 6430 9715
rect 5603 9678 5659 9712
rect 5693 9678 6430 9712
rect 5603 9677 6430 9678
rect 5603 9643 6361 9677
rect 6395 9643 6430 9677
rect 5603 9621 6430 9643
rect 4921 9497 5019 9526
rect 4921 9463 4954 9497
rect 4988 9463 5019 9497
rect 4921 9425 5019 9463
rect 4921 9391 4954 9425
rect 4988 9391 5019 9425
rect 4921 9362 5019 9391
rect 6833 4440 7096 4504
rect 370 4215 685 4272
rect -17839 783 -17703 798
rect -17839 677 -17826 783
rect -17720 677 -17703 783
rect -17839 662 -17703 677
rect 370 546 570 4215
rect 6968 798 7096 4440
rect 6963 782 7096 798
rect 6963 676 6977 782
rect 7083 676 7096 782
rect 6963 662 7096 676
rect 370 440 421 546
rect 527 440 570 546
rect 370 425 570 440
use 3_INPUT_NOR_MAG  3_INPUT_NOR_MAG_0
timestamp 1717691374
transform 1 0 -32501 0 1 5775
box -80 -736 945 956
use 3AND_MAGIC  3AND_MAGIC_0
timestamp 1717691374
transform -1 0 -31386 0 -1 3692
box -48 -929 1456 459
use 3AND_MAGIC  3AND_MAGIC_1
timestamp 1717691374
transform 1 0 -30797 0 1 9475
box -48 -929 1456 459
use 3AND_MAGIC  3AND_MAGIC_2
timestamp 1717691374
transform 1 0 -32627 0 1 11411
box -48 -929 1456 459
use 7b_counter_new  7b_counter_new_0
timestamp 1717691374
transform 1 0 15673 0 1 4170
box -15678 -4161 62341 11526
use AND_1  AND_1_0
timestamp 1717691374
transform 1 0 -32630 0 1 8683
box -204 -132 1711 1174
use AND_1  AND_1_1
timestamp 1717691374
transform 1 0 -30688 0 1 10592
box -204 -132 1711 1174
use DFF_MAG  DFF_MAG_0
timestamp 1717691374
transform 1 0 3249 0 1 4592
box -2652 -1119 3660 811
use DivideBy2_magic  DivideBy2_magic_0
timestamp 1717691374
transform -1 0 -21649 0 -1 6620
box -2642 -1119 3660 811
use DivideBy2_magic  DivideBy2_magic_1
timestamp 1717691374
transform -1 0 -21649 0 -1 11547
box -2642 -1119 3660 811
use divider_magic  divider_magic_0
timestamp 1717691374
transform 1 0 815 0 1 -5504
box -18550 8609 -2256 18169
use MUX_1  MUX_1_0
timestamp 1717691374
transform 1 0 -29352 0 -1 6248
box -88 -416 3361 2650
use MUX_1  MUX_1_1
timestamp 1717691374
transform 1 0 -24363 0 -1 10272
box -88 -416 3361 2650
use MUX_1  MUX_1_2
timestamp 1717691374
transform 1 0 -29352 0 -1 11248
box -88 -416 3361 2650
use NOR_MAGIC  NOR_MAGIC_0
timestamp 1717691374
transform 1 0 -30394 0 1 6056
box -13 -652 636 681
use NOR_MAGIC  NOR_MAGIC_1
timestamp 1717691374
transform 1 0 -31299 0 1 6057
box -13 -652 636 681
use OR_MAGIC  OR_MAGIC_0
timestamp 1717691374
transform -1 0 -19953 0 1 10306
box -2036 715 -1189 2359
use OR_MAGIC  OR_MAGIC_1
timestamp 1717691374
transform -1 0 -19926 0 1 5372
box -2036 715 -1189 2359
<< labels >>
flabel locali s 2705 735 2705 735 0 FreeSans 4000 0 0 0 P0
flabel locali s -17559 9584 -17559 9584 0 FreeSans 2000 0 0 0 P3
flabel locali s -1654 965 -1654 965 0 FreeSans 4000 0 0 0 CLK
flabel locali s -20972 2881 -20972 2881 0 FreeSans 2000 0 0 0 D2_1
flabel locali s -20420 2656 -20420 2656 0 FreeSans 2000 0 0 0 D2_2
flabel locali s -20056 2417 -20056 2417 0 FreeSans 2000 0 0 0 D2_3
flabel locali s -19654 2167 -19654 2167 0 FreeSans 2000 0 0 0 D2_4
flabel locali s -19393 1879 -19393 1879 0 FreeSans 2000 0 0 0 D2_5
flabel locali s -19051 1591 -19051 1591 0 FreeSans 2000 0 0 0 D2_6
flabel locali s -18643 1211 -18643 1211 0 FreeSans 2000 0 0 0 D2_7
flabel locali s -18758 477 -18758 477 0 FreeSans 2000 0 0 0 LD
flabel locali s -2013 13443 -2013 13443 0 FreeSans 4000 0 0 0 VSS
flabel locali s -3203 14207 -3203 14207 0 FreeSans 4000 0 0 0 VDD
flabel metal1 s 18937 12148 18937 12148 0 FreeSans 4000 0 0 0 Q1
flabel metal1 s 13523 12586 13523 12586 0 FreeSans 4000 0 0 0 Q2
flabel metal1 s 13016 13046 13016 13046 0 FreeSans 4000 0 0 0 Q3
flabel metal1 s 12417 13576 12417 13576 0 FreeSans 4000 0 0 0 Q4
flabel metal1 s 18384 14060 18384 14060 0 FreeSans 4000 0 0 0 Q5
flabel metal1 s 18775 14682 18775 14682 0 FreeSans 4000 0 0 0 Q6
flabel metal1 s 20203 15626 20203 15626 0 FreeSans 4000 0 0 0 Q7
flabel locali s -17649 6672 -17649 6672 0 FreeSans 2000 0 0 0 P2
flabel locali s -31383 7763 -31383 7763 0 FreeSans 2000 0 0 0 OUT1
<< end >>
