magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect -223 -982 -159 -975
rect -3 -998 1159 483
<< pwell >>
rect -90 -2389 1154 -2157
<< psubdiff >>
rect -64 -2222 1128 -2183
rect -64 -2324 22 -2222
rect 1008 -2324 1128 -2222
rect -64 -2363 1128 -2324
<< nsubdiff >>
rect 49 401 1099 447
rect 49 367 124 401
rect 158 367 192 401
rect 226 367 260 401
rect 294 367 328 401
rect 362 367 396 401
rect 430 367 464 401
rect 498 367 532 401
rect 566 367 600 401
rect 634 367 668 401
rect 702 367 736 401
rect 770 367 804 401
rect 838 367 872 401
rect 906 367 940 401
rect 974 367 1099 401
rect 49 315 1099 367
<< psubdiffcont >>
rect 22 -2324 1008 -2222
<< nsubdiffcont >>
rect 124 367 158 401
rect 192 367 226 401
rect 260 367 294 401
rect 328 367 362 401
rect 396 367 430 401
rect 464 367 498 401
rect 532 367 566 401
rect 600 367 634 401
rect 668 367 702 401
rect 736 367 770 401
rect 804 367 838 401
rect 872 367 906 401
rect 940 367 974 401
<< poly >>
rect 91 -69 291 -35
rect 349 -69 549 -36
rect 607 -69 807 -36
rect 865 -69 1065 -36
rect 91 -85 1065 -69
rect 91 -119 109 -85
rect 143 -109 1065 -85
rect 143 -119 560 -109
rect 91 -143 560 -119
rect 594 -113 1065 -109
rect 594 -143 974 -113
rect 91 -147 974 -143
rect 1008 -147 1065 -113
rect 91 -181 1065 -147
rect 91 -237 291 -181
rect 349 -238 549 -181
rect 607 -238 807 -181
rect 865 -238 1065 -181
rect 91 -555 291 -540
rect 91 -589 167 -555
rect 201 -589 291 -555
rect 91 -610 291 -589
rect 90 -957 1065 -862
rect -156 -975 -96 -960
rect -232 -991 -96 -975
rect -232 -1025 -208 -991
rect -174 -1025 -96 -991
rect -232 -1054 -96 -1025
rect -156 -1055 -96 -1054
rect 96 -1323 296 -1292
rect 353 -1323 554 -1292
rect 612 -1323 812 -1292
rect 870 -1323 1070 -1292
rect 96 -1351 1070 -1323
rect 96 -1352 960 -1351
rect 96 -1357 679 -1352
rect 96 -1391 398 -1357
rect 432 -1386 679 -1357
rect 713 -1385 960 -1352
rect 994 -1385 1070 -1351
rect 713 -1386 1070 -1385
rect 432 -1391 1070 -1386
rect 96 -1397 1070 -1391
rect 96 -1440 296 -1397
rect 353 -1440 554 -1397
rect 612 -1440 813 -1397
rect 870 -1440 1070 -1397
rect 96 -1782 1071 -1770
rect 96 -1816 168 -1782
rect 202 -1812 1071 -1782
rect 202 -1816 296 -1812
rect 96 -1840 296 -1816
rect 354 -1840 555 -1812
rect 612 -1840 813 -1812
rect 870 -1840 1071 -1812
<< polycont >>
rect 109 -119 143 -85
rect 560 -143 594 -109
rect 974 -147 1008 -113
rect 167 -589 201 -555
rect -208 -1025 -174 -991
rect 398 -1391 432 -1357
rect 679 -1386 713 -1352
rect 960 -1385 994 -1351
rect 168 -1816 202 -1782
<< locali >>
rect 1751 14982 3341 15029
rect 1751 14876 1950 14982
rect 3280 14876 3341 14982
rect 1751 14839 3341 14876
rect -3 401 1159 483
rect -3 367 124 401
rect 158 367 192 401
rect 226 367 260 401
rect 294 367 328 401
rect 362 367 396 401
rect 430 367 464 401
rect 498 367 532 401
rect 566 367 600 401
rect 634 367 668 401
rect 702 367 736 401
rect 770 367 804 401
rect 838 367 872 401
rect 906 367 940 401
rect 974 367 1159 401
rect -3 355 1159 367
rect -3 321 1235 355
rect -3 290 1159 321
rect 303 171 337 290
rect 819 171 853 290
rect 44 -66 79 -36
rect -317 -85 162 -66
rect -317 -119 109 -85
rect 143 -119 162 -85
rect 561 -88 595 -37
rect 91 -136 162 -119
rect 537 -109 618 -88
rect 537 -143 560 -109
rect 594 -143 618 -109
rect 537 -163 618 -143
rect 951 -107 1032 -92
rect 1077 -107 1111 -36
rect 951 -113 1111 -107
rect 951 -147 974 -113
rect 1008 -141 1111 -113
rect 1008 -147 1032 -141
rect 951 -167 1032 -147
rect 303 -485 337 -439
rect 819 -485 853 -440
rect 150 -552 217 -542
rect -202 -555 217 -552
rect -202 -586 167 -555
rect -202 -770 -168 -586
rect 150 -589 167 -586
rect 201 -589 217 -555
rect 150 -609 217 -589
rect 303 -590 853 -485
rect 303 -632 337 -590
rect 819 -632 853 -590
rect 45 -881 79 -840
rect 561 -881 595 -839
rect 1077 -881 1111 -840
rect 1201 -881 1235 321
rect -84 -915 1235 -881
rect -223 -990 -159 -975
rect -297 -991 -159 -990
rect -297 -1025 -208 -991
rect -174 -1025 -159 -991
rect -297 -1026 -159 -1025
rect -223 -1043 -159 -1026
rect 308 -998 858 -964
rect 308 -1075 342 -998
rect 824 -1062 858 -998
rect 308 -1352 342 -1270
rect -404 -1355 342 -1352
rect 380 -1355 453 -1336
rect 661 -1352 734 -1331
rect 661 -1355 679 -1352
rect -404 -1357 679 -1355
rect -404 -1386 398 -1357
rect 308 -1389 398 -1386
rect 380 -1391 398 -1389
rect 432 -1386 679 -1357
rect 713 -1355 734 -1352
rect 942 -1351 1015 -1330
rect 942 -1355 960 -1351
rect 713 -1385 960 -1355
rect 994 -1385 1015 -1351
rect 713 -1386 1015 -1385
rect 432 -1389 1015 -1386
rect 432 -1391 453 -1389
rect 380 -1414 453 -1391
rect 661 -1409 734 -1389
rect 942 -1408 1015 -1389
rect 308 -1717 342 -1669
rect 824 -1717 858 -1669
rect 308 -1751 858 -1717
rect 152 -1770 218 -1764
rect -430 -1782 218 -1770
rect -430 -1816 168 -1782
rect 202 -1816 218 -1782
rect -430 -1823 218 -1816
rect 152 -1832 218 -1823
rect 308 -1865 342 -1751
rect 824 -1876 858 -1751
rect 50 -2166 84 -2069
rect 566 -2166 600 -2070
rect 1082 -2166 1116 -2069
rect 2294 -2075 7783 -1997
rect -148 -2173 1194 -2166
rect 2294 -2173 2404 -2075
rect -905 -2222 2404 -2173
rect -905 -2324 22 -2222
rect 1008 -2253 2404 -2222
rect 7694 -2253 7783 -2075
rect 1008 -2324 7783 -2253
rect -905 -2330 7783 -2324
rect -905 -2363 3949 -2330
rect -905 -2719 -715 -2363
rect -148 -2385 1194 -2363
rect -1410 -71383 -178 -2719
rect 3404 -79274 29439 -78979
rect 3404 -80028 3772 -79274
rect 29078 -80028 29439 -79274
rect 3404 -80200 29439 -80028
<< viali >>
rect 1950 14876 3280 14982
rect 2404 -2253 7694 -2075
rect 34 -2301 68 -2267
rect 3772 -80028 29078 -79274
<< metal1 >>
rect 1866 14987 3401 15069
rect 1866 14978 1949 14987
rect 1364 14925 1949 14978
rect 1364 -117 1417 14925
rect 1866 14871 1949 14925
rect 3281 14871 3401 14987
rect 1866 14825 3401 14871
rect 39 -127 1443 -117
rect -3766 -163 1443 -127
rect -3766 -173 85 -163
rect -3766 -899 -1443 -173
rect 39 -244 85 -173
rect 555 -236 601 -163
rect 1071 -170 1443 -163
rect 1071 -236 1117 -170
rect -3766 -71546 -2997 -899
rect -208 -1081 -162 -933
rect 44 -1027 1123 -981
rect 44 -1066 90 -1027
rect 560 -1066 607 -1027
rect 1076 -1066 1123 -1027
rect -52 -1149 54 -1091
rect -90 -2179 -44 -1164
rect 44 -1352 1122 -1347
rect 1232 -1352 1278 -170
rect 44 -1393 1278 -1352
rect 44 -1469 90 -1393
rect 560 -1466 606 -1393
rect 1076 -1398 1278 -1393
rect 1076 -1466 1122 -1398
rect 2294 -2042 7783 -1997
rect -90 -2250 125 -2179
rect -100 -2267 125 -2250
rect -100 -2301 34 -2267
rect 68 -2301 125 -2267
rect -100 -2366 125 -2301
rect 2294 -2286 2399 -2042
rect 7699 -2286 7783 -2042
rect 2294 -2330 7783 -2286
rect -3766 -71854 -2429 -71546
rect -2248 -71803 -2120 -71722
rect -1928 -71784 -1755 -71712
rect -1262 -71734 -1089 -71662
rect -1595 -71806 -1422 -71734
rect -942 -71794 -769 -71722
rect -595 -71741 -422 -71669
rect -270 -71795 -97 -71723
rect 70 -71750 243 -71678
rect 385 -71750 558 -71678
rect -3766 -71957 -2997 -71854
rect -2411 -72368 -2283 -72287
rect -2085 -72334 -1957 -72253
rect -1774 -72315 -1601 -72243
rect -1422 -72309 -1249 -72237
rect -1117 -72334 -944 -72262
rect -764 -72348 -591 -72276
rect -440 -72355 -267 -72283
rect -103 -72343 70 -72271
rect 234 -72299 407 -72227
rect 529 -72644 579 -72525
rect -2424 -72857 -2262 -72781
rect -2089 -72833 -1927 -72757
rect -1757 -72826 -1595 -72750
rect -1426 -72809 -1264 -72733
rect -1097 -72812 -935 -72736
rect -766 -72743 -604 -72667
rect -427 -72785 -265 -72709
rect -102 -72726 60 -72650
rect 219 -72740 381 -72664
rect -2265 -73541 -2103 -73465
rect -1937 -73559 -1775 -73483
rect -1585 -73573 -1423 -73497
rect -1284 -73604 -1122 -73528
rect -942 -73600 -780 -73524
rect -589 -73631 -427 -73555
rect -285 -73631 -123 -73555
rect 64 -73614 226 -73538
rect 395 -73624 557 -73548
rect -2459 -73779 -2409 -73662
rect -2254 -73879 -2103 -73806
rect -1913 -73877 -1762 -73804
rect -1597 -73875 -1446 -73802
rect -1261 -73868 -1110 -73795
rect -926 -73877 -775 -73804
rect -594 -73890 -443 -73817
rect -262 -73886 -111 -73813
rect 65 -73870 216 -73797
rect 403 -73866 554 -73793
rect -2418 -74791 -2267 -74718
rect -2086 -74756 -1935 -74683
rect -1763 -74771 -1612 -74698
rect -1437 -74764 -1286 -74691
rect -1090 -74764 -939 -74691
rect -774 -74773 -623 -74700
rect -424 -74773 -273 -74700
rect -97 -74766 54 -74693
rect 222 -74746 373 -74673
rect 529 -74915 579 -74798
rect -2415 -75010 -2235 -74930
rect -2109 -75006 -1929 -74926
rect -1765 -75022 -1585 -74942
rect -1436 -75026 -1256 -74946
rect -1115 -75018 -935 -74938
rect -764 -75022 -584 -74942
rect -439 -75018 -259 -74938
rect -106 -75022 74 -74942
rect 207 -75037 387 -74957
rect -2258 -75874 -2078 -75794
rect -1941 -75870 -1761 -75790
rect -1597 -75874 -1417 -75794
rect -1280 -75885 -1100 -75805
rect -932 -75885 -752 -75805
rect -611 -75889 -431 -75809
rect -290 -75885 -110 -75805
rect 54 -75839 234 -75759
rect 375 -75889 562 -75805
rect -2459 -76051 -2409 -75934
rect -2277 -76180 -2109 -76108
rect -1931 -76180 -1763 -76108
rect -1598 -76192 -1430 -76120
rect -1268 -76168 -1100 -76096
rect -947 -76160 -779 -76088
rect -625 -76156 -457 -76084
rect -268 -76180 -100 -76108
rect 54 -76172 222 -76100
rect 383 -76148 551 -76076
rect -2104 -76971 -1936 -76899
rect -2433 -77047 -2265 -76975
rect -1758 -76999 -1590 -76927
rect -1437 -77003 -1269 -76931
rect -1111 -76975 -943 -76903
rect -778 -76979 -610 -76907
rect -453 -76995 -285 -76923
rect -123 -77023 45 -76951
rect 214 -77011 382 -76939
rect 514 -79178 593 -77031
rect 3404 -79178 29439 -78979
rect 409 -79273 29439 -79178
rect 409 -79274 3791 -79273
rect 29059 -79274 29439 -79273
rect 409 -80028 3772 -79274
rect 29078 -80028 29439 -79274
rect 409 -80029 3791 -80028
rect 29059 -80029 29439 -80028
rect 409 -80046 29439 -80029
rect 3404 -80200 29439 -80046
<< via1 >>
rect 1949 14982 3281 14987
rect 1949 14876 1950 14982
rect 1950 14876 3280 14982
rect 3280 14876 3281 14982
rect 1949 14871 3281 14876
rect 2399 -2075 7699 -2042
rect 2399 -2253 2404 -2075
rect 2404 -2253 7694 -2075
rect 7694 -2253 7699 -2075
rect 2399 -2286 7699 -2253
rect 3791 -79274 29059 -79273
rect 3791 -80028 29059 -79274
rect 3791 -80029 29059 -80028
<< metal2 >>
rect 1866 14997 3401 15069
rect 1866 14861 1947 14997
rect 3283 14861 3401 14997
rect 1866 14825 3401 14861
rect 2294 -2042 7783 -1997
rect 2294 -2286 2399 -2042
rect 7699 -2286 7783 -2042
rect 2294 -2330 7783 -2286
rect 3404 -79263 29439 -78979
rect 3404 -79273 3797 -79263
rect 29053 -79273 29439 -79263
rect 3404 -80029 3791 -79273
rect 29059 -80029 29439 -79273
rect 3404 -80039 3797 -80029
rect 29053 -80039 29439 -80029
rect 3404 -80200 29439 -80039
<< via2 >>
rect 1947 14987 3283 14997
rect 1947 14871 1949 14987
rect 1949 14871 3281 14987
rect 3281 14871 3283 14987
rect 1947 14861 3283 14871
rect 2421 -2272 7677 -2056
rect 3797 -79273 29053 -79263
rect 3797 -80029 29053 -79273
rect 3797 -80039 29053 -80029
<< metal3 >>
rect 1866 15001 3401 15069
rect 1866 14857 1943 15001
rect 3287 14857 3401 15001
rect 1866 14825 3401 14857
rect 2294 -2052 7783 -1997
rect 2294 -2276 2417 -2052
rect 7681 -2276 7783 -2052
rect 2294 -2330 7783 -2276
rect 3404 -79259 29439 -78979
rect 3404 -80043 3793 -79259
rect 29057 -80043 29439 -79259
rect 3404 -80200 29439 -80043
<< via3 >>
rect 1943 14997 3287 15001
rect 1943 14861 1947 14997
rect 1947 14861 3283 14997
rect 3283 14861 3287 14997
rect 1943 14857 3287 14861
rect 2417 -2056 7681 -2052
rect 2417 -2272 2421 -2056
rect 2421 -2272 7677 -2056
rect 7677 -2272 7681 -2056
rect 2417 -2276 7681 -2272
rect 3793 -79263 29057 -79259
rect 3793 -80039 3797 -79263
rect 3797 -80039 29053 -79263
rect 29053 -80039 29057 -79263
rect 3793 -80043 29057 -80039
<< metal4 >>
rect 1809 15001 19858 15106
rect 1809 14857 1943 15001
rect 3287 14857 19858 15001
rect 1809 14815 19858 14857
rect 2747 14651 2851 14815
rect 5359 14651 5463 14815
rect 7971 14651 8075 14815
rect 10583 14651 10687 14815
rect 13195 14651 13299 14815
rect 15807 14651 15911 14815
rect 18419 14651 18523 14815
rect 4027 -1860 4131 -1374
rect 6639 -1860 6743 -1381
rect 9251 -1860 9355 -1381
rect 11863 -1860 11967 -1381
rect 14475 -1860 14579 -1381
rect 17087 -1860 17191 -1372
rect 19699 -1860 19803 -1381
rect 2189 -2052 19803 -1860
rect 2189 -2276 2417 -2052
rect 7681 -2222 19803 -2052
rect 7681 -2276 80252 -2222
rect 2189 -2440 80252 -2276
rect 2453 -3078 80252 -2440
rect 7120 -3292 7224 -3078
rect 12732 -3292 12836 -3078
rect 18344 -3292 18448 -3078
rect 23956 -3292 24060 -3078
rect 29568 -3292 29672 -3078
rect 35180 -3292 35284 -3078
rect 40792 -3292 40896 -3078
rect 46404 -3292 46508 -3078
rect 52016 -3292 52120 -3078
rect 57628 -3292 57732 -3078
rect 63240 -3313 63344 -3078
rect 68852 -3292 68956 -3078
rect 74464 -3292 74568 -3078
rect 80076 -3292 80180 -3078
rect 4340 -78625 4444 -77564
rect 9952 -78625 10056 -77559
rect 15564 -78625 15668 -77537
rect 21176 -78625 21280 -77559
rect 26788 -78625 26892 -77537
rect 32400 -78625 32504 -77564
rect 38012 -78625 38116 -77537
rect 43624 -78625 43728 -77564
rect 49236 -78625 49340 -77559
rect 54848 -78625 54952 -77564
rect 60460 -78625 60564 -77559
rect 66072 -78625 66176 -77563
rect 71684 -78625 71788 -77552
rect 77296 -78625 77400 -77564
rect 1721 -79259 80012 -78625
rect 1721 -80043 3793 -79259
rect 29057 -80043 80012 -79259
rect 1721 -80648 80012 -80043
use sky130_fd_pr__cap_mim_m3_1_6V5NNB  sky130_fd_pr__cap_mim_m3_1_6V5NNB_0
timestamp 1717691374
transform 1 0 10781 0 -1 6635
box -9022 -8120 9022 8120
use sky130_fd_pr__cap_mim_m3_1_FDLZWY  sky130_fd_pr__cap_mim_m3_1_FDLZWY_0
timestamp 1717691374
transform 1 0 41016 0 1 -40428
box -39164 -37240 39164 37240
use sky130_fd_pr__nfet_01v8_lvt_N79YZL  sky130_fd_pr__nfet_01v8_lvt_N79YZL_0
timestamp 1717691374
transform 1 0 583 0 1 -1166
box -571 -126 571 126
use sky130_fd_pr__nfet_01v8_lvt_N79YZL  sky130_fd_pr__nfet_01v8_lvt_N79YZL_1
timestamp 1717691374
transform 1 0 583 0 1 -1566
box -571 -126 571 126
use sky130_fd_pr__nfet_01v8_lvt_N79YZL  sky130_fd_pr__nfet_01v8_lvt_N79YZL_2
timestamp 1717691374
transform 1 0 583 0 1 -1966
box -571 -126 571 126
use sky130_fd_pr__nfet_01v8_Z3KAEG  sky130_fd_pr__nfet_01v8_Z3KAEG_0
timestamp 1717691374
transform 1 0 -126 0 1 -1123
box -114 -68 114 68
use sky130_fd_pr__pfet_01v8_AHD6SB  sky130_fd_pr__pfet_01v8_AHD6SB_0
timestamp 1717691374
transform 1 0 -126 0 1 -854
box -124 -142 124 142
use sky130_fd_pr__pfet_01v8_lvt_KNF787  sky130_fd_pr__pfet_01v8_lvt_KNF787_0
timestamp 1717691374
transform 1 0 578 0 1 67
box -581 -162 581 162
use sky130_fd_pr__pfet_01v8_lvt_KNF787  sky130_fd_pr__pfet_01v8_lvt_KNF787_1
timestamp 1717691374
transform 1 0 578 0 1 -336
box -581 -162 581 162
use sky130_fd_pr__pfet_01v8_lvt_KNF787  sky130_fd_pr__pfet_01v8_lvt_KNF787_2
timestamp 1717691374
transform 1 0 578 0 1 -736
box -581 -162 581 162
use sky130_fd_pr__res_xhigh_po_0p35_APUJRU  sky130_fd_pr__res_xhigh_po_0p35_APUJRU_0
timestamp 1717691374
transform 1 0 -940 0 1 -74289
box -1685 -2944 1685 2944
<< labels >>
flabel locali s 125 -100 125 -100 0 FreeSans 2000 0 0 0 ITAIL
flabel metal1 s -193 -154 -193 -154 0 FreeSans 1000 0 0 0 VCTRL
flabel locali s -275 -1005 -275 -1005 0 FreeSans 1000 0 0 0 UP
flabel locali s -377 -1366 -377 -1366 0 FreeSans 1000 0 0 0 ITAIL1
flabel locali s 523 -2273 523 -2273 0 FreeSans 1000 0 0 0 VSS
flabel locali s 546 385 546 385 0 FreeSans 1000 0 0 0 VDD
flabel locali s -420 -1800 -420 -1800 0 FreeSans 1000 0 0 0 down
<< end >>
