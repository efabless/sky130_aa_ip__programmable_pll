magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< pwell >>
rect -1685 2858 1685 2944
rect -1685 -2858 -1599 2858
rect 1599 -2858 1685 2858
rect -1685 -2944 1685 -2858
<< psubdiff >>
rect -1659 2884 -1547 2918
rect -1513 2884 -1479 2918
rect -1445 2884 -1411 2918
rect -1377 2884 -1343 2918
rect -1309 2884 -1275 2918
rect -1241 2884 -1207 2918
rect -1173 2884 -1139 2918
rect -1105 2884 -1071 2918
rect -1037 2884 -1003 2918
rect -969 2884 -935 2918
rect -901 2884 -867 2918
rect -833 2884 -799 2918
rect -765 2884 -731 2918
rect -697 2884 -663 2918
rect -629 2884 -595 2918
rect -561 2884 -527 2918
rect -493 2884 -459 2918
rect -425 2884 -391 2918
rect -357 2884 -323 2918
rect -289 2884 -255 2918
rect -221 2884 -187 2918
rect -153 2884 -119 2918
rect -85 2884 -51 2918
rect -17 2884 17 2918
rect 51 2884 85 2918
rect 119 2884 153 2918
rect 187 2884 221 2918
rect 255 2884 289 2918
rect 323 2884 357 2918
rect 391 2884 425 2918
rect 459 2884 493 2918
rect 527 2884 561 2918
rect 595 2884 629 2918
rect 663 2884 697 2918
rect 731 2884 765 2918
rect 799 2884 833 2918
rect 867 2884 901 2918
rect 935 2884 969 2918
rect 1003 2884 1037 2918
rect 1071 2884 1105 2918
rect 1139 2884 1173 2918
rect 1207 2884 1241 2918
rect 1275 2884 1309 2918
rect 1343 2884 1377 2918
rect 1411 2884 1445 2918
rect 1479 2884 1513 2918
rect 1547 2884 1659 2918
rect -1659 2805 -1625 2884
rect 1625 2805 1659 2884
rect -1659 2737 -1625 2771
rect -1659 2669 -1625 2703
rect -1659 2601 -1625 2635
rect -1659 2533 -1625 2567
rect -1659 2465 -1625 2499
rect -1659 2397 -1625 2431
rect -1659 2329 -1625 2363
rect -1659 2261 -1625 2295
rect -1659 2193 -1625 2227
rect -1659 2125 -1625 2159
rect -1659 2057 -1625 2091
rect -1659 1989 -1625 2023
rect -1659 1921 -1625 1955
rect -1659 1853 -1625 1887
rect -1659 1785 -1625 1819
rect 1625 2737 1659 2771
rect 1625 2669 1659 2703
rect 1625 2601 1659 2635
rect 1625 2533 1659 2567
rect 1625 2465 1659 2499
rect 1625 2397 1659 2431
rect 1625 2329 1659 2363
rect 1625 2261 1659 2295
rect 1625 2193 1659 2227
rect 1625 2125 1659 2159
rect 1625 2057 1659 2091
rect 1625 1989 1659 2023
rect 1625 1921 1659 1955
rect 1625 1853 1659 1887
rect 1625 1785 1659 1819
rect -1659 1717 -1625 1751
rect -1659 1649 -1625 1683
rect 1625 1717 1659 1751
rect -1659 1581 -1625 1615
rect -1659 1513 -1625 1547
rect -1659 1445 -1625 1479
rect -1659 1377 -1625 1411
rect -1659 1309 -1625 1343
rect -1659 1241 -1625 1275
rect -1659 1173 -1625 1207
rect -1659 1105 -1625 1139
rect -1659 1037 -1625 1071
rect -1659 969 -1625 1003
rect -1659 901 -1625 935
rect -1659 833 -1625 867
rect -1659 765 -1625 799
rect -1659 697 -1625 731
rect -1659 629 -1625 663
rect 1625 1649 1659 1683
rect 1625 1581 1659 1615
rect 1625 1513 1659 1547
rect 1625 1445 1659 1479
rect 1625 1377 1659 1411
rect 1625 1309 1659 1343
rect 1625 1241 1659 1275
rect 1625 1173 1659 1207
rect 1625 1105 1659 1139
rect 1625 1037 1659 1071
rect 1625 969 1659 1003
rect 1625 901 1659 935
rect 1625 833 1659 867
rect 1625 765 1659 799
rect 1625 697 1659 731
rect 1625 629 1659 663
rect -1659 561 -1625 595
rect -1659 493 -1625 527
rect 1625 561 1659 595
rect -1659 425 -1625 459
rect -1659 357 -1625 391
rect -1659 289 -1625 323
rect -1659 221 -1625 255
rect -1659 153 -1625 187
rect -1659 85 -1625 119
rect -1659 17 -1625 51
rect -1659 -51 -1625 -17
rect -1659 -119 -1625 -85
rect -1659 -187 -1625 -153
rect -1659 -255 -1625 -221
rect -1659 -323 -1625 -289
rect -1659 -391 -1625 -357
rect -1659 -459 -1625 -425
rect -1659 -527 -1625 -493
rect 1625 493 1659 527
rect 1625 425 1659 459
rect 1625 357 1659 391
rect 1625 289 1659 323
rect 1625 221 1659 255
rect 1625 153 1659 187
rect 1625 85 1659 119
rect 1625 17 1659 51
rect 1625 -51 1659 -17
rect 1625 -119 1659 -85
rect 1625 -187 1659 -153
rect 1625 -255 1659 -221
rect 1625 -323 1659 -289
rect 1625 -391 1659 -357
rect 1625 -459 1659 -425
rect -1659 -595 -1625 -561
rect 1625 -527 1659 -493
rect 1625 -595 1659 -561
rect -1659 -663 -1625 -629
rect -1659 -731 -1625 -697
rect -1659 -799 -1625 -765
rect -1659 -867 -1625 -833
rect -1659 -935 -1625 -901
rect -1659 -1003 -1625 -969
rect -1659 -1071 -1625 -1037
rect -1659 -1139 -1625 -1105
rect -1659 -1207 -1625 -1173
rect -1659 -1275 -1625 -1241
rect -1659 -1343 -1625 -1309
rect -1659 -1411 -1625 -1377
rect -1659 -1479 -1625 -1445
rect -1659 -1547 -1625 -1513
rect -1659 -1615 -1625 -1581
rect -1659 -1683 -1625 -1649
rect 1625 -663 1659 -629
rect 1625 -731 1659 -697
rect 1625 -799 1659 -765
rect 1625 -867 1659 -833
rect 1625 -935 1659 -901
rect 1625 -1003 1659 -969
rect 1625 -1071 1659 -1037
rect 1625 -1139 1659 -1105
rect 1625 -1207 1659 -1173
rect 1625 -1275 1659 -1241
rect 1625 -1343 1659 -1309
rect 1625 -1411 1659 -1377
rect 1625 -1479 1659 -1445
rect 1625 -1547 1659 -1513
rect 1625 -1615 1659 -1581
rect -1659 -1751 -1625 -1717
rect 1625 -1683 1659 -1649
rect 1625 -1751 1659 -1717
rect -1659 -1819 -1625 -1785
rect -1659 -1887 -1625 -1853
rect -1659 -1955 -1625 -1921
rect -1659 -2023 -1625 -1989
rect -1659 -2091 -1625 -2057
rect -1659 -2159 -1625 -2125
rect -1659 -2227 -1625 -2193
rect -1659 -2295 -1625 -2261
rect -1659 -2363 -1625 -2329
rect -1659 -2431 -1625 -2397
rect -1659 -2499 -1625 -2465
rect -1659 -2567 -1625 -2533
rect -1659 -2635 -1625 -2601
rect -1659 -2703 -1625 -2669
rect -1659 -2771 -1625 -2737
rect 1625 -1819 1659 -1785
rect 1625 -1887 1659 -1853
rect 1625 -1955 1659 -1921
rect 1625 -2023 1659 -1989
rect 1625 -2091 1659 -2057
rect 1625 -2159 1659 -2125
rect 1625 -2227 1659 -2193
rect 1625 -2295 1659 -2261
rect 1625 -2363 1659 -2329
rect 1625 -2431 1659 -2397
rect 1625 -2499 1659 -2465
rect 1625 -2567 1659 -2533
rect 1625 -2635 1659 -2601
rect 1625 -2703 1659 -2669
rect 1625 -2771 1659 -2737
rect -1659 -2884 -1625 -2805
rect 1625 -2884 1659 -2805
rect -1659 -2918 -1547 -2884
rect -1513 -2918 -1479 -2884
rect -1445 -2918 -1411 -2884
rect -1377 -2918 -1343 -2884
rect -1309 -2918 -1275 -2884
rect -1241 -2918 -1207 -2884
rect -1173 -2918 -1139 -2884
rect -1105 -2918 -1071 -2884
rect -1037 -2918 -1003 -2884
rect -969 -2918 -935 -2884
rect -901 -2918 -867 -2884
rect -833 -2918 -799 -2884
rect -765 -2918 -731 -2884
rect -697 -2918 -663 -2884
rect -629 -2918 -595 -2884
rect -561 -2918 -527 -2884
rect -493 -2918 -459 -2884
rect -425 -2918 -391 -2884
rect -357 -2918 -323 -2884
rect -289 -2918 -255 -2884
rect -221 -2918 -187 -2884
rect -153 -2918 -119 -2884
rect -85 -2918 -51 -2884
rect -17 -2918 17 -2884
rect 51 -2918 85 -2884
rect 119 -2918 153 -2884
rect 187 -2918 221 -2884
rect 255 -2918 289 -2884
rect 323 -2918 357 -2884
rect 391 -2918 425 -2884
rect 459 -2918 493 -2884
rect 527 -2918 561 -2884
rect 595 -2918 629 -2884
rect 663 -2918 697 -2884
rect 731 -2918 765 -2884
rect 799 -2918 833 -2884
rect 867 -2918 901 -2884
rect 935 -2918 969 -2884
rect 1003 -2918 1037 -2884
rect 1071 -2918 1105 -2884
rect 1139 -2918 1173 -2884
rect 1207 -2918 1241 -2884
rect 1275 -2918 1309 -2884
rect 1343 -2918 1377 -2884
rect 1411 -2918 1445 -2884
rect 1479 -2918 1513 -2884
rect 1547 -2918 1659 -2884
<< psubdiffcont >>
rect -1547 2884 -1513 2918
rect -1479 2884 -1445 2918
rect -1411 2884 -1377 2918
rect -1343 2884 -1309 2918
rect -1275 2884 -1241 2918
rect -1207 2884 -1173 2918
rect -1139 2884 -1105 2918
rect -1071 2884 -1037 2918
rect -1003 2884 -969 2918
rect -935 2884 -901 2918
rect -867 2884 -833 2918
rect -799 2884 -765 2918
rect -731 2884 -697 2918
rect -663 2884 -629 2918
rect -595 2884 -561 2918
rect -527 2884 -493 2918
rect -459 2884 -425 2918
rect -391 2884 -357 2918
rect -323 2884 -289 2918
rect -255 2884 -221 2918
rect -187 2884 -153 2918
rect -119 2884 -85 2918
rect -51 2884 -17 2918
rect 17 2884 51 2918
rect 85 2884 119 2918
rect 153 2884 187 2918
rect 221 2884 255 2918
rect 289 2884 323 2918
rect 357 2884 391 2918
rect 425 2884 459 2918
rect 493 2884 527 2918
rect 561 2884 595 2918
rect 629 2884 663 2918
rect 697 2884 731 2918
rect 765 2884 799 2918
rect 833 2884 867 2918
rect 901 2884 935 2918
rect 969 2884 1003 2918
rect 1037 2884 1071 2918
rect 1105 2884 1139 2918
rect 1173 2884 1207 2918
rect 1241 2884 1275 2918
rect 1309 2884 1343 2918
rect 1377 2884 1411 2918
rect 1445 2884 1479 2918
rect 1513 2884 1547 2918
rect -1659 2771 -1625 2805
rect -1659 2703 -1625 2737
rect -1659 2635 -1625 2669
rect -1659 2567 -1625 2601
rect -1659 2499 -1625 2533
rect -1659 2431 -1625 2465
rect -1659 2363 -1625 2397
rect -1659 2295 -1625 2329
rect -1659 2227 -1625 2261
rect -1659 2159 -1625 2193
rect -1659 2091 -1625 2125
rect -1659 2023 -1625 2057
rect -1659 1955 -1625 1989
rect -1659 1887 -1625 1921
rect -1659 1819 -1625 1853
rect -1659 1751 -1625 1785
rect 1625 2771 1659 2805
rect 1625 2703 1659 2737
rect 1625 2635 1659 2669
rect 1625 2567 1659 2601
rect 1625 2499 1659 2533
rect 1625 2431 1659 2465
rect 1625 2363 1659 2397
rect 1625 2295 1659 2329
rect 1625 2227 1659 2261
rect 1625 2159 1659 2193
rect 1625 2091 1659 2125
rect 1625 2023 1659 2057
rect 1625 1955 1659 1989
rect 1625 1887 1659 1921
rect 1625 1819 1659 1853
rect -1659 1683 -1625 1717
rect 1625 1751 1659 1785
rect 1625 1683 1659 1717
rect -1659 1615 -1625 1649
rect -1659 1547 -1625 1581
rect -1659 1479 -1625 1513
rect -1659 1411 -1625 1445
rect -1659 1343 -1625 1377
rect -1659 1275 -1625 1309
rect -1659 1207 -1625 1241
rect -1659 1139 -1625 1173
rect -1659 1071 -1625 1105
rect -1659 1003 -1625 1037
rect -1659 935 -1625 969
rect -1659 867 -1625 901
rect -1659 799 -1625 833
rect -1659 731 -1625 765
rect -1659 663 -1625 697
rect -1659 595 -1625 629
rect 1625 1615 1659 1649
rect 1625 1547 1659 1581
rect 1625 1479 1659 1513
rect 1625 1411 1659 1445
rect 1625 1343 1659 1377
rect 1625 1275 1659 1309
rect 1625 1207 1659 1241
rect 1625 1139 1659 1173
rect 1625 1071 1659 1105
rect 1625 1003 1659 1037
rect 1625 935 1659 969
rect 1625 867 1659 901
rect 1625 799 1659 833
rect 1625 731 1659 765
rect 1625 663 1659 697
rect -1659 527 -1625 561
rect 1625 595 1659 629
rect 1625 527 1659 561
rect -1659 459 -1625 493
rect -1659 391 -1625 425
rect -1659 323 -1625 357
rect -1659 255 -1625 289
rect -1659 187 -1625 221
rect -1659 119 -1625 153
rect -1659 51 -1625 85
rect -1659 -17 -1625 17
rect -1659 -85 -1625 -51
rect -1659 -153 -1625 -119
rect -1659 -221 -1625 -187
rect -1659 -289 -1625 -255
rect -1659 -357 -1625 -323
rect -1659 -425 -1625 -391
rect -1659 -493 -1625 -459
rect 1625 459 1659 493
rect 1625 391 1659 425
rect 1625 323 1659 357
rect 1625 255 1659 289
rect 1625 187 1659 221
rect 1625 119 1659 153
rect 1625 51 1659 85
rect 1625 -17 1659 17
rect 1625 -85 1659 -51
rect 1625 -153 1659 -119
rect 1625 -221 1659 -187
rect 1625 -289 1659 -255
rect 1625 -357 1659 -323
rect 1625 -425 1659 -391
rect 1625 -493 1659 -459
rect -1659 -561 -1625 -527
rect -1659 -629 -1625 -595
rect 1625 -561 1659 -527
rect -1659 -697 -1625 -663
rect -1659 -765 -1625 -731
rect -1659 -833 -1625 -799
rect -1659 -901 -1625 -867
rect -1659 -969 -1625 -935
rect -1659 -1037 -1625 -1003
rect -1659 -1105 -1625 -1071
rect -1659 -1173 -1625 -1139
rect -1659 -1241 -1625 -1207
rect -1659 -1309 -1625 -1275
rect -1659 -1377 -1625 -1343
rect -1659 -1445 -1625 -1411
rect -1659 -1513 -1625 -1479
rect -1659 -1581 -1625 -1547
rect -1659 -1649 -1625 -1615
rect 1625 -629 1659 -595
rect 1625 -697 1659 -663
rect 1625 -765 1659 -731
rect 1625 -833 1659 -799
rect 1625 -901 1659 -867
rect 1625 -969 1659 -935
rect 1625 -1037 1659 -1003
rect 1625 -1105 1659 -1071
rect 1625 -1173 1659 -1139
rect 1625 -1241 1659 -1207
rect 1625 -1309 1659 -1275
rect 1625 -1377 1659 -1343
rect 1625 -1445 1659 -1411
rect 1625 -1513 1659 -1479
rect 1625 -1581 1659 -1547
rect 1625 -1649 1659 -1615
rect -1659 -1717 -1625 -1683
rect -1659 -1785 -1625 -1751
rect 1625 -1717 1659 -1683
rect -1659 -1853 -1625 -1819
rect -1659 -1921 -1625 -1887
rect -1659 -1989 -1625 -1955
rect -1659 -2057 -1625 -2023
rect -1659 -2125 -1625 -2091
rect -1659 -2193 -1625 -2159
rect -1659 -2261 -1625 -2227
rect -1659 -2329 -1625 -2295
rect -1659 -2397 -1625 -2363
rect -1659 -2465 -1625 -2431
rect -1659 -2533 -1625 -2499
rect -1659 -2601 -1625 -2567
rect -1659 -2669 -1625 -2635
rect -1659 -2737 -1625 -2703
rect -1659 -2805 -1625 -2771
rect 1625 -1785 1659 -1751
rect 1625 -1853 1659 -1819
rect 1625 -1921 1659 -1887
rect 1625 -1989 1659 -1955
rect 1625 -2057 1659 -2023
rect 1625 -2125 1659 -2091
rect 1625 -2193 1659 -2159
rect 1625 -2261 1659 -2227
rect 1625 -2329 1659 -2295
rect 1625 -2397 1659 -2363
rect 1625 -2465 1659 -2431
rect 1625 -2533 1659 -2499
rect 1625 -2601 1659 -2567
rect 1625 -2669 1659 -2635
rect 1625 -2737 1659 -2703
rect 1625 -2805 1659 -2771
rect -1547 -2918 -1513 -2884
rect -1479 -2918 -1445 -2884
rect -1411 -2918 -1377 -2884
rect -1343 -2918 -1309 -2884
rect -1275 -2918 -1241 -2884
rect -1207 -2918 -1173 -2884
rect -1139 -2918 -1105 -2884
rect -1071 -2918 -1037 -2884
rect -1003 -2918 -969 -2884
rect -935 -2918 -901 -2884
rect -867 -2918 -833 -2884
rect -799 -2918 -765 -2884
rect -731 -2918 -697 -2884
rect -663 -2918 -629 -2884
rect -595 -2918 -561 -2884
rect -527 -2918 -493 -2884
rect -459 -2918 -425 -2884
rect -391 -2918 -357 -2884
rect -323 -2918 -289 -2884
rect -255 -2918 -221 -2884
rect -187 -2918 -153 -2884
rect -119 -2918 -85 -2884
rect -51 -2918 -17 -2884
rect 17 -2918 51 -2884
rect 85 -2918 119 -2884
rect 153 -2918 187 -2884
rect 221 -2918 255 -2884
rect 289 -2918 323 -2884
rect 357 -2918 391 -2884
rect 425 -2918 459 -2884
rect 493 -2918 527 -2884
rect 561 -2918 595 -2884
rect 629 -2918 663 -2884
rect 697 -2918 731 -2884
rect 765 -2918 799 -2884
rect 833 -2918 867 -2884
rect 901 -2918 935 -2884
rect 969 -2918 1003 -2884
rect 1037 -2918 1071 -2884
rect 1105 -2918 1139 -2884
rect 1173 -2918 1207 -2884
rect 1241 -2918 1275 -2884
rect 1309 -2918 1343 -2884
rect 1377 -2918 1411 -2884
rect 1445 -2918 1479 -2884
rect 1513 -2918 1547 -2884
<< xpolycontact >>
rect -1529 2356 -1459 2788
rect -1529 1756 -1459 2188
rect -1363 2356 -1293 2788
rect -1363 1756 -1293 2188
rect -1197 2356 -1127 2788
rect -1197 1756 -1127 2188
rect -1031 2356 -961 2788
rect -1031 1756 -961 2188
rect -865 2356 -795 2788
rect -865 1756 -795 2188
rect -699 2356 -629 2788
rect -699 1756 -629 2188
rect -533 2356 -463 2788
rect -533 1756 -463 2188
rect -367 2356 -297 2788
rect -367 1756 -297 2188
rect -201 2356 -131 2788
rect -201 1756 -131 2188
rect -35 2356 35 2788
rect -35 1756 35 2188
rect 131 2356 201 2788
rect 131 1756 201 2188
rect 297 2356 367 2788
rect 297 1756 367 2188
rect 463 2356 533 2788
rect 463 1756 533 2188
rect 629 2356 699 2788
rect 629 1756 699 2188
rect 795 2356 865 2788
rect 795 1756 865 2188
rect 961 2356 1031 2788
rect 961 1756 1031 2188
rect 1127 2356 1197 2788
rect 1127 1756 1197 2188
rect 1293 2356 1363 2788
rect 1293 1756 1363 2188
rect 1459 2356 1529 2788
rect 1459 1756 1529 2188
rect -1529 1220 -1459 1652
rect -1529 620 -1459 1052
rect -1363 1220 -1293 1652
rect -1363 620 -1293 1052
rect -1197 1220 -1127 1652
rect -1197 620 -1127 1052
rect -1031 1220 -961 1652
rect -1031 620 -961 1052
rect -865 1220 -795 1652
rect -865 620 -795 1052
rect -699 1220 -629 1652
rect -699 620 -629 1052
rect -533 1220 -463 1652
rect -533 620 -463 1052
rect -367 1220 -297 1652
rect -367 620 -297 1052
rect -201 1220 -131 1652
rect -201 620 -131 1052
rect -35 1220 35 1652
rect -35 620 35 1052
rect 131 1220 201 1652
rect 131 620 201 1052
rect 297 1220 367 1652
rect 297 620 367 1052
rect 463 1220 533 1652
rect 463 620 533 1052
rect 629 1220 699 1652
rect 629 620 699 1052
rect 795 1220 865 1652
rect 795 620 865 1052
rect 961 1220 1031 1652
rect 961 620 1031 1052
rect 1127 1220 1197 1652
rect 1127 620 1197 1052
rect 1293 1220 1363 1652
rect 1293 620 1363 1052
rect 1459 1220 1529 1652
rect 1459 620 1529 1052
rect -1529 84 -1459 516
rect -1529 -516 -1459 -84
rect -1363 84 -1293 516
rect -1363 -516 -1293 -84
rect -1197 84 -1127 516
rect -1197 -516 -1127 -84
rect -1031 84 -961 516
rect -1031 -516 -961 -84
rect -865 84 -795 516
rect -865 -516 -795 -84
rect -699 84 -629 516
rect -699 -516 -629 -84
rect -533 84 -463 516
rect -533 -516 -463 -84
rect -367 84 -297 516
rect -367 -516 -297 -84
rect -201 84 -131 516
rect -201 -516 -131 -84
rect -35 84 35 516
rect -35 -516 35 -84
rect 131 84 201 516
rect 131 -516 201 -84
rect 297 84 367 516
rect 297 -516 367 -84
rect 463 84 533 516
rect 463 -516 533 -84
rect 629 84 699 516
rect 629 -516 699 -84
rect 795 84 865 516
rect 795 -516 865 -84
rect 961 84 1031 516
rect 961 -516 1031 -84
rect 1127 84 1197 516
rect 1127 -516 1197 -84
rect 1293 84 1363 516
rect 1293 -516 1363 -84
rect 1459 84 1529 516
rect 1459 -516 1529 -84
rect -1529 -1052 -1459 -620
rect -1529 -1652 -1459 -1220
rect -1363 -1052 -1293 -620
rect -1363 -1652 -1293 -1220
rect -1197 -1052 -1127 -620
rect -1197 -1652 -1127 -1220
rect -1031 -1052 -961 -620
rect -1031 -1652 -961 -1220
rect -865 -1052 -795 -620
rect -865 -1652 -795 -1220
rect -699 -1052 -629 -620
rect -699 -1652 -629 -1220
rect -533 -1052 -463 -620
rect -533 -1652 -463 -1220
rect -367 -1052 -297 -620
rect -367 -1652 -297 -1220
rect -201 -1052 -131 -620
rect -201 -1652 -131 -1220
rect -35 -1052 35 -620
rect -35 -1652 35 -1220
rect 131 -1052 201 -620
rect 131 -1652 201 -1220
rect 297 -1052 367 -620
rect 297 -1652 367 -1220
rect 463 -1052 533 -620
rect 463 -1652 533 -1220
rect 629 -1052 699 -620
rect 629 -1652 699 -1220
rect 795 -1052 865 -620
rect 795 -1652 865 -1220
rect 961 -1052 1031 -620
rect 961 -1652 1031 -1220
rect 1127 -1052 1197 -620
rect 1127 -1652 1197 -1220
rect 1293 -1052 1363 -620
rect 1293 -1652 1363 -1220
rect 1459 -1052 1529 -620
rect 1459 -1652 1529 -1220
rect -1529 -2188 -1459 -1756
rect -1529 -2788 -1459 -2356
rect -1363 -2188 -1293 -1756
rect -1363 -2788 -1293 -2356
rect -1197 -2188 -1127 -1756
rect -1197 -2788 -1127 -2356
rect -1031 -2188 -961 -1756
rect -1031 -2788 -961 -2356
rect -865 -2188 -795 -1756
rect -865 -2788 -795 -2356
rect -699 -2188 -629 -1756
rect -699 -2788 -629 -2356
rect -533 -2188 -463 -1756
rect -533 -2788 -463 -2356
rect -367 -2188 -297 -1756
rect -367 -2788 -297 -2356
rect -201 -2188 -131 -1756
rect -201 -2788 -131 -2356
rect -35 -2188 35 -1756
rect -35 -2788 35 -2356
rect 131 -2188 201 -1756
rect 131 -2788 201 -2356
rect 297 -2188 367 -1756
rect 297 -2788 367 -2356
rect 463 -2188 533 -1756
rect 463 -2788 533 -2356
rect 629 -2188 699 -1756
rect 629 -2788 699 -2356
rect 795 -2188 865 -1756
rect 795 -2788 865 -2356
rect 961 -2188 1031 -1756
rect 961 -2788 1031 -2356
rect 1127 -2188 1197 -1756
rect 1127 -2788 1197 -2356
rect 1293 -2188 1363 -1756
rect 1293 -2788 1363 -2356
rect 1459 -2188 1529 -1756
rect 1459 -2788 1529 -2356
<< xpolyres >>
rect -1529 2188 -1459 2356
rect -1363 2188 -1293 2356
rect -1197 2188 -1127 2356
rect -1031 2188 -961 2356
rect -865 2188 -795 2356
rect -699 2188 -629 2356
rect -533 2188 -463 2356
rect -367 2188 -297 2356
rect -201 2188 -131 2356
rect -35 2188 35 2356
rect 131 2188 201 2356
rect 297 2188 367 2356
rect 463 2188 533 2356
rect 629 2188 699 2356
rect 795 2188 865 2356
rect 961 2188 1031 2356
rect 1127 2188 1197 2356
rect 1293 2188 1363 2356
rect 1459 2188 1529 2356
rect -1529 1052 -1459 1220
rect -1363 1052 -1293 1220
rect -1197 1052 -1127 1220
rect -1031 1052 -961 1220
rect -865 1052 -795 1220
rect -699 1052 -629 1220
rect -533 1052 -463 1220
rect -367 1052 -297 1220
rect -201 1052 -131 1220
rect -35 1052 35 1220
rect 131 1052 201 1220
rect 297 1052 367 1220
rect 463 1052 533 1220
rect 629 1052 699 1220
rect 795 1052 865 1220
rect 961 1052 1031 1220
rect 1127 1052 1197 1220
rect 1293 1052 1363 1220
rect 1459 1052 1529 1220
rect -1529 -84 -1459 84
rect -1363 -84 -1293 84
rect -1197 -84 -1127 84
rect -1031 -84 -961 84
rect -865 -84 -795 84
rect -699 -84 -629 84
rect -533 -84 -463 84
rect -367 -84 -297 84
rect -201 -84 -131 84
rect -35 -84 35 84
rect 131 -84 201 84
rect 297 -84 367 84
rect 463 -84 533 84
rect 629 -84 699 84
rect 795 -84 865 84
rect 961 -84 1031 84
rect 1127 -84 1197 84
rect 1293 -84 1363 84
rect 1459 -84 1529 84
rect -1529 -1220 -1459 -1052
rect -1363 -1220 -1293 -1052
rect -1197 -1220 -1127 -1052
rect -1031 -1220 -961 -1052
rect -865 -1220 -795 -1052
rect -699 -1220 -629 -1052
rect -533 -1220 -463 -1052
rect -367 -1220 -297 -1052
rect -201 -1220 -131 -1052
rect -35 -1220 35 -1052
rect 131 -1220 201 -1052
rect 297 -1220 367 -1052
rect 463 -1220 533 -1052
rect 629 -1220 699 -1052
rect 795 -1220 865 -1052
rect 961 -1220 1031 -1052
rect 1127 -1220 1197 -1052
rect 1293 -1220 1363 -1052
rect 1459 -1220 1529 -1052
rect -1529 -2356 -1459 -2188
rect -1363 -2356 -1293 -2188
rect -1197 -2356 -1127 -2188
rect -1031 -2356 -961 -2188
rect -865 -2356 -795 -2188
rect -699 -2356 -629 -2188
rect -533 -2356 -463 -2188
rect -367 -2356 -297 -2188
rect -201 -2356 -131 -2188
rect -35 -2356 35 -2188
rect 131 -2356 201 -2188
rect 297 -2356 367 -2188
rect 463 -2356 533 -2188
rect 629 -2356 699 -2188
rect 795 -2356 865 -2188
rect 961 -2356 1031 -2188
rect 1127 -2356 1197 -2188
rect 1293 -2356 1363 -2188
rect 1459 -2356 1529 -2188
<< locali >>
rect -1659 2884 -1547 2918
rect -1513 2884 -1479 2918
rect -1445 2884 -1411 2918
rect -1377 2884 -1343 2918
rect -1309 2884 -1275 2918
rect -1241 2884 -1207 2918
rect -1173 2884 -1139 2918
rect -1105 2884 -1071 2918
rect -1037 2884 -1003 2918
rect -969 2884 -935 2918
rect -901 2884 -867 2918
rect -833 2884 -799 2918
rect -765 2884 -731 2918
rect -697 2884 -663 2918
rect -629 2884 -595 2918
rect -561 2884 -527 2918
rect -493 2884 -459 2918
rect -425 2884 -391 2918
rect -357 2884 -323 2918
rect -289 2884 -255 2918
rect -221 2884 -187 2918
rect -153 2884 -119 2918
rect -85 2884 -51 2918
rect -17 2884 17 2918
rect 51 2884 85 2918
rect 119 2884 153 2918
rect 187 2884 221 2918
rect 255 2884 289 2918
rect 323 2884 357 2918
rect 391 2884 425 2918
rect 459 2884 493 2918
rect 527 2884 561 2918
rect 595 2884 629 2918
rect 663 2884 697 2918
rect 731 2884 765 2918
rect 799 2884 833 2918
rect 867 2884 901 2918
rect 935 2884 969 2918
rect 1003 2884 1037 2918
rect 1071 2884 1105 2918
rect 1139 2884 1173 2918
rect 1207 2884 1241 2918
rect 1275 2884 1309 2918
rect 1343 2884 1377 2918
rect 1411 2884 1445 2918
rect 1479 2884 1513 2918
rect 1547 2884 1659 2918
rect -1659 2805 -1625 2884
rect 1625 2805 1659 2884
rect -1659 2737 -1625 2771
rect -1659 2669 -1625 2703
rect -1659 2601 -1625 2635
rect -1659 2533 -1625 2567
rect -1659 2465 -1625 2499
rect -1659 2397 -1625 2431
rect -1659 2329 -1625 2363
rect 1625 2737 1659 2771
rect 1625 2669 1659 2703
rect 1625 2601 1659 2635
rect 1625 2533 1659 2567
rect 1625 2465 1659 2499
rect 1625 2397 1659 2431
rect -1659 2261 -1625 2295
rect -1659 2193 -1625 2227
rect 1625 2329 1659 2363
rect 1625 2261 1659 2295
rect 1625 2193 1659 2227
rect -1659 2125 -1625 2159
rect -1659 2057 -1625 2091
rect -1659 1989 -1625 2023
rect -1659 1921 -1625 1955
rect -1659 1853 -1625 1887
rect -1659 1785 -1625 1819
rect 1625 2125 1659 2159
rect 1625 2057 1659 2091
rect 1625 1989 1659 2023
rect 1625 1921 1659 1955
rect 1625 1853 1659 1887
rect 1625 1785 1659 1819
rect -1659 1717 -1625 1751
rect -1659 1649 -1625 1683
rect 1625 1717 1659 1751
rect -1659 1581 -1625 1615
rect -1659 1513 -1625 1547
rect -1659 1445 -1625 1479
rect -1659 1377 -1625 1411
rect -1659 1309 -1625 1343
rect -1659 1241 -1625 1275
rect 1625 1649 1659 1683
rect 1625 1581 1659 1615
rect 1625 1513 1659 1547
rect 1625 1445 1659 1479
rect 1625 1377 1659 1411
rect 1625 1309 1659 1343
rect 1625 1241 1659 1275
rect -1659 1173 -1625 1207
rect -1659 1105 -1625 1139
rect -1659 1037 -1625 1071
rect 1625 1173 1659 1207
rect 1625 1105 1659 1139
rect -1659 969 -1625 1003
rect -1659 901 -1625 935
rect -1659 833 -1625 867
rect -1659 765 -1625 799
rect -1659 697 -1625 731
rect -1659 629 -1625 663
rect 1625 1037 1659 1071
rect 1625 969 1659 1003
rect 1625 901 1659 935
rect 1625 833 1659 867
rect 1625 765 1659 799
rect 1625 697 1659 731
rect 1625 629 1659 663
rect -1659 561 -1625 595
rect -1659 493 -1625 527
rect 1625 561 1659 595
rect -1659 425 -1625 459
rect -1659 357 -1625 391
rect -1659 289 -1625 323
rect -1659 221 -1625 255
rect -1659 153 -1625 187
rect -1659 85 -1625 119
rect 1625 493 1659 527
rect 1625 425 1659 459
rect 1625 357 1659 391
rect 1625 289 1659 323
rect 1625 221 1659 255
rect 1625 153 1659 187
rect 1625 85 1659 119
rect -1659 17 -1625 51
rect -1659 -51 -1625 -17
rect 1625 17 1659 51
rect 1625 -51 1659 -17
rect -1659 -119 -1625 -85
rect -1659 -187 -1625 -153
rect -1659 -255 -1625 -221
rect -1659 -323 -1625 -289
rect -1659 -391 -1625 -357
rect -1659 -459 -1625 -425
rect -1659 -527 -1625 -493
rect 1625 -119 1659 -85
rect 1625 -187 1659 -153
rect 1625 -255 1659 -221
rect 1625 -323 1659 -289
rect 1625 -391 1659 -357
rect 1625 -459 1659 -425
rect -1659 -595 -1625 -561
rect 1625 -527 1659 -493
rect 1625 -595 1659 -561
rect -1659 -663 -1625 -629
rect -1659 -731 -1625 -697
rect -1659 -799 -1625 -765
rect -1659 -867 -1625 -833
rect -1659 -935 -1625 -901
rect -1659 -1003 -1625 -969
rect -1659 -1071 -1625 -1037
rect 1625 -663 1659 -629
rect 1625 -731 1659 -697
rect 1625 -799 1659 -765
rect 1625 -867 1659 -833
rect 1625 -935 1659 -901
rect 1625 -1003 1659 -969
rect -1659 -1139 -1625 -1105
rect -1659 -1207 -1625 -1173
rect 1625 -1071 1659 -1037
rect 1625 -1139 1659 -1105
rect 1625 -1207 1659 -1173
rect -1659 -1275 -1625 -1241
rect -1659 -1343 -1625 -1309
rect -1659 -1411 -1625 -1377
rect -1659 -1479 -1625 -1445
rect -1659 -1547 -1625 -1513
rect -1659 -1615 -1625 -1581
rect -1659 -1683 -1625 -1649
rect 1625 -1275 1659 -1241
rect 1625 -1343 1659 -1309
rect 1625 -1411 1659 -1377
rect 1625 -1479 1659 -1445
rect 1625 -1547 1659 -1513
rect 1625 -1615 1659 -1581
rect -1659 -1751 -1625 -1717
rect 1625 -1683 1659 -1649
rect 1625 -1751 1659 -1717
rect -1659 -1819 -1625 -1785
rect -1659 -1887 -1625 -1853
rect -1659 -1955 -1625 -1921
rect -1659 -2023 -1625 -1989
rect -1659 -2091 -1625 -2057
rect -1659 -2159 -1625 -2125
rect 1625 -1819 1659 -1785
rect 1625 -1887 1659 -1853
rect 1625 -1955 1659 -1921
rect 1625 -2023 1659 -1989
rect 1625 -2091 1659 -2057
rect 1625 -2159 1659 -2125
rect -1659 -2227 -1625 -2193
rect -1659 -2295 -1625 -2261
rect -1659 -2363 -1625 -2329
rect 1625 -2227 1659 -2193
rect 1625 -2295 1659 -2261
rect -1659 -2431 -1625 -2397
rect -1659 -2499 -1625 -2465
rect -1659 -2567 -1625 -2533
rect -1659 -2635 -1625 -2601
rect -1659 -2703 -1625 -2669
rect -1659 -2771 -1625 -2737
rect 1625 -2363 1659 -2329
rect 1625 -2431 1659 -2397
rect 1625 -2499 1659 -2465
rect 1625 -2567 1659 -2533
rect 1625 -2635 1659 -2601
rect 1625 -2703 1659 -2669
rect 1625 -2771 1659 -2737
rect -1659 -2884 -1625 -2805
rect 1625 -2884 1659 -2805
rect -1659 -2918 -1547 -2884
rect -1513 -2918 -1479 -2884
rect -1445 -2918 -1411 -2884
rect -1377 -2918 -1343 -2884
rect -1309 -2918 -1275 -2884
rect -1241 -2918 -1207 -2884
rect -1173 -2918 -1139 -2884
rect -1105 -2918 -1071 -2884
rect -1037 -2918 -1003 -2884
rect -969 -2918 -935 -2884
rect -901 -2918 -867 -2884
rect -833 -2918 -799 -2884
rect -765 -2918 -731 -2884
rect -697 -2918 -663 -2884
rect -629 -2918 -595 -2884
rect -561 -2918 -527 -2884
rect -493 -2918 -459 -2884
rect -425 -2918 -391 -2884
rect -357 -2918 -323 -2884
rect -289 -2918 -255 -2884
rect -221 -2918 -187 -2884
rect -153 -2918 -119 -2884
rect -85 -2918 -51 -2884
rect -17 -2918 17 -2884
rect 51 -2918 85 -2884
rect 119 -2918 153 -2884
rect 187 -2918 221 -2884
rect 255 -2918 289 -2884
rect 323 -2918 357 -2884
rect 391 -2918 425 -2884
rect 459 -2918 493 -2884
rect 527 -2918 561 -2884
rect 595 -2918 629 -2884
rect 663 -2918 697 -2884
rect 731 -2918 765 -2884
rect 799 -2918 833 -2884
rect 867 -2918 901 -2884
rect 935 -2918 969 -2884
rect 1003 -2918 1037 -2884
rect 1071 -2918 1105 -2884
rect 1139 -2918 1173 -2884
rect 1207 -2918 1241 -2884
rect 1275 -2918 1309 -2884
rect 1343 -2918 1377 -2884
rect 1411 -2918 1445 -2884
rect 1479 -2918 1513 -2884
rect 1547 -2918 1659 -2884
<< viali >>
rect -1511 2734 -1477 2768
rect -1511 2662 -1477 2696
rect -1511 2590 -1477 2624
rect -1511 2518 -1477 2552
rect -1511 2446 -1477 2480
rect -1511 2374 -1477 2408
rect -1345 2734 -1311 2768
rect -1345 2662 -1311 2696
rect -1345 2590 -1311 2624
rect -1345 2518 -1311 2552
rect -1345 2446 -1311 2480
rect -1345 2374 -1311 2408
rect -1179 2734 -1145 2768
rect -1179 2662 -1145 2696
rect -1179 2590 -1145 2624
rect -1179 2518 -1145 2552
rect -1179 2446 -1145 2480
rect -1179 2374 -1145 2408
rect -1013 2734 -979 2768
rect -1013 2662 -979 2696
rect -1013 2590 -979 2624
rect -1013 2518 -979 2552
rect -1013 2446 -979 2480
rect -1013 2374 -979 2408
rect -847 2734 -813 2768
rect -847 2662 -813 2696
rect -847 2590 -813 2624
rect -847 2518 -813 2552
rect -847 2446 -813 2480
rect -847 2374 -813 2408
rect -681 2734 -647 2768
rect -681 2662 -647 2696
rect -681 2590 -647 2624
rect -681 2518 -647 2552
rect -681 2446 -647 2480
rect -681 2374 -647 2408
rect -515 2734 -481 2768
rect -515 2662 -481 2696
rect -515 2590 -481 2624
rect -515 2518 -481 2552
rect -515 2446 -481 2480
rect -515 2374 -481 2408
rect -349 2734 -315 2768
rect -349 2662 -315 2696
rect -349 2590 -315 2624
rect -349 2518 -315 2552
rect -349 2446 -315 2480
rect -349 2374 -315 2408
rect -183 2734 -149 2768
rect -183 2662 -149 2696
rect -183 2590 -149 2624
rect -183 2518 -149 2552
rect -183 2446 -149 2480
rect -183 2374 -149 2408
rect -17 2734 17 2768
rect -17 2662 17 2696
rect -17 2590 17 2624
rect -17 2518 17 2552
rect -17 2446 17 2480
rect -17 2374 17 2408
rect 149 2734 183 2768
rect 149 2662 183 2696
rect 149 2590 183 2624
rect 149 2518 183 2552
rect 149 2446 183 2480
rect 149 2374 183 2408
rect 315 2734 349 2768
rect 315 2662 349 2696
rect 315 2590 349 2624
rect 315 2518 349 2552
rect 315 2446 349 2480
rect 315 2374 349 2408
rect 481 2734 515 2768
rect 481 2662 515 2696
rect 481 2590 515 2624
rect 481 2518 515 2552
rect 481 2446 515 2480
rect 481 2374 515 2408
rect 647 2734 681 2768
rect 647 2662 681 2696
rect 647 2590 681 2624
rect 647 2518 681 2552
rect 647 2446 681 2480
rect 647 2374 681 2408
rect 813 2734 847 2768
rect 813 2662 847 2696
rect 813 2590 847 2624
rect 813 2518 847 2552
rect 813 2446 847 2480
rect 813 2374 847 2408
rect 979 2734 1013 2768
rect 979 2662 1013 2696
rect 979 2590 1013 2624
rect 979 2518 1013 2552
rect 979 2446 1013 2480
rect 979 2374 1013 2408
rect 1145 2734 1179 2768
rect 1145 2662 1179 2696
rect 1145 2590 1179 2624
rect 1145 2518 1179 2552
rect 1145 2446 1179 2480
rect 1145 2374 1179 2408
rect 1311 2734 1345 2768
rect 1311 2662 1345 2696
rect 1311 2590 1345 2624
rect 1311 2518 1345 2552
rect 1311 2446 1345 2480
rect 1311 2374 1345 2408
rect 1477 2734 1511 2768
rect 1477 2662 1511 2696
rect 1477 2590 1511 2624
rect 1477 2518 1511 2552
rect 1477 2446 1511 2480
rect 1477 2374 1511 2408
rect -1511 2135 -1477 2169
rect -1511 2063 -1477 2097
rect -1511 1991 -1477 2025
rect -1511 1919 -1477 1953
rect -1511 1847 -1477 1881
rect -1511 1775 -1477 1809
rect -1345 2135 -1311 2169
rect -1345 2063 -1311 2097
rect -1345 1991 -1311 2025
rect -1345 1919 -1311 1953
rect -1345 1847 -1311 1881
rect -1345 1775 -1311 1809
rect -1179 2135 -1145 2169
rect -1179 2063 -1145 2097
rect -1179 1991 -1145 2025
rect -1179 1919 -1145 1953
rect -1179 1847 -1145 1881
rect -1179 1775 -1145 1809
rect -1013 2135 -979 2169
rect -1013 2063 -979 2097
rect -1013 1991 -979 2025
rect -1013 1919 -979 1953
rect -1013 1847 -979 1881
rect -1013 1775 -979 1809
rect -847 2135 -813 2169
rect -847 2063 -813 2097
rect -847 1991 -813 2025
rect -847 1919 -813 1953
rect -847 1847 -813 1881
rect -847 1775 -813 1809
rect -681 2135 -647 2169
rect -681 2063 -647 2097
rect -681 1991 -647 2025
rect -681 1919 -647 1953
rect -681 1847 -647 1881
rect -681 1775 -647 1809
rect -515 2135 -481 2169
rect -515 2063 -481 2097
rect -515 1991 -481 2025
rect -515 1919 -481 1953
rect -515 1847 -481 1881
rect -515 1775 -481 1809
rect -349 2135 -315 2169
rect -349 2063 -315 2097
rect -349 1991 -315 2025
rect -349 1919 -315 1953
rect -349 1847 -315 1881
rect -349 1775 -315 1809
rect -183 2135 -149 2169
rect -183 2063 -149 2097
rect -183 1991 -149 2025
rect -183 1919 -149 1953
rect -183 1847 -149 1881
rect -183 1775 -149 1809
rect -17 2135 17 2169
rect -17 2063 17 2097
rect -17 1991 17 2025
rect -17 1919 17 1953
rect -17 1847 17 1881
rect -17 1775 17 1809
rect 149 2135 183 2169
rect 149 2063 183 2097
rect 149 1991 183 2025
rect 149 1919 183 1953
rect 149 1847 183 1881
rect 149 1775 183 1809
rect 315 2135 349 2169
rect 315 2063 349 2097
rect 315 1991 349 2025
rect 315 1919 349 1953
rect 315 1847 349 1881
rect 315 1775 349 1809
rect 481 2135 515 2169
rect 481 2063 515 2097
rect 481 1991 515 2025
rect 481 1919 515 1953
rect 481 1847 515 1881
rect 481 1775 515 1809
rect 647 2135 681 2169
rect 647 2063 681 2097
rect 647 1991 681 2025
rect 647 1919 681 1953
rect 647 1847 681 1881
rect 647 1775 681 1809
rect 813 2135 847 2169
rect 813 2063 847 2097
rect 813 1991 847 2025
rect 813 1919 847 1953
rect 813 1847 847 1881
rect 813 1775 847 1809
rect 979 2135 1013 2169
rect 979 2063 1013 2097
rect 979 1991 1013 2025
rect 979 1919 1013 1953
rect 979 1847 1013 1881
rect 979 1775 1013 1809
rect 1145 2135 1179 2169
rect 1145 2063 1179 2097
rect 1145 1991 1179 2025
rect 1145 1919 1179 1953
rect 1145 1847 1179 1881
rect 1145 1775 1179 1809
rect 1311 2135 1345 2169
rect 1311 2063 1345 2097
rect 1311 1991 1345 2025
rect 1311 1919 1345 1953
rect 1311 1847 1345 1881
rect 1311 1775 1345 1809
rect 1477 2135 1511 2169
rect 1477 2063 1511 2097
rect 1477 1991 1511 2025
rect 1477 1919 1511 1953
rect 1477 1847 1511 1881
rect 1477 1775 1511 1809
rect -1511 1598 -1477 1632
rect -1511 1526 -1477 1560
rect -1511 1454 -1477 1488
rect -1511 1382 -1477 1416
rect -1511 1310 -1477 1344
rect -1511 1238 -1477 1272
rect -1345 1598 -1311 1632
rect -1345 1526 -1311 1560
rect -1345 1454 -1311 1488
rect -1345 1382 -1311 1416
rect -1345 1310 -1311 1344
rect -1345 1238 -1311 1272
rect -1179 1598 -1145 1632
rect -1179 1526 -1145 1560
rect -1179 1454 -1145 1488
rect -1179 1382 -1145 1416
rect -1179 1310 -1145 1344
rect -1179 1238 -1145 1272
rect -1013 1598 -979 1632
rect -1013 1526 -979 1560
rect -1013 1454 -979 1488
rect -1013 1382 -979 1416
rect -1013 1310 -979 1344
rect -1013 1238 -979 1272
rect -847 1598 -813 1632
rect -847 1526 -813 1560
rect -847 1454 -813 1488
rect -847 1382 -813 1416
rect -847 1310 -813 1344
rect -847 1238 -813 1272
rect -681 1598 -647 1632
rect -681 1526 -647 1560
rect -681 1454 -647 1488
rect -681 1382 -647 1416
rect -681 1310 -647 1344
rect -681 1238 -647 1272
rect -515 1598 -481 1632
rect -515 1526 -481 1560
rect -515 1454 -481 1488
rect -515 1382 -481 1416
rect -515 1310 -481 1344
rect -515 1238 -481 1272
rect -349 1598 -315 1632
rect -349 1526 -315 1560
rect -349 1454 -315 1488
rect -349 1382 -315 1416
rect -349 1310 -315 1344
rect -349 1238 -315 1272
rect -183 1598 -149 1632
rect -183 1526 -149 1560
rect -183 1454 -149 1488
rect -183 1382 -149 1416
rect -183 1310 -149 1344
rect -183 1238 -149 1272
rect -17 1598 17 1632
rect -17 1526 17 1560
rect -17 1454 17 1488
rect -17 1382 17 1416
rect -17 1310 17 1344
rect -17 1238 17 1272
rect 149 1598 183 1632
rect 149 1526 183 1560
rect 149 1454 183 1488
rect 149 1382 183 1416
rect 149 1310 183 1344
rect 149 1238 183 1272
rect 315 1598 349 1632
rect 315 1526 349 1560
rect 315 1454 349 1488
rect 315 1382 349 1416
rect 315 1310 349 1344
rect 315 1238 349 1272
rect 481 1598 515 1632
rect 481 1526 515 1560
rect 481 1454 515 1488
rect 481 1382 515 1416
rect 481 1310 515 1344
rect 481 1238 515 1272
rect 647 1598 681 1632
rect 647 1526 681 1560
rect 647 1454 681 1488
rect 647 1382 681 1416
rect 647 1310 681 1344
rect 647 1238 681 1272
rect 813 1598 847 1632
rect 813 1526 847 1560
rect 813 1454 847 1488
rect 813 1382 847 1416
rect 813 1310 847 1344
rect 813 1238 847 1272
rect 979 1598 1013 1632
rect 979 1526 1013 1560
rect 979 1454 1013 1488
rect 979 1382 1013 1416
rect 979 1310 1013 1344
rect 979 1238 1013 1272
rect 1145 1598 1179 1632
rect 1145 1526 1179 1560
rect 1145 1454 1179 1488
rect 1145 1382 1179 1416
rect 1145 1310 1179 1344
rect 1145 1238 1179 1272
rect 1311 1598 1345 1632
rect 1311 1526 1345 1560
rect 1311 1454 1345 1488
rect 1311 1382 1345 1416
rect 1311 1310 1345 1344
rect 1311 1238 1345 1272
rect 1477 1598 1511 1632
rect 1477 1526 1511 1560
rect 1477 1454 1511 1488
rect 1477 1382 1511 1416
rect 1477 1310 1511 1344
rect 1477 1238 1511 1272
rect -1511 999 -1477 1033
rect -1511 927 -1477 961
rect -1511 855 -1477 889
rect -1511 783 -1477 817
rect -1511 711 -1477 745
rect -1511 639 -1477 673
rect -1345 999 -1311 1033
rect -1345 927 -1311 961
rect -1345 855 -1311 889
rect -1345 783 -1311 817
rect -1345 711 -1311 745
rect -1345 639 -1311 673
rect -1179 999 -1145 1033
rect -1179 927 -1145 961
rect -1179 855 -1145 889
rect -1179 783 -1145 817
rect -1179 711 -1145 745
rect -1179 639 -1145 673
rect -1013 999 -979 1033
rect -1013 927 -979 961
rect -1013 855 -979 889
rect -1013 783 -979 817
rect -1013 711 -979 745
rect -1013 639 -979 673
rect -847 999 -813 1033
rect -847 927 -813 961
rect -847 855 -813 889
rect -847 783 -813 817
rect -847 711 -813 745
rect -847 639 -813 673
rect -681 999 -647 1033
rect -681 927 -647 961
rect -681 855 -647 889
rect -681 783 -647 817
rect -681 711 -647 745
rect -681 639 -647 673
rect -515 999 -481 1033
rect -515 927 -481 961
rect -515 855 -481 889
rect -515 783 -481 817
rect -515 711 -481 745
rect -515 639 -481 673
rect -349 999 -315 1033
rect -349 927 -315 961
rect -349 855 -315 889
rect -349 783 -315 817
rect -349 711 -315 745
rect -349 639 -315 673
rect -183 999 -149 1033
rect -183 927 -149 961
rect -183 855 -149 889
rect -183 783 -149 817
rect -183 711 -149 745
rect -183 639 -149 673
rect -17 999 17 1033
rect -17 927 17 961
rect -17 855 17 889
rect -17 783 17 817
rect -17 711 17 745
rect -17 639 17 673
rect 149 999 183 1033
rect 149 927 183 961
rect 149 855 183 889
rect 149 783 183 817
rect 149 711 183 745
rect 149 639 183 673
rect 315 999 349 1033
rect 315 927 349 961
rect 315 855 349 889
rect 315 783 349 817
rect 315 711 349 745
rect 315 639 349 673
rect 481 999 515 1033
rect 481 927 515 961
rect 481 855 515 889
rect 481 783 515 817
rect 481 711 515 745
rect 481 639 515 673
rect 647 999 681 1033
rect 647 927 681 961
rect 647 855 681 889
rect 647 783 681 817
rect 647 711 681 745
rect 647 639 681 673
rect 813 999 847 1033
rect 813 927 847 961
rect 813 855 847 889
rect 813 783 847 817
rect 813 711 847 745
rect 813 639 847 673
rect 979 999 1013 1033
rect 979 927 1013 961
rect 979 855 1013 889
rect 979 783 1013 817
rect 979 711 1013 745
rect 979 639 1013 673
rect 1145 999 1179 1033
rect 1145 927 1179 961
rect 1145 855 1179 889
rect 1145 783 1179 817
rect 1145 711 1179 745
rect 1145 639 1179 673
rect 1311 999 1345 1033
rect 1311 927 1345 961
rect 1311 855 1345 889
rect 1311 783 1345 817
rect 1311 711 1345 745
rect 1311 639 1345 673
rect 1477 999 1511 1033
rect 1477 927 1511 961
rect 1477 855 1511 889
rect 1477 783 1511 817
rect 1477 711 1511 745
rect 1477 639 1511 673
rect -1511 462 -1477 496
rect -1511 390 -1477 424
rect -1511 318 -1477 352
rect -1511 246 -1477 280
rect -1511 174 -1477 208
rect -1511 102 -1477 136
rect -1345 462 -1311 496
rect -1345 390 -1311 424
rect -1345 318 -1311 352
rect -1345 246 -1311 280
rect -1345 174 -1311 208
rect -1345 102 -1311 136
rect -1179 462 -1145 496
rect -1179 390 -1145 424
rect -1179 318 -1145 352
rect -1179 246 -1145 280
rect -1179 174 -1145 208
rect -1179 102 -1145 136
rect -1013 462 -979 496
rect -1013 390 -979 424
rect -1013 318 -979 352
rect -1013 246 -979 280
rect -1013 174 -979 208
rect -1013 102 -979 136
rect -847 462 -813 496
rect -847 390 -813 424
rect -847 318 -813 352
rect -847 246 -813 280
rect -847 174 -813 208
rect -847 102 -813 136
rect -681 462 -647 496
rect -681 390 -647 424
rect -681 318 -647 352
rect -681 246 -647 280
rect -681 174 -647 208
rect -681 102 -647 136
rect -515 462 -481 496
rect -515 390 -481 424
rect -515 318 -481 352
rect -515 246 -481 280
rect -515 174 -481 208
rect -515 102 -481 136
rect -349 462 -315 496
rect -349 390 -315 424
rect -349 318 -315 352
rect -349 246 -315 280
rect -349 174 -315 208
rect -349 102 -315 136
rect -183 462 -149 496
rect -183 390 -149 424
rect -183 318 -149 352
rect -183 246 -149 280
rect -183 174 -149 208
rect -183 102 -149 136
rect -17 462 17 496
rect -17 390 17 424
rect -17 318 17 352
rect -17 246 17 280
rect -17 174 17 208
rect -17 102 17 136
rect 149 462 183 496
rect 149 390 183 424
rect 149 318 183 352
rect 149 246 183 280
rect 149 174 183 208
rect 149 102 183 136
rect 315 462 349 496
rect 315 390 349 424
rect 315 318 349 352
rect 315 246 349 280
rect 315 174 349 208
rect 315 102 349 136
rect 481 462 515 496
rect 481 390 515 424
rect 481 318 515 352
rect 481 246 515 280
rect 481 174 515 208
rect 481 102 515 136
rect 647 462 681 496
rect 647 390 681 424
rect 647 318 681 352
rect 647 246 681 280
rect 647 174 681 208
rect 647 102 681 136
rect 813 462 847 496
rect 813 390 847 424
rect 813 318 847 352
rect 813 246 847 280
rect 813 174 847 208
rect 813 102 847 136
rect 979 462 1013 496
rect 979 390 1013 424
rect 979 318 1013 352
rect 979 246 1013 280
rect 979 174 1013 208
rect 979 102 1013 136
rect 1145 462 1179 496
rect 1145 390 1179 424
rect 1145 318 1179 352
rect 1145 246 1179 280
rect 1145 174 1179 208
rect 1145 102 1179 136
rect 1311 462 1345 496
rect 1311 390 1345 424
rect 1311 318 1345 352
rect 1311 246 1345 280
rect 1311 174 1345 208
rect 1311 102 1345 136
rect 1477 462 1511 496
rect 1477 390 1511 424
rect 1477 318 1511 352
rect 1477 246 1511 280
rect 1477 174 1511 208
rect 1477 102 1511 136
rect -1511 -137 -1477 -103
rect -1511 -209 -1477 -175
rect -1511 -281 -1477 -247
rect -1511 -353 -1477 -319
rect -1511 -425 -1477 -391
rect -1511 -497 -1477 -463
rect -1345 -137 -1311 -103
rect -1345 -209 -1311 -175
rect -1345 -281 -1311 -247
rect -1345 -353 -1311 -319
rect -1345 -425 -1311 -391
rect -1345 -497 -1311 -463
rect -1179 -137 -1145 -103
rect -1179 -209 -1145 -175
rect -1179 -281 -1145 -247
rect -1179 -353 -1145 -319
rect -1179 -425 -1145 -391
rect -1179 -497 -1145 -463
rect -1013 -137 -979 -103
rect -1013 -209 -979 -175
rect -1013 -281 -979 -247
rect -1013 -353 -979 -319
rect -1013 -425 -979 -391
rect -1013 -497 -979 -463
rect -847 -137 -813 -103
rect -847 -209 -813 -175
rect -847 -281 -813 -247
rect -847 -353 -813 -319
rect -847 -425 -813 -391
rect -847 -497 -813 -463
rect -681 -137 -647 -103
rect -681 -209 -647 -175
rect -681 -281 -647 -247
rect -681 -353 -647 -319
rect -681 -425 -647 -391
rect -681 -497 -647 -463
rect -515 -137 -481 -103
rect -515 -209 -481 -175
rect -515 -281 -481 -247
rect -515 -353 -481 -319
rect -515 -425 -481 -391
rect -515 -497 -481 -463
rect -349 -137 -315 -103
rect -349 -209 -315 -175
rect -349 -281 -315 -247
rect -349 -353 -315 -319
rect -349 -425 -315 -391
rect -349 -497 -315 -463
rect -183 -137 -149 -103
rect -183 -209 -149 -175
rect -183 -281 -149 -247
rect -183 -353 -149 -319
rect -183 -425 -149 -391
rect -183 -497 -149 -463
rect -17 -137 17 -103
rect -17 -209 17 -175
rect -17 -281 17 -247
rect -17 -353 17 -319
rect -17 -425 17 -391
rect -17 -497 17 -463
rect 149 -137 183 -103
rect 149 -209 183 -175
rect 149 -281 183 -247
rect 149 -353 183 -319
rect 149 -425 183 -391
rect 149 -497 183 -463
rect 315 -137 349 -103
rect 315 -209 349 -175
rect 315 -281 349 -247
rect 315 -353 349 -319
rect 315 -425 349 -391
rect 315 -497 349 -463
rect 481 -137 515 -103
rect 481 -209 515 -175
rect 481 -281 515 -247
rect 481 -353 515 -319
rect 481 -425 515 -391
rect 481 -497 515 -463
rect 647 -137 681 -103
rect 647 -209 681 -175
rect 647 -281 681 -247
rect 647 -353 681 -319
rect 647 -425 681 -391
rect 647 -497 681 -463
rect 813 -137 847 -103
rect 813 -209 847 -175
rect 813 -281 847 -247
rect 813 -353 847 -319
rect 813 -425 847 -391
rect 813 -497 847 -463
rect 979 -137 1013 -103
rect 979 -209 1013 -175
rect 979 -281 1013 -247
rect 979 -353 1013 -319
rect 979 -425 1013 -391
rect 979 -497 1013 -463
rect 1145 -137 1179 -103
rect 1145 -209 1179 -175
rect 1145 -281 1179 -247
rect 1145 -353 1179 -319
rect 1145 -425 1179 -391
rect 1145 -497 1179 -463
rect 1311 -137 1345 -103
rect 1311 -209 1345 -175
rect 1311 -281 1345 -247
rect 1311 -353 1345 -319
rect 1311 -425 1345 -391
rect 1311 -497 1345 -463
rect 1477 -137 1511 -103
rect 1477 -209 1511 -175
rect 1477 -281 1511 -247
rect 1477 -353 1511 -319
rect 1477 -425 1511 -391
rect 1477 -497 1511 -463
rect -1511 -674 -1477 -640
rect -1511 -746 -1477 -712
rect -1511 -818 -1477 -784
rect -1511 -890 -1477 -856
rect -1511 -962 -1477 -928
rect -1511 -1034 -1477 -1000
rect -1345 -674 -1311 -640
rect -1345 -746 -1311 -712
rect -1345 -818 -1311 -784
rect -1345 -890 -1311 -856
rect -1345 -962 -1311 -928
rect -1345 -1034 -1311 -1000
rect -1179 -674 -1145 -640
rect -1179 -746 -1145 -712
rect -1179 -818 -1145 -784
rect -1179 -890 -1145 -856
rect -1179 -962 -1145 -928
rect -1179 -1034 -1145 -1000
rect -1013 -674 -979 -640
rect -1013 -746 -979 -712
rect -1013 -818 -979 -784
rect -1013 -890 -979 -856
rect -1013 -962 -979 -928
rect -1013 -1034 -979 -1000
rect -847 -674 -813 -640
rect -847 -746 -813 -712
rect -847 -818 -813 -784
rect -847 -890 -813 -856
rect -847 -962 -813 -928
rect -847 -1034 -813 -1000
rect -681 -674 -647 -640
rect -681 -746 -647 -712
rect -681 -818 -647 -784
rect -681 -890 -647 -856
rect -681 -962 -647 -928
rect -681 -1034 -647 -1000
rect -515 -674 -481 -640
rect -515 -746 -481 -712
rect -515 -818 -481 -784
rect -515 -890 -481 -856
rect -515 -962 -481 -928
rect -515 -1034 -481 -1000
rect -349 -674 -315 -640
rect -349 -746 -315 -712
rect -349 -818 -315 -784
rect -349 -890 -315 -856
rect -349 -962 -315 -928
rect -349 -1034 -315 -1000
rect -183 -674 -149 -640
rect -183 -746 -149 -712
rect -183 -818 -149 -784
rect -183 -890 -149 -856
rect -183 -962 -149 -928
rect -183 -1034 -149 -1000
rect -17 -674 17 -640
rect -17 -746 17 -712
rect -17 -818 17 -784
rect -17 -890 17 -856
rect -17 -962 17 -928
rect -17 -1034 17 -1000
rect 149 -674 183 -640
rect 149 -746 183 -712
rect 149 -818 183 -784
rect 149 -890 183 -856
rect 149 -962 183 -928
rect 149 -1034 183 -1000
rect 315 -674 349 -640
rect 315 -746 349 -712
rect 315 -818 349 -784
rect 315 -890 349 -856
rect 315 -962 349 -928
rect 315 -1034 349 -1000
rect 481 -674 515 -640
rect 481 -746 515 -712
rect 481 -818 515 -784
rect 481 -890 515 -856
rect 481 -962 515 -928
rect 481 -1034 515 -1000
rect 647 -674 681 -640
rect 647 -746 681 -712
rect 647 -818 681 -784
rect 647 -890 681 -856
rect 647 -962 681 -928
rect 647 -1034 681 -1000
rect 813 -674 847 -640
rect 813 -746 847 -712
rect 813 -818 847 -784
rect 813 -890 847 -856
rect 813 -962 847 -928
rect 813 -1034 847 -1000
rect 979 -674 1013 -640
rect 979 -746 1013 -712
rect 979 -818 1013 -784
rect 979 -890 1013 -856
rect 979 -962 1013 -928
rect 979 -1034 1013 -1000
rect 1145 -674 1179 -640
rect 1145 -746 1179 -712
rect 1145 -818 1179 -784
rect 1145 -890 1179 -856
rect 1145 -962 1179 -928
rect 1145 -1034 1179 -1000
rect 1311 -674 1345 -640
rect 1311 -746 1345 -712
rect 1311 -818 1345 -784
rect 1311 -890 1345 -856
rect 1311 -962 1345 -928
rect 1311 -1034 1345 -1000
rect 1477 -674 1511 -640
rect 1477 -746 1511 -712
rect 1477 -818 1511 -784
rect 1477 -890 1511 -856
rect 1477 -962 1511 -928
rect 1477 -1034 1511 -1000
rect -1511 -1273 -1477 -1239
rect -1511 -1345 -1477 -1311
rect -1511 -1417 -1477 -1383
rect -1511 -1489 -1477 -1455
rect -1511 -1561 -1477 -1527
rect -1511 -1633 -1477 -1599
rect -1345 -1273 -1311 -1239
rect -1345 -1345 -1311 -1311
rect -1345 -1417 -1311 -1383
rect -1345 -1489 -1311 -1455
rect -1345 -1561 -1311 -1527
rect -1345 -1633 -1311 -1599
rect -1179 -1273 -1145 -1239
rect -1179 -1345 -1145 -1311
rect -1179 -1417 -1145 -1383
rect -1179 -1489 -1145 -1455
rect -1179 -1561 -1145 -1527
rect -1179 -1633 -1145 -1599
rect -1013 -1273 -979 -1239
rect -1013 -1345 -979 -1311
rect -1013 -1417 -979 -1383
rect -1013 -1489 -979 -1455
rect -1013 -1561 -979 -1527
rect -1013 -1633 -979 -1599
rect -847 -1273 -813 -1239
rect -847 -1345 -813 -1311
rect -847 -1417 -813 -1383
rect -847 -1489 -813 -1455
rect -847 -1561 -813 -1527
rect -847 -1633 -813 -1599
rect -681 -1273 -647 -1239
rect -681 -1345 -647 -1311
rect -681 -1417 -647 -1383
rect -681 -1489 -647 -1455
rect -681 -1561 -647 -1527
rect -681 -1633 -647 -1599
rect -515 -1273 -481 -1239
rect -515 -1345 -481 -1311
rect -515 -1417 -481 -1383
rect -515 -1489 -481 -1455
rect -515 -1561 -481 -1527
rect -515 -1633 -481 -1599
rect -349 -1273 -315 -1239
rect -349 -1345 -315 -1311
rect -349 -1417 -315 -1383
rect -349 -1489 -315 -1455
rect -349 -1561 -315 -1527
rect -349 -1633 -315 -1599
rect -183 -1273 -149 -1239
rect -183 -1345 -149 -1311
rect -183 -1417 -149 -1383
rect -183 -1489 -149 -1455
rect -183 -1561 -149 -1527
rect -183 -1633 -149 -1599
rect -17 -1273 17 -1239
rect -17 -1345 17 -1311
rect -17 -1417 17 -1383
rect -17 -1489 17 -1455
rect -17 -1561 17 -1527
rect -17 -1633 17 -1599
rect 149 -1273 183 -1239
rect 149 -1345 183 -1311
rect 149 -1417 183 -1383
rect 149 -1489 183 -1455
rect 149 -1561 183 -1527
rect 149 -1633 183 -1599
rect 315 -1273 349 -1239
rect 315 -1345 349 -1311
rect 315 -1417 349 -1383
rect 315 -1489 349 -1455
rect 315 -1561 349 -1527
rect 315 -1633 349 -1599
rect 481 -1273 515 -1239
rect 481 -1345 515 -1311
rect 481 -1417 515 -1383
rect 481 -1489 515 -1455
rect 481 -1561 515 -1527
rect 481 -1633 515 -1599
rect 647 -1273 681 -1239
rect 647 -1345 681 -1311
rect 647 -1417 681 -1383
rect 647 -1489 681 -1455
rect 647 -1561 681 -1527
rect 647 -1633 681 -1599
rect 813 -1273 847 -1239
rect 813 -1345 847 -1311
rect 813 -1417 847 -1383
rect 813 -1489 847 -1455
rect 813 -1561 847 -1527
rect 813 -1633 847 -1599
rect 979 -1273 1013 -1239
rect 979 -1345 1013 -1311
rect 979 -1417 1013 -1383
rect 979 -1489 1013 -1455
rect 979 -1561 1013 -1527
rect 979 -1633 1013 -1599
rect 1145 -1273 1179 -1239
rect 1145 -1345 1179 -1311
rect 1145 -1417 1179 -1383
rect 1145 -1489 1179 -1455
rect 1145 -1561 1179 -1527
rect 1145 -1633 1179 -1599
rect 1311 -1273 1345 -1239
rect 1311 -1345 1345 -1311
rect 1311 -1417 1345 -1383
rect 1311 -1489 1345 -1455
rect 1311 -1561 1345 -1527
rect 1311 -1633 1345 -1599
rect 1477 -1273 1511 -1239
rect 1477 -1345 1511 -1311
rect 1477 -1417 1511 -1383
rect 1477 -1489 1511 -1455
rect 1477 -1561 1511 -1527
rect 1477 -1633 1511 -1599
rect -1511 -1810 -1477 -1776
rect -1511 -1882 -1477 -1848
rect -1511 -1954 -1477 -1920
rect -1511 -2026 -1477 -1992
rect -1511 -2098 -1477 -2064
rect -1511 -2170 -1477 -2136
rect -1345 -1810 -1311 -1776
rect -1345 -1882 -1311 -1848
rect -1345 -1954 -1311 -1920
rect -1345 -2026 -1311 -1992
rect -1345 -2098 -1311 -2064
rect -1345 -2170 -1311 -2136
rect -1179 -1810 -1145 -1776
rect -1179 -1882 -1145 -1848
rect -1179 -1954 -1145 -1920
rect -1179 -2026 -1145 -1992
rect -1179 -2098 -1145 -2064
rect -1179 -2170 -1145 -2136
rect -1013 -1810 -979 -1776
rect -1013 -1882 -979 -1848
rect -1013 -1954 -979 -1920
rect -1013 -2026 -979 -1992
rect -1013 -2098 -979 -2064
rect -1013 -2170 -979 -2136
rect -847 -1810 -813 -1776
rect -847 -1882 -813 -1848
rect -847 -1954 -813 -1920
rect -847 -2026 -813 -1992
rect -847 -2098 -813 -2064
rect -847 -2170 -813 -2136
rect -681 -1810 -647 -1776
rect -681 -1882 -647 -1848
rect -681 -1954 -647 -1920
rect -681 -2026 -647 -1992
rect -681 -2098 -647 -2064
rect -681 -2170 -647 -2136
rect -515 -1810 -481 -1776
rect -515 -1882 -481 -1848
rect -515 -1954 -481 -1920
rect -515 -2026 -481 -1992
rect -515 -2098 -481 -2064
rect -515 -2170 -481 -2136
rect -349 -1810 -315 -1776
rect -349 -1882 -315 -1848
rect -349 -1954 -315 -1920
rect -349 -2026 -315 -1992
rect -349 -2098 -315 -2064
rect -349 -2170 -315 -2136
rect -183 -1810 -149 -1776
rect -183 -1882 -149 -1848
rect -183 -1954 -149 -1920
rect -183 -2026 -149 -1992
rect -183 -2098 -149 -2064
rect -183 -2170 -149 -2136
rect -17 -1810 17 -1776
rect -17 -1882 17 -1848
rect -17 -1954 17 -1920
rect -17 -2026 17 -1992
rect -17 -2098 17 -2064
rect -17 -2170 17 -2136
rect 149 -1810 183 -1776
rect 149 -1882 183 -1848
rect 149 -1954 183 -1920
rect 149 -2026 183 -1992
rect 149 -2098 183 -2064
rect 149 -2170 183 -2136
rect 315 -1810 349 -1776
rect 315 -1882 349 -1848
rect 315 -1954 349 -1920
rect 315 -2026 349 -1992
rect 315 -2098 349 -2064
rect 315 -2170 349 -2136
rect 481 -1810 515 -1776
rect 481 -1882 515 -1848
rect 481 -1954 515 -1920
rect 481 -2026 515 -1992
rect 481 -2098 515 -2064
rect 481 -2170 515 -2136
rect 647 -1810 681 -1776
rect 647 -1882 681 -1848
rect 647 -1954 681 -1920
rect 647 -2026 681 -1992
rect 647 -2098 681 -2064
rect 647 -2170 681 -2136
rect 813 -1810 847 -1776
rect 813 -1882 847 -1848
rect 813 -1954 847 -1920
rect 813 -2026 847 -1992
rect 813 -2098 847 -2064
rect 813 -2170 847 -2136
rect 979 -1810 1013 -1776
rect 979 -1882 1013 -1848
rect 979 -1954 1013 -1920
rect 979 -2026 1013 -1992
rect 979 -2098 1013 -2064
rect 979 -2170 1013 -2136
rect 1145 -1810 1179 -1776
rect 1145 -1882 1179 -1848
rect 1145 -1954 1179 -1920
rect 1145 -2026 1179 -1992
rect 1145 -2098 1179 -2064
rect 1145 -2170 1179 -2136
rect 1311 -1810 1345 -1776
rect 1311 -1882 1345 -1848
rect 1311 -1954 1345 -1920
rect 1311 -2026 1345 -1992
rect 1311 -2098 1345 -2064
rect 1311 -2170 1345 -2136
rect 1477 -1810 1511 -1776
rect 1477 -1882 1511 -1848
rect 1477 -1954 1511 -1920
rect 1477 -2026 1511 -1992
rect 1477 -2098 1511 -2064
rect 1477 -2170 1511 -2136
rect -1511 -2409 -1477 -2375
rect -1511 -2481 -1477 -2447
rect -1511 -2553 -1477 -2519
rect -1511 -2625 -1477 -2591
rect -1511 -2697 -1477 -2663
rect -1511 -2769 -1477 -2735
rect -1345 -2409 -1311 -2375
rect -1345 -2481 -1311 -2447
rect -1345 -2553 -1311 -2519
rect -1345 -2625 -1311 -2591
rect -1345 -2697 -1311 -2663
rect -1345 -2769 -1311 -2735
rect -1179 -2409 -1145 -2375
rect -1179 -2481 -1145 -2447
rect -1179 -2553 -1145 -2519
rect -1179 -2625 -1145 -2591
rect -1179 -2697 -1145 -2663
rect -1179 -2769 -1145 -2735
rect -1013 -2409 -979 -2375
rect -1013 -2481 -979 -2447
rect -1013 -2553 -979 -2519
rect -1013 -2625 -979 -2591
rect -1013 -2697 -979 -2663
rect -1013 -2769 -979 -2735
rect -847 -2409 -813 -2375
rect -847 -2481 -813 -2447
rect -847 -2553 -813 -2519
rect -847 -2625 -813 -2591
rect -847 -2697 -813 -2663
rect -847 -2769 -813 -2735
rect -681 -2409 -647 -2375
rect -681 -2481 -647 -2447
rect -681 -2553 -647 -2519
rect -681 -2625 -647 -2591
rect -681 -2697 -647 -2663
rect -681 -2769 -647 -2735
rect -515 -2409 -481 -2375
rect -515 -2481 -481 -2447
rect -515 -2553 -481 -2519
rect -515 -2625 -481 -2591
rect -515 -2697 -481 -2663
rect -515 -2769 -481 -2735
rect -349 -2409 -315 -2375
rect -349 -2481 -315 -2447
rect -349 -2553 -315 -2519
rect -349 -2625 -315 -2591
rect -349 -2697 -315 -2663
rect -349 -2769 -315 -2735
rect -183 -2409 -149 -2375
rect -183 -2481 -149 -2447
rect -183 -2553 -149 -2519
rect -183 -2625 -149 -2591
rect -183 -2697 -149 -2663
rect -183 -2769 -149 -2735
rect -17 -2409 17 -2375
rect -17 -2481 17 -2447
rect -17 -2553 17 -2519
rect -17 -2625 17 -2591
rect -17 -2697 17 -2663
rect -17 -2769 17 -2735
rect 149 -2409 183 -2375
rect 149 -2481 183 -2447
rect 149 -2553 183 -2519
rect 149 -2625 183 -2591
rect 149 -2697 183 -2663
rect 149 -2769 183 -2735
rect 315 -2409 349 -2375
rect 315 -2481 349 -2447
rect 315 -2553 349 -2519
rect 315 -2625 349 -2591
rect 315 -2697 349 -2663
rect 315 -2769 349 -2735
rect 481 -2409 515 -2375
rect 481 -2481 515 -2447
rect 481 -2553 515 -2519
rect 481 -2625 515 -2591
rect 481 -2697 515 -2663
rect 481 -2769 515 -2735
rect 647 -2409 681 -2375
rect 647 -2481 681 -2447
rect 647 -2553 681 -2519
rect 647 -2625 681 -2591
rect 647 -2697 681 -2663
rect 647 -2769 681 -2735
rect 813 -2409 847 -2375
rect 813 -2481 847 -2447
rect 813 -2553 847 -2519
rect 813 -2625 847 -2591
rect 813 -2697 847 -2663
rect 813 -2769 847 -2735
rect 979 -2409 1013 -2375
rect 979 -2481 1013 -2447
rect 979 -2553 1013 -2519
rect 979 -2625 1013 -2591
rect 979 -2697 1013 -2663
rect 979 -2769 1013 -2735
rect 1145 -2409 1179 -2375
rect 1145 -2481 1179 -2447
rect 1145 -2553 1179 -2519
rect 1145 -2625 1179 -2591
rect 1145 -2697 1179 -2663
rect 1145 -2769 1179 -2735
rect 1311 -2409 1345 -2375
rect 1311 -2481 1345 -2447
rect 1311 -2553 1345 -2519
rect 1311 -2625 1345 -2591
rect 1311 -2697 1345 -2663
rect 1311 -2769 1345 -2735
rect 1477 -2409 1511 -2375
rect 1477 -2481 1511 -2447
rect 1477 -2553 1511 -2519
rect 1477 -2625 1511 -2591
rect 1477 -2697 1511 -2663
rect 1477 -2769 1511 -2735
<< metal1 >>
rect -1519 2768 -1469 2782
rect -1519 2734 -1511 2768
rect -1477 2734 -1469 2768
rect -1519 2696 -1469 2734
rect -1519 2662 -1511 2696
rect -1477 2662 -1469 2696
rect -1519 2624 -1469 2662
rect -1519 2590 -1511 2624
rect -1477 2590 -1469 2624
rect -1519 2552 -1469 2590
rect -1519 2518 -1511 2552
rect -1477 2518 -1469 2552
rect -1519 2480 -1469 2518
rect -1519 2446 -1511 2480
rect -1477 2446 -1469 2480
rect -1519 2408 -1469 2446
rect -1519 2374 -1511 2408
rect -1477 2374 -1469 2408
rect -1519 2361 -1469 2374
rect -1353 2768 -1303 2782
rect -1353 2734 -1345 2768
rect -1311 2734 -1303 2768
rect -1353 2696 -1303 2734
rect -1353 2662 -1345 2696
rect -1311 2662 -1303 2696
rect -1353 2624 -1303 2662
rect -1353 2590 -1345 2624
rect -1311 2590 -1303 2624
rect -1353 2552 -1303 2590
rect -1353 2518 -1345 2552
rect -1311 2518 -1303 2552
rect -1353 2480 -1303 2518
rect -1353 2446 -1345 2480
rect -1311 2446 -1303 2480
rect -1353 2408 -1303 2446
rect -1353 2374 -1345 2408
rect -1311 2374 -1303 2408
rect -1353 2361 -1303 2374
rect -1187 2768 -1137 2782
rect -1187 2734 -1179 2768
rect -1145 2734 -1137 2768
rect -1187 2696 -1137 2734
rect -1187 2662 -1179 2696
rect -1145 2662 -1137 2696
rect -1187 2624 -1137 2662
rect -1187 2590 -1179 2624
rect -1145 2590 -1137 2624
rect -1187 2552 -1137 2590
rect -1187 2518 -1179 2552
rect -1145 2518 -1137 2552
rect -1187 2480 -1137 2518
rect -1187 2446 -1179 2480
rect -1145 2446 -1137 2480
rect -1187 2408 -1137 2446
rect -1187 2374 -1179 2408
rect -1145 2374 -1137 2408
rect -1187 2361 -1137 2374
rect -1021 2768 -971 2782
rect -1021 2734 -1013 2768
rect -979 2734 -971 2768
rect -1021 2696 -971 2734
rect -1021 2662 -1013 2696
rect -979 2662 -971 2696
rect -1021 2624 -971 2662
rect -1021 2590 -1013 2624
rect -979 2590 -971 2624
rect -1021 2552 -971 2590
rect -1021 2518 -1013 2552
rect -979 2518 -971 2552
rect -1021 2480 -971 2518
rect -1021 2446 -1013 2480
rect -979 2446 -971 2480
rect -1021 2408 -971 2446
rect -1021 2374 -1013 2408
rect -979 2374 -971 2408
rect -1021 2361 -971 2374
rect -855 2768 -805 2782
rect -855 2734 -847 2768
rect -813 2734 -805 2768
rect -855 2696 -805 2734
rect -855 2662 -847 2696
rect -813 2662 -805 2696
rect -855 2624 -805 2662
rect -855 2590 -847 2624
rect -813 2590 -805 2624
rect -855 2552 -805 2590
rect -855 2518 -847 2552
rect -813 2518 -805 2552
rect -855 2480 -805 2518
rect -855 2446 -847 2480
rect -813 2446 -805 2480
rect -855 2408 -805 2446
rect -855 2374 -847 2408
rect -813 2374 -805 2408
rect -855 2361 -805 2374
rect -689 2768 -639 2782
rect -689 2734 -681 2768
rect -647 2734 -639 2768
rect -689 2696 -639 2734
rect -689 2662 -681 2696
rect -647 2662 -639 2696
rect -689 2624 -639 2662
rect -689 2590 -681 2624
rect -647 2590 -639 2624
rect -689 2552 -639 2590
rect -689 2518 -681 2552
rect -647 2518 -639 2552
rect -689 2480 -639 2518
rect -689 2446 -681 2480
rect -647 2446 -639 2480
rect -689 2408 -639 2446
rect -689 2374 -681 2408
rect -647 2374 -639 2408
rect -689 2361 -639 2374
rect -523 2768 -473 2782
rect -523 2734 -515 2768
rect -481 2734 -473 2768
rect -523 2696 -473 2734
rect -523 2662 -515 2696
rect -481 2662 -473 2696
rect -523 2624 -473 2662
rect -523 2590 -515 2624
rect -481 2590 -473 2624
rect -523 2552 -473 2590
rect -523 2518 -515 2552
rect -481 2518 -473 2552
rect -523 2480 -473 2518
rect -523 2446 -515 2480
rect -481 2446 -473 2480
rect -523 2408 -473 2446
rect -523 2374 -515 2408
rect -481 2374 -473 2408
rect -523 2361 -473 2374
rect -357 2768 -307 2782
rect -357 2734 -349 2768
rect -315 2734 -307 2768
rect -357 2696 -307 2734
rect -357 2662 -349 2696
rect -315 2662 -307 2696
rect -357 2624 -307 2662
rect -357 2590 -349 2624
rect -315 2590 -307 2624
rect -357 2552 -307 2590
rect -357 2518 -349 2552
rect -315 2518 -307 2552
rect -357 2480 -307 2518
rect -357 2446 -349 2480
rect -315 2446 -307 2480
rect -357 2408 -307 2446
rect -357 2374 -349 2408
rect -315 2374 -307 2408
rect -357 2361 -307 2374
rect -191 2768 -141 2782
rect -191 2734 -183 2768
rect -149 2734 -141 2768
rect -191 2696 -141 2734
rect -191 2662 -183 2696
rect -149 2662 -141 2696
rect -191 2624 -141 2662
rect -191 2590 -183 2624
rect -149 2590 -141 2624
rect -191 2552 -141 2590
rect -191 2518 -183 2552
rect -149 2518 -141 2552
rect -191 2480 -141 2518
rect -191 2446 -183 2480
rect -149 2446 -141 2480
rect -191 2408 -141 2446
rect -191 2374 -183 2408
rect -149 2374 -141 2408
rect -191 2361 -141 2374
rect -25 2768 25 2782
rect -25 2734 -17 2768
rect 17 2734 25 2768
rect -25 2696 25 2734
rect -25 2662 -17 2696
rect 17 2662 25 2696
rect -25 2624 25 2662
rect -25 2590 -17 2624
rect 17 2590 25 2624
rect -25 2552 25 2590
rect -25 2518 -17 2552
rect 17 2518 25 2552
rect -25 2480 25 2518
rect -25 2446 -17 2480
rect 17 2446 25 2480
rect -25 2408 25 2446
rect -25 2374 -17 2408
rect 17 2374 25 2408
rect -25 2361 25 2374
rect 141 2768 191 2782
rect 141 2734 149 2768
rect 183 2734 191 2768
rect 141 2696 191 2734
rect 141 2662 149 2696
rect 183 2662 191 2696
rect 141 2624 191 2662
rect 141 2590 149 2624
rect 183 2590 191 2624
rect 141 2552 191 2590
rect 141 2518 149 2552
rect 183 2518 191 2552
rect 141 2480 191 2518
rect 141 2446 149 2480
rect 183 2446 191 2480
rect 141 2408 191 2446
rect 141 2374 149 2408
rect 183 2374 191 2408
rect 141 2361 191 2374
rect 307 2768 357 2782
rect 307 2734 315 2768
rect 349 2734 357 2768
rect 307 2696 357 2734
rect 307 2662 315 2696
rect 349 2662 357 2696
rect 307 2624 357 2662
rect 307 2590 315 2624
rect 349 2590 357 2624
rect 307 2552 357 2590
rect 307 2518 315 2552
rect 349 2518 357 2552
rect 307 2480 357 2518
rect 307 2446 315 2480
rect 349 2446 357 2480
rect 307 2408 357 2446
rect 307 2374 315 2408
rect 349 2374 357 2408
rect 307 2361 357 2374
rect 473 2768 523 2782
rect 473 2734 481 2768
rect 515 2734 523 2768
rect 473 2696 523 2734
rect 473 2662 481 2696
rect 515 2662 523 2696
rect 473 2624 523 2662
rect 473 2590 481 2624
rect 515 2590 523 2624
rect 473 2552 523 2590
rect 473 2518 481 2552
rect 515 2518 523 2552
rect 473 2480 523 2518
rect 473 2446 481 2480
rect 515 2446 523 2480
rect 473 2408 523 2446
rect 473 2374 481 2408
rect 515 2374 523 2408
rect 473 2361 523 2374
rect 639 2768 689 2782
rect 639 2734 647 2768
rect 681 2734 689 2768
rect 639 2696 689 2734
rect 639 2662 647 2696
rect 681 2662 689 2696
rect 639 2624 689 2662
rect 639 2590 647 2624
rect 681 2590 689 2624
rect 639 2552 689 2590
rect 639 2518 647 2552
rect 681 2518 689 2552
rect 639 2480 689 2518
rect 639 2446 647 2480
rect 681 2446 689 2480
rect 639 2408 689 2446
rect 639 2374 647 2408
rect 681 2374 689 2408
rect 639 2361 689 2374
rect 805 2768 855 2782
rect 805 2734 813 2768
rect 847 2734 855 2768
rect 805 2696 855 2734
rect 805 2662 813 2696
rect 847 2662 855 2696
rect 805 2624 855 2662
rect 805 2590 813 2624
rect 847 2590 855 2624
rect 805 2552 855 2590
rect 805 2518 813 2552
rect 847 2518 855 2552
rect 805 2480 855 2518
rect 805 2446 813 2480
rect 847 2446 855 2480
rect 805 2408 855 2446
rect 805 2374 813 2408
rect 847 2374 855 2408
rect 805 2361 855 2374
rect 971 2768 1021 2782
rect 971 2734 979 2768
rect 1013 2734 1021 2768
rect 971 2696 1021 2734
rect 971 2662 979 2696
rect 1013 2662 1021 2696
rect 971 2624 1021 2662
rect 971 2590 979 2624
rect 1013 2590 1021 2624
rect 971 2552 1021 2590
rect 971 2518 979 2552
rect 1013 2518 1021 2552
rect 971 2480 1021 2518
rect 971 2446 979 2480
rect 1013 2446 1021 2480
rect 971 2408 1021 2446
rect 971 2374 979 2408
rect 1013 2374 1021 2408
rect 971 2361 1021 2374
rect 1137 2768 1187 2782
rect 1137 2734 1145 2768
rect 1179 2734 1187 2768
rect 1137 2696 1187 2734
rect 1137 2662 1145 2696
rect 1179 2662 1187 2696
rect 1137 2624 1187 2662
rect 1137 2590 1145 2624
rect 1179 2590 1187 2624
rect 1137 2552 1187 2590
rect 1137 2518 1145 2552
rect 1179 2518 1187 2552
rect 1137 2480 1187 2518
rect 1137 2446 1145 2480
rect 1179 2446 1187 2480
rect 1137 2408 1187 2446
rect 1137 2374 1145 2408
rect 1179 2374 1187 2408
rect 1137 2361 1187 2374
rect 1303 2768 1353 2782
rect 1303 2734 1311 2768
rect 1345 2734 1353 2768
rect 1303 2696 1353 2734
rect 1303 2662 1311 2696
rect 1345 2662 1353 2696
rect 1303 2624 1353 2662
rect 1303 2590 1311 2624
rect 1345 2590 1353 2624
rect 1303 2552 1353 2590
rect 1303 2518 1311 2552
rect 1345 2518 1353 2552
rect 1303 2480 1353 2518
rect 1303 2446 1311 2480
rect 1345 2446 1353 2480
rect 1303 2408 1353 2446
rect 1303 2374 1311 2408
rect 1345 2374 1353 2408
rect 1303 2361 1353 2374
rect 1469 2768 1519 2782
rect 1469 2734 1477 2768
rect 1511 2734 1519 2768
rect 1469 2696 1519 2734
rect 1469 2662 1477 2696
rect 1511 2662 1519 2696
rect 1469 2624 1519 2662
rect 1469 2590 1477 2624
rect 1511 2590 1519 2624
rect 1469 2552 1519 2590
rect 1469 2518 1477 2552
rect 1511 2518 1519 2552
rect 1469 2480 1519 2518
rect 1469 2446 1477 2480
rect 1511 2446 1519 2480
rect 1469 2408 1519 2446
rect 1469 2374 1477 2408
rect 1511 2374 1519 2408
rect 1469 2361 1519 2374
rect -1519 2169 -1469 2183
rect -1519 2135 -1511 2169
rect -1477 2135 -1469 2169
rect -1519 2097 -1469 2135
rect -1519 2063 -1511 2097
rect -1477 2063 -1469 2097
rect -1519 2025 -1469 2063
rect -1519 1991 -1511 2025
rect -1477 1991 -1469 2025
rect -1519 1953 -1469 1991
rect -1519 1919 -1511 1953
rect -1477 1919 -1469 1953
rect -1519 1881 -1469 1919
rect -1519 1847 -1511 1881
rect -1477 1847 -1469 1881
rect -1519 1809 -1469 1847
rect -1519 1775 -1511 1809
rect -1477 1775 -1469 1809
rect -1519 1762 -1469 1775
rect -1353 2169 -1303 2183
rect -1353 2135 -1345 2169
rect -1311 2135 -1303 2169
rect -1353 2097 -1303 2135
rect -1353 2063 -1345 2097
rect -1311 2063 -1303 2097
rect -1353 2025 -1303 2063
rect -1353 1991 -1345 2025
rect -1311 1991 -1303 2025
rect -1353 1953 -1303 1991
rect -1353 1919 -1345 1953
rect -1311 1919 -1303 1953
rect -1353 1881 -1303 1919
rect -1353 1847 -1345 1881
rect -1311 1847 -1303 1881
rect -1353 1809 -1303 1847
rect -1353 1775 -1345 1809
rect -1311 1775 -1303 1809
rect -1353 1762 -1303 1775
rect -1187 2169 -1137 2183
rect -1187 2135 -1179 2169
rect -1145 2135 -1137 2169
rect -1187 2097 -1137 2135
rect -1187 2063 -1179 2097
rect -1145 2063 -1137 2097
rect -1187 2025 -1137 2063
rect -1187 1991 -1179 2025
rect -1145 1991 -1137 2025
rect -1187 1953 -1137 1991
rect -1187 1919 -1179 1953
rect -1145 1919 -1137 1953
rect -1187 1881 -1137 1919
rect -1187 1847 -1179 1881
rect -1145 1847 -1137 1881
rect -1187 1809 -1137 1847
rect -1187 1775 -1179 1809
rect -1145 1775 -1137 1809
rect -1187 1762 -1137 1775
rect -1021 2169 -971 2183
rect -1021 2135 -1013 2169
rect -979 2135 -971 2169
rect -1021 2097 -971 2135
rect -1021 2063 -1013 2097
rect -979 2063 -971 2097
rect -1021 2025 -971 2063
rect -1021 1991 -1013 2025
rect -979 1991 -971 2025
rect -1021 1953 -971 1991
rect -1021 1919 -1013 1953
rect -979 1919 -971 1953
rect -1021 1881 -971 1919
rect -1021 1847 -1013 1881
rect -979 1847 -971 1881
rect -1021 1809 -971 1847
rect -1021 1775 -1013 1809
rect -979 1775 -971 1809
rect -1021 1762 -971 1775
rect -855 2169 -805 2183
rect -855 2135 -847 2169
rect -813 2135 -805 2169
rect -855 2097 -805 2135
rect -855 2063 -847 2097
rect -813 2063 -805 2097
rect -855 2025 -805 2063
rect -855 1991 -847 2025
rect -813 1991 -805 2025
rect -855 1953 -805 1991
rect -855 1919 -847 1953
rect -813 1919 -805 1953
rect -855 1881 -805 1919
rect -855 1847 -847 1881
rect -813 1847 -805 1881
rect -855 1809 -805 1847
rect -855 1775 -847 1809
rect -813 1775 -805 1809
rect -855 1762 -805 1775
rect -689 2169 -639 2183
rect -689 2135 -681 2169
rect -647 2135 -639 2169
rect -689 2097 -639 2135
rect -689 2063 -681 2097
rect -647 2063 -639 2097
rect -689 2025 -639 2063
rect -689 1991 -681 2025
rect -647 1991 -639 2025
rect -689 1953 -639 1991
rect -689 1919 -681 1953
rect -647 1919 -639 1953
rect -689 1881 -639 1919
rect -689 1847 -681 1881
rect -647 1847 -639 1881
rect -689 1809 -639 1847
rect -689 1775 -681 1809
rect -647 1775 -639 1809
rect -689 1762 -639 1775
rect -523 2169 -473 2183
rect -523 2135 -515 2169
rect -481 2135 -473 2169
rect -523 2097 -473 2135
rect -523 2063 -515 2097
rect -481 2063 -473 2097
rect -523 2025 -473 2063
rect -523 1991 -515 2025
rect -481 1991 -473 2025
rect -523 1953 -473 1991
rect -523 1919 -515 1953
rect -481 1919 -473 1953
rect -523 1881 -473 1919
rect -523 1847 -515 1881
rect -481 1847 -473 1881
rect -523 1809 -473 1847
rect -523 1775 -515 1809
rect -481 1775 -473 1809
rect -523 1762 -473 1775
rect -357 2169 -307 2183
rect -357 2135 -349 2169
rect -315 2135 -307 2169
rect -357 2097 -307 2135
rect -357 2063 -349 2097
rect -315 2063 -307 2097
rect -357 2025 -307 2063
rect -357 1991 -349 2025
rect -315 1991 -307 2025
rect -357 1953 -307 1991
rect -357 1919 -349 1953
rect -315 1919 -307 1953
rect -357 1881 -307 1919
rect -357 1847 -349 1881
rect -315 1847 -307 1881
rect -357 1809 -307 1847
rect -357 1775 -349 1809
rect -315 1775 -307 1809
rect -357 1762 -307 1775
rect -191 2169 -141 2183
rect -191 2135 -183 2169
rect -149 2135 -141 2169
rect -191 2097 -141 2135
rect -191 2063 -183 2097
rect -149 2063 -141 2097
rect -191 2025 -141 2063
rect -191 1991 -183 2025
rect -149 1991 -141 2025
rect -191 1953 -141 1991
rect -191 1919 -183 1953
rect -149 1919 -141 1953
rect -191 1881 -141 1919
rect -191 1847 -183 1881
rect -149 1847 -141 1881
rect -191 1809 -141 1847
rect -191 1775 -183 1809
rect -149 1775 -141 1809
rect -191 1762 -141 1775
rect -25 2169 25 2183
rect -25 2135 -17 2169
rect 17 2135 25 2169
rect -25 2097 25 2135
rect -25 2063 -17 2097
rect 17 2063 25 2097
rect -25 2025 25 2063
rect -25 1991 -17 2025
rect 17 1991 25 2025
rect -25 1953 25 1991
rect -25 1919 -17 1953
rect 17 1919 25 1953
rect -25 1881 25 1919
rect -25 1847 -17 1881
rect 17 1847 25 1881
rect -25 1809 25 1847
rect -25 1775 -17 1809
rect 17 1775 25 1809
rect -25 1762 25 1775
rect 141 2169 191 2183
rect 141 2135 149 2169
rect 183 2135 191 2169
rect 141 2097 191 2135
rect 141 2063 149 2097
rect 183 2063 191 2097
rect 141 2025 191 2063
rect 141 1991 149 2025
rect 183 1991 191 2025
rect 141 1953 191 1991
rect 141 1919 149 1953
rect 183 1919 191 1953
rect 141 1881 191 1919
rect 141 1847 149 1881
rect 183 1847 191 1881
rect 141 1809 191 1847
rect 141 1775 149 1809
rect 183 1775 191 1809
rect 141 1762 191 1775
rect 307 2169 357 2183
rect 307 2135 315 2169
rect 349 2135 357 2169
rect 307 2097 357 2135
rect 307 2063 315 2097
rect 349 2063 357 2097
rect 307 2025 357 2063
rect 307 1991 315 2025
rect 349 1991 357 2025
rect 307 1953 357 1991
rect 307 1919 315 1953
rect 349 1919 357 1953
rect 307 1881 357 1919
rect 307 1847 315 1881
rect 349 1847 357 1881
rect 307 1809 357 1847
rect 307 1775 315 1809
rect 349 1775 357 1809
rect 307 1762 357 1775
rect 473 2169 523 2183
rect 473 2135 481 2169
rect 515 2135 523 2169
rect 473 2097 523 2135
rect 473 2063 481 2097
rect 515 2063 523 2097
rect 473 2025 523 2063
rect 473 1991 481 2025
rect 515 1991 523 2025
rect 473 1953 523 1991
rect 473 1919 481 1953
rect 515 1919 523 1953
rect 473 1881 523 1919
rect 473 1847 481 1881
rect 515 1847 523 1881
rect 473 1809 523 1847
rect 473 1775 481 1809
rect 515 1775 523 1809
rect 473 1762 523 1775
rect 639 2169 689 2183
rect 639 2135 647 2169
rect 681 2135 689 2169
rect 639 2097 689 2135
rect 639 2063 647 2097
rect 681 2063 689 2097
rect 639 2025 689 2063
rect 639 1991 647 2025
rect 681 1991 689 2025
rect 639 1953 689 1991
rect 639 1919 647 1953
rect 681 1919 689 1953
rect 639 1881 689 1919
rect 639 1847 647 1881
rect 681 1847 689 1881
rect 639 1809 689 1847
rect 639 1775 647 1809
rect 681 1775 689 1809
rect 639 1762 689 1775
rect 805 2169 855 2183
rect 805 2135 813 2169
rect 847 2135 855 2169
rect 805 2097 855 2135
rect 805 2063 813 2097
rect 847 2063 855 2097
rect 805 2025 855 2063
rect 805 1991 813 2025
rect 847 1991 855 2025
rect 805 1953 855 1991
rect 805 1919 813 1953
rect 847 1919 855 1953
rect 805 1881 855 1919
rect 805 1847 813 1881
rect 847 1847 855 1881
rect 805 1809 855 1847
rect 805 1775 813 1809
rect 847 1775 855 1809
rect 805 1762 855 1775
rect 971 2169 1021 2183
rect 971 2135 979 2169
rect 1013 2135 1021 2169
rect 971 2097 1021 2135
rect 971 2063 979 2097
rect 1013 2063 1021 2097
rect 971 2025 1021 2063
rect 971 1991 979 2025
rect 1013 1991 1021 2025
rect 971 1953 1021 1991
rect 971 1919 979 1953
rect 1013 1919 1021 1953
rect 971 1881 1021 1919
rect 971 1847 979 1881
rect 1013 1847 1021 1881
rect 971 1809 1021 1847
rect 971 1775 979 1809
rect 1013 1775 1021 1809
rect 971 1762 1021 1775
rect 1137 2169 1187 2183
rect 1137 2135 1145 2169
rect 1179 2135 1187 2169
rect 1137 2097 1187 2135
rect 1137 2063 1145 2097
rect 1179 2063 1187 2097
rect 1137 2025 1187 2063
rect 1137 1991 1145 2025
rect 1179 1991 1187 2025
rect 1137 1953 1187 1991
rect 1137 1919 1145 1953
rect 1179 1919 1187 1953
rect 1137 1881 1187 1919
rect 1137 1847 1145 1881
rect 1179 1847 1187 1881
rect 1137 1809 1187 1847
rect 1137 1775 1145 1809
rect 1179 1775 1187 1809
rect 1137 1762 1187 1775
rect 1303 2169 1353 2183
rect 1303 2135 1311 2169
rect 1345 2135 1353 2169
rect 1303 2097 1353 2135
rect 1303 2063 1311 2097
rect 1345 2063 1353 2097
rect 1303 2025 1353 2063
rect 1303 1991 1311 2025
rect 1345 1991 1353 2025
rect 1303 1953 1353 1991
rect 1303 1919 1311 1953
rect 1345 1919 1353 1953
rect 1303 1881 1353 1919
rect 1303 1847 1311 1881
rect 1345 1847 1353 1881
rect 1303 1809 1353 1847
rect 1303 1775 1311 1809
rect 1345 1775 1353 1809
rect 1303 1762 1353 1775
rect 1469 2169 1519 2183
rect 1469 2135 1477 2169
rect 1511 2135 1519 2169
rect 1469 2097 1519 2135
rect 1469 2063 1477 2097
rect 1511 2063 1519 2097
rect 1469 2025 1519 2063
rect 1469 1991 1477 2025
rect 1511 1991 1519 2025
rect 1469 1953 1519 1991
rect 1469 1919 1477 1953
rect 1511 1919 1519 1953
rect 1469 1881 1519 1919
rect 1469 1847 1477 1881
rect 1511 1847 1519 1881
rect 1469 1809 1519 1847
rect 1469 1775 1477 1809
rect 1511 1775 1519 1809
rect 1469 1762 1519 1775
rect -1519 1632 -1469 1646
rect -1519 1598 -1511 1632
rect -1477 1598 -1469 1632
rect -1519 1560 -1469 1598
rect -1519 1526 -1511 1560
rect -1477 1526 -1469 1560
rect -1519 1488 -1469 1526
rect -1519 1454 -1511 1488
rect -1477 1454 -1469 1488
rect -1519 1416 -1469 1454
rect -1519 1382 -1511 1416
rect -1477 1382 -1469 1416
rect -1519 1344 -1469 1382
rect -1519 1310 -1511 1344
rect -1477 1310 -1469 1344
rect -1519 1272 -1469 1310
rect -1519 1238 -1511 1272
rect -1477 1238 -1469 1272
rect -1519 1225 -1469 1238
rect -1353 1632 -1303 1646
rect -1353 1598 -1345 1632
rect -1311 1598 -1303 1632
rect -1353 1560 -1303 1598
rect -1353 1526 -1345 1560
rect -1311 1526 -1303 1560
rect -1353 1488 -1303 1526
rect -1353 1454 -1345 1488
rect -1311 1454 -1303 1488
rect -1353 1416 -1303 1454
rect -1353 1382 -1345 1416
rect -1311 1382 -1303 1416
rect -1353 1344 -1303 1382
rect -1353 1310 -1345 1344
rect -1311 1310 -1303 1344
rect -1353 1272 -1303 1310
rect -1353 1238 -1345 1272
rect -1311 1238 -1303 1272
rect -1353 1225 -1303 1238
rect -1187 1632 -1137 1646
rect -1187 1598 -1179 1632
rect -1145 1598 -1137 1632
rect -1187 1560 -1137 1598
rect -1187 1526 -1179 1560
rect -1145 1526 -1137 1560
rect -1187 1488 -1137 1526
rect -1187 1454 -1179 1488
rect -1145 1454 -1137 1488
rect -1187 1416 -1137 1454
rect -1187 1382 -1179 1416
rect -1145 1382 -1137 1416
rect -1187 1344 -1137 1382
rect -1187 1310 -1179 1344
rect -1145 1310 -1137 1344
rect -1187 1272 -1137 1310
rect -1187 1238 -1179 1272
rect -1145 1238 -1137 1272
rect -1187 1225 -1137 1238
rect -1021 1632 -971 1646
rect -1021 1598 -1013 1632
rect -979 1598 -971 1632
rect -1021 1560 -971 1598
rect -1021 1526 -1013 1560
rect -979 1526 -971 1560
rect -1021 1488 -971 1526
rect -1021 1454 -1013 1488
rect -979 1454 -971 1488
rect -1021 1416 -971 1454
rect -1021 1382 -1013 1416
rect -979 1382 -971 1416
rect -1021 1344 -971 1382
rect -1021 1310 -1013 1344
rect -979 1310 -971 1344
rect -1021 1272 -971 1310
rect -1021 1238 -1013 1272
rect -979 1238 -971 1272
rect -1021 1225 -971 1238
rect -855 1632 -805 1646
rect -855 1598 -847 1632
rect -813 1598 -805 1632
rect -855 1560 -805 1598
rect -855 1526 -847 1560
rect -813 1526 -805 1560
rect -855 1488 -805 1526
rect -855 1454 -847 1488
rect -813 1454 -805 1488
rect -855 1416 -805 1454
rect -855 1382 -847 1416
rect -813 1382 -805 1416
rect -855 1344 -805 1382
rect -855 1310 -847 1344
rect -813 1310 -805 1344
rect -855 1272 -805 1310
rect -855 1238 -847 1272
rect -813 1238 -805 1272
rect -855 1225 -805 1238
rect -689 1632 -639 1646
rect -689 1598 -681 1632
rect -647 1598 -639 1632
rect -689 1560 -639 1598
rect -689 1526 -681 1560
rect -647 1526 -639 1560
rect -689 1488 -639 1526
rect -689 1454 -681 1488
rect -647 1454 -639 1488
rect -689 1416 -639 1454
rect -689 1382 -681 1416
rect -647 1382 -639 1416
rect -689 1344 -639 1382
rect -689 1310 -681 1344
rect -647 1310 -639 1344
rect -689 1272 -639 1310
rect -689 1238 -681 1272
rect -647 1238 -639 1272
rect -689 1225 -639 1238
rect -523 1632 -473 1646
rect -523 1598 -515 1632
rect -481 1598 -473 1632
rect -523 1560 -473 1598
rect -523 1526 -515 1560
rect -481 1526 -473 1560
rect -523 1488 -473 1526
rect -523 1454 -515 1488
rect -481 1454 -473 1488
rect -523 1416 -473 1454
rect -523 1382 -515 1416
rect -481 1382 -473 1416
rect -523 1344 -473 1382
rect -523 1310 -515 1344
rect -481 1310 -473 1344
rect -523 1272 -473 1310
rect -523 1238 -515 1272
rect -481 1238 -473 1272
rect -523 1225 -473 1238
rect -357 1632 -307 1646
rect -357 1598 -349 1632
rect -315 1598 -307 1632
rect -357 1560 -307 1598
rect -357 1526 -349 1560
rect -315 1526 -307 1560
rect -357 1488 -307 1526
rect -357 1454 -349 1488
rect -315 1454 -307 1488
rect -357 1416 -307 1454
rect -357 1382 -349 1416
rect -315 1382 -307 1416
rect -357 1344 -307 1382
rect -357 1310 -349 1344
rect -315 1310 -307 1344
rect -357 1272 -307 1310
rect -357 1238 -349 1272
rect -315 1238 -307 1272
rect -357 1225 -307 1238
rect -191 1632 -141 1646
rect -191 1598 -183 1632
rect -149 1598 -141 1632
rect -191 1560 -141 1598
rect -191 1526 -183 1560
rect -149 1526 -141 1560
rect -191 1488 -141 1526
rect -191 1454 -183 1488
rect -149 1454 -141 1488
rect -191 1416 -141 1454
rect -191 1382 -183 1416
rect -149 1382 -141 1416
rect -191 1344 -141 1382
rect -191 1310 -183 1344
rect -149 1310 -141 1344
rect -191 1272 -141 1310
rect -191 1238 -183 1272
rect -149 1238 -141 1272
rect -191 1225 -141 1238
rect -25 1632 25 1646
rect -25 1598 -17 1632
rect 17 1598 25 1632
rect -25 1560 25 1598
rect -25 1526 -17 1560
rect 17 1526 25 1560
rect -25 1488 25 1526
rect -25 1454 -17 1488
rect 17 1454 25 1488
rect -25 1416 25 1454
rect -25 1382 -17 1416
rect 17 1382 25 1416
rect -25 1344 25 1382
rect -25 1310 -17 1344
rect 17 1310 25 1344
rect -25 1272 25 1310
rect -25 1238 -17 1272
rect 17 1238 25 1272
rect -25 1225 25 1238
rect 141 1632 191 1646
rect 141 1598 149 1632
rect 183 1598 191 1632
rect 141 1560 191 1598
rect 141 1526 149 1560
rect 183 1526 191 1560
rect 141 1488 191 1526
rect 141 1454 149 1488
rect 183 1454 191 1488
rect 141 1416 191 1454
rect 141 1382 149 1416
rect 183 1382 191 1416
rect 141 1344 191 1382
rect 141 1310 149 1344
rect 183 1310 191 1344
rect 141 1272 191 1310
rect 141 1238 149 1272
rect 183 1238 191 1272
rect 141 1225 191 1238
rect 307 1632 357 1646
rect 307 1598 315 1632
rect 349 1598 357 1632
rect 307 1560 357 1598
rect 307 1526 315 1560
rect 349 1526 357 1560
rect 307 1488 357 1526
rect 307 1454 315 1488
rect 349 1454 357 1488
rect 307 1416 357 1454
rect 307 1382 315 1416
rect 349 1382 357 1416
rect 307 1344 357 1382
rect 307 1310 315 1344
rect 349 1310 357 1344
rect 307 1272 357 1310
rect 307 1238 315 1272
rect 349 1238 357 1272
rect 307 1225 357 1238
rect 473 1632 523 1646
rect 473 1598 481 1632
rect 515 1598 523 1632
rect 473 1560 523 1598
rect 473 1526 481 1560
rect 515 1526 523 1560
rect 473 1488 523 1526
rect 473 1454 481 1488
rect 515 1454 523 1488
rect 473 1416 523 1454
rect 473 1382 481 1416
rect 515 1382 523 1416
rect 473 1344 523 1382
rect 473 1310 481 1344
rect 515 1310 523 1344
rect 473 1272 523 1310
rect 473 1238 481 1272
rect 515 1238 523 1272
rect 473 1225 523 1238
rect 639 1632 689 1646
rect 639 1598 647 1632
rect 681 1598 689 1632
rect 639 1560 689 1598
rect 639 1526 647 1560
rect 681 1526 689 1560
rect 639 1488 689 1526
rect 639 1454 647 1488
rect 681 1454 689 1488
rect 639 1416 689 1454
rect 639 1382 647 1416
rect 681 1382 689 1416
rect 639 1344 689 1382
rect 639 1310 647 1344
rect 681 1310 689 1344
rect 639 1272 689 1310
rect 639 1238 647 1272
rect 681 1238 689 1272
rect 639 1225 689 1238
rect 805 1632 855 1646
rect 805 1598 813 1632
rect 847 1598 855 1632
rect 805 1560 855 1598
rect 805 1526 813 1560
rect 847 1526 855 1560
rect 805 1488 855 1526
rect 805 1454 813 1488
rect 847 1454 855 1488
rect 805 1416 855 1454
rect 805 1382 813 1416
rect 847 1382 855 1416
rect 805 1344 855 1382
rect 805 1310 813 1344
rect 847 1310 855 1344
rect 805 1272 855 1310
rect 805 1238 813 1272
rect 847 1238 855 1272
rect 805 1225 855 1238
rect 971 1632 1021 1646
rect 971 1598 979 1632
rect 1013 1598 1021 1632
rect 971 1560 1021 1598
rect 971 1526 979 1560
rect 1013 1526 1021 1560
rect 971 1488 1021 1526
rect 971 1454 979 1488
rect 1013 1454 1021 1488
rect 971 1416 1021 1454
rect 971 1382 979 1416
rect 1013 1382 1021 1416
rect 971 1344 1021 1382
rect 971 1310 979 1344
rect 1013 1310 1021 1344
rect 971 1272 1021 1310
rect 971 1238 979 1272
rect 1013 1238 1021 1272
rect 971 1225 1021 1238
rect 1137 1632 1187 1646
rect 1137 1598 1145 1632
rect 1179 1598 1187 1632
rect 1137 1560 1187 1598
rect 1137 1526 1145 1560
rect 1179 1526 1187 1560
rect 1137 1488 1187 1526
rect 1137 1454 1145 1488
rect 1179 1454 1187 1488
rect 1137 1416 1187 1454
rect 1137 1382 1145 1416
rect 1179 1382 1187 1416
rect 1137 1344 1187 1382
rect 1137 1310 1145 1344
rect 1179 1310 1187 1344
rect 1137 1272 1187 1310
rect 1137 1238 1145 1272
rect 1179 1238 1187 1272
rect 1137 1225 1187 1238
rect 1303 1632 1353 1646
rect 1303 1598 1311 1632
rect 1345 1598 1353 1632
rect 1303 1560 1353 1598
rect 1303 1526 1311 1560
rect 1345 1526 1353 1560
rect 1303 1488 1353 1526
rect 1303 1454 1311 1488
rect 1345 1454 1353 1488
rect 1303 1416 1353 1454
rect 1303 1382 1311 1416
rect 1345 1382 1353 1416
rect 1303 1344 1353 1382
rect 1303 1310 1311 1344
rect 1345 1310 1353 1344
rect 1303 1272 1353 1310
rect 1303 1238 1311 1272
rect 1345 1238 1353 1272
rect 1303 1225 1353 1238
rect 1469 1632 1519 1646
rect 1469 1598 1477 1632
rect 1511 1598 1519 1632
rect 1469 1560 1519 1598
rect 1469 1526 1477 1560
rect 1511 1526 1519 1560
rect 1469 1488 1519 1526
rect 1469 1454 1477 1488
rect 1511 1454 1519 1488
rect 1469 1416 1519 1454
rect 1469 1382 1477 1416
rect 1511 1382 1519 1416
rect 1469 1344 1519 1382
rect 1469 1310 1477 1344
rect 1511 1310 1519 1344
rect 1469 1272 1519 1310
rect 1469 1238 1477 1272
rect 1511 1238 1519 1272
rect 1469 1225 1519 1238
rect -1519 1033 -1469 1047
rect -1519 999 -1511 1033
rect -1477 999 -1469 1033
rect -1519 961 -1469 999
rect -1519 927 -1511 961
rect -1477 927 -1469 961
rect -1519 889 -1469 927
rect -1519 855 -1511 889
rect -1477 855 -1469 889
rect -1519 817 -1469 855
rect -1519 783 -1511 817
rect -1477 783 -1469 817
rect -1519 745 -1469 783
rect -1519 711 -1511 745
rect -1477 711 -1469 745
rect -1519 673 -1469 711
rect -1519 639 -1511 673
rect -1477 639 -1469 673
rect -1519 626 -1469 639
rect -1353 1033 -1303 1047
rect -1353 999 -1345 1033
rect -1311 999 -1303 1033
rect -1353 961 -1303 999
rect -1353 927 -1345 961
rect -1311 927 -1303 961
rect -1353 889 -1303 927
rect -1353 855 -1345 889
rect -1311 855 -1303 889
rect -1353 817 -1303 855
rect -1353 783 -1345 817
rect -1311 783 -1303 817
rect -1353 745 -1303 783
rect -1353 711 -1345 745
rect -1311 711 -1303 745
rect -1353 673 -1303 711
rect -1353 639 -1345 673
rect -1311 639 -1303 673
rect -1353 626 -1303 639
rect -1187 1033 -1137 1047
rect -1187 999 -1179 1033
rect -1145 999 -1137 1033
rect -1187 961 -1137 999
rect -1187 927 -1179 961
rect -1145 927 -1137 961
rect -1187 889 -1137 927
rect -1187 855 -1179 889
rect -1145 855 -1137 889
rect -1187 817 -1137 855
rect -1187 783 -1179 817
rect -1145 783 -1137 817
rect -1187 745 -1137 783
rect -1187 711 -1179 745
rect -1145 711 -1137 745
rect -1187 673 -1137 711
rect -1187 639 -1179 673
rect -1145 639 -1137 673
rect -1187 626 -1137 639
rect -1021 1033 -971 1047
rect -1021 999 -1013 1033
rect -979 999 -971 1033
rect -1021 961 -971 999
rect -1021 927 -1013 961
rect -979 927 -971 961
rect -1021 889 -971 927
rect -1021 855 -1013 889
rect -979 855 -971 889
rect -1021 817 -971 855
rect -1021 783 -1013 817
rect -979 783 -971 817
rect -1021 745 -971 783
rect -1021 711 -1013 745
rect -979 711 -971 745
rect -1021 673 -971 711
rect -1021 639 -1013 673
rect -979 639 -971 673
rect -1021 626 -971 639
rect -855 1033 -805 1047
rect -855 999 -847 1033
rect -813 999 -805 1033
rect -855 961 -805 999
rect -855 927 -847 961
rect -813 927 -805 961
rect -855 889 -805 927
rect -855 855 -847 889
rect -813 855 -805 889
rect -855 817 -805 855
rect -855 783 -847 817
rect -813 783 -805 817
rect -855 745 -805 783
rect -855 711 -847 745
rect -813 711 -805 745
rect -855 673 -805 711
rect -855 639 -847 673
rect -813 639 -805 673
rect -855 626 -805 639
rect -689 1033 -639 1047
rect -689 999 -681 1033
rect -647 999 -639 1033
rect -689 961 -639 999
rect -689 927 -681 961
rect -647 927 -639 961
rect -689 889 -639 927
rect -689 855 -681 889
rect -647 855 -639 889
rect -689 817 -639 855
rect -689 783 -681 817
rect -647 783 -639 817
rect -689 745 -639 783
rect -689 711 -681 745
rect -647 711 -639 745
rect -689 673 -639 711
rect -689 639 -681 673
rect -647 639 -639 673
rect -689 626 -639 639
rect -523 1033 -473 1047
rect -523 999 -515 1033
rect -481 999 -473 1033
rect -523 961 -473 999
rect -523 927 -515 961
rect -481 927 -473 961
rect -523 889 -473 927
rect -523 855 -515 889
rect -481 855 -473 889
rect -523 817 -473 855
rect -523 783 -515 817
rect -481 783 -473 817
rect -523 745 -473 783
rect -523 711 -515 745
rect -481 711 -473 745
rect -523 673 -473 711
rect -523 639 -515 673
rect -481 639 -473 673
rect -523 626 -473 639
rect -357 1033 -307 1047
rect -357 999 -349 1033
rect -315 999 -307 1033
rect -357 961 -307 999
rect -357 927 -349 961
rect -315 927 -307 961
rect -357 889 -307 927
rect -357 855 -349 889
rect -315 855 -307 889
rect -357 817 -307 855
rect -357 783 -349 817
rect -315 783 -307 817
rect -357 745 -307 783
rect -357 711 -349 745
rect -315 711 -307 745
rect -357 673 -307 711
rect -357 639 -349 673
rect -315 639 -307 673
rect -357 626 -307 639
rect -191 1033 -141 1047
rect -191 999 -183 1033
rect -149 999 -141 1033
rect -191 961 -141 999
rect -191 927 -183 961
rect -149 927 -141 961
rect -191 889 -141 927
rect -191 855 -183 889
rect -149 855 -141 889
rect -191 817 -141 855
rect -191 783 -183 817
rect -149 783 -141 817
rect -191 745 -141 783
rect -191 711 -183 745
rect -149 711 -141 745
rect -191 673 -141 711
rect -191 639 -183 673
rect -149 639 -141 673
rect -191 626 -141 639
rect -25 1033 25 1047
rect -25 999 -17 1033
rect 17 999 25 1033
rect -25 961 25 999
rect -25 927 -17 961
rect 17 927 25 961
rect -25 889 25 927
rect -25 855 -17 889
rect 17 855 25 889
rect -25 817 25 855
rect -25 783 -17 817
rect 17 783 25 817
rect -25 745 25 783
rect -25 711 -17 745
rect 17 711 25 745
rect -25 673 25 711
rect -25 639 -17 673
rect 17 639 25 673
rect -25 626 25 639
rect 141 1033 191 1047
rect 141 999 149 1033
rect 183 999 191 1033
rect 141 961 191 999
rect 141 927 149 961
rect 183 927 191 961
rect 141 889 191 927
rect 141 855 149 889
rect 183 855 191 889
rect 141 817 191 855
rect 141 783 149 817
rect 183 783 191 817
rect 141 745 191 783
rect 141 711 149 745
rect 183 711 191 745
rect 141 673 191 711
rect 141 639 149 673
rect 183 639 191 673
rect 141 626 191 639
rect 307 1033 357 1047
rect 307 999 315 1033
rect 349 999 357 1033
rect 307 961 357 999
rect 307 927 315 961
rect 349 927 357 961
rect 307 889 357 927
rect 307 855 315 889
rect 349 855 357 889
rect 307 817 357 855
rect 307 783 315 817
rect 349 783 357 817
rect 307 745 357 783
rect 307 711 315 745
rect 349 711 357 745
rect 307 673 357 711
rect 307 639 315 673
rect 349 639 357 673
rect 307 626 357 639
rect 473 1033 523 1047
rect 473 999 481 1033
rect 515 999 523 1033
rect 473 961 523 999
rect 473 927 481 961
rect 515 927 523 961
rect 473 889 523 927
rect 473 855 481 889
rect 515 855 523 889
rect 473 817 523 855
rect 473 783 481 817
rect 515 783 523 817
rect 473 745 523 783
rect 473 711 481 745
rect 515 711 523 745
rect 473 673 523 711
rect 473 639 481 673
rect 515 639 523 673
rect 473 626 523 639
rect 639 1033 689 1047
rect 639 999 647 1033
rect 681 999 689 1033
rect 639 961 689 999
rect 639 927 647 961
rect 681 927 689 961
rect 639 889 689 927
rect 639 855 647 889
rect 681 855 689 889
rect 639 817 689 855
rect 639 783 647 817
rect 681 783 689 817
rect 639 745 689 783
rect 639 711 647 745
rect 681 711 689 745
rect 639 673 689 711
rect 639 639 647 673
rect 681 639 689 673
rect 639 626 689 639
rect 805 1033 855 1047
rect 805 999 813 1033
rect 847 999 855 1033
rect 805 961 855 999
rect 805 927 813 961
rect 847 927 855 961
rect 805 889 855 927
rect 805 855 813 889
rect 847 855 855 889
rect 805 817 855 855
rect 805 783 813 817
rect 847 783 855 817
rect 805 745 855 783
rect 805 711 813 745
rect 847 711 855 745
rect 805 673 855 711
rect 805 639 813 673
rect 847 639 855 673
rect 805 626 855 639
rect 971 1033 1021 1047
rect 971 999 979 1033
rect 1013 999 1021 1033
rect 971 961 1021 999
rect 971 927 979 961
rect 1013 927 1021 961
rect 971 889 1021 927
rect 971 855 979 889
rect 1013 855 1021 889
rect 971 817 1021 855
rect 971 783 979 817
rect 1013 783 1021 817
rect 971 745 1021 783
rect 971 711 979 745
rect 1013 711 1021 745
rect 971 673 1021 711
rect 971 639 979 673
rect 1013 639 1021 673
rect 971 626 1021 639
rect 1137 1033 1187 1047
rect 1137 999 1145 1033
rect 1179 999 1187 1033
rect 1137 961 1187 999
rect 1137 927 1145 961
rect 1179 927 1187 961
rect 1137 889 1187 927
rect 1137 855 1145 889
rect 1179 855 1187 889
rect 1137 817 1187 855
rect 1137 783 1145 817
rect 1179 783 1187 817
rect 1137 745 1187 783
rect 1137 711 1145 745
rect 1179 711 1187 745
rect 1137 673 1187 711
rect 1137 639 1145 673
rect 1179 639 1187 673
rect 1137 626 1187 639
rect 1303 1033 1353 1047
rect 1303 999 1311 1033
rect 1345 999 1353 1033
rect 1303 961 1353 999
rect 1303 927 1311 961
rect 1345 927 1353 961
rect 1303 889 1353 927
rect 1303 855 1311 889
rect 1345 855 1353 889
rect 1303 817 1353 855
rect 1303 783 1311 817
rect 1345 783 1353 817
rect 1303 745 1353 783
rect 1303 711 1311 745
rect 1345 711 1353 745
rect 1303 673 1353 711
rect 1303 639 1311 673
rect 1345 639 1353 673
rect 1303 626 1353 639
rect 1469 1033 1519 1047
rect 1469 999 1477 1033
rect 1511 999 1519 1033
rect 1469 961 1519 999
rect 1469 927 1477 961
rect 1511 927 1519 961
rect 1469 889 1519 927
rect 1469 855 1477 889
rect 1511 855 1519 889
rect 1469 817 1519 855
rect 1469 783 1477 817
rect 1511 783 1519 817
rect 1469 745 1519 783
rect 1469 711 1477 745
rect 1511 711 1519 745
rect 1469 673 1519 711
rect 1469 639 1477 673
rect 1511 639 1519 673
rect 1469 626 1519 639
rect -1519 496 -1469 510
rect -1519 462 -1511 496
rect -1477 462 -1469 496
rect -1519 424 -1469 462
rect -1519 390 -1511 424
rect -1477 390 -1469 424
rect -1519 352 -1469 390
rect -1519 318 -1511 352
rect -1477 318 -1469 352
rect -1519 280 -1469 318
rect -1519 246 -1511 280
rect -1477 246 -1469 280
rect -1519 208 -1469 246
rect -1519 174 -1511 208
rect -1477 174 -1469 208
rect -1519 136 -1469 174
rect -1519 102 -1511 136
rect -1477 102 -1469 136
rect -1519 89 -1469 102
rect -1353 496 -1303 510
rect -1353 462 -1345 496
rect -1311 462 -1303 496
rect -1353 424 -1303 462
rect -1353 390 -1345 424
rect -1311 390 -1303 424
rect -1353 352 -1303 390
rect -1353 318 -1345 352
rect -1311 318 -1303 352
rect -1353 280 -1303 318
rect -1353 246 -1345 280
rect -1311 246 -1303 280
rect -1353 208 -1303 246
rect -1353 174 -1345 208
rect -1311 174 -1303 208
rect -1353 136 -1303 174
rect -1353 102 -1345 136
rect -1311 102 -1303 136
rect -1353 89 -1303 102
rect -1187 496 -1137 510
rect -1187 462 -1179 496
rect -1145 462 -1137 496
rect -1187 424 -1137 462
rect -1187 390 -1179 424
rect -1145 390 -1137 424
rect -1187 352 -1137 390
rect -1187 318 -1179 352
rect -1145 318 -1137 352
rect -1187 280 -1137 318
rect -1187 246 -1179 280
rect -1145 246 -1137 280
rect -1187 208 -1137 246
rect -1187 174 -1179 208
rect -1145 174 -1137 208
rect -1187 136 -1137 174
rect -1187 102 -1179 136
rect -1145 102 -1137 136
rect -1187 89 -1137 102
rect -1021 496 -971 510
rect -1021 462 -1013 496
rect -979 462 -971 496
rect -1021 424 -971 462
rect -1021 390 -1013 424
rect -979 390 -971 424
rect -1021 352 -971 390
rect -1021 318 -1013 352
rect -979 318 -971 352
rect -1021 280 -971 318
rect -1021 246 -1013 280
rect -979 246 -971 280
rect -1021 208 -971 246
rect -1021 174 -1013 208
rect -979 174 -971 208
rect -1021 136 -971 174
rect -1021 102 -1013 136
rect -979 102 -971 136
rect -1021 89 -971 102
rect -855 496 -805 510
rect -855 462 -847 496
rect -813 462 -805 496
rect -855 424 -805 462
rect -855 390 -847 424
rect -813 390 -805 424
rect -855 352 -805 390
rect -855 318 -847 352
rect -813 318 -805 352
rect -855 280 -805 318
rect -855 246 -847 280
rect -813 246 -805 280
rect -855 208 -805 246
rect -855 174 -847 208
rect -813 174 -805 208
rect -855 136 -805 174
rect -855 102 -847 136
rect -813 102 -805 136
rect -855 89 -805 102
rect -689 496 -639 510
rect -689 462 -681 496
rect -647 462 -639 496
rect -689 424 -639 462
rect -689 390 -681 424
rect -647 390 -639 424
rect -689 352 -639 390
rect -689 318 -681 352
rect -647 318 -639 352
rect -689 280 -639 318
rect -689 246 -681 280
rect -647 246 -639 280
rect -689 208 -639 246
rect -689 174 -681 208
rect -647 174 -639 208
rect -689 136 -639 174
rect -689 102 -681 136
rect -647 102 -639 136
rect -689 89 -639 102
rect -523 496 -473 510
rect -523 462 -515 496
rect -481 462 -473 496
rect -523 424 -473 462
rect -523 390 -515 424
rect -481 390 -473 424
rect -523 352 -473 390
rect -523 318 -515 352
rect -481 318 -473 352
rect -523 280 -473 318
rect -523 246 -515 280
rect -481 246 -473 280
rect -523 208 -473 246
rect -523 174 -515 208
rect -481 174 -473 208
rect -523 136 -473 174
rect -523 102 -515 136
rect -481 102 -473 136
rect -523 89 -473 102
rect -357 496 -307 510
rect -357 462 -349 496
rect -315 462 -307 496
rect -357 424 -307 462
rect -357 390 -349 424
rect -315 390 -307 424
rect -357 352 -307 390
rect -357 318 -349 352
rect -315 318 -307 352
rect -357 280 -307 318
rect -357 246 -349 280
rect -315 246 -307 280
rect -357 208 -307 246
rect -357 174 -349 208
rect -315 174 -307 208
rect -357 136 -307 174
rect -357 102 -349 136
rect -315 102 -307 136
rect -357 89 -307 102
rect -191 496 -141 510
rect -191 462 -183 496
rect -149 462 -141 496
rect -191 424 -141 462
rect -191 390 -183 424
rect -149 390 -141 424
rect -191 352 -141 390
rect -191 318 -183 352
rect -149 318 -141 352
rect -191 280 -141 318
rect -191 246 -183 280
rect -149 246 -141 280
rect -191 208 -141 246
rect -191 174 -183 208
rect -149 174 -141 208
rect -191 136 -141 174
rect -191 102 -183 136
rect -149 102 -141 136
rect -191 89 -141 102
rect -25 496 25 510
rect -25 462 -17 496
rect 17 462 25 496
rect -25 424 25 462
rect -25 390 -17 424
rect 17 390 25 424
rect -25 352 25 390
rect -25 318 -17 352
rect 17 318 25 352
rect -25 280 25 318
rect -25 246 -17 280
rect 17 246 25 280
rect -25 208 25 246
rect -25 174 -17 208
rect 17 174 25 208
rect -25 136 25 174
rect -25 102 -17 136
rect 17 102 25 136
rect -25 89 25 102
rect 141 496 191 510
rect 141 462 149 496
rect 183 462 191 496
rect 141 424 191 462
rect 141 390 149 424
rect 183 390 191 424
rect 141 352 191 390
rect 141 318 149 352
rect 183 318 191 352
rect 141 280 191 318
rect 141 246 149 280
rect 183 246 191 280
rect 141 208 191 246
rect 141 174 149 208
rect 183 174 191 208
rect 141 136 191 174
rect 141 102 149 136
rect 183 102 191 136
rect 141 89 191 102
rect 307 496 357 510
rect 307 462 315 496
rect 349 462 357 496
rect 307 424 357 462
rect 307 390 315 424
rect 349 390 357 424
rect 307 352 357 390
rect 307 318 315 352
rect 349 318 357 352
rect 307 280 357 318
rect 307 246 315 280
rect 349 246 357 280
rect 307 208 357 246
rect 307 174 315 208
rect 349 174 357 208
rect 307 136 357 174
rect 307 102 315 136
rect 349 102 357 136
rect 307 89 357 102
rect 473 496 523 510
rect 473 462 481 496
rect 515 462 523 496
rect 473 424 523 462
rect 473 390 481 424
rect 515 390 523 424
rect 473 352 523 390
rect 473 318 481 352
rect 515 318 523 352
rect 473 280 523 318
rect 473 246 481 280
rect 515 246 523 280
rect 473 208 523 246
rect 473 174 481 208
rect 515 174 523 208
rect 473 136 523 174
rect 473 102 481 136
rect 515 102 523 136
rect 473 89 523 102
rect 639 496 689 510
rect 639 462 647 496
rect 681 462 689 496
rect 639 424 689 462
rect 639 390 647 424
rect 681 390 689 424
rect 639 352 689 390
rect 639 318 647 352
rect 681 318 689 352
rect 639 280 689 318
rect 639 246 647 280
rect 681 246 689 280
rect 639 208 689 246
rect 639 174 647 208
rect 681 174 689 208
rect 639 136 689 174
rect 639 102 647 136
rect 681 102 689 136
rect 639 89 689 102
rect 805 496 855 510
rect 805 462 813 496
rect 847 462 855 496
rect 805 424 855 462
rect 805 390 813 424
rect 847 390 855 424
rect 805 352 855 390
rect 805 318 813 352
rect 847 318 855 352
rect 805 280 855 318
rect 805 246 813 280
rect 847 246 855 280
rect 805 208 855 246
rect 805 174 813 208
rect 847 174 855 208
rect 805 136 855 174
rect 805 102 813 136
rect 847 102 855 136
rect 805 89 855 102
rect 971 496 1021 510
rect 971 462 979 496
rect 1013 462 1021 496
rect 971 424 1021 462
rect 971 390 979 424
rect 1013 390 1021 424
rect 971 352 1021 390
rect 971 318 979 352
rect 1013 318 1021 352
rect 971 280 1021 318
rect 971 246 979 280
rect 1013 246 1021 280
rect 971 208 1021 246
rect 971 174 979 208
rect 1013 174 1021 208
rect 971 136 1021 174
rect 971 102 979 136
rect 1013 102 1021 136
rect 971 89 1021 102
rect 1137 496 1187 510
rect 1137 462 1145 496
rect 1179 462 1187 496
rect 1137 424 1187 462
rect 1137 390 1145 424
rect 1179 390 1187 424
rect 1137 352 1187 390
rect 1137 318 1145 352
rect 1179 318 1187 352
rect 1137 280 1187 318
rect 1137 246 1145 280
rect 1179 246 1187 280
rect 1137 208 1187 246
rect 1137 174 1145 208
rect 1179 174 1187 208
rect 1137 136 1187 174
rect 1137 102 1145 136
rect 1179 102 1187 136
rect 1137 89 1187 102
rect 1303 496 1353 510
rect 1303 462 1311 496
rect 1345 462 1353 496
rect 1303 424 1353 462
rect 1303 390 1311 424
rect 1345 390 1353 424
rect 1303 352 1353 390
rect 1303 318 1311 352
rect 1345 318 1353 352
rect 1303 280 1353 318
rect 1303 246 1311 280
rect 1345 246 1353 280
rect 1303 208 1353 246
rect 1303 174 1311 208
rect 1345 174 1353 208
rect 1303 136 1353 174
rect 1303 102 1311 136
rect 1345 102 1353 136
rect 1303 89 1353 102
rect 1469 496 1519 510
rect 1469 462 1477 496
rect 1511 462 1519 496
rect 1469 424 1519 462
rect 1469 390 1477 424
rect 1511 390 1519 424
rect 1469 352 1519 390
rect 1469 318 1477 352
rect 1511 318 1519 352
rect 1469 280 1519 318
rect 1469 246 1477 280
rect 1511 246 1519 280
rect 1469 208 1519 246
rect 1469 174 1477 208
rect 1511 174 1519 208
rect 1469 136 1519 174
rect 1469 102 1477 136
rect 1511 102 1519 136
rect 1469 89 1519 102
rect -1519 -103 -1469 -89
rect -1519 -137 -1511 -103
rect -1477 -137 -1469 -103
rect -1519 -175 -1469 -137
rect -1519 -209 -1511 -175
rect -1477 -209 -1469 -175
rect -1519 -247 -1469 -209
rect -1519 -281 -1511 -247
rect -1477 -281 -1469 -247
rect -1519 -319 -1469 -281
rect -1519 -353 -1511 -319
rect -1477 -353 -1469 -319
rect -1519 -391 -1469 -353
rect -1519 -425 -1511 -391
rect -1477 -425 -1469 -391
rect -1519 -463 -1469 -425
rect -1519 -497 -1511 -463
rect -1477 -497 -1469 -463
rect -1519 -510 -1469 -497
rect -1353 -103 -1303 -89
rect -1353 -137 -1345 -103
rect -1311 -137 -1303 -103
rect -1353 -175 -1303 -137
rect -1353 -209 -1345 -175
rect -1311 -209 -1303 -175
rect -1353 -247 -1303 -209
rect -1353 -281 -1345 -247
rect -1311 -281 -1303 -247
rect -1353 -319 -1303 -281
rect -1353 -353 -1345 -319
rect -1311 -353 -1303 -319
rect -1353 -391 -1303 -353
rect -1353 -425 -1345 -391
rect -1311 -425 -1303 -391
rect -1353 -463 -1303 -425
rect -1353 -497 -1345 -463
rect -1311 -497 -1303 -463
rect -1353 -510 -1303 -497
rect -1187 -103 -1137 -89
rect -1187 -137 -1179 -103
rect -1145 -137 -1137 -103
rect -1187 -175 -1137 -137
rect -1187 -209 -1179 -175
rect -1145 -209 -1137 -175
rect -1187 -247 -1137 -209
rect -1187 -281 -1179 -247
rect -1145 -281 -1137 -247
rect -1187 -319 -1137 -281
rect -1187 -353 -1179 -319
rect -1145 -353 -1137 -319
rect -1187 -391 -1137 -353
rect -1187 -425 -1179 -391
rect -1145 -425 -1137 -391
rect -1187 -463 -1137 -425
rect -1187 -497 -1179 -463
rect -1145 -497 -1137 -463
rect -1187 -510 -1137 -497
rect -1021 -103 -971 -89
rect -1021 -137 -1013 -103
rect -979 -137 -971 -103
rect -1021 -175 -971 -137
rect -1021 -209 -1013 -175
rect -979 -209 -971 -175
rect -1021 -247 -971 -209
rect -1021 -281 -1013 -247
rect -979 -281 -971 -247
rect -1021 -319 -971 -281
rect -1021 -353 -1013 -319
rect -979 -353 -971 -319
rect -1021 -391 -971 -353
rect -1021 -425 -1013 -391
rect -979 -425 -971 -391
rect -1021 -463 -971 -425
rect -1021 -497 -1013 -463
rect -979 -497 -971 -463
rect -1021 -510 -971 -497
rect -855 -103 -805 -89
rect -855 -137 -847 -103
rect -813 -137 -805 -103
rect -855 -175 -805 -137
rect -855 -209 -847 -175
rect -813 -209 -805 -175
rect -855 -247 -805 -209
rect -855 -281 -847 -247
rect -813 -281 -805 -247
rect -855 -319 -805 -281
rect -855 -353 -847 -319
rect -813 -353 -805 -319
rect -855 -391 -805 -353
rect -855 -425 -847 -391
rect -813 -425 -805 -391
rect -855 -463 -805 -425
rect -855 -497 -847 -463
rect -813 -497 -805 -463
rect -855 -510 -805 -497
rect -689 -103 -639 -89
rect -689 -137 -681 -103
rect -647 -137 -639 -103
rect -689 -175 -639 -137
rect -689 -209 -681 -175
rect -647 -209 -639 -175
rect -689 -247 -639 -209
rect -689 -281 -681 -247
rect -647 -281 -639 -247
rect -689 -319 -639 -281
rect -689 -353 -681 -319
rect -647 -353 -639 -319
rect -689 -391 -639 -353
rect -689 -425 -681 -391
rect -647 -425 -639 -391
rect -689 -463 -639 -425
rect -689 -497 -681 -463
rect -647 -497 -639 -463
rect -689 -510 -639 -497
rect -523 -103 -473 -89
rect -523 -137 -515 -103
rect -481 -137 -473 -103
rect -523 -175 -473 -137
rect -523 -209 -515 -175
rect -481 -209 -473 -175
rect -523 -247 -473 -209
rect -523 -281 -515 -247
rect -481 -281 -473 -247
rect -523 -319 -473 -281
rect -523 -353 -515 -319
rect -481 -353 -473 -319
rect -523 -391 -473 -353
rect -523 -425 -515 -391
rect -481 -425 -473 -391
rect -523 -463 -473 -425
rect -523 -497 -515 -463
rect -481 -497 -473 -463
rect -523 -510 -473 -497
rect -357 -103 -307 -89
rect -357 -137 -349 -103
rect -315 -137 -307 -103
rect -357 -175 -307 -137
rect -357 -209 -349 -175
rect -315 -209 -307 -175
rect -357 -247 -307 -209
rect -357 -281 -349 -247
rect -315 -281 -307 -247
rect -357 -319 -307 -281
rect -357 -353 -349 -319
rect -315 -353 -307 -319
rect -357 -391 -307 -353
rect -357 -425 -349 -391
rect -315 -425 -307 -391
rect -357 -463 -307 -425
rect -357 -497 -349 -463
rect -315 -497 -307 -463
rect -357 -510 -307 -497
rect -191 -103 -141 -89
rect -191 -137 -183 -103
rect -149 -137 -141 -103
rect -191 -175 -141 -137
rect -191 -209 -183 -175
rect -149 -209 -141 -175
rect -191 -247 -141 -209
rect -191 -281 -183 -247
rect -149 -281 -141 -247
rect -191 -319 -141 -281
rect -191 -353 -183 -319
rect -149 -353 -141 -319
rect -191 -391 -141 -353
rect -191 -425 -183 -391
rect -149 -425 -141 -391
rect -191 -463 -141 -425
rect -191 -497 -183 -463
rect -149 -497 -141 -463
rect -191 -510 -141 -497
rect -25 -103 25 -89
rect -25 -137 -17 -103
rect 17 -137 25 -103
rect -25 -175 25 -137
rect -25 -209 -17 -175
rect 17 -209 25 -175
rect -25 -247 25 -209
rect -25 -281 -17 -247
rect 17 -281 25 -247
rect -25 -319 25 -281
rect -25 -353 -17 -319
rect 17 -353 25 -319
rect -25 -391 25 -353
rect -25 -425 -17 -391
rect 17 -425 25 -391
rect -25 -463 25 -425
rect -25 -497 -17 -463
rect 17 -497 25 -463
rect -25 -510 25 -497
rect 141 -103 191 -89
rect 141 -137 149 -103
rect 183 -137 191 -103
rect 141 -175 191 -137
rect 141 -209 149 -175
rect 183 -209 191 -175
rect 141 -247 191 -209
rect 141 -281 149 -247
rect 183 -281 191 -247
rect 141 -319 191 -281
rect 141 -353 149 -319
rect 183 -353 191 -319
rect 141 -391 191 -353
rect 141 -425 149 -391
rect 183 -425 191 -391
rect 141 -463 191 -425
rect 141 -497 149 -463
rect 183 -497 191 -463
rect 141 -510 191 -497
rect 307 -103 357 -89
rect 307 -137 315 -103
rect 349 -137 357 -103
rect 307 -175 357 -137
rect 307 -209 315 -175
rect 349 -209 357 -175
rect 307 -247 357 -209
rect 307 -281 315 -247
rect 349 -281 357 -247
rect 307 -319 357 -281
rect 307 -353 315 -319
rect 349 -353 357 -319
rect 307 -391 357 -353
rect 307 -425 315 -391
rect 349 -425 357 -391
rect 307 -463 357 -425
rect 307 -497 315 -463
rect 349 -497 357 -463
rect 307 -510 357 -497
rect 473 -103 523 -89
rect 473 -137 481 -103
rect 515 -137 523 -103
rect 473 -175 523 -137
rect 473 -209 481 -175
rect 515 -209 523 -175
rect 473 -247 523 -209
rect 473 -281 481 -247
rect 515 -281 523 -247
rect 473 -319 523 -281
rect 473 -353 481 -319
rect 515 -353 523 -319
rect 473 -391 523 -353
rect 473 -425 481 -391
rect 515 -425 523 -391
rect 473 -463 523 -425
rect 473 -497 481 -463
rect 515 -497 523 -463
rect 473 -510 523 -497
rect 639 -103 689 -89
rect 639 -137 647 -103
rect 681 -137 689 -103
rect 639 -175 689 -137
rect 639 -209 647 -175
rect 681 -209 689 -175
rect 639 -247 689 -209
rect 639 -281 647 -247
rect 681 -281 689 -247
rect 639 -319 689 -281
rect 639 -353 647 -319
rect 681 -353 689 -319
rect 639 -391 689 -353
rect 639 -425 647 -391
rect 681 -425 689 -391
rect 639 -463 689 -425
rect 639 -497 647 -463
rect 681 -497 689 -463
rect 639 -510 689 -497
rect 805 -103 855 -89
rect 805 -137 813 -103
rect 847 -137 855 -103
rect 805 -175 855 -137
rect 805 -209 813 -175
rect 847 -209 855 -175
rect 805 -247 855 -209
rect 805 -281 813 -247
rect 847 -281 855 -247
rect 805 -319 855 -281
rect 805 -353 813 -319
rect 847 -353 855 -319
rect 805 -391 855 -353
rect 805 -425 813 -391
rect 847 -425 855 -391
rect 805 -463 855 -425
rect 805 -497 813 -463
rect 847 -497 855 -463
rect 805 -510 855 -497
rect 971 -103 1021 -89
rect 971 -137 979 -103
rect 1013 -137 1021 -103
rect 971 -175 1021 -137
rect 971 -209 979 -175
rect 1013 -209 1021 -175
rect 971 -247 1021 -209
rect 971 -281 979 -247
rect 1013 -281 1021 -247
rect 971 -319 1021 -281
rect 971 -353 979 -319
rect 1013 -353 1021 -319
rect 971 -391 1021 -353
rect 971 -425 979 -391
rect 1013 -425 1021 -391
rect 971 -463 1021 -425
rect 971 -497 979 -463
rect 1013 -497 1021 -463
rect 971 -510 1021 -497
rect 1137 -103 1187 -89
rect 1137 -137 1145 -103
rect 1179 -137 1187 -103
rect 1137 -175 1187 -137
rect 1137 -209 1145 -175
rect 1179 -209 1187 -175
rect 1137 -247 1187 -209
rect 1137 -281 1145 -247
rect 1179 -281 1187 -247
rect 1137 -319 1187 -281
rect 1137 -353 1145 -319
rect 1179 -353 1187 -319
rect 1137 -391 1187 -353
rect 1137 -425 1145 -391
rect 1179 -425 1187 -391
rect 1137 -463 1187 -425
rect 1137 -497 1145 -463
rect 1179 -497 1187 -463
rect 1137 -510 1187 -497
rect 1303 -103 1353 -89
rect 1303 -137 1311 -103
rect 1345 -137 1353 -103
rect 1303 -175 1353 -137
rect 1303 -209 1311 -175
rect 1345 -209 1353 -175
rect 1303 -247 1353 -209
rect 1303 -281 1311 -247
rect 1345 -281 1353 -247
rect 1303 -319 1353 -281
rect 1303 -353 1311 -319
rect 1345 -353 1353 -319
rect 1303 -391 1353 -353
rect 1303 -425 1311 -391
rect 1345 -425 1353 -391
rect 1303 -463 1353 -425
rect 1303 -497 1311 -463
rect 1345 -497 1353 -463
rect 1303 -510 1353 -497
rect 1469 -103 1519 -89
rect 1469 -137 1477 -103
rect 1511 -137 1519 -103
rect 1469 -175 1519 -137
rect 1469 -209 1477 -175
rect 1511 -209 1519 -175
rect 1469 -247 1519 -209
rect 1469 -281 1477 -247
rect 1511 -281 1519 -247
rect 1469 -319 1519 -281
rect 1469 -353 1477 -319
rect 1511 -353 1519 -319
rect 1469 -391 1519 -353
rect 1469 -425 1477 -391
rect 1511 -425 1519 -391
rect 1469 -463 1519 -425
rect 1469 -497 1477 -463
rect 1511 -497 1519 -463
rect 1469 -510 1519 -497
rect -1519 -640 -1469 -626
rect -1519 -674 -1511 -640
rect -1477 -674 -1469 -640
rect -1519 -712 -1469 -674
rect -1519 -746 -1511 -712
rect -1477 -746 -1469 -712
rect -1519 -784 -1469 -746
rect -1519 -818 -1511 -784
rect -1477 -818 -1469 -784
rect -1519 -856 -1469 -818
rect -1519 -890 -1511 -856
rect -1477 -890 -1469 -856
rect -1519 -928 -1469 -890
rect -1519 -962 -1511 -928
rect -1477 -962 -1469 -928
rect -1519 -1000 -1469 -962
rect -1519 -1034 -1511 -1000
rect -1477 -1034 -1469 -1000
rect -1519 -1047 -1469 -1034
rect -1353 -640 -1303 -626
rect -1353 -674 -1345 -640
rect -1311 -674 -1303 -640
rect -1353 -712 -1303 -674
rect -1353 -746 -1345 -712
rect -1311 -746 -1303 -712
rect -1353 -784 -1303 -746
rect -1353 -818 -1345 -784
rect -1311 -818 -1303 -784
rect -1353 -856 -1303 -818
rect -1353 -890 -1345 -856
rect -1311 -890 -1303 -856
rect -1353 -928 -1303 -890
rect -1353 -962 -1345 -928
rect -1311 -962 -1303 -928
rect -1353 -1000 -1303 -962
rect -1353 -1034 -1345 -1000
rect -1311 -1034 -1303 -1000
rect -1353 -1047 -1303 -1034
rect -1187 -640 -1137 -626
rect -1187 -674 -1179 -640
rect -1145 -674 -1137 -640
rect -1187 -712 -1137 -674
rect -1187 -746 -1179 -712
rect -1145 -746 -1137 -712
rect -1187 -784 -1137 -746
rect -1187 -818 -1179 -784
rect -1145 -818 -1137 -784
rect -1187 -856 -1137 -818
rect -1187 -890 -1179 -856
rect -1145 -890 -1137 -856
rect -1187 -928 -1137 -890
rect -1187 -962 -1179 -928
rect -1145 -962 -1137 -928
rect -1187 -1000 -1137 -962
rect -1187 -1034 -1179 -1000
rect -1145 -1034 -1137 -1000
rect -1187 -1047 -1137 -1034
rect -1021 -640 -971 -626
rect -1021 -674 -1013 -640
rect -979 -674 -971 -640
rect -1021 -712 -971 -674
rect -1021 -746 -1013 -712
rect -979 -746 -971 -712
rect -1021 -784 -971 -746
rect -1021 -818 -1013 -784
rect -979 -818 -971 -784
rect -1021 -856 -971 -818
rect -1021 -890 -1013 -856
rect -979 -890 -971 -856
rect -1021 -928 -971 -890
rect -1021 -962 -1013 -928
rect -979 -962 -971 -928
rect -1021 -1000 -971 -962
rect -1021 -1034 -1013 -1000
rect -979 -1034 -971 -1000
rect -1021 -1047 -971 -1034
rect -855 -640 -805 -626
rect -855 -674 -847 -640
rect -813 -674 -805 -640
rect -855 -712 -805 -674
rect -855 -746 -847 -712
rect -813 -746 -805 -712
rect -855 -784 -805 -746
rect -855 -818 -847 -784
rect -813 -818 -805 -784
rect -855 -856 -805 -818
rect -855 -890 -847 -856
rect -813 -890 -805 -856
rect -855 -928 -805 -890
rect -855 -962 -847 -928
rect -813 -962 -805 -928
rect -855 -1000 -805 -962
rect -855 -1034 -847 -1000
rect -813 -1034 -805 -1000
rect -855 -1047 -805 -1034
rect -689 -640 -639 -626
rect -689 -674 -681 -640
rect -647 -674 -639 -640
rect -689 -712 -639 -674
rect -689 -746 -681 -712
rect -647 -746 -639 -712
rect -689 -784 -639 -746
rect -689 -818 -681 -784
rect -647 -818 -639 -784
rect -689 -856 -639 -818
rect -689 -890 -681 -856
rect -647 -890 -639 -856
rect -689 -928 -639 -890
rect -689 -962 -681 -928
rect -647 -962 -639 -928
rect -689 -1000 -639 -962
rect -689 -1034 -681 -1000
rect -647 -1034 -639 -1000
rect -689 -1047 -639 -1034
rect -523 -640 -473 -626
rect -523 -674 -515 -640
rect -481 -674 -473 -640
rect -523 -712 -473 -674
rect -523 -746 -515 -712
rect -481 -746 -473 -712
rect -523 -784 -473 -746
rect -523 -818 -515 -784
rect -481 -818 -473 -784
rect -523 -856 -473 -818
rect -523 -890 -515 -856
rect -481 -890 -473 -856
rect -523 -928 -473 -890
rect -523 -962 -515 -928
rect -481 -962 -473 -928
rect -523 -1000 -473 -962
rect -523 -1034 -515 -1000
rect -481 -1034 -473 -1000
rect -523 -1047 -473 -1034
rect -357 -640 -307 -626
rect -357 -674 -349 -640
rect -315 -674 -307 -640
rect -357 -712 -307 -674
rect -357 -746 -349 -712
rect -315 -746 -307 -712
rect -357 -784 -307 -746
rect -357 -818 -349 -784
rect -315 -818 -307 -784
rect -357 -856 -307 -818
rect -357 -890 -349 -856
rect -315 -890 -307 -856
rect -357 -928 -307 -890
rect -357 -962 -349 -928
rect -315 -962 -307 -928
rect -357 -1000 -307 -962
rect -357 -1034 -349 -1000
rect -315 -1034 -307 -1000
rect -357 -1047 -307 -1034
rect -191 -640 -141 -626
rect -191 -674 -183 -640
rect -149 -674 -141 -640
rect -191 -712 -141 -674
rect -191 -746 -183 -712
rect -149 -746 -141 -712
rect -191 -784 -141 -746
rect -191 -818 -183 -784
rect -149 -818 -141 -784
rect -191 -856 -141 -818
rect -191 -890 -183 -856
rect -149 -890 -141 -856
rect -191 -928 -141 -890
rect -191 -962 -183 -928
rect -149 -962 -141 -928
rect -191 -1000 -141 -962
rect -191 -1034 -183 -1000
rect -149 -1034 -141 -1000
rect -191 -1047 -141 -1034
rect -25 -640 25 -626
rect -25 -674 -17 -640
rect 17 -674 25 -640
rect -25 -712 25 -674
rect -25 -746 -17 -712
rect 17 -746 25 -712
rect -25 -784 25 -746
rect -25 -818 -17 -784
rect 17 -818 25 -784
rect -25 -856 25 -818
rect -25 -890 -17 -856
rect 17 -890 25 -856
rect -25 -928 25 -890
rect -25 -962 -17 -928
rect 17 -962 25 -928
rect -25 -1000 25 -962
rect -25 -1034 -17 -1000
rect 17 -1034 25 -1000
rect -25 -1047 25 -1034
rect 141 -640 191 -626
rect 141 -674 149 -640
rect 183 -674 191 -640
rect 141 -712 191 -674
rect 141 -746 149 -712
rect 183 -746 191 -712
rect 141 -784 191 -746
rect 141 -818 149 -784
rect 183 -818 191 -784
rect 141 -856 191 -818
rect 141 -890 149 -856
rect 183 -890 191 -856
rect 141 -928 191 -890
rect 141 -962 149 -928
rect 183 -962 191 -928
rect 141 -1000 191 -962
rect 141 -1034 149 -1000
rect 183 -1034 191 -1000
rect 141 -1047 191 -1034
rect 307 -640 357 -626
rect 307 -674 315 -640
rect 349 -674 357 -640
rect 307 -712 357 -674
rect 307 -746 315 -712
rect 349 -746 357 -712
rect 307 -784 357 -746
rect 307 -818 315 -784
rect 349 -818 357 -784
rect 307 -856 357 -818
rect 307 -890 315 -856
rect 349 -890 357 -856
rect 307 -928 357 -890
rect 307 -962 315 -928
rect 349 -962 357 -928
rect 307 -1000 357 -962
rect 307 -1034 315 -1000
rect 349 -1034 357 -1000
rect 307 -1047 357 -1034
rect 473 -640 523 -626
rect 473 -674 481 -640
rect 515 -674 523 -640
rect 473 -712 523 -674
rect 473 -746 481 -712
rect 515 -746 523 -712
rect 473 -784 523 -746
rect 473 -818 481 -784
rect 515 -818 523 -784
rect 473 -856 523 -818
rect 473 -890 481 -856
rect 515 -890 523 -856
rect 473 -928 523 -890
rect 473 -962 481 -928
rect 515 -962 523 -928
rect 473 -1000 523 -962
rect 473 -1034 481 -1000
rect 515 -1034 523 -1000
rect 473 -1047 523 -1034
rect 639 -640 689 -626
rect 639 -674 647 -640
rect 681 -674 689 -640
rect 639 -712 689 -674
rect 639 -746 647 -712
rect 681 -746 689 -712
rect 639 -784 689 -746
rect 639 -818 647 -784
rect 681 -818 689 -784
rect 639 -856 689 -818
rect 639 -890 647 -856
rect 681 -890 689 -856
rect 639 -928 689 -890
rect 639 -962 647 -928
rect 681 -962 689 -928
rect 639 -1000 689 -962
rect 639 -1034 647 -1000
rect 681 -1034 689 -1000
rect 639 -1047 689 -1034
rect 805 -640 855 -626
rect 805 -674 813 -640
rect 847 -674 855 -640
rect 805 -712 855 -674
rect 805 -746 813 -712
rect 847 -746 855 -712
rect 805 -784 855 -746
rect 805 -818 813 -784
rect 847 -818 855 -784
rect 805 -856 855 -818
rect 805 -890 813 -856
rect 847 -890 855 -856
rect 805 -928 855 -890
rect 805 -962 813 -928
rect 847 -962 855 -928
rect 805 -1000 855 -962
rect 805 -1034 813 -1000
rect 847 -1034 855 -1000
rect 805 -1047 855 -1034
rect 971 -640 1021 -626
rect 971 -674 979 -640
rect 1013 -674 1021 -640
rect 971 -712 1021 -674
rect 971 -746 979 -712
rect 1013 -746 1021 -712
rect 971 -784 1021 -746
rect 971 -818 979 -784
rect 1013 -818 1021 -784
rect 971 -856 1021 -818
rect 971 -890 979 -856
rect 1013 -890 1021 -856
rect 971 -928 1021 -890
rect 971 -962 979 -928
rect 1013 -962 1021 -928
rect 971 -1000 1021 -962
rect 971 -1034 979 -1000
rect 1013 -1034 1021 -1000
rect 971 -1047 1021 -1034
rect 1137 -640 1187 -626
rect 1137 -674 1145 -640
rect 1179 -674 1187 -640
rect 1137 -712 1187 -674
rect 1137 -746 1145 -712
rect 1179 -746 1187 -712
rect 1137 -784 1187 -746
rect 1137 -818 1145 -784
rect 1179 -818 1187 -784
rect 1137 -856 1187 -818
rect 1137 -890 1145 -856
rect 1179 -890 1187 -856
rect 1137 -928 1187 -890
rect 1137 -962 1145 -928
rect 1179 -962 1187 -928
rect 1137 -1000 1187 -962
rect 1137 -1034 1145 -1000
rect 1179 -1034 1187 -1000
rect 1137 -1047 1187 -1034
rect 1303 -640 1353 -626
rect 1303 -674 1311 -640
rect 1345 -674 1353 -640
rect 1303 -712 1353 -674
rect 1303 -746 1311 -712
rect 1345 -746 1353 -712
rect 1303 -784 1353 -746
rect 1303 -818 1311 -784
rect 1345 -818 1353 -784
rect 1303 -856 1353 -818
rect 1303 -890 1311 -856
rect 1345 -890 1353 -856
rect 1303 -928 1353 -890
rect 1303 -962 1311 -928
rect 1345 -962 1353 -928
rect 1303 -1000 1353 -962
rect 1303 -1034 1311 -1000
rect 1345 -1034 1353 -1000
rect 1303 -1047 1353 -1034
rect 1469 -640 1519 -626
rect 1469 -674 1477 -640
rect 1511 -674 1519 -640
rect 1469 -712 1519 -674
rect 1469 -746 1477 -712
rect 1511 -746 1519 -712
rect 1469 -784 1519 -746
rect 1469 -818 1477 -784
rect 1511 -818 1519 -784
rect 1469 -856 1519 -818
rect 1469 -890 1477 -856
rect 1511 -890 1519 -856
rect 1469 -928 1519 -890
rect 1469 -962 1477 -928
rect 1511 -962 1519 -928
rect 1469 -1000 1519 -962
rect 1469 -1034 1477 -1000
rect 1511 -1034 1519 -1000
rect 1469 -1047 1519 -1034
rect -1519 -1239 -1469 -1225
rect -1519 -1273 -1511 -1239
rect -1477 -1273 -1469 -1239
rect -1519 -1311 -1469 -1273
rect -1519 -1345 -1511 -1311
rect -1477 -1345 -1469 -1311
rect -1519 -1383 -1469 -1345
rect -1519 -1417 -1511 -1383
rect -1477 -1417 -1469 -1383
rect -1519 -1455 -1469 -1417
rect -1519 -1489 -1511 -1455
rect -1477 -1489 -1469 -1455
rect -1519 -1527 -1469 -1489
rect -1519 -1561 -1511 -1527
rect -1477 -1561 -1469 -1527
rect -1519 -1599 -1469 -1561
rect -1519 -1633 -1511 -1599
rect -1477 -1633 -1469 -1599
rect -1519 -1646 -1469 -1633
rect -1353 -1239 -1303 -1225
rect -1353 -1273 -1345 -1239
rect -1311 -1273 -1303 -1239
rect -1353 -1311 -1303 -1273
rect -1353 -1345 -1345 -1311
rect -1311 -1345 -1303 -1311
rect -1353 -1383 -1303 -1345
rect -1353 -1417 -1345 -1383
rect -1311 -1417 -1303 -1383
rect -1353 -1455 -1303 -1417
rect -1353 -1489 -1345 -1455
rect -1311 -1489 -1303 -1455
rect -1353 -1527 -1303 -1489
rect -1353 -1561 -1345 -1527
rect -1311 -1561 -1303 -1527
rect -1353 -1599 -1303 -1561
rect -1353 -1633 -1345 -1599
rect -1311 -1633 -1303 -1599
rect -1353 -1646 -1303 -1633
rect -1187 -1239 -1137 -1225
rect -1187 -1273 -1179 -1239
rect -1145 -1273 -1137 -1239
rect -1187 -1311 -1137 -1273
rect -1187 -1345 -1179 -1311
rect -1145 -1345 -1137 -1311
rect -1187 -1383 -1137 -1345
rect -1187 -1417 -1179 -1383
rect -1145 -1417 -1137 -1383
rect -1187 -1455 -1137 -1417
rect -1187 -1489 -1179 -1455
rect -1145 -1489 -1137 -1455
rect -1187 -1527 -1137 -1489
rect -1187 -1561 -1179 -1527
rect -1145 -1561 -1137 -1527
rect -1187 -1599 -1137 -1561
rect -1187 -1633 -1179 -1599
rect -1145 -1633 -1137 -1599
rect -1187 -1646 -1137 -1633
rect -1021 -1239 -971 -1225
rect -1021 -1273 -1013 -1239
rect -979 -1273 -971 -1239
rect -1021 -1311 -971 -1273
rect -1021 -1345 -1013 -1311
rect -979 -1345 -971 -1311
rect -1021 -1383 -971 -1345
rect -1021 -1417 -1013 -1383
rect -979 -1417 -971 -1383
rect -1021 -1455 -971 -1417
rect -1021 -1489 -1013 -1455
rect -979 -1489 -971 -1455
rect -1021 -1527 -971 -1489
rect -1021 -1561 -1013 -1527
rect -979 -1561 -971 -1527
rect -1021 -1599 -971 -1561
rect -1021 -1633 -1013 -1599
rect -979 -1633 -971 -1599
rect -1021 -1646 -971 -1633
rect -855 -1239 -805 -1225
rect -855 -1273 -847 -1239
rect -813 -1273 -805 -1239
rect -855 -1311 -805 -1273
rect -855 -1345 -847 -1311
rect -813 -1345 -805 -1311
rect -855 -1383 -805 -1345
rect -855 -1417 -847 -1383
rect -813 -1417 -805 -1383
rect -855 -1455 -805 -1417
rect -855 -1489 -847 -1455
rect -813 -1489 -805 -1455
rect -855 -1527 -805 -1489
rect -855 -1561 -847 -1527
rect -813 -1561 -805 -1527
rect -855 -1599 -805 -1561
rect -855 -1633 -847 -1599
rect -813 -1633 -805 -1599
rect -855 -1646 -805 -1633
rect -689 -1239 -639 -1225
rect -689 -1273 -681 -1239
rect -647 -1273 -639 -1239
rect -689 -1311 -639 -1273
rect -689 -1345 -681 -1311
rect -647 -1345 -639 -1311
rect -689 -1383 -639 -1345
rect -689 -1417 -681 -1383
rect -647 -1417 -639 -1383
rect -689 -1455 -639 -1417
rect -689 -1489 -681 -1455
rect -647 -1489 -639 -1455
rect -689 -1527 -639 -1489
rect -689 -1561 -681 -1527
rect -647 -1561 -639 -1527
rect -689 -1599 -639 -1561
rect -689 -1633 -681 -1599
rect -647 -1633 -639 -1599
rect -689 -1646 -639 -1633
rect -523 -1239 -473 -1225
rect -523 -1273 -515 -1239
rect -481 -1273 -473 -1239
rect -523 -1311 -473 -1273
rect -523 -1345 -515 -1311
rect -481 -1345 -473 -1311
rect -523 -1383 -473 -1345
rect -523 -1417 -515 -1383
rect -481 -1417 -473 -1383
rect -523 -1455 -473 -1417
rect -523 -1489 -515 -1455
rect -481 -1489 -473 -1455
rect -523 -1527 -473 -1489
rect -523 -1561 -515 -1527
rect -481 -1561 -473 -1527
rect -523 -1599 -473 -1561
rect -523 -1633 -515 -1599
rect -481 -1633 -473 -1599
rect -523 -1646 -473 -1633
rect -357 -1239 -307 -1225
rect -357 -1273 -349 -1239
rect -315 -1273 -307 -1239
rect -357 -1311 -307 -1273
rect -357 -1345 -349 -1311
rect -315 -1345 -307 -1311
rect -357 -1383 -307 -1345
rect -357 -1417 -349 -1383
rect -315 -1417 -307 -1383
rect -357 -1455 -307 -1417
rect -357 -1489 -349 -1455
rect -315 -1489 -307 -1455
rect -357 -1527 -307 -1489
rect -357 -1561 -349 -1527
rect -315 -1561 -307 -1527
rect -357 -1599 -307 -1561
rect -357 -1633 -349 -1599
rect -315 -1633 -307 -1599
rect -357 -1646 -307 -1633
rect -191 -1239 -141 -1225
rect -191 -1273 -183 -1239
rect -149 -1273 -141 -1239
rect -191 -1311 -141 -1273
rect -191 -1345 -183 -1311
rect -149 -1345 -141 -1311
rect -191 -1383 -141 -1345
rect -191 -1417 -183 -1383
rect -149 -1417 -141 -1383
rect -191 -1455 -141 -1417
rect -191 -1489 -183 -1455
rect -149 -1489 -141 -1455
rect -191 -1527 -141 -1489
rect -191 -1561 -183 -1527
rect -149 -1561 -141 -1527
rect -191 -1599 -141 -1561
rect -191 -1633 -183 -1599
rect -149 -1633 -141 -1599
rect -191 -1646 -141 -1633
rect -25 -1239 25 -1225
rect -25 -1273 -17 -1239
rect 17 -1273 25 -1239
rect -25 -1311 25 -1273
rect -25 -1345 -17 -1311
rect 17 -1345 25 -1311
rect -25 -1383 25 -1345
rect -25 -1417 -17 -1383
rect 17 -1417 25 -1383
rect -25 -1455 25 -1417
rect -25 -1489 -17 -1455
rect 17 -1489 25 -1455
rect -25 -1527 25 -1489
rect -25 -1561 -17 -1527
rect 17 -1561 25 -1527
rect -25 -1599 25 -1561
rect -25 -1633 -17 -1599
rect 17 -1633 25 -1599
rect -25 -1646 25 -1633
rect 141 -1239 191 -1225
rect 141 -1273 149 -1239
rect 183 -1273 191 -1239
rect 141 -1311 191 -1273
rect 141 -1345 149 -1311
rect 183 -1345 191 -1311
rect 141 -1383 191 -1345
rect 141 -1417 149 -1383
rect 183 -1417 191 -1383
rect 141 -1455 191 -1417
rect 141 -1489 149 -1455
rect 183 -1489 191 -1455
rect 141 -1527 191 -1489
rect 141 -1561 149 -1527
rect 183 -1561 191 -1527
rect 141 -1599 191 -1561
rect 141 -1633 149 -1599
rect 183 -1633 191 -1599
rect 141 -1646 191 -1633
rect 307 -1239 357 -1225
rect 307 -1273 315 -1239
rect 349 -1273 357 -1239
rect 307 -1311 357 -1273
rect 307 -1345 315 -1311
rect 349 -1345 357 -1311
rect 307 -1383 357 -1345
rect 307 -1417 315 -1383
rect 349 -1417 357 -1383
rect 307 -1455 357 -1417
rect 307 -1489 315 -1455
rect 349 -1489 357 -1455
rect 307 -1527 357 -1489
rect 307 -1561 315 -1527
rect 349 -1561 357 -1527
rect 307 -1599 357 -1561
rect 307 -1633 315 -1599
rect 349 -1633 357 -1599
rect 307 -1646 357 -1633
rect 473 -1239 523 -1225
rect 473 -1273 481 -1239
rect 515 -1273 523 -1239
rect 473 -1311 523 -1273
rect 473 -1345 481 -1311
rect 515 -1345 523 -1311
rect 473 -1383 523 -1345
rect 473 -1417 481 -1383
rect 515 -1417 523 -1383
rect 473 -1455 523 -1417
rect 473 -1489 481 -1455
rect 515 -1489 523 -1455
rect 473 -1527 523 -1489
rect 473 -1561 481 -1527
rect 515 -1561 523 -1527
rect 473 -1599 523 -1561
rect 473 -1633 481 -1599
rect 515 -1633 523 -1599
rect 473 -1646 523 -1633
rect 639 -1239 689 -1225
rect 639 -1273 647 -1239
rect 681 -1273 689 -1239
rect 639 -1311 689 -1273
rect 639 -1345 647 -1311
rect 681 -1345 689 -1311
rect 639 -1383 689 -1345
rect 639 -1417 647 -1383
rect 681 -1417 689 -1383
rect 639 -1455 689 -1417
rect 639 -1489 647 -1455
rect 681 -1489 689 -1455
rect 639 -1527 689 -1489
rect 639 -1561 647 -1527
rect 681 -1561 689 -1527
rect 639 -1599 689 -1561
rect 639 -1633 647 -1599
rect 681 -1633 689 -1599
rect 639 -1646 689 -1633
rect 805 -1239 855 -1225
rect 805 -1273 813 -1239
rect 847 -1273 855 -1239
rect 805 -1311 855 -1273
rect 805 -1345 813 -1311
rect 847 -1345 855 -1311
rect 805 -1383 855 -1345
rect 805 -1417 813 -1383
rect 847 -1417 855 -1383
rect 805 -1455 855 -1417
rect 805 -1489 813 -1455
rect 847 -1489 855 -1455
rect 805 -1527 855 -1489
rect 805 -1561 813 -1527
rect 847 -1561 855 -1527
rect 805 -1599 855 -1561
rect 805 -1633 813 -1599
rect 847 -1633 855 -1599
rect 805 -1646 855 -1633
rect 971 -1239 1021 -1225
rect 971 -1273 979 -1239
rect 1013 -1273 1021 -1239
rect 971 -1311 1021 -1273
rect 971 -1345 979 -1311
rect 1013 -1345 1021 -1311
rect 971 -1383 1021 -1345
rect 971 -1417 979 -1383
rect 1013 -1417 1021 -1383
rect 971 -1455 1021 -1417
rect 971 -1489 979 -1455
rect 1013 -1489 1021 -1455
rect 971 -1527 1021 -1489
rect 971 -1561 979 -1527
rect 1013 -1561 1021 -1527
rect 971 -1599 1021 -1561
rect 971 -1633 979 -1599
rect 1013 -1633 1021 -1599
rect 971 -1646 1021 -1633
rect 1137 -1239 1187 -1225
rect 1137 -1273 1145 -1239
rect 1179 -1273 1187 -1239
rect 1137 -1311 1187 -1273
rect 1137 -1345 1145 -1311
rect 1179 -1345 1187 -1311
rect 1137 -1383 1187 -1345
rect 1137 -1417 1145 -1383
rect 1179 -1417 1187 -1383
rect 1137 -1455 1187 -1417
rect 1137 -1489 1145 -1455
rect 1179 -1489 1187 -1455
rect 1137 -1527 1187 -1489
rect 1137 -1561 1145 -1527
rect 1179 -1561 1187 -1527
rect 1137 -1599 1187 -1561
rect 1137 -1633 1145 -1599
rect 1179 -1633 1187 -1599
rect 1137 -1646 1187 -1633
rect 1303 -1239 1353 -1225
rect 1303 -1273 1311 -1239
rect 1345 -1273 1353 -1239
rect 1303 -1311 1353 -1273
rect 1303 -1345 1311 -1311
rect 1345 -1345 1353 -1311
rect 1303 -1383 1353 -1345
rect 1303 -1417 1311 -1383
rect 1345 -1417 1353 -1383
rect 1303 -1455 1353 -1417
rect 1303 -1489 1311 -1455
rect 1345 -1489 1353 -1455
rect 1303 -1527 1353 -1489
rect 1303 -1561 1311 -1527
rect 1345 -1561 1353 -1527
rect 1303 -1599 1353 -1561
rect 1303 -1633 1311 -1599
rect 1345 -1633 1353 -1599
rect 1303 -1646 1353 -1633
rect 1469 -1239 1519 -1225
rect 1469 -1273 1477 -1239
rect 1511 -1273 1519 -1239
rect 1469 -1311 1519 -1273
rect 1469 -1345 1477 -1311
rect 1511 -1345 1519 -1311
rect 1469 -1383 1519 -1345
rect 1469 -1417 1477 -1383
rect 1511 -1417 1519 -1383
rect 1469 -1455 1519 -1417
rect 1469 -1489 1477 -1455
rect 1511 -1489 1519 -1455
rect 1469 -1527 1519 -1489
rect 1469 -1561 1477 -1527
rect 1511 -1561 1519 -1527
rect 1469 -1599 1519 -1561
rect 1469 -1633 1477 -1599
rect 1511 -1633 1519 -1599
rect 1469 -1646 1519 -1633
rect -1519 -1776 -1469 -1762
rect -1519 -1810 -1511 -1776
rect -1477 -1810 -1469 -1776
rect -1519 -1848 -1469 -1810
rect -1519 -1882 -1511 -1848
rect -1477 -1882 -1469 -1848
rect -1519 -1920 -1469 -1882
rect -1519 -1954 -1511 -1920
rect -1477 -1954 -1469 -1920
rect -1519 -1992 -1469 -1954
rect -1519 -2026 -1511 -1992
rect -1477 -2026 -1469 -1992
rect -1519 -2064 -1469 -2026
rect -1519 -2098 -1511 -2064
rect -1477 -2098 -1469 -2064
rect -1519 -2136 -1469 -2098
rect -1519 -2170 -1511 -2136
rect -1477 -2170 -1469 -2136
rect -1519 -2183 -1469 -2170
rect -1353 -1776 -1303 -1762
rect -1353 -1810 -1345 -1776
rect -1311 -1810 -1303 -1776
rect -1353 -1848 -1303 -1810
rect -1353 -1882 -1345 -1848
rect -1311 -1882 -1303 -1848
rect -1353 -1920 -1303 -1882
rect -1353 -1954 -1345 -1920
rect -1311 -1954 -1303 -1920
rect -1353 -1992 -1303 -1954
rect -1353 -2026 -1345 -1992
rect -1311 -2026 -1303 -1992
rect -1353 -2064 -1303 -2026
rect -1353 -2098 -1345 -2064
rect -1311 -2098 -1303 -2064
rect -1353 -2136 -1303 -2098
rect -1353 -2170 -1345 -2136
rect -1311 -2170 -1303 -2136
rect -1353 -2183 -1303 -2170
rect -1187 -1776 -1137 -1762
rect -1187 -1810 -1179 -1776
rect -1145 -1810 -1137 -1776
rect -1187 -1848 -1137 -1810
rect -1187 -1882 -1179 -1848
rect -1145 -1882 -1137 -1848
rect -1187 -1920 -1137 -1882
rect -1187 -1954 -1179 -1920
rect -1145 -1954 -1137 -1920
rect -1187 -1992 -1137 -1954
rect -1187 -2026 -1179 -1992
rect -1145 -2026 -1137 -1992
rect -1187 -2064 -1137 -2026
rect -1187 -2098 -1179 -2064
rect -1145 -2098 -1137 -2064
rect -1187 -2136 -1137 -2098
rect -1187 -2170 -1179 -2136
rect -1145 -2170 -1137 -2136
rect -1187 -2183 -1137 -2170
rect -1021 -1776 -971 -1762
rect -1021 -1810 -1013 -1776
rect -979 -1810 -971 -1776
rect -1021 -1848 -971 -1810
rect -1021 -1882 -1013 -1848
rect -979 -1882 -971 -1848
rect -1021 -1920 -971 -1882
rect -1021 -1954 -1013 -1920
rect -979 -1954 -971 -1920
rect -1021 -1992 -971 -1954
rect -1021 -2026 -1013 -1992
rect -979 -2026 -971 -1992
rect -1021 -2064 -971 -2026
rect -1021 -2098 -1013 -2064
rect -979 -2098 -971 -2064
rect -1021 -2136 -971 -2098
rect -1021 -2170 -1013 -2136
rect -979 -2170 -971 -2136
rect -1021 -2183 -971 -2170
rect -855 -1776 -805 -1762
rect -855 -1810 -847 -1776
rect -813 -1810 -805 -1776
rect -855 -1848 -805 -1810
rect -855 -1882 -847 -1848
rect -813 -1882 -805 -1848
rect -855 -1920 -805 -1882
rect -855 -1954 -847 -1920
rect -813 -1954 -805 -1920
rect -855 -1992 -805 -1954
rect -855 -2026 -847 -1992
rect -813 -2026 -805 -1992
rect -855 -2064 -805 -2026
rect -855 -2098 -847 -2064
rect -813 -2098 -805 -2064
rect -855 -2136 -805 -2098
rect -855 -2170 -847 -2136
rect -813 -2170 -805 -2136
rect -855 -2183 -805 -2170
rect -689 -1776 -639 -1762
rect -689 -1810 -681 -1776
rect -647 -1810 -639 -1776
rect -689 -1848 -639 -1810
rect -689 -1882 -681 -1848
rect -647 -1882 -639 -1848
rect -689 -1920 -639 -1882
rect -689 -1954 -681 -1920
rect -647 -1954 -639 -1920
rect -689 -1992 -639 -1954
rect -689 -2026 -681 -1992
rect -647 -2026 -639 -1992
rect -689 -2064 -639 -2026
rect -689 -2098 -681 -2064
rect -647 -2098 -639 -2064
rect -689 -2136 -639 -2098
rect -689 -2170 -681 -2136
rect -647 -2170 -639 -2136
rect -689 -2183 -639 -2170
rect -523 -1776 -473 -1762
rect -523 -1810 -515 -1776
rect -481 -1810 -473 -1776
rect -523 -1848 -473 -1810
rect -523 -1882 -515 -1848
rect -481 -1882 -473 -1848
rect -523 -1920 -473 -1882
rect -523 -1954 -515 -1920
rect -481 -1954 -473 -1920
rect -523 -1992 -473 -1954
rect -523 -2026 -515 -1992
rect -481 -2026 -473 -1992
rect -523 -2064 -473 -2026
rect -523 -2098 -515 -2064
rect -481 -2098 -473 -2064
rect -523 -2136 -473 -2098
rect -523 -2170 -515 -2136
rect -481 -2170 -473 -2136
rect -523 -2183 -473 -2170
rect -357 -1776 -307 -1762
rect -357 -1810 -349 -1776
rect -315 -1810 -307 -1776
rect -357 -1848 -307 -1810
rect -357 -1882 -349 -1848
rect -315 -1882 -307 -1848
rect -357 -1920 -307 -1882
rect -357 -1954 -349 -1920
rect -315 -1954 -307 -1920
rect -357 -1992 -307 -1954
rect -357 -2026 -349 -1992
rect -315 -2026 -307 -1992
rect -357 -2064 -307 -2026
rect -357 -2098 -349 -2064
rect -315 -2098 -307 -2064
rect -357 -2136 -307 -2098
rect -357 -2170 -349 -2136
rect -315 -2170 -307 -2136
rect -357 -2183 -307 -2170
rect -191 -1776 -141 -1762
rect -191 -1810 -183 -1776
rect -149 -1810 -141 -1776
rect -191 -1848 -141 -1810
rect -191 -1882 -183 -1848
rect -149 -1882 -141 -1848
rect -191 -1920 -141 -1882
rect -191 -1954 -183 -1920
rect -149 -1954 -141 -1920
rect -191 -1992 -141 -1954
rect -191 -2026 -183 -1992
rect -149 -2026 -141 -1992
rect -191 -2064 -141 -2026
rect -191 -2098 -183 -2064
rect -149 -2098 -141 -2064
rect -191 -2136 -141 -2098
rect -191 -2170 -183 -2136
rect -149 -2170 -141 -2136
rect -191 -2183 -141 -2170
rect -25 -1776 25 -1762
rect -25 -1810 -17 -1776
rect 17 -1810 25 -1776
rect -25 -1848 25 -1810
rect -25 -1882 -17 -1848
rect 17 -1882 25 -1848
rect -25 -1920 25 -1882
rect -25 -1954 -17 -1920
rect 17 -1954 25 -1920
rect -25 -1992 25 -1954
rect -25 -2026 -17 -1992
rect 17 -2026 25 -1992
rect -25 -2064 25 -2026
rect -25 -2098 -17 -2064
rect 17 -2098 25 -2064
rect -25 -2136 25 -2098
rect -25 -2170 -17 -2136
rect 17 -2170 25 -2136
rect -25 -2183 25 -2170
rect 141 -1776 191 -1762
rect 141 -1810 149 -1776
rect 183 -1810 191 -1776
rect 141 -1848 191 -1810
rect 141 -1882 149 -1848
rect 183 -1882 191 -1848
rect 141 -1920 191 -1882
rect 141 -1954 149 -1920
rect 183 -1954 191 -1920
rect 141 -1992 191 -1954
rect 141 -2026 149 -1992
rect 183 -2026 191 -1992
rect 141 -2064 191 -2026
rect 141 -2098 149 -2064
rect 183 -2098 191 -2064
rect 141 -2136 191 -2098
rect 141 -2170 149 -2136
rect 183 -2170 191 -2136
rect 141 -2183 191 -2170
rect 307 -1776 357 -1762
rect 307 -1810 315 -1776
rect 349 -1810 357 -1776
rect 307 -1848 357 -1810
rect 307 -1882 315 -1848
rect 349 -1882 357 -1848
rect 307 -1920 357 -1882
rect 307 -1954 315 -1920
rect 349 -1954 357 -1920
rect 307 -1992 357 -1954
rect 307 -2026 315 -1992
rect 349 -2026 357 -1992
rect 307 -2064 357 -2026
rect 307 -2098 315 -2064
rect 349 -2098 357 -2064
rect 307 -2136 357 -2098
rect 307 -2170 315 -2136
rect 349 -2170 357 -2136
rect 307 -2183 357 -2170
rect 473 -1776 523 -1762
rect 473 -1810 481 -1776
rect 515 -1810 523 -1776
rect 473 -1848 523 -1810
rect 473 -1882 481 -1848
rect 515 -1882 523 -1848
rect 473 -1920 523 -1882
rect 473 -1954 481 -1920
rect 515 -1954 523 -1920
rect 473 -1992 523 -1954
rect 473 -2026 481 -1992
rect 515 -2026 523 -1992
rect 473 -2064 523 -2026
rect 473 -2098 481 -2064
rect 515 -2098 523 -2064
rect 473 -2136 523 -2098
rect 473 -2170 481 -2136
rect 515 -2170 523 -2136
rect 473 -2183 523 -2170
rect 639 -1776 689 -1762
rect 639 -1810 647 -1776
rect 681 -1810 689 -1776
rect 639 -1848 689 -1810
rect 639 -1882 647 -1848
rect 681 -1882 689 -1848
rect 639 -1920 689 -1882
rect 639 -1954 647 -1920
rect 681 -1954 689 -1920
rect 639 -1992 689 -1954
rect 639 -2026 647 -1992
rect 681 -2026 689 -1992
rect 639 -2064 689 -2026
rect 639 -2098 647 -2064
rect 681 -2098 689 -2064
rect 639 -2136 689 -2098
rect 639 -2170 647 -2136
rect 681 -2170 689 -2136
rect 639 -2183 689 -2170
rect 805 -1776 855 -1762
rect 805 -1810 813 -1776
rect 847 -1810 855 -1776
rect 805 -1848 855 -1810
rect 805 -1882 813 -1848
rect 847 -1882 855 -1848
rect 805 -1920 855 -1882
rect 805 -1954 813 -1920
rect 847 -1954 855 -1920
rect 805 -1992 855 -1954
rect 805 -2026 813 -1992
rect 847 -2026 855 -1992
rect 805 -2064 855 -2026
rect 805 -2098 813 -2064
rect 847 -2098 855 -2064
rect 805 -2136 855 -2098
rect 805 -2170 813 -2136
rect 847 -2170 855 -2136
rect 805 -2183 855 -2170
rect 971 -1776 1021 -1762
rect 971 -1810 979 -1776
rect 1013 -1810 1021 -1776
rect 971 -1848 1021 -1810
rect 971 -1882 979 -1848
rect 1013 -1882 1021 -1848
rect 971 -1920 1021 -1882
rect 971 -1954 979 -1920
rect 1013 -1954 1021 -1920
rect 971 -1992 1021 -1954
rect 971 -2026 979 -1992
rect 1013 -2026 1021 -1992
rect 971 -2064 1021 -2026
rect 971 -2098 979 -2064
rect 1013 -2098 1021 -2064
rect 971 -2136 1021 -2098
rect 971 -2170 979 -2136
rect 1013 -2170 1021 -2136
rect 971 -2183 1021 -2170
rect 1137 -1776 1187 -1762
rect 1137 -1810 1145 -1776
rect 1179 -1810 1187 -1776
rect 1137 -1848 1187 -1810
rect 1137 -1882 1145 -1848
rect 1179 -1882 1187 -1848
rect 1137 -1920 1187 -1882
rect 1137 -1954 1145 -1920
rect 1179 -1954 1187 -1920
rect 1137 -1992 1187 -1954
rect 1137 -2026 1145 -1992
rect 1179 -2026 1187 -1992
rect 1137 -2064 1187 -2026
rect 1137 -2098 1145 -2064
rect 1179 -2098 1187 -2064
rect 1137 -2136 1187 -2098
rect 1137 -2170 1145 -2136
rect 1179 -2170 1187 -2136
rect 1137 -2183 1187 -2170
rect 1303 -1776 1353 -1762
rect 1303 -1810 1311 -1776
rect 1345 -1810 1353 -1776
rect 1303 -1848 1353 -1810
rect 1303 -1882 1311 -1848
rect 1345 -1882 1353 -1848
rect 1303 -1920 1353 -1882
rect 1303 -1954 1311 -1920
rect 1345 -1954 1353 -1920
rect 1303 -1992 1353 -1954
rect 1303 -2026 1311 -1992
rect 1345 -2026 1353 -1992
rect 1303 -2064 1353 -2026
rect 1303 -2098 1311 -2064
rect 1345 -2098 1353 -2064
rect 1303 -2136 1353 -2098
rect 1303 -2170 1311 -2136
rect 1345 -2170 1353 -2136
rect 1303 -2183 1353 -2170
rect 1469 -1776 1519 -1762
rect 1469 -1810 1477 -1776
rect 1511 -1810 1519 -1776
rect 1469 -1848 1519 -1810
rect 1469 -1882 1477 -1848
rect 1511 -1882 1519 -1848
rect 1469 -1920 1519 -1882
rect 1469 -1954 1477 -1920
rect 1511 -1954 1519 -1920
rect 1469 -1992 1519 -1954
rect 1469 -2026 1477 -1992
rect 1511 -2026 1519 -1992
rect 1469 -2064 1519 -2026
rect 1469 -2098 1477 -2064
rect 1511 -2098 1519 -2064
rect 1469 -2136 1519 -2098
rect 1469 -2170 1477 -2136
rect 1511 -2170 1519 -2136
rect 1469 -2183 1519 -2170
rect -1519 -2375 -1469 -2361
rect -1519 -2409 -1511 -2375
rect -1477 -2409 -1469 -2375
rect -1519 -2447 -1469 -2409
rect -1519 -2481 -1511 -2447
rect -1477 -2481 -1469 -2447
rect -1519 -2519 -1469 -2481
rect -1519 -2553 -1511 -2519
rect -1477 -2553 -1469 -2519
rect -1519 -2591 -1469 -2553
rect -1519 -2625 -1511 -2591
rect -1477 -2625 -1469 -2591
rect -1519 -2663 -1469 -2625
rect -1519 -2697 -1511 -2663
rect -1477 -2697 -1469 -2663
rect -1519 -2735 -1469 -2697
rect -1519 -2769 -1511 -2735
rect -1477 -2769 -1469 -2735
rect -1519 -2782 -1469 -2769
rect -1353 -2375 -1303 -2361
rect -1353 -2409 -1345 -2375
rect -1311 -2409 -1303 -2375
rect -1353 -2447 -1303 -2409
rect -1353 -2481 -1345 -2447
rect -1311 -2481 -1303 -2447
rect -1353 -2519 -1303 -2481
rect -1353 -2553 -1345 -2519
rect -1311 -2553 -1303 -2519
rect -1353 -2591 -1303 -2553
rect -1353 -2625 -1345 -2591
rect -1311 -2625 -1303 -2591
rect -1353 -2663 -1303 -2625
rect -1353 -2697 -1345 -2663
rect -1311 -2697 -1303 -2663
rect -1353 -2735 -1303 -2697
rect -1353 -2769 -1345 -2735
rect -1311 -2769 -1303 -2735
rect -1353 -2782 -1303 -2769
rect -1187 -2375 -1137 -2361
rect -1187 -2409 -1179 -2375
rect -1145 -2409 -1137 -2375
rect -1187 -2447 -1137 -2409
rect -1187 -2481 -1179 -2447
rect -1145 -2481 -1137 -2447
rect -1187 -2519 -1137 -2481
rect -1187 -2553 -1179 -2519
rect -1145 -2553 -1137 -2519
rect -1187 -2591 -1137 -2553
rect -1187 -2625 -1179 -2591
rect -1145 -2625 -1137 -2591
rect -1187 -2663 -1137 -2625
rect -1187 -2697 -1179 -2663
rect -1145 -2697 -1137 -2663
rect -1187 -2735 -1137 -2697
rect -1187 -2769 -1179 -2735
rect -1145 -2769 -1137 -2735
rect -1187 -2782 -1137 -2769
rect -1021 -2375 -971 -2361
rect -1021 -2409 -1013 -2375
rect -979 -2409 -971 -2375
rect -1021 -2447 -971 -2409
rect -1021 -2481 -1013 -2447
rect -979 -2481 -971 -2447
rect -1021 -2519 -971 -2481
rect -1021 -2553 -1013 -2519
rect -979 -2553 -971 -2519
rect -1021 -2591 -971 -2553
rect -1021 -2625 -1013 -2591
rect -979 -2625 -971 -2591
rect -1021 -2663 -971 -2625
rect -1021 -2697 -1013 -2663
rect -979 -2697 -971 -2663
rect -1021 -2735 -971 -2697
rect -1021 -2769 -1013 -2735
rect -979 -2769 -971 -2735
rect -1021 -2782 -971 -2769
rect -855 -2375 -805 -2361
rect -855 -2409 -847 -2375
rect -813 -2409 -805 -2375
rect -855 -2447 -805 -2409
rect -855 -2481 -847 -2447
rect -813 -2481 -805 -2447
rect -855 -2519 -805 -2481
rect -855 -2553 -847 -2519
rect -813 -2553 -805 -2519
rect -855 -2591 -805 -2553
rect -855 -2625 -847 -2591
rect -813 -2625 -805 -2591
rect -855 -2663 -805 -2625
rect -855 -2697 -847 -2663
rect -813 -2697 -805 -2663
rect -855 -2735 -805 -2697
rect -855 -2769 -847 -2735
rect -813 -2769 -805 -2735
rect -855 -2782 -805 -2769
rect -689 -2375 -639 -2361
rect -689 -2409 -681 -2375
rect -647 -2409 -639 -2375
rect -689 -2447 -639 -2409
rect -689 -2481 -681 -2447
rect -647 -2481 -639 -2447
rect -689 -2519 -639 -2481
rect -689 -2553 -681 -2519
rect -647 -2553 -639 -2519
rect -689 -2591 -639 -2553
rect -689 -2625 -681 -2591
rect -647 -2625 -639 -2591
rect -689 -2663 -639 -2625
rect -689 -2697 -681 -2663
rect -647 -2697 -639 -2663
rect -689 -2735 -639 -2697
rect -689 -2769 -681 -2735
rect -647 -2769 -639 -2735
rect -689 -2782 -639 -2769
rect -523 -2375 -473 -2361
rect -523 -2409 -515 -2375
rect -481 -2409 -473 -2375
rect -523 -2447 -473 -2409
rect -523 -2481 -515 -2447
rect -481 -2481 -473 -2447
rect -523 -2519 -473 -2481
rect -523 -2553 -515 -2519
rect -481 -2553 -473 -2519
rect -523 -2591 -473 -2553
rect -523 -2625 -515 -2591
rect -481 -2625 -473 -2591
rect -523 -2663 -473 -2625
rect -523 -2697 -515 -2663
rect -481 -2697 -473 -2663
rect -523 -2735 -473 -2697
rect -523 -2769 -515 -2735
rect -481 -2769 -473 -2735
rect -523 -2782 -473 -2769
rect -357 -2375 -307 -2361
rect -357 -2409 -349 -2375
rect -315 -2409 -307 -2375
rect -357 -2447 -307 -2409
rect -357 -2481 -349 -2447
rect -315 -2481 -307 -2447
rect -357 -2519 -307 -2481
rect -357 -2553 -349 -2519
rect -315 -2553 -307 -2519
rect -357 -2591 -307 -2553
rect -357 -2625 -349 -2591
rect -315 -2625 -307 -2591
rect -357 -2663 -307 -2625
rect -357 -2697 -349 -2663
rect -315 -2697 -307 -2663
rect -357 -2735 -307 -2697
rect -357 -2769 -349 -2735
rect -315 -2769 -307 -2735
rect -357 -2782 -307 -2769
rect -191 -2375 -141 -2361
rect -191 -2409 -183 -2375
rect -149 -2409 -141 -2375
rect -191 -2447 -141 -2409
rect -191 -2481 -183 -2447
rect -149 -2481 -141 -2447
rect -191 -2519 -141 -2481
rect -191 -2553 -183 -2519
rect -149 -2553 -141 -2519
rect -191 -2591 -141 -2553
rect -191 -2625 -183 -2591
rect -149 -2625 -141 -2591
rect -191 -2663 -141 -2625
rect -191 -2697 -183 -2663
rect -149 -2697 -141 -2663
rect -191 -2735 -141 -2697
rect -191 -2769 -183 -2735
rect -149 -2769 -141 -2735
rect -191 -2782 -141 -2769
rect -25 -2375 25 -2361
rect -25 -2409 -17 -2375
rect 17 -2409 25 -2375
rect -25 -2447 25 -2409
rect -25 -2481 -17 -2447
rect 17 -2481 25 -2447
rect -25 -2519 25 -2481
rect -25 -2553 -17 -2519
rect 17 -2553 25 -2519
rect -25 -2591 25 -2553
rect -25 -2625 -17 -2591
rect 17 -2625 25 -2591
rect -25 -2663 25 -2625
rect -25 -2697 -17 -2663
rect 17 -2697 25 -2663
rect -25 -2735 25 -2697
rect -25 -2769 -17 -2735
rect 17 -2769 25 -2735
rect -25 -2782 25 -2769
rect 141 -2375 191 -2361
rect 141 -2409 149 -2375
rect 183 -2409 191 -2375
rect 141 -2447 191 -2409
rect 141 -2481 149 -2447
rect 183 -2481 191 -2447
rect 141 -2519 191 -2481
rect 141 -2553 149 -2519
rect 183 -2553 191 -2519
rect 141 -2591 191 -2553
rect 141 -2625 149 -2591
rect 183 -2625 191 -2591
rect 141 -2663 191 -2625
rect 141 -2697 149 -2663
rect 183 -2697 191 -2663
rect 141 -2735 191 -2697
rect 141 -2769 149 -2735
rect 183 -2769 191 -2735
rect 141 -2782 191 -2769
rect 307 -2375 357 -2361
rect 307 -2409 315 -2375
rect 349 -2409 357 -2375
rect 307 -2447 357 -2409
rect 307 -2481 315 -2447
rect 349 -2481 357 -2447
rect 307 -2519 357 -2481
rect 307 -2553 315 -2519
rect 349 -2553 357 -2519
rect 307 -2591 357 -2553
rect 307 -2625 315 -2591
rect 349 -2625 357 -2591
rect 307 -2663 357 -2625
rect 307 -2697 315 -2663
rect 349 -2697 357 -2663
rect 307 -2735 357 -2697
rect 307 -2769 315 -2735
rect 349 -2769 357 -2735
rect 307 -2782 357 -2769
rect 473 -2375 523 -2361
rect 473 -2409 481 -2375
rect 515 -2409 523 -2375
rect 473 -2447 523 -2409
rect 473 -2481 481 -2447
rect 515 -2481 523 -2447
rect 473 -2519 523 -2481
rect 473 -2553 481 -2519
rect 515 -2553 523 -2519
rect 473 -2591 523 -2553
rect 473 -2625 481 -2591
rect 515 -2625 523 -2591
rect 473 -2663 523 -2625
rect 473 -2697 481 -2663
rect 515 -2697 523 -2663
rect 473 -2735 523 -2697
rect 473 -2769 481 -2735
rect 515 -2769 523 -2735
rect 473 -2782 523 -2769
rect 639 -2375 689 -2361
rect 639 -2409 647 -2375
rect 681 -2409 689 -2375
rect 639 -2447 689 -2409
rect 639 -2481 647 -2447
rect 681 -2481 689 -2447
rect 639 -2519 689 -2481
rect 639 -2553 647 -2519
rect 681 -2553 689 -2519
rect 639 -2591 689 -2553
rect 639 -2625 647 -2591
rect 681 -2625 689 -2591
rect 639 -2663 689 -2625
rect 639 -2697 647 -2663
rect 681 -2697 689 -2663
rect 639 -2735 689 -2697
rect 639 -2769 647 -2735
rect 681 -2769 689 -2735
rect 639 -2782 689 -2769
rect 805 -2375 855 -2361
rect 805 -2409 813 -2375
rect 847 -2409 855 -2375
rect 805 -2447 855 -2409
rect 805 -2481 813 -2447
rect 847 -2481 855 -2447
rect 805 -2519 855 -2481
rect 805 -2553 813 -2519
rect 847 -2553 855 -2519
rect 805 -2591 855 -2553
rect 805 -2625 813 -2591
rect 847 -2625 855 -2591
rect 805 -2663 855 -2625
rect 805 -2697 813 -2663
rect 847 -2697 855 -2663
rect 805 -2735 855 -2697
rect 805 -2769 813 -2735
rect 847 -2769 855 -2735
rect 805 -2782 855 -2769
rect 971 -2375 1021 -2361
rect 971 -2409 979 -2375
rect 1013 -2409 1021 -2375
rect 971 -2447 1021 -2409
rect 971 -2481 979 -2447
rect 1013 -2481 1021 -2447
rect 971 -2519 1021 -2481
rect 971 -2553 979 -2519
rect 1013 -2553 1021 -2519
rect 971 -2591 1021 -2553
rect 971 -2625 979 -2591
rect 1013 -2625 1021 -2591
rect 971 -2663 1021 -2625
rect 971 -2697 979 -2663
rect 1013 -2697 1021 -2663
rect 971 -2735 1021 -2697
rect 971 -2769 979 -2735
rect 1013 -2769 1021 -2735
rect 971 -2782 1021 -2769
rect 1137 -2375 1187 -2361
rect 1137 -2409 1145 -2375
rect 1179 -2409 1187 -2375
rect 1137 -2447 1187 -2409
rect 1137 -2481 1145 -2447
rect 1179 -2481 1187 -2447
rect 1137 -2519 1187 -2481
rect 1137 -2553 1145 -2519
rect 1179 -2553 1187 -2519
rect 1137 -2591 1187 -2553
rect 1137 -2625 1145 -2591
rect 1179 -2625 1187 -2591
rect 1137 -2663 1187 -2625
rect 1137 -2697 1145 -2663
rect 1179 -2697 1187 -2663
rect 1137 -2735 1187 -2697
rect 1137 -2769 1145 -2735
rect 1179 -2769 1187 -2735
rect 1137 -2782 1187 -2769
rect 1303 -2375 1353 -2361
rect 1303 -2409 1311 -2375
rect 1345 -2409 1353 -2375
rect 1303 -2447 1353 -2409
rect 1303 -2481 1311 -2447
rect 1345 -2481 1353 -2447
rect 1303 -2519 1353 -2481
rect 1303 -2553 1311 -2519
rect 1345 -2553 1353 -2519
rect 1303 -2591 1353 -2553
rect 1303 -2625 1311 -2591
rect 1345 -2625 1353 -2591
rect 1303 -2663 1353 -2625
rect 1303 -2697 1311 -2663
rect 1345 -2697 1353 -2663
rect 1303 -2735 1353 -2697
rect 1303 -2769 1311 -2735
rect 1345 -2769 1353 -2735
rect 1303 -2782 1353 -2769
rect 1469 -2375 1519 -2361
rect 1469 -2409 1477 -2375
rect 1511 -2409 1519 -2375
rect 1469 -2447 1519 -2409
rect 1469 -2481 1477 -2447
rect 1511 -2481 1519 -2447
rect 1469 -2519 1519 -2481
rect 1469 -2553 1477 -2519
rect 1511 -2553 1519 -2519
rect 1469 -2591 1519 -2553
rect 1469 -2625 1477 -2591
rect 1511 -2625 1519 -2591
rect 1469 -2663 1519 -2625
rect 1469 -2697 1477 -2663
rect 1511 -2697 1519 -2663
rect 1469 -2735 1519 -2697
rect 1469 -2769 1477 -2735
rect 1511 -2769 1519 -2735
rect 1469 -2782 1519 -2769
<< properties >>
string FIXED_BBOX -1642 -2901 1642 2901
<< end >>
