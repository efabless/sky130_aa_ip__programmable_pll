magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< metal3 >>
rect -39164 37092 -33792 37120
rect -39164 37028 -33876 37092
rect -33812 37028 -33792 37092
rect -39164 37012 -33792 37028
rect -39164 36948 -33876 37012
rect -33812 36948 -33792 37012
rect -39164 36932 -33792 36948
rect -39164 36868 -33876 36932
rect -33812 36868 -33792 36932
rect -39164 36852 -33792 36868
rect -39164 36788 -33876 36852
rect -33812 36788 -33792 36852
rect -39164 36772 -33792 36788
rect -39164 36708 -33876 36772
rect -33812 36708 -33792 36772
rect -39164 36692 -33792 36708
rect -39164 36628 -33876 36692
rect -33812 36628 -33792 36692
rect -39164 36612 -33792 36628
rect -39164 36548 -33876 36612
rect -33812 36548 -33792 36612
rect -39164 36532 -33792 36548
rect -39164 36468 -33876 36532
rect -33812 36468 -33792 36532
rect -39164 36452 -33792 36468
rect -39164 36388 -33876 36452
rect -33812 36388 -33792 36452
rect -39164 36372 -33792 36388
rect -39164 36308 -33876 36372
rect -33812 36308 -33792 36372
rect -39164 36292 -33792 36308
rect -39164 36228 -33876 36292
rect -33812 36228 -33792 36292
rect -39164 36212 -33792 36228
rect -39164 36148 -33876 36212
rect -33812 36148 -33792 36212
rect -39164 36132 -33792 36148
rect -39164 36068 -33876 36132
rect -33812 36068 -33792 36132
rect -39164 36052 -33792 36068
rect -39164 35988 -33876 36052
rect -33812 35988 -33792 36052
rect -39164 35972 -33792 35988
rect -39164 35908 -33876 35972
rect -33812 35908 -33792 35972
rect -39164 35892 -33792 35908
rect -39164 35828 -33876 35892
rect -33812 35828 -33792 35892
rect -39164 35812 -33792 35828
rect -39164 35748 -33876 35812
rect -33812 35748 -33792 35812
rect -39164 35732 -33792 35748
rect -39164 35668 -33876 35732
rect -33812 35668 -33792 35732
rect -39164 35652 -33792 35668
rect -39164 35588 -33876 35652
rect -33812 35588 -33792 35652
rect -39164 35572 -33792 35588
rect -39164 35508 -33876 35572
rect -33812 35508 -33792 35572
rect -39164 35492 -33792 35508
rect -39164 35428 -33876 35492
rect -33812 35428 -33792 35492
rect -39164 35412 -33792 35428
rect -39164 35348 -33876 35412
rect -33812 35348 -33792 35412
rect -39164 35332 -33792 35348
rect -39164 35268 -33876 35332
rect -33812 35268 -33792 35332
rect -39164 35252 -33792 35268
rect -39164 35188 -33876 35252
rect -33812 35188 -33792 35252
rect -39164 35172 -33792 35188
rect -39164 35108 -33876 35172
rect -33812 35108 -33792 35172
rect -39164 35092 -33792 35108
rect -39164 35028 -33876 35092
rect -33812 35028 -33792 35092
rect -39164 35012 -33792 35028
rect -39164 34948 -33876 35012
rect -33812 34948 -33792 35012
rect -39164 34932 -33792 34948
rect -39164 34868 -33876 34932
rect -33812 34868 -33792 34932
rect -39164 34852 -33792 34868
rect -39164 34788 -33876 34852
rect -33812 34788 -33792 34852
rect -39164 34772 -33792 34788
rect -39164 34708 -33876 34772
rect -33812 34708 -33792 34772
rect -39164 34692 -33792 34708
rect -39164 34628 -33876 34692
rect -33812 34628 -33792 34692
rect -39164 34612 -33792 34628
rect -39164 34548 -33876 34612
rect -33812 34548 -33792 34612
rect -39164 34532 -33792 34548
rect -39164 34468 -33876 34532
rect -33812 34468 -33792 34532
rect -39164 34452 -33792 34468
rect -39164 34388 -33876 34452
rect -33812 34388 -33792 34452
rect -39164 34372 -33792 34388
rect -39164 34308 -33876 34372
rect -33812 34308 -33792 34372
rect -39164 34292 -33792 34308
rect -39164 34228 -33876 34292
rect -33812 34228 -33792 34292
rect -39164 34212 -33792 34228
rect -39164 34148 -33876 34212
rect -33812 34148 -33792 34212
rect -39164 34132 -33792 34148
rect -39164 34068 -33876 34132
rect -33812 34068 -33792 34132
rect -39164 34052 -33792 34068
rect -39164 33988 -33876 34052
rect -33812 33988 -33792 34052
rect -39164 33972 -33792 33988
rect -39164 33908 -33876 33972
rect -33812 33908 -33792 33972
rect -39164 33892 -33792 33908
rect -39164 33828 -33876 33892
rect -33812 33828 -33792 33892
rect -39164 33812 -33792 33828
rect -39164 33748 -33876 33812
rect -33812 33748 -33792 33812
rect -39164 33732 -33792 33748
rect -39164 33668 -33876 33732
rect -33812 33668 -33792 33732
rect -39164 33652 -33792 33668
rect -39164 33588 -33876 33652
rect -33812 33588 -33792 33652
rect -39164 33572 -33792 33588
rect -39164 33508 -33876 33572
rect -33812 33508 -33792 33572
rect -39164 33492 -33792 33508
rect -39164 33428 -33876 33492
rect -33812 33428 -33792 33492
rect -39164 33412 -33792 33428
rect -39164 33348 -33876 33412
rect -33812 33348 -33792 33412
rect -39164 33332 -33792 33348
rect -39164 33268 -33876 33332
rect -33812 33268 -33792 33332
rect -39164 33252 -33792 33268
rect -39164 33188 -33876 33252
rect -33812 33188 -33792 33252
rect -39164 33172 -33792 33188
rect -39164 33108 -33876 33172
rect -33812 33108 -33792 33172
rect -39164 33092 -33792 33108
rect -39164 33028 -33876 33092
rect -33812 33028 -33792 33092
rect -39164 33012 -33792 33028
rect -39164 32948 -33876 33012
rect -33812 32948 -33792 33012
rect -39164 32932 -33792 32948
rect -39164 32868 -33876 32932
rect -33812 32868 -33792 32932
rect -39164 32852 -33792 32868
rect -39164 32788 -33876 32852
rect -33812 32788 -33792 32852
rect -39164 32772 -33792 32788
rect -39164 32708 -33876 32772
rect -33812 32708 -33792 32772
rect -39164 32692 -33792 32708
rect -39164 32628 -33876 32692
rect -33812 32628 -33792 32692
rect -39164 32612 -33792 32628
rect -39164 32548 -33876 32612
rect -33812 32548 -33792 32612
rect -39164 32532 -33792 32548
rect -39164 32468 -33876 32532
rect -33812 32468 -33792 32532
rect -39164 32452 -33792 32468
rect -39164 32388 -33876 32452
rect -33812 32388 -33792 32452
rect -39164 32372 -33792 32388
rect -39164 32308 -33876 32372
rect -33812 32308 -33792 32372
rect -39164 32292 -33792 32308
rect -39164 32228 -33876 32292
rect -33812 32228 -33792 32292
rect -39164 32212 -33792 32228
rect -39164 32148 -33876 32212
rect -33812 32148 -33792 32212
rect -39164 32132 -33792 32148
rect -39164 32068 -33876 32132
rect -33812 32068 -33792 32132
rect -39164 32040 -33792 32068
rect -33552 37092 -28180 37120
rect -33552 37028 -28264 37092
rect -28200 37028 -28180 37092
rect -33552 37012 -28180 37028
rect -33552 36948 -28264 37012
rect -28200 36948 -28180 37012
rect -33552 36932 -28180 36948
rect -33552 36868 -28264 36932
rect -28200 36868 -28180 36932
rect -33552 36852 -28180 36868
rect -33552 36788 -28264 36852
rect -28200 36788 -28180 36852
rect -33552 36772 -28180 36788
rect -33552 36708 -28264 36772
rect -28200 36708 -28180 36772
rect -33552 36692 -28180 36708
rect -33552 36628 -28264 36692
rect -28200 36628 -28180 36692
rect -33552 36612 -28180 36628
rect -33552 36548 -28264 36612
rect -28200 36548 -28180 36612
rect -33552 36532 -28180 36548
rect -33552 36468 -28264 36532
rect -28200 36468 -28180 36532
rect -33552 36452 -28180 36468
rect -33552 36388 -28264 36452
rect -28200 36388 -28180 36452
rect -33552 36372 -28180 36388
rect -33552 36308 -28264 36372
rect -28200 36308 -28180 36372
rect -33552 36292 -28180 36308
rect -33552 36228 -28264 36292
rect -28200 36228 -28180 36292
rect -33552 36212 -28180 36228
rect -33552 36148 -28264 36212
rect -28200 36148 -28180 36212
rect -33552 36132 -28180 36148
rect -33552 36068 -28264 36132
rect -28200 36068 -28180 36132
rect -33552 36052 -28180 36068
rect -33552 35988 -28264 36052
rect -28200 35988 -28180 36052
rect -33552 35972 -28180 35988
rect -33552 35908 -28264 35972
rect -28200 35908 -28180 35972
rect -33552 35892 -28180 35908
rect -33552 35828 -28264 35892
rect -28200 35828 -28180 35892
rect -33552 35812 -28180 35828
rect -33552 35748 -28264 35812
rect -28200 35748 -28180 35812
rect -33552 35732 -28180 35748
rect -33552 35668 -28264 35732
rect -28200 35668 -28180 35732
rect -33552 35652 -28180 35668
rect -33552 35588 -28264 35652
rect -28200 35588 -28180 35652
rect -33552 35572 -28180 35588
rect -33552 35508 -28264 35572
rect -28200 35508 -28180 35572
rect -33552 35492 -28180 35508
rect -33552 35428 -28264 35492
rect -28200 35428 -28180 35492
rect -33552 35412 -28180 35428
rect -33552 35348 -28264 35412
rect -28200 35348 -28180 35412
rect -33552 35332 -28180 35348
rect -33552 35268 -28264 35332
rect -28200 35268 -28180 35332
rect -33552 35252 -28180 35268
rect -33552 35188 -28264 35252
rect -28200 35188 -28180 35252
rect -33552 35172 -28180 35188
rect -33552 35108 -28264 35172
rect -28200 35108 -28180 35172
rect -33552 35092 -28180 35108
rect -33552 35028 -28264 35092
rect -28200 35028 -28180 35092
rect -33552 35012 -28180 35028
rect -33552 34948 -28264 35012
rect -28200 34948 -28180 35012
rect -33552 34932 -28180 34948
rect -33552 34868 -28264 34932
rect -28200 34868 -28180 34932
rect -33552 34852 -28180 34868
rect -33552 34788 -28264 34852
rect -28200 34788 -28180 34852
rect -33552 34772 -28180 34788
rect -33552 34708 -28264 34772
rect -28200 34708 -28180 34772
rect -33552 34692 -28180 34708
rect -33552 34628 -28264 34692
rect -28200 34628 -28180 34692
rect -33552 34612 -28180 34628
rect -33552 34548 -28264 34612
rect -28200 34548 -28180 34612
rect -33552 34532 -28180 34548
rect -33552 34468 -28264 34532
rect -28200 34468 -28180 34532
rect -33552 34452 -28180 34468
rect -33552 34388 -28264 34452
rect -28200 34388 -28180 34452
rect -33552 34372 -28180 34388
rect -33552 34308 -28264 34372
rect -28200 34308 -28180 34372
rect -33552 34292 -28180 34308
rect -33552 34228 -28264 34292
rect -28200 34228 -28180 34292
rect -33552 34212 -28180 34228
rect -33552 34148 -28264 34212
rect -28200 34148 -28180 34212
rect -33552 34132 -28180 34148
rect -33552 34068 -28264 34132
rect -28200 34068 -28180 34132
rect -33552 34052 -28180 34068
rect -33552 33988 -28264 34052
rect -28200 33988 -28180 34052
rect -33552 33972 -28180 33988
rect -33552 33908 -28264 33972
rect -28200 33908 -28180 33972
rect -33552 33892 -28180 33908
rect -33552 33828 -28264 33892
rect -28200 33828 -28180 33892
rect -33552 33812 -28180 33828
rect -33552 33748 -28264 33812
rect -28200 33748 -28180 33812
rect -33552 33732 -28180 33748
rect -33552 33668 -28264 33732
rect -28200 33668 -28180 33732
rect -33552 33652 -28180 33668
rect -33552 33588 -28264 33652
rect -28200 33588 -28180 33652
rect -33552 33572 -28180 33588
rect -33552 33508 -28264 33572
rect -28200 33508 -28180 33572
rect -33552 33492 -28180 33508
rect -33552 33428 -28264 33492
rect -28200 33428 -28180 33492
rect -33552 33412 -28180 33428
rect -33552 33348 -28264 33412
rect -28200 33348 -28180 33412
rect -33552 33332 -28180 33348
rect -33552 33268 -28264 33332
rect -28200 33268 -28180 33332
rect -33552 33252 -28180 33268
rect -33552 33188 -28264 33252
rect -28200 33188 -28180 33252
rect -33552 33172 -28180 33188
rect -33552 33108 -28264 33172
rect -28200 33108 -28180 33172
rect -33552 33092 -28180 33108
rect -33552 33028 -28264 33092
rect -28200 33028 -28180 33092
rect -33552 33012 -28180 33028
rect -33552 32948 -28264 33012
rect -28200 32948 -28180 33012
rect -33552 32932 -28180 32948
rect -33552 32868 -28264 32932
rect -28200 32868 -28180 32932
rect -33552 32852 -28180 32868
rect -33552 32788 -28264 32852
rect -28200 32788 -28180 32852
rect -33552 32772 -28180 32788
rect -33552 32708 -28264 32772
rect -28200 32708 -28180 32772
rect -33552 32692 -28180 32708
rect -33552 32628 -28264 32692
rect -28200 32628 -28180 32692
rect -33552 32612 -28180 32628
rect -33552 32548 -28264 32612
rect -28200 32548 -28180 32612
rect -33552 32532 -28180 32548
rect -33552 32468 -28264 32532
rect -28200 32468 -28180 32532
rect -33552 32452 -28180 32468
rect -33552 32388 -28264 32452
rect -28200 32388 -28180 32452
rect -33552 32372 -28180 32388
rect -33552 32308 -28264 32372
rect -28200 32308 -28180 32372
rect -33552 32292 -28180 32308
rect -33552 32228 -28264 32292
rect -28200 32228 -28180 32292
rect -33552 32212 -28180 32228
rect -33552 32148 -28264 32212
rect -28200 32148 -28180 32212
rect -33552 32132 -28180 32148
rect -33552 32068 -28264 32132
rect -28200 32068 -28180 32132
rect -33552 32040 -28180 32068
rect -27940 37092 -22568 37120
rect -27940 37028 -22652 37092
rect -22588 37028 -22568 37092
rect -27940 37012 -22568 37028
rect -27940 36948 -22652 37012
rect -22588 36948 -22568 37012
rect -27940 36932 -22568 36948
rect -27940 36868 -22652 36932
rect -22588 36868 -22568 36932
rect -27940 36852 -22568 36868
rect -27940 36788 -22652 36852
rect -22588 36788 -22568 36852
rect -27940 36772 -22568 36788
rect -27940 36708 -22652 36772
rect -22588 36708 -22568 36772
rect -27940 36692 -22568 36708
rect -27940 36628 -22652 36692
rect -22588 36628 -22568 36692
rect -27940 36612 -22568 36628
rect -27940 36548 -22652 36612
rect -22588 36548 -22568 36612
rect -27940 36532 -22568 36548
rect -27940 36468 -22652 36532
rect -22588 36468 -22568 36532
rect -27940 36452 -22568 36468
rect -27940 36388 -22652 36452
rect -22588 36388 -22568 36452
rect -27940 36372 -22568 36388
rect -27940 36308 -22652 36372
rect -22588 36308 -22568 36372
rect -27940 36292 -22568 36308
rect -27940 36228 -22652 36292
rect -22588 36228 -22568 36292
rect -27940 36212 -22568 36228
rect -27940 36148 -22652 36212
rect -22588 36148 -22568 36212
rect -27940 36132 -22568 36148
rect -27940 36068 -22652 36132
rect -22588 36068 -22568 36132
rect -27940 36052 -22568 36068
rect -27940 35988 -22652 36052
rect -22588 35988 -22568 36052
rect -27940 35972 -22568 35988
rect -27940 35908 -22652 35972
rect -22588 35908 -22568 35972
rect -27940 35892 -22568 35908
rect -27940 35828 -22652 35892
rect -22588 35828 -22568 35892
rect -27940 35812 -22568 35828
rect -27940 35748 -22652 35812
rect -22588 35748 -22568 35812
rect -27940 35732 -22568 35748
rect -27940 35668 -22652 35732
rect -22588 35668 -22568 35732
rect -27940 35652 -22568 35668
rect -27940 35588 -22652 35652
rect -22588 35588 -22568 35652
rect -27940 35572 -22568 35588
rect -27940 35508 -22652 35572
rect -22588 35508 -22568 35572
rect -27940 35492 -22568 35508
rect -27940 35428 -22652 35492
rect -22588 35428 -22568 35492
rect -27940 35412 -22568 35428
rect -27940 35348 -22652 35412
rect -22588 35348 -22568 35412
rect -27940 35332 -22568 35348
rect -27940 35268 -22652 35332
rect -22588 35268 -22568 35332
rect -27940 35252 -22568 35268
rect -27940 35188 -22652 35252
rect -22588 35188 -22568 35252
rect -27940 35172 -22568 35188
rect -27940 35108 -22652 35172
rect -22588 35108 -22568 35172
rect -27940 35092 -22568 35108
rect -27940 35028 -22652 35092
rect -22588 35028 -22568 35092
rect -27940 35012 -22568 35028
rect -27940 34948 -22652 35012
rect -22588 34948 -22568 35012
rect -27940 34932 -22568 34948
rect -27940 34868 -22652 34932
rect -22588 34868 -22568 34932
rect -27940 34852 -22568 34868
rect -27940 34788 -22652 34852
rect -22588 34788 -22568 34852
rect -27940 34772 -22568 34788
rect -27940 34708 -22652 34772
rect -22588 34708 -22568 34772
rect -27940 34692 -22568 34708
rect -27940 34628 -22652 34692
rect -22588 34628 -22568 34692
rect -27940 34612 -22568 34628
rect -27940 34548 -22652 34612
rect -22588 34548 -22568 34612
rect -27940 34532 -22568 34548
rect -27940 34468 -22652 34532
rect -22588 34468 -22568 34532
rect -27940 34452 -22568 34468
rect -27940 34388 -22652 34452
rect -22588 34388 -22568 34452
rect -27940 34372 -22568 34388
rect -27940 34308 -22652 34372
rect -22588 34308 -22568 34372
rect -27940 34292 -22568 34308
rect -27940 34228 -22652 34292
rect -22588 34228 -22568 34292
rect -27940 34212 -22568 34228
rect -27940 34148 -22652 34212
rect -22588 34148 -22568 34212
rect -27940 34132 -22568 34148
rect -27940 34068 -22652 34132
rect -22588 34068 -22568 34132
rect -27940 34052 -22568 34068
rect -27940 33988 -22652 34052
rect -22588 33988 -22568 34052
rect -27940 33972 -22568 33988
rect -27940 33908 -22652 33972
rect -22588 33908 -22568 33972
rect -27940 33892 -22568 33908
rect -27940 33828 -22652 33892
rect -22588 33828 -22568 33892
rect -27940 33812 -22568 33828
rect -27940 33748 -22652 33812
rect -22588 33748 -22568 33812
rect -27940 33732 -22568 33748
rect -27940 33668 -22652 33732
rect -22588 33668 -22568 33732
rect -27940 33652 -22568 33668
rect -27940 33588 -22652 33652
rect -22588 33588 -22568 33652
rect -27940 33572 -22568 33588
rect -27940 33508 -22652 33572
rect -22588 33508 -22568 33572
rect -27940 33492 -22568 33508
rect -27940 33428 -22652 33492
rect -22588 33428 -22568 33492
rect -27940 33412 -22568 33428
rect -27940 33348 -22652 33412
rect -22588 33348 -22568 33412
rect -27940 33332 -22568 33348
rect -27940 33268 -22652 33332
rect -22588 33268 -22568 33332
rect -27940 33252 -22568 33268
rect -27940 33188 -22652 33252
rect -22588 33188 -22568 33252
rect -27940 33172 -22568 33188
rect -27940 33108 -22652 33172
rect -22588 33108 -22568 33172
rect -27940 33092 -22568 33108
rect -27940 33028 -22652 33092
rect -22588 33028 -22568 33092
rect -27940 33012 -22568 33028
rect -27940 32948 -22652 33012
rect -22588 32948 -22568 33012
rect -27940 32932 -22568 32948
rect -27940 32868 -22652 32932
rect -22588 32868 -22568 32932
rect -27940 32852 -22568 32868
rect -27940 32788 -22652 32852
rect -22588 32788 -22568 32852
rect -27940 32772 -22568 32788
rect -27940 32708 -22652 32772
rect -22588 32708 -22568 32772
rect -27940 32692 -22568 32708
rect -27940 32628 -22652 32692
rect -22588 32628 -22568 32692
rect -27940 32612 -22568 32628
rect -27940 32548 -22652 32612
rect -22588 32548 -22568 32612
rect -27940 32532 -22568 32548
rect -27940 32468 -22652 32532
rect -22588 32468 -22568 32532
rect -27940 32452 -22568 32468
rect -27940 32388 -22652 32452
rect -22588 32388 -22568 32452
rect -27940 32372 -22568 32388
rect -27940 32308 -22652 32372
rect -22588 32308 -22568 32372
rect -27940 32292 -22568 32308
rect -27940 32228 -22652 32292
rect -22588 32228 -22568 32292
rect -27940 32212 -22568 32228
rect -27940 32148 -22652 32212
rect -22588 32148 -22568 32212
rect -27940 32132 -22568 32148
rect -27940 32068 -22652 32132
rect -22588 32068 -22568 32132
rect -27940 32040 -22568 32068
rect -22328 37092 -16956 37120
rect -22328 37028 -17040 37092
rect -16976 37028 -16956 37092
rect -22328 37012 -16956 37028
rect -22328 36948 -17040 37012
rect -16976 36948 -16956 37012
rect -22328 36932 -16956 36948
rect -22328 36868 -17040 36932
rect -16976 36868 -16956 36932
rect -22328 36852 -16956 36868
rect -22328 36788 -17040 36852
rect -16976 36788 -16956 36852
rect -22328 36772 -16956 36788
rect -22328 36708 -17040 36772
rect -16976 36708 -16956 36772
rect -22328 36692 -16956 36708
rect -22328 36628 -17040 36692
rect -16976 36628 -16956 36692
rect -22328 36612 -16956 36628
rect -22328 36548 -17040 36612
rect -16976 36548 -16956 36612
rect -22328 36532 -16956 36548
rect -22328 36468 -17040 36532
rect -16976 36468 -16956 36532
rect -22328 36452 -16956 36468
rect -22328 36388 -17040 36452
rect -16976 36388 -16956 36452
rect -22328 36372 -16956 36388
rect -22328 36308 -17040 36372
rect -16976 36308 -16956 36372
rect -22328 36292 -16956 36308
rect -22328 36228 -17040 36292
rect -16976 36228 -16956 36292
rect -22328 36212 -16956 36228
rect -22328 36148 -17040 36212
rect -16976 36148 -16956 36212
rect -22328 36132 -16956 36148
rect -22328 36068 -17040 36132
rect -16976 36068 -16956 36132
rect -22328 36052 -16956 36068
rect -22328 35988 -17040 36052
rect -16976 35988 -16956 36052
rect -22328 35972 -16956 35988
rect -22328 35908 -17040 35972
rect -16976 35908 -16956 35972
rect -22328 35892 -16956 35908
rect -22328 35828 -17040 35892
rect -16976 35828 -16956 35892
rect -22328 35812 -16956 35828
rect -22328 35748 -17040 35812
rect -16976 35748 -16956 35812
rect -22328 35732 -16956 35748
rect -22328 35668 -17040 35732
rect -16976 35668 -16956 35732
rect -22328 35652 -16956 35668
rect -22328 35588 -17040 35652
rect -16976 35588 -16956 35652
rect -22328 35572 -16956 35588
rect -22328 35508 -17040 35572
rect -16976 35508 -16956 35572
rect -22328 35492 -16956 35508
rect -22328 35428 -17040 35492
rect -16976 35428 -16956 35492
rect -22328 35412 -16956 35428
rect -22328 35348 -17040 35412
rect -16976 35348 -16956 35412
rect -22328 35332 -16956 35348
rect -22328 35268 -17040 35332
rect -16976 35268 -16956 35332
rect -22328 35252 -16956 35268
rect -22328 35188 -17040 35252
rect -16976 35188 -16956 35252
rect -22328 35172 -16956 35188
rect -22328 35108 -17040 35172
rect -16976 35108 -16956 35172
rect -22328 35092 -16956 35108
rect -22328 35028 -17040 35092
rect -16976 35028 -16956 35092
rect -22328 35012 -16956 35028
rect -22328 34948 -17040 35012
rect -16976 34948 -16956 35012
rect -22328 34932 -16956 34948
rect -22328 34868 -17040 34932
rect -16976 34868 -16956 34932
rect -22328 34852 -16956 34868
rect -22328 34788 -17040 34852
rect -16976 34788 -16956 34852
rect -22328 34772 -16956 34788
rect -22328 34708 -17040 34772
rect -16976 34708 -16956 34772
rect -22328 34692 -16956 34708
rect -22328 34628 -17040 34692
rect -16976 34628 -16956 34692
rect -22328 34612 -16956 34628
rect -22328 34548 -17040 34612
rect -16976 34548 -16956 34612
rect -22328 34532 -16956 34548
rect -22328 34468 -17040 34532
rect -16976 34468 -16956 34532
rect -22328 34452 -16956 34468
rect -22328 34388 -17040 34452
rect -16976 34388 -16956 34452
rect -22328 34372 -16956 34388
rect -22328 34308 -17040 34372
rect -16976 34308 -16956 34372
rect -22328 34292 -16956 34308
rect -22328 34228 -17040 34292
rect -16976 34228 -16956 34292
rect -22328 34212 -16956 34228
rect -22328 34148 -17040 34212
rect -16976 34148 -16956 34212
rect -22328 34132 -16956 34148
rect -22328 34068 -17040 34132
rect -16976 34068 -16956 34132
rect -22328 34052 -16956 34068
rect -22328 33988 -17040 34052
rect -16976 33988 -16956 34052
rect -22328 33972 -16956 33988
rect -22328 33908 -17040 33972
rect -16976 33908 -16956 33972
rect -22328 33892 -16956 33908
rect -22328 33828 -17040 33892
rect -16976 33828 -16956 33892
rect -22328 33812 -16956 33828
rect -22328 33748 -17040 33812
rect -16976 33748 -16956 33812
rect -22328 33732 -16956 33748
rect -22328 33668 -17040 33732
rect -16976 33668 -16956 33732
rect -22328 33652 -16956 33668
rect -22328 33588 -17040 33652
rect -16976 33588 -16956 33652
rect -22328 33572 -16956 33588
rect -22328 33508 -17040 33572
rect -16976 33508 -16956 33572
rect -22328 33492 -16956 33508
rect -22328 33428 -17040 33492
rect -16976 33428 -16956 33492
rect -22328 33412 -16956 33428
rect -22328 33348 -17040 33412
rect -16976 33348 -16956 33412
rect -22328 33332 -16956 33348
rect -22328 33268 -17040 33332
rect -16976 33268 -16956 33332
rect -22328 33252 -16956 33268
rect -22328 33188 -17040 33252
rect -16976 33188 -16956 33252
rect -22328 33172 -16956 33188
rect -22328 33108 -17040 33172
rect -16976 33108 -16956 33172
rect -22328 33092 -16956 33108
rect -22328 33028 -17040 33092
rect -16976 33028 -16956 33092
rect -22328 33012 -16956 33028
rect -22328 32948 -17040 33012
rect -16976 32948 -16956 33012
rect -22328 32932 -16956 32948
rect -22328 32868 -17040 32932
rect -16976 32868 -16956 32932
rect -22328 32852 -16956 32868
rect -22328 32788 -17040 32852
rect -16976 32788 -16956 32852
rect -22328 32772 -16956 32788
rect -22328 32708 -17040 32772
rect -16976 32708 -16956 32772
rect -22328 32692 -16956 32708
rect -22328 32628 -17040 32692
rect -16976 32628 -16956 32692
rect -22328 32612 -16956 32628
rect -22328 32548 -17040 32612
rect -16976 32548 -16956 32612
rect -22328 32532 -16956 32548
rect -22328 32468 -17040 32532
rect -16976 32468 -16956 32532
rect -22328 32452 -16956 32468
rect -22328 32388 -17040 32452
rect -16976 32388 -16956 32452
rect -22328 32372 -16956 32388
rect -22328 32308 -17040 32372
rect -16976 32308 -16956 32372
rect -22328 32292 -16956 32308
rect -22328 32228 -17040 32292
rect -16976 32228 -16956 32292
rect -22328 32212 -16956 32228
rect -22328 32148 -17040 32212
rect -16976 32148 -16956 32212
rect -22328 32132 -16956 32148
rect -22328 32068 -17040 32132
rect -16976 32068 -16956 32132
rect -22328 32040 -16956 32068
rect -16716 37092 -11344 37120
rect -16716 37028 -11428 37092
rect -11364 37028 -11344 37092
rect -16716 37012 -11344 37028
rect -16716 36948 -11428 37012
rect -11364 36948 -11344 37012
rect -16716 36932 -11344 36948
rect -16716 36868 -11428 36932
rect -11364 36868 -11344 36932
rect -16716 36852 -11344 36868
rect -16716 36788 -11428 36852
rect -11364 36788 -11344 36852
rect -16716 36772 -11344 36788
rect -16716 36708 -11428 36772
rect -11364 36708 -11344 36772
rect -16716 36692 -11344 36708
rect -16716 36628 -11428 36692
rect -11364 36628 -11344 36692
rect -16716 36612 -11344 36628
rect -16716 36548 -11428 36612
rect -11364 36548 -11344 36612
rect -16716 36532 -11344 36548
rect -16716 36468 -11428 36532
rect -11364 36468 -11344 36532
rect -16716 36452 -11344 36468
rect -16716 36388 -11428 36452
rect -11364 36388 -11344 36452
rect -16716 36372 -11344 36388
rect -16716 36308 -11428 36372
rect -11364 36308 -11344 36372
rect -16716 36292 -11344 36308
rect -16716 36228 -11428 36292
rect -11364 36228 -11344 36292
rect -16716 36212 -11344 36228
rect -16716 36148 -11428 36212
rect -11364 36148 -11344 36212
rect -16716 36132 -11344 36148
rect -16716 36068 -11428 36132
rect -11364 36068 -11344 36132
rect -16716 36052 -11344 36068
rect -16716 35988 -11428 36052
rect -11364 35988 -11344 36052
rect -16716 35972 -11344 35988
rect -16716 35908 -11428 35972
rect -11364 35908 -11344 35972
rect -16716 35892 -11344 35908
rect -16716 35828 -11428 35892
rect -11364 35828 -11344 35892
rect -16716 35812 -11344 35828
rect -16716 35748 -11428 35812
rect -11364 35748 -11344 35812
rect -16716 35732 -11344 35748
rect -16716 35668 -11428 35732
rect -11364 35668 -11344 35732
rect -16716 35652 -11344 35668
rect -16716 35588 -11428 35652
rect -11364 35588 -11344 35652
rect -16716 35572 -11344 35588
rect -16716 35508 -11428 35572
rect -11364 35508 -11344 35572
rect -16716 35492 -11344 35508
rect -16716 35428 -11428 35492
rect -11364 35428 -11344 35492
rect -16716 35412 -11344 35428
rect -16716 35348 -11428 35412
rect -11364 35348 -11344 35412
rect -16716 35332 -11344 35348
rect -16716 35268 -11428 35332
rect -11364 35268 -11344 35332
rect -16716 35252 -11344 35268
rect -16716 35188 -11428 35252
rect -11364 35188 -11344 35252
rect -16716 35172 -11344 35188
rect -16716 35108 -11428 35172
rect -11364 35108 -11344 35172
rect -16716 35092 -11344 35108
rect -16716 35028 -11428 35092
rect -11364 35028 -11344 35092
rect -16716 35012 -11344 35028
rect -16716 34948 -11428 35012
rect -11364 34948 -11344 35012
rect -16716 34932 -11344 34948
rect -16716 34868 -11428 34932
rect -11364 34868 -11344 34932
rect -16716 34852 -11344 34868
rect -16716 34788 -11428 34852
rect -11364 34788 -11344 34852
rect -16716 34772 -11344 34788
rect -16716 34708 -11428 34772
rect -11364 34708 -11344 34772
rect -16716 34692 -11344 34708
rect -16716 34628 -11428 34692
rect -11364 34628 -11344 34692
rect -16716 34612 -11344 34628
rect -16716 34548 -11428 34612
rect -11364 34548 -11344 34612
rect -16716 34532 -11344 34548
rect -16716 34468 -11428 34532
rect -11364 34468 -11344 34532
rect -16716 34452 -11344 34468
rect -16716 34388 -11428 34452
rect -11364 34388 -11344 34452
rect -16716 34372 -11344 34388
rect -16716 34308 -11428 34372
rect -11364 34308 -11344 34372
rect -16716 34292 -11344 34308
rect -16716 34228 -11428 34292
rect -11364 34228 -11344 34292
rect -16716 34212 -11344 34228
rect -16716 34148 -11428 34212
rect -11364 34148 -11344 34212
rect -16716 34132 -11344 34148
rect -16716 34068 -11428 34132
rect -11364 34068 -11344 34132
rect -16716 34052 -11344 34068
rect -16716 33988 -11428 34052
rect -11364 33988 -11344 34052
rect -16716 33972 -11344 33988
rect -16716 33908 -11428 33972
rect -11364 33908 -11344 33972
rect -16716 33892 -11344 33908
rect -16716 33828 -11428 33892
rect -11364 33828 -11344 33892
rect -16716 33812 -11344 33828
rect -16716 33748 -11428 33812
rect -11364 33748 -11344 33812
rect -16716 33732 -11344 33748
rect -16716 33668 -11428 33732
rect -11364 33668 -11344 33732
rect -16716 33652 -11344 33668
rect -16716 33588 -11428 33652
rect -11364 33588 -11344 33652
rect -16716 33572 -11344 33588
rect -16716 33508 -11428 33572
rect -11364 33508 -11344 33572
rect -16716 33492 -11344 33508
rect -16716 33428 -11428 33492
rect -11364 33428 -11344 33492
rect -16716 33412 -11344 33428
rect -16716 33348 -11428 33412
rect -11364 33348 -11344 33412
rect -16716 33332 -11344 33348
rect -16716 33268 -11428 33332
rect -11364 33268 -11344 33332
rect -16716 33252 -11344 33268
rect -16716 33188 -11428 33252
rect -11364 33188 -11344 33252
rect -16716 33172 -11344 33188
rect -16716 33108 -11428 33172
rect -11364 33108 -11344 33172
rect -16716 33092 -11344 33108
rect -16716 33028 -11428 33092
rect -11364 33028 -11344 33092
rect -16716 33012 -11344 33028
rect -16716 32948 -11428 33012
rect -11364 32948 -11344 33012
rect -16716 32932 -11344 32948
rect -16716 32868 -11428 32932
rect -11364 32868 -11344 32932
rect -16716 32852 -11344 32868
rect -16716 32788 -11428 32852
rect -11364 32788 -11344 32852
rect -16716 32772 -11344 32788
rect -16716 32708 -11428 32772
rect -11364 32708 -11344 32772
rect -16716 32692 -11344 32708
rect -16716 32628 -11428 32692
rect -11364 32628 -11344 32692
rect -16716 32612 -11344 32628
rect -16716 32548 -11428 32612
rect -11364 32548 -11344 32612
rect -16716 32532 -11344 32548
rect -16716 32468 -11428 32532
rect -11364 32468 -11344 32532
rect -16716 32452 -11344 32468
rect -16716 32388 -11428 32452
rect -11364 32388 -11344 32452
rect -16716 32372 -11344 32388
rect -16716 32308 -11428 32372
rect -11364 32308 -11344 32372
rect -16716 32292 -11344 32308
rect -16716 32228 -11428 32292
rect -11364 32228 -11344 32292
rect -16716 32212 -11344 32228
rect -16716 32148 -11428 32212
rect -11364 32148 -11344 32212
rect -16716 32132 -11344 32148
rect -16716 32068 -11428 32132
rect -11364 32068 -11344 32132
rect -16716 32040 -11344 32068
rect -11104 37092 -5732 37120
rect -11104 37028 -5816 37092
rect -5752 37028 -5732 37092
rect -11104 37012 -5732 37028
rect -11104 36948 -5816 37012
rect -5752 36948 -5732 37012
rect -11104 36932 -5732 36948
rect -11104 36868 -5816 36932
rect -5752 36868 -5732 36932
rect -11104 36852 -5732 36868
rect -11104 36788 -5816 36852
rect -5752 36788 -5732 36852
rect -11104 36772 -5732 36788
rect -11104 36708 -5816 36772
rect -5752 36708 -5732 36772
rect -11104 36692 -5732 36708
rect -11104 36628 -5816 36692
rect -5752 36628 -5732 36692
rect -11104 36612 -5732 36628
rect -11104 36548 -5816 36612
rect -5752 36548 -5732 36612
rect -11104 36532 -5732 36548
rect -11104 36468 -5816 36532
rect -5752 36468 -5732 36532
rect -11104 36452 -5732 36468
rect -11104 36388 -5816 36452
rect -5752 36388 -5732 36452
rect -11104 36372 -5732 36388
rect -11104 36308 -5816 36372
rect -5752 36308 -5732 36372
rect -11104 36292 -5732 36308
rect -11104 36228 -5816 36292
rect -5752 36228 -5732 36292
rect -11104 36212 -5732 36228
rect -11104 36148 -5816 36212
rect -5752 36148 -5732 36212
rect -11104 36132 -5732 36148
rect -11104 36068 -5816 36132
rect -5752 36068 -5732 36132
rect -11104 36052 -5732 36068
rect -11104 35988 -5816 36052
rect -5752 35988 -5732 36052
rect -11104 35972 -5732 35988
rect -11104 35908 -5816 35972
rect -5752 35908 -5732 35972
rect -11104 35892 -5732 35908
rect -11104 35828 -5816 35892
rect -5752 35828 -5732 35892
rect -11104 35812 -5732 35828
rect -11104 35748 -5816 35812
rect -5752 35748 -5732 35812
rect -11104 35732 -5732 35748
rect -11104 35668 -5816 35732
rect -5752 35668 -5732 35732
rect -11104 35652 -5732 35668
rect -11104 35588 -5816 35652
rect -5752 35588 -5732 35652
rect -11104 35572 -5732 35588
rect -11104 35508 -5816 35572
rect -5752 35508 -5732 35572
rect -11104 35492 -5732 35508
rect -11104 35428 -5816 35492
rect -5752 35428 -5732 35492
rect -11104 35412 -5732 35428
rect -11104 35348 -5816 35412
rect -5752 35348 -5732 35412
rect -11104 35332 -5732 35348
rect -11104 35268 -5816 35332
rect -5752 35268 -5732 35332
rect -11104 35252 -5732 35268
rect -11104 35188 -5816 35252
rect -5752 35188 -5732 35252
rect -11104 35172 -5732 35188
rect -11104 35108 -5816 35172
rect -5752 35108 -5732 35172
rect -11104 35092 -5732 35108
rect -11104 35028 -5816 35092
rect -5752 35028 -5732 35092
rect -11104 35012 -5732 35028
rect -11104 34948 -5816 35012
rect -5752 34948 -5732 35012
rect -11104 34932 -5732 34948
rect -11104 34868 -5816 34932
rect -5752 34868 -5732 34932
rect -11104 34852 -5732 34868
rect -11104 34788 -5816 34852
rect -5752 34788 -5732 34852
rect -11104 34772 -5732 34788
rect -11104 34708 -5816 34772
rect -5752 34708 -5732 34772
rect -11104 34692 -5732 34708
rect -11104 34628 -5816 34692
rect -5752 34628 -5732 34692
rect -11104 34612 -5732 34628
rect -11104 34548 -5816 34612
rect -5752 34548 -5732 34612
rect -11104 34532 -5732 34548
rect -11104 34468 -5816 34532
rect -5752 34468 -5732 34532
rect -11104 34452 -5732 34468
rect -11104 34388 -5816 34452
rect -5752 34388 -5732 34452
rect -11104 34372 -5732 34388
rect -11104 34308 -5816 34372
rect -5752 34308 -5732 34372
rect -11104 34292 -5732 34308
rect -11104 34228 -5816 34292
rect -5752 34228 -5732 34292
rect -11104 34212 -5732 34228
rect -11104 34148 -5816 34212
rect -5752 34148 -5732 34212
rect -11104 34132 -5732 34148
rect -11104 34068 -5816 34132
rect -5752 34068 -5732 34132
rect -11104 34052 -5732 34068
rect -11104 33988 -5816 34052
rect -5752 33988 -5732 34052
rect -11104 33972 -5732 33988
rect -11104 33908 -5816 33972
rect -5752 33908 -5732 33972
rect -11104 33892 -5732 33908
rect -11104 33828 -5816 33892
rect -5752 33828 -5732 33892
rect -11104 33812 -5732 33828
rect -11104 33748 -5816 33812
rect -5752 33748 -5732 33812
rect -11104 33732 -5732 33748
rect -11104 33668 -5816 33732
rect -5752 33668 -5732 33732
rect -11104 33652 -5732 33668
rect -11104 33588 -5816 33652
rect -5752 33588 -5732 33652
rect -11104 33572 -5732 33588
rect -11104 33508 -5816 33572
rect -5752 33508 -5732 33572
rect -11104 33492 -5732 33508
rect -11104 33428 -5816 33492
rect -5752 33428 -5732 33492
rect -11104 33412 -5732 33428
rect -11104 33348 -5816 33412
rect -5752 33348 -5732 33412
rect -11104 33332 -5732 33348
rect -11104 33268 -5816 33332
rect -5752 33268 -5732 33332
rect -11104 33252 -5732 33268
rect -11104 33188 -5816 33252
rect -5752 33188 -5732 33252
rect -11104 33172 -5732 33188
rect -11104 33108 -5816 33172
rect -5752 33108 -5732 33172
rect -11104 33092 -5732 33108
rect -11104 33028 -5816 33092
rect -5752 33028 -5732 33092
rect -11104 33012 -5732 33028
rect -11104 32948 -5816 33012
rect -5752 32948 -5732 33012
rect -11104 32932 -5732 32948
rect -11104 32868 -5816 32932
rect -5752 32868 -5732 32932
rect -11104 32852 -5732 32868
rect -11104 32788 -5816 32852
rect -5752 32788 -5732 32852
rect -11104 32772 -5732 32788
rect -11104 32708 -5816 32772
rect -5752 32708 -5732 32772
rect -11104 32692 -5732 32708
rect -11104 32628 -5816 32692
rect -5752 32628 -5732 32692
rect -11104 32612 -5732 32628
rect -11104 32548 -5816 32612
rect -5752 32548 -5732 32612
rect -11104 32532 -5732 32548
rect -11104 32468 -5816 32532
rect -5752 32468 -5732 32532
rect -11104 32452 -5732 32468
rect -11104 32388 -5816 32452
rect -5752 32388 -5732 32452
rect -11104 32372 -5732 32388
rect -11104 32308 -5816 32372
rect -5752 32308 -5732 32372
rect -11104 32292 -5732 32308
rect -11104 32228 -5816 32292
rect -5752 32228 -5732 32292
rect -11104 32212 -5732 32228
rect -11104 32148 -5816 32212
rect -5752 32148 -5732 32212
rect -11104 32132 -5732 32148
rect -11104 32068 -5816 32132
rect -5752 32068 -5732 32132
rect -11104 32040 -5732 32068
rect -5492 37092 -120 37120
rect -5492 37028 -204 37092
rect -140 37028 -120 37092
rect -5492 37012 -120 37028
rect -5492 36948 -204 37012
rect -140 36948 -120 37012
rect -5492 36932 -120 36948
rect -5492 36868 -204 36932
rect -140 36868 -120 36932
rect -5492 36852 -120 36868
rect -5492 36788 -204 36852
rect -140 36788 -120 36852
rect -5492 36772 -120 36788
rect -5492 36708 -204 36772
rect -140 36708 -120 36772
rect -5492 36692 -120 36708
rect -5492 36628 -204 36692
rect -140 36628 -120 36692
rect -5492 36612 -120 36628
rect -5492 36548 -204 36612
rect -140 36548 -120 36612
rect -5492 36532 -120 36548
rect -5492 36468 -204 36532
rect -140 36468 -120 36532
rect -5492 36452 -120 36468
rect -5492 36388 -204 36452
rect -140 36388 -120 36452
rect -5492 36372 -120 36388
rect -5492 36308 -204 36372
rect -140 36308 -120 36372
rect -5492 36292 -120 36308
rect -5492 36228 -204 36292
rect -140 36228 -120 36292
rect -5492 36212 -120 36228
rect -5492 36148 -204 36212
rect -140 36148 -120 36212
rect -5492 36132 -120 36148
rect -5492 36068 -204 36132
rect -140 36068 -120 36132
rect -5492 36052 -120 36068
rect -5492 35988 -204 36052
rect -140 35988 -120 36052
rect -5492 35972 -120 35988
rect -5492 35908 -204 35972
rect -140 35908 -120 35972
rect -5492 35892 -120 35908
rect -5492 35828 -204 35892
rect -140 35828 -120 35892
rect -5492 35812 -120 35828
rect -5492 35748 -204 35812
rect -140 35748 -120 35812
rect -5492 35732 -120 35748
rect -5492 35668 -204 35732
rect -140 35668 -120 35732
rect -5492 35652 -120 35668
rect -5492 35588 -204 35652
rect -140 35588 -120 35652
rect -5492 35572 -120 35588
rect -5492 35508 -204 35572
rect -140 35508 -120 35572
rect -5492 35492 -120 35508
rect -5492 35428 -204 35492
rect -140 35428 -120 35492
rect -5492 35412 -120 35428
rect -5492 35348 -204 35412
rect -140 35348 -120 35412
rect -5492 35332 -120 35348
rect -5492 35268 -204 35332
rect -140 35268 -120 35332
rect -5492 35252 -120 35268
rect -5492 35188 -204 35252
rect -140 35188 -120 35252
rect -5492 35172 -120 35188
rect -5492 35108 -204 35172
rect -140 35108 -120 35172
rect -5492 35092 -120 35108
rect -5492 35028 -204 35092
rect -140 35028 -120 35092
rect -5492 35012 -120 35028
rect -5492 34948 -204 35012
rect -140 34948 -120 35012
rect -5492 34932 -120 34948
rect -5492 34868 -204 34932
rect -140 34868 -120 34932
rect -5492 34852 -120 34868
rect -5492 34788 -204 34852
rect -140 34788 -120 34852
rect -5492 34772 -120 34788
rect -5492 34708 -204 34772
rect -140 34708 -120 34772
rect -5492 34692 -120 34708
rect -5492 34628 -204 34692
rect -140 34628 -120 34692
rect -5492 34612 -120 34628
rect -5492 34548 -204 34612
rect -140 34548 -120 34612
rect -5492 34532 -120 34548
rect -5492 34468 -204 34532
rect -140 34468 -120 34532
rect -5492 34452 -120 34468
rect -5492 34388 -204 34452
rect -140 34388 -120 34452
rect -5492 34372 -120 34388
rect -5492 34308 -204 34372
rect -140 34308 -120 34372
rect -5492 34292 -120 34308
rect -5492 34228 -204 34292
rect -140 34228 -120 34292
rect -5492 34212 -120 34228
rect -5492 34148 -204 34212
rect -140 34148 -120 34212
rect -5492 34132 -120 34148
rect -5492 34068 -204 34132
rect -140 34068 -120 34132
rect -5492 34052 -120 34068
rect -5492 33988 -204 34052
rect -140 33988 -120 34052
rect -5492 33972 -120 33988
rect -5492 33908 -204 33972
rect -140 33908 -120 33972
rect -5492 33892 -120 33908
rect -5492 33828 -204 33892
rect -140 33828 -120 33892
rect -5492 33812 -120 33828
rect -5492 33748 -204 33812
rect -140 33748 -120 33812
rect -5492 33732 -120 33748
rect -5492 33668 -204 33732
rect -140 33668 -120 33732
rect -5492 33652 -120 33668
rect -5492 33588 -204 33652
rect -140 33588 -120 33652
rect -5492 33572 -120 33588
rect -5492 33508 -204 33572
rect -140 33508 -120 33572
rect -5492 33492 -120 33508
rect -5492 33428 -204 33492
rect -140 33428 -120 33492
rect -5492 33412 -120 33428
rect -5492 33348 -204 33412
rect -140 33348 -120 33412
rect -5492 33332 -120 33348
rect -5492 33268 -204 33332
rect -140 33268 -120 33332
rect -5492 33252 -120 33268
rect -5492 33188 -204 33252
rect -140 33188 -120 33252
rect -5492 33172 -120 33188
rect -5492 33108 -204 33172
rect -140 33108 -120 33172
rect -5492 33092 -120 33108
rect -5492 33028 -204 33092
rect -140 33028 -120 33092
rect -5492 33012 -120 33028
rect -5492 32948 -204 33012
rect -140 32948 -120 33012
rect -5492 32932 -120 32948
rect -5492 32868 -204 32932
rect -140 32868 -120 32932
rect -5492 32852 -120 32868
rect -5492 32788 -204 32852
rect -140 32788 -120 32852
rect -5492 32772 -120 32788
rect -5492 32708 -204 32772
rect -140 32708 -120 32772
rect -5492 32692 -120 32708
rect -5492 32628 -204 32692
rect -140 32628 -120 32692
rect -5492 32612 -120 32628
rect -5492 32548 -204 32612
rect -140 32548 -120 32612
rect -5492 32532 -120 32548
rect -5492 32468 -204 32532
rect -140 32468 -120 32532
rect -5492 32452 -120 32468
rect -5492 32388 -204 32452
rect -140 32388 -120 32452
rect -5492 32372 -120 32388
rect -5492 32308 -204 32372
rect -140 32308 -120 32372
rect -5492 32292 -120 32308
rect -5492 32228 -204 32292
rect -140 32228 -120 32292
rect -5492 32212 -120 32228
rect -5492 32148 -204 32212
rect -140 32148 -120 32212
rect -5492 32132 -120 32148
rect -5492 32068 -204 32132
rect -140 32068 -120 32132
rect -5492 32040 -120 32068
rect 120 37092 5492 37120
rect 120 37028 5408 37092
rect 5472 37028 5492 37092
rect 120 37012 5492 37028
rect 120 36948 5408 37012
rect 5472 36948 5492 37012
rect 120 36932 5492 36948
rect 120 36868 5408 36932
rect 5472 36868 5492 36932
rect 120 36852 5492 36868
rect 120 36788 5408 36852
rect 5472 36788 5492 36852
rect 120 36772 5492 36788
rect 120 36708 5408 36772
rect 5472 36708 5492 36772
rect 120 36692 5492 36708
rect 120 36628 5408 36692
rect 5472 36628 5492 36692
rect 120 36612 5492 36628
rect 120 36548 5408 36612
rect 5472 36548 5492 36612
rect 120 36532 5492 36548
rect 120 36468 5408 36532
rect 5472 36468 5492 36532
rect 120 36452 5492 36468
rect 120 36388 5408 36452
rect 5472 36388 5492 36452
rect 120 36372 5492 36388
rect 120 36308 5408 36372
rect 5472 36308 5492 36372
rect 120 36292 5492 36308
rect 120 36228 5408 36292
rect 5472 36228 5492 36292
rect 120 36212 5492 36228
rect 120 36148 5408 36212
rect 5472 36148 5492 36212
rect 120 36132 5492 36148
rect 120 36068 5408 36132
rect 5472 36068 5492 36132
rect 120 36052 5492 36068
rect 120 35988 5408 36052
rect 5472 35988 5492 36052
rect 120 35972 5492 35988
rect 120 35908 5408 35972
rect 5472 35908 5492 35972
rect 120 35892 5492 35908
rect 120 35828 5408 35892
rect 5472 35828 5492 35892
rect 120 35812 5492 35828
rect 120 35748 5408 35812
rect 5472 35748 5492 35812
rect 120 35732 5492 35748
rect 120 35668 5408 35732
rect 5472 35668 5492 35732
rect 120 35652 5492 35668
rect 120 35588 5408 35652
rect 5472 35588 5492 35652
rect 120 35572 5492 35588
rect 120 35508 5408 35572
rect 5472 35508 5492 35572
rect 120 35492 5492 35508
rect 120 35428 5408 35492
rect 5472 35428 5492 35492
rect 120 35412 5492 35428
rect 120 35348 5408 35412
rect 5472 35348 5492 35412
rect 120 35332 5492 35348
rect 120 35268 5408 35332
rect 5472 35268 5492 35332
rect 120 35252 5492 35268
rect 120 35188 5408 35252
rect 5472 35188 5492 35252
rect 120 35172 5492 35188
rect 120 35108 5408 35172
rect 5472 35108 5492 35172
rect 120 35092 5492 35108
rect 120 35028 5408 35092
rect 5472 35028 5492 35092
rect 120 35012 5492 35028
rect 120 34948 5408 35012
rect 5472 34948 5492 35012
rect 120 34932 5492 34948
rect 120 34868 5408 34932
rect 5472 34868 5492 34932
rect 120 34852 5492 34868
rect 120 34788 5408 34852
rect 5472 34788 5492 34852
rect 120 34772 5492 34788
rect 120 34708 5408 34772
rect 5472 34708 5492 34772
rect 120 34692 5492 34708
rect 120 34628 5408 34692
rect 5472 34628 5492 34692
rect 120 34612 5492 34628
rect 120 34548 5408 34612
rect 5472 34548 5492 34612
rect 120 34532 5492 34548
rect 120 34468 5408 34532
rect 5472 34468 5492 34532
rect 120 34452 5492 34468
rect 120 34388 5408 34452
rect 5472 34388 5492 34452
rect 120 34372 5492 34388
rect 120 34308 5408 34372
rect 5472 34308 5492 34372
rect 120 34292 5492 34308
rect 120 34228 5408 34292
rect 5472 34228 5492 34292
rect 120 34212 5492 34228
rect 120 34148 5408 34212
rect 5472 34148 5492 34212
rect 120 34132 5492 34148
rect 120 34068 5408 34132
rect 5472 34068 5492 34132
rect 120 34052 5492 34068
rect 120 33988 5408 34052
rect 5472 33988 5492 34052
rect 120 33972 5492 33988
rect 120 33908 5408 33972
rect 5472 33908 5492 33972
rect 120 33892 5492 33908
rect 120 33828 5408 33892
rect 5472 33828 5492 33892
rect 120 33812 5492 33828
rect 120 33748 5408 33812
rect 5472 33748 5492 33812
rect 120 33732 5492 33748
rect 120 33668 5408 33732
rect 5472 33668 5492 33732
rect 120 33652 5492 33668
rect 120 33588 5408 33652
rect 5472 33588 5492 33652
rect 120 33572 5492 33588
rect 120 33508 5408 33572
rect 5472 33508 5492 33572
rect 120 33492 5492 33508
rect 120 33428 5408 33492
rect 5472 33428 5492 33492
rect 120 33412 5492 33428
rect 120 33348 5408 33412
rect 5472 33348 5492 33412
rect 120 33332 5492 33348
rect 120 33268 5408 33332
rect 5472 33268 5492 33332
rect 120 33252 5492 33268
rect 120 33188 5408 33252
rect 5472 33188 5492 33252
rect 120 33172 5492 33188
rect 120 33108 5408 33172
rect 5472 33108 5492 33172
rect 120 33092 5492 33108
rect 120 33028 5408 33092
rect 5472 33028 5492 33092
rect 120 33012 5492 33028
rect 120 32948 5408 33012
rect 5472 32948 5492 33012
rect 120 32932 5492 32948
rect 120 32868 5408 32932
rect 5472 32868 5492 32932
rect 120 32852 5492 32868
rect 120 32788 5408 32852
rect 5472 32788 5492 32852
rect 120 32772 5492 32788
rect 120 32708 5408 32772
rect 5472 32708 5492 32772
rect 120 32692 5492 32708
rect 120 32628 5408 32692
rect 5472 32628 5492 32692
rect 120 32612 5492 32628
rect 120 32548 5408 32612
rect 5472 32548 5492 32612
rect 120 32532 5492 32548
rect 120 32468 5408 32532
rect 5472 32468 5492 32532
rect 120 32452 5492 32468
rect 120 32388 5408 32452
rect 5472 32388 5492 32452
rect 120 32372 5492 32388
rect 120 32308 5408 32372
rect 5472 32308 5492 32372
rect 120 32292 5492 32308
rect 120 32228 5408 32292
rect 5472 32228 5492 32292
rect 120 32212 5492 32228
rect 120 32148 5408 32212
rect 5472 32148 5492 32212
rect 120 32132 5492 32148
rect 120 32068 5408 32132
rect 5472 32068 5492 32132
rect 120 32040 5492 32068
rect 5732 37092 11104 37120
rect 5732 37028 11020 37092
rect 11084 37028 11104 37092
rect 5732 37012 11104 37028
rect 5732 36948 11020 37012
rect 11084 36948 11104 37012
rect 5732 36932 11104 36948
rect 5732 36868 11020 36932
rect 11084 36868 11104 36932
rect 5732 36852 11104 36868
rect 5732 36788 11020 36852
rect 11084 36788 11104 36852
rect 5732 36772 11104 36788
rect 5732 36708 11020 36772
rect 11084 36708 11104 36772
rect 5732 36692 11104 36708
rect 5732 36628 11020 36692
rect 11084 36628 11104 36692
rect 5732 36612 11104 36628
rect 5732 36548 11020 36612
rect 11084 36548 11104 36612
rect 5732 36532 11104 36548
rect 5732 36468 11020 36532
rect 11084 36468 11104 36532
rect 5732 36452 11104 36468
rect 5732 36388 11020 36452
rect 11084 36388 11104 36452
rect 5732 36372 11104 36388
rect 5732 36308 11020 36372
rect 11084 36308 11104 36372
rect 5732 36292 11104 36308
rect 5732 36228 11020 36292
rect 11084 36228 11104 36292
rect 5732 36212 11104 36228
rect 5732 36148 11020 36212
rect 11084 36148 11104 36212
rect 5732 36132 11104 36148
rect 5732 36068 11020 36132
rect 11084 36068 11104 36132
rect 5732 36052 11104 36068
rect 5732 35988 11020 36052
rect 11084 35988 11104 36052
rect 5732 35972 11104 35988
rect 5732 35908 11020 35972
rect 11084 35908 11104 35972
rect 5732 35892 11104 35908
rect 5732 35828 11020 35892
rect 11084 35828 11104 35892
rect 5732 35812 11104 35828
rect 5732 35748 11020 35812
rect 11084 35748 11104 35812
rect 5732 35732 11104 35748
rect 5732 35668 11020 35732
rect 11084 35668 11104 35732
rect 5732 35652 11104 35668
rect 5732 35588 11020 35652
rect 11084 35588 11104 35652
rect 5732 35572 11104 35588
rect 5732 35508 11020 35572
rect 11084 35508 11104 35572
rect 5732 35492 11104 35508
rect 5732 35428 11020 35492
rect 11084 35428 11104 35492
rect 5732 35412 11104 35428
rect 5732 35348 11020 35412
rect 11084 35348 11104 35412
rect 5732 35332 11104 35348
rect 5732 35268 11020 35332
rect 11084 35268 11104 35332
rect 5732 35252 11104 35268
rect 5732 35188 11020 35252
rect 11084 35188 11104 35252
rect 5732 35172 11104 35188
rect 5732 35108 11020 35172
rect 11084 35108 11104 35172
rect 5732 35092 11104 35108
rect 5732 35028 11020 35092
rect 11084 35028 11104 35092
rect 5732 35012 11104 35028
rect 5732 34948 11020 35012
rect 11084 34948 11104 35012
rect 5732 34932 11104 34948
rect 5732 34868 11020 34932
rect 11084 34868 11104 34932
rect 5732 34852 11104 34868
rect 5732 34788 11020 34852
rect 11084 34788 11104 34852
rect 5732 34772 11104 34788
rect 5732 34708 11020 34772
rect 11084 34708 11104 34772
rect 5732 34692 11104 34708
rect 5732 34628 11020 34692
rect 11084 34628 11104 34692
rect 5732 34612 11104 34628
rect 5732 34548 11020 34612
rect 11084 34548 11104 34612
rect 5732 34532 11104 34548
rect 5732 34468 11020 34532
rect 11084 34468 11104 34532
rect 5732 34452 11104 34468
rect 5732 34388 11020 34452
rect 11084 34388 11104 34452
rect 5732 34372 11104 34388
rect 5732 34308 11020 34372
rect 11084 34308 11104 34372
rect 5732 34292 11104 34308
rect 5732 34228 11020 34292
rect 11084 34228 11104 34292
rect 5732 34212 11104 34228
rect 5732 34148 11020 34212
rect 11084 34148 11104 34212
rect 5732 34132 11104 34148
rect 5732 34068 11020 34132
rect 11084 34068 11104 34132
rect 5732 34052 11104 34068
rect 5732 33988 11020 34052
rect 11084 33988 11104 34052
rect 5732 33972 11104 33988
rect 5732 33908 11020 33972
rect 11084 33908 11104 33972
rect 5732 33892 11104 33908
rect 5732 33828 11020 33892
rect 11084 33828 11104 33892
rect 5732 33812 11104 33828
rect 5732 33748 11020 33812
rect 11084 33748 11104 33812
rect 5732 33732 11104 33748
rect 5732 33668 11020 33732
rect 11084 33668 11104 33732
rect 5732 33652 11104 33668
rect 5732 33588 11020 33652
rect 11084 33588 11104 33652
rect 5732 33572 11104 33588
rect 5732 33508 11020 33572
rect 11084 33508 11104 33572
rect 5732 33492 11104 33508
rect 5732 33428 11020 33492
rect 11084 33428 11104 33492
rect 5732 33412 11104 33428
rect 5732 33348 11020 33412
rect 11084 33348 11104 33412
rect 5732 33332 11104 33348
rect 5732 33268 11020 33332
rect 11084 33268 11104 33332
rect 5732 33252 11104 33268
rect 5732 33188 11020 33252
rect 11084 33188 11104 33252
rect 5732 33172 11104 33188
rect 5732 33108 11020 33172
rect 11084 33108 11104 33172
rect 5732 33092 11104 33108
rect 5732 33028 11020 33092
rect 11084 33028 11104 33092
rect 5732 33012 11104 33028
rect 5732 32948 11020 33012
rect 11084 32948 11104 33012
rect 5732 32932 11104 32948
rect 5732 32868 11020 32932
rect 11084 32868 11104 32932
rect 5732 32852 11104 32868
rect 5732 32788 11020 32852
rect 11084 32788 11104 32852
rect 5732 32772 11104 32788
rect 5732 32708 11020 32772
rect 11084 32708 11104 32772
rect 5732 32692 11104 32708
rect 5732 32628 11020 32692
rect 11084 32628 11104 32692
rect 5732 32612 11104 32628
rect 5732 32548 11020 32612
rect 11084 32548 11104 32612
rect 5732 32532 11104 32548
rect 5732 32468 11020 32532
rect 11084 32468 11104 32532
rect 5732 32452 11104 32468
rect 5732 32388 11020 32452
rect 11084 32388 11104 32452
rect 5732 32372 11104 32388
rect 5732 32308 11020 32372
rect 11084 32308 11104 32372
rect 5732 32292 11104 32308
rect 5732 32228 11020 32292
rect 11084 32228 11104 32292
rect 5732 32212 11104 32228
rect 5732 32148 11020 32212
rect 11084 32148 11104 32212
rect 5732 32132 11104 32148
rect 5732 32068 11020 32132
rect 11084 32068 11104 32132
rect 5732 32040 11104 32068
rect 11344 37092 16716 37120
rect 11344 37028 16632 37092
rect 16696 37028 16716 37092
rect 11344 37012 16716 37028
rect 11344 36948 16632 37012
rect 16696 36948 16716 37012
rect 11344 36932 16716 36948
rect 11344 36868 16632 36932
rect 16696 36868 16716 36932
rect 11344 36852 16716 36868
rect 11344 36788 16632 36852
rect 16696 36788 16716 36852
rect 11344 36772 16716 36788
rect 11344 36708 16632 36772
rect 16696 36708 16716 36772
rect 11344 36692 16716 36708
rect 11344 36628 16632 36692
rect 16696 36628 16716 36692
rect 11344 36612 16716 36628
rect 11344 36548 16632 36612
rect 16696 36548 16716 36612
rect 11344 36532 16716 36548
rect 11344 36468 16632 36532
rect 16696 36468 16716 36532
rect 11344 36452 16716 36468
rect 11344 36388 16632 36452
rect 16696 36388 16716 36452
rect 11344 36372 16716 36388
rect 11344 36308 16632 36372
rect 16696 36308 16716 36372
rect 11344 36292 16716 36308
rect 11344 36228 16632 36292
rect 16696 36228 16716 36292
rect 11344 36212 16716 36228
rect 11344 36148 16632 36212
rect 16696 36148 16716 36212
rect 11344 36132 16716 36148
rect 11344 36068 16632 36132
rect 16696 36068 16716 36132
rect 11344 36052 16716 36068
rect 11344 35988 16632 36052
rect 16696 35988 16716 36052
rect 11344 35972 16716 35988
rect 11344 35908 16632 35972
rect 16696 35908 16716 35972
rect 11344 35892 16716 35908
rect 11344 35828 16632 35892
rect 16696 35828 16716 35892
rect 11344 35812 16716 35828
rect 11344 35748 16632 35812
rect 16696 35748 16716 35812
rect 11344 35732 16716 35748
rect 11344 35668 16632 35732
rect 16696 35668 16716 35732
rect 11344 35652 16716 35668
rect 11344 35588 16632 35652
rect 16696 35588 16716 35652
rect 11344 35572 16716 35588
rect 11344 35508 16632 35572
rect 16696 35508 16716 35572
rect 11344 35492 16716 35508
rect 11344 35428 16632 35492
rect 16696 35428 16716 35492
rect 11344 35412 16716 35428
rect 11344 35348 16632 35412
rect 16696 35348 16716 35412
rect 11344 35332 16716 35348
rect 11344 35268 16632 35332
rect 16696 35268 16716 35332
rect 11344 35252 16716 35268
rect 11344 35188 16632 35252
rect 16696 35188 16716 35252
rect 11344 35172 16716 35188
rect 11344 35108 16632 35172
rect 16696 35108 16716 35172
rect 11344 35092 16716 35108
rect 11344 35028 16632 35092
rect 16696 35028 16716 35092
rect 11344 35012 16716 35028
rect 11344 34948 16632 35012
rect 16696 34948 16716 35012
rect 11344 34932 16716 34948
rect 11344 34868 16632 34932
rect 16696 34868 16716 34932
rect 11344 34852 16716 34868
rect 11344 34788 16632 34852
rect 16696 34788 16716 34852
rect 11344 34772 16716 34788
rect 11344 34708 16632 34772
rect 16696 34708 16716 34772
rect 11344 34692 16716 34708
rect 11344 34628 16632 34692
rect 16696 34628 16716 34692
rect 11344 34612 16716 34628
rect 11344 34548 16632 34612
rect 16696 34548 16716 34612
rect 11344 34532 16716 34548
rect 11344 34468 16632 34532
rect 16696 34468 16716 34532
rect 11344 34452 16716 34468
rect 11344 34388 16632 34452
rect 16696 34388 16716 34452
rect 11344 34372 16716 34388
rect 11344 34308 16632 34372
rect 16696 34308 16716 34372
rect 11344 34292 16716 34308
rect 11344 34228 16632 34292
rect 16696 34228 16716 34292
rect 11344 34212 16716 34228
rect 11344 34148 16632 34212
rect 16696 34148 16716 34212
rect 11344 34132 16716 34148
rect 11344 34068 16632 34132
rect 16696 34068 16716 34132
rect 11344 34052 16716 34068
rect 11344 33988 16632 34052
rect 16696 33988 16716 34052
rect 11344 33972 16716 33988
rect 11344 33908 16632 33972
rect 16696 33908 16716 33972
rect 11344 33892 16716 33908
rect 11344 33828 16632 33892
rect 16696 33828 16716 33892
rect 11344 33812 16716 33828
rect 11344 33748 16632 33812
rect 16696 33748 16716 33812
rect 11344 33732 16716 33748
rect 11344 33668 16632 33732
rect 16696 33668 16716 33732
rect 11344 33652 16716 33668
rect 11344 33588 16632 33652
rect 16696 33588 16716 33652
rect 11344 33572 16716 33588
rect 11344 33508 16632 33572
rect 16696 33508 16716 33572
rect 11344 33492 16716 33508
rect 11344 33428 16632 33492
rect 16696 33428 16716 33492
rect 11344 33412 16716 33428
rect 11344 33348 16632 33412
rect 16696 33348 16716 33412
rect 11344 33332 16716 33348
rect 11344 33268 16632 33332
rect 16696 33268 16716 33332
rect 11344 33252 16716 33268
rect 11344 33188 16632 33252
rect 16696 33188 16716 33252
rect 11344 33172 16716 33188
rect 11344 33108 16632 33172
rect 16696 33108 16716 33172
rect 11344 33092 16716 33108
rect 11344 33028 16632 33092
rect 16696 33028 16716 33092
rect 11344 33012 16716 33028
rect 11344 32948 16632 33012
rect 16696 32948 16716 33012
rect 11344 32932 16716 32948
rect 11344 32868 16632 32932
rect 16696 32868 16716 32932
rect 11344 32852 16716 32868
rect 11344 32788 16632 32852
rect 16696 32788 16716 32852
rect 11344 32772 16716 32788
rect 11344 32708 16632 32772
rect 16696 32708 16716 32772
rect 11344 32692 16716 32708
rect 11344 32628 16632 32692
rect 16696 32628 16716 32692
rect 11344 32612 16716 32628
rect 11344 32548 16632 32612
rect 16696 32548 16716 32612
rect 11344 32532 16716 32548
rect 11344 32468 16632 32532
rect 16696 32468 16716 32532
rect 11344 32452 16716 32468
rect 11344 32388 16632 32452
rect 16696 32388 16716 32452
rect 11344 32372 16716 32388
rect 11344 32308 16632 32372
rect 16696 32308 16716 32372
rect 11344 32292 16716 32308
rect 11344 32228 16632 32292
rect 16696 32228 16716 32292
rect 11344 32212 16716 32228
rect 11344 32148 16632 32212
rect 16696 32148 16716 32212
rect 11344 32132 16716 32148
rect 11344 32068 16632 32132
rect 16696 32068 16716 32132
rect 11344 32040 16716 32068
rect 16956 37092 22328 37120
rect 16956 37028 22244 37092
rect 22308 37028 22328 37092
rect 16956 37012 22328 37028
rect 16956 36948 22244 37012
rect 22308 36948 22328 37012
rect 16956 36932 22328 36948
rect 16956 36868 22244 36932
rect 22308 36868 22328 36932
rect 16956 36852 22328 36868
rect 16956 36788 22244 36852
rect 22308 36788 22328 36852
rect 16956 36772 22328 36788
rect 16956 36708 22244 36772
rect 22308 36708 22328 36772
rect 16956 36692 22328 36708
rect 16956 36628 22244 36692
rect 22308 36628 22328 36692
rect 16956 36612 22328 36628
rect 16956 36548 22244 36612
rect 22308 36548 22328 36612
rect 16956 36532 22328 36548
rect 16956 36468 22244 36532
rect 22308 36468 22328 36532
rect 16956 36452 22328 36468
rect 16956 36388 22244 36452
rect 22308 36388 22328 36452
rect 16956 36372 22328 36388
rect 16956 36308 22244 36372
rect 22308 36308 22328 36372
rect 16956 36292 22328 36308
rect 16956 36228 22244 36292
rect 22308 36228 22328 36292
rect 16956 36212 22328 36228
rect 16956 36148 22244 36212
rect 22308 36148 22328 36212
rect 16956 36132 22328 36148
rect 16956 36068 22244 36132
rect 22308 36068 22328 36132
rect 16956 36052 22328 36068
rect 16956 35988 22244 36052
rect 22308 35988 22328 36052
rect 16956 35972 22328 35988
rect 16956 35908 22244 35972
rect 22308 35908 22328 35972
rect 16956 35892 22328 35908
rect 16956 35828 22244 35892
rect 22308 35828 22328 35892
rect 16956 35812 22328 35828
rect 16956 35748 22244 35812
rect 22308 35748 22328 35812
rect 16956 35732 22328 35748
rect 16956 35668 22244 35732
rect 22308 35668 22328 35732
rect 16956 35652 22328 35668
rect 16956 35588 22244 35652
rect 22308 35588 22328 35652
rect 16956 35572 22328 35588
rect 16956 35508 22244 35572
rect 22308 35508 22328 35572
rect 16956 35492 22328 35508
rect 16956 35428 22244 35492
rect 22308 35428 22328 35492
rect 16956 35412 22328 35428
rect 16956 35348 22244 35412
rect 22308 35348 22328 35412
rect 16956 35332 22328 35348
rect 16956 35268 22244 35332
rect 22308 35268 22328 35332
rect 16956 35252 22328 35268
rect 16956 35188 22244 35252
rect 22308 35188 22328 35252
rect 16956 35172 22328 35188
rect 16956 35108 22244 35172
rect 22308 35108 22328 35172
rect 16956 35092 22328 35108
rect 16956 35028 22244 35092
rect 22308 35028 22328 35092
rect 16956 35012 22328 35028
rect 16956 34948 22244 35012
rect 22308 34948 22328 35012
rect 16956 34932 22328 34948
rect 16956 34868 22244 34932
rect 22308 34868 22328 34932
rect 16956 34852 22328 34868
rect 16956 34788 22244 34852
rect 22308 34788 22328 34852
rect 16956 34772 22328 34788
rect 16956 34708 22244 34772
rect 22308 34708 22328 34772
rect 16956 34692 22328 34708
rect 16956 34628 22244 34692
rect 22308 34628 22328 34692
rect 16956 34612 22328 34628
rect 16956 34548 22244 34612
rect 22308 34548 22328 34612
rect 16956 34532 22328 34548
rect 16956 34468 22244 34532
rect 22308 34468 22328 34532
rect 16956 34452 22328 34468
rect 16956 34388 22244 34452
rect 22308 34388 22328 34452
rect 16956 34372 22328 34388
rect 16956 34308 22244 34372
rect 22308 34308 22328 34372
rect 16956 34292 22328 34308
rect 16956 34228 22244 34292
rect 22308 34228 22328 34292
rect 16956 34212 22328 34228
rect 16956 34148 22244 34212
rect 22308 34148 22328 34212
rect 16956 34132 22328 34148
rect 16956 34068 22244 34132
rect 22308 34068 22328 34132
rect 16956 34052 22328 34068
rect 16956 33988 22244 34052
rect 22308 33988 22328 34052
rect 16956 33972 22328 33988
rect 16956 33908 22244 33972
rect 22308 33908 22328 33972
rect 16956 33892 22328 33908
rect 16956 33828 22244 33892
rect 22308 33828 22328 33892
rect 16956 33812 22328 33828
rect 16956 33748 22244 33812
rect 22308 33748 22328 33812
rect 16956 33732 22328 33748
rect 16956 33668 22244 33732
rect 22308 33668 22328 33732
rect 16956 33652 22328 33668
rect 16956 33588 22244 33652
rect 22308 33588 22328 33652
rect 16956 33572 22328 33588
rect 16956 33508 22244 33572
rect 22308 33508 22328 33572
rect 16956 33492 22328 33508
rect 16956 33428 22244 33492
rect 22308 33428 22328 33492
rect 16956 33412 22328 33428
rect 16956 33348 22244 33412
rect 22308 33348 22328 33412
rect 16956 33332 22328 33348
rect 16956 33268 22244 33332
rect 22308 33268 22328 33332
rect 16956 33252 22328 33268
rect 16956 33188 22244 33252
rect 22308 33188 22328 33252
rect 16956 33172 22328 33188
rect 16956 33108 22244 33172
rect 22308 33108 22328 33172
rect 16956 33092 22328 33108
rect 16956 33028 22244 33092
rect 22308 33028 22328 33092
rect 16956 33012 22328 33028
rect 16956 32948 22244 33012
rect 22308 32948 22328 33012
rect 16956 32932 22328 32948
rect 16956 32868 22244 32932
rect 22308 32868 22328 32932
rect 16956 32852 22328 32868
rect 16956 32788 22244 32852
rect 22308 32788 22328 32852
rect 16956 32772 22328 32788
rect 16956 32708 22244 32772
rect 22308 32708 22328 32772
rect 16956 32692 22328 32708
rect 16956 32628 22244 32692
rect 22308 32628 22328 32692
rect 16956 32612 22328 32628
rect 16956 32548 22244 32612
rect 22308 32548 22328 32612
rect 16956 32532 22328 32548
rect 16956 32468 22244 32532
rect 22308 32468 22328 32532
rect 16956 32452 22328 32468
rect 16956 32388 22244 32452
rect 22308 32388 22328 32452
rect 16956 32372 22328 32388
rect 16956 32308 22244 32372
rect 22308 32308 22328 32372
rect 16956 32292 22328 32308
rect 16956 32228 22244 32292
rect 22308 32228 22328 32292
rect 16956 32212 22328 32228
rect 16956 32148 22244 32212
rect 22308 32148 22328 32212
rect 16956 32132 22328 32148
rect 16956 32068 22244 32132
rect 22308 32068 22328 32132
rect 16956 32040 22328 32068
rect 22568 37092 27940 37120
rect 22568 37028 27856 37092
rect 27920 37028 27940 37092
rect 22568 37012 27940 37028
rect 22568 36948 27856 37012
rect 27920 36948 27940 37012
rect 22568 36932 27940 36948
rect 22568 36868 27856 36932
rect 27920 36868 27940 36932
rect 22568 36852 27940 36868
rect 22568 36788 27856 36852
rect 27920 36788 27940 36852
rect 22568 36772 27940 36788
rect 22568 36708 27856 36772
rect 27920 36708 27940 36772
rect 22568 36692 27940 36708
rect 22568 36628 27856 36692
rect 27920 36628 27940 36692
rect 22568 36612 27940 36628
rect 22568 36548 27856 36612
rect 27920 36548 27940 36612
rect 22568 36532 27940 36548
rect 22568 36468 27856 36532
rect 27920 36468 27940 36532
rect 22568 36452 27940 36468
rect 22568 36388 27856 36452
rect 27920 36388 27940 36452
rect 22568 36372 27940 36388
rect 22568 36308 27856 36372
rect 27920 36308 27940 36372
rect 22568 36292 27940 36308
rect 22568 36228 27856 36292
rect 27920 36228 27940 36292
rect 22568 36212 27940 36228
rect 22568 36148 27856 36212
rect 27920 36148 27940 36212
rect 22568 36132 27940 36148
rect 22568 36068 27856 36132
rect 27920 36068 27940 36132
rect 22568 36052 27940 36068
rect 22568 35988 27856 36052
rect 27920 35988 27940 36052
rect 22568 35972 27940 35988
rect 22568 35908 27856 35972
rect 27920 35908 27940 35972
rect 22568 35892 27940 35908
rect 22568 35828 27856 35892
rect 27920 35828 27940 35892
rect 22568 35812 27940 35828
rect 22568 35748 27856 35812
rect 27920 35748 27940 35812
rect 22568 35732 27940 35748
rect 22568 35668 27856 35732
rect 27920 35668 27940 35732
rect 22568 35652 27940 35668
rect 22568 35588 27856 35652
rect 27920 35588 27940 35652
rect 22568 35572 27940 35588
rect 22568 35508 27856 35572
rect 27920 35508 27940 35572
rect 22568 35492 27940 35508
rect 22568 35428 27856 35492
rect 27920 35428 27940 35492
rect 22568 35412 27940 35428
rect 22568 35348 27856 35412
rect 27920 35348 27940 35412
rect 22568 35332 27940 35348
rect 22568 35268 27856 35332
rect 27920 35268 27940 35332
rect 22568 35252 27940 35268
rect 22568 35188 27856 35252
rect 27920 35188 27940 35252
rect 22568 35172 27940 35188
rect 22568 35108 27856 35172
rect 27920 35108 27940 35172
rect 22568 35092 27940 35108
rect 22568 35028 27856 35092
rect 27920 35028 27940 35092
rect 22568 35012 27940 35028
rect 22568 34948 27856 35012
rect 27920 34948 27940 35012
rect 22568 34932 27940 34948
rect 22568 34868 27856 34932
rect 27920 34868 27940 34932
rect 22568 34852 27940 34868
rect 22568 34788 27856 34852
rect 27920 34788 27940 34852
rect 22568 34772 27940 34788
rect 22568 34708 27856 34772
rect 27920 34708 27940 34772
rect 22568 34692 27940 34708
rect 22568 34628 27856 34692
rect 27920 34628 27940 34692
rect 22568 34612 27940 34628
rect 22568 34548 27856 34612
rect 27920 34548 27940 34612
rect 22568 34532 27940 34548
rect 22568 34468 27856 34532
rect 27920 34468 27940 34532
rect 22568 34452 27940 34468
rect 22568 34388 27856 34452
rect 27920 34388 27940 34452
rect 22568 34372 27940 34388
rect 22568 34308 27856 34372
rect 27920 34308 27940 34372
rect 22568 34292 27940 34308
rect 22568 34228 27856 34292
rect 27920 34228 27940 34292
rect 22568 34212 27940 34228
rect 22568 34148 27856 34212
rect 27920 34148 27940 34212
rect 22568 34132 27940 34148
rect 22568 34068 27856 34132
rect 27920 34068 27940 34132
rect 22568 34052 27940 34068
rect 22568 33988 27856 34052
rect 27920 33988 27940 34052
rect 22568 33972 27940 33988
rect 22568 33908 27856 33972
rect 27920 33908 27940 33972
rect 22568 33892 27940 33908
rect 22568 33828 27856 33892
rect 27920 33828 27940 33892
rect 22568 33812 27940 33828
rect 22568 33748 27856 33812
rect 27920 33748 27940 33812
rect 22568 33732 27940 33748
rect 22568 33668 27856 33732
rect 27920 33668 27940 33732
rect 22568 33652 27940 33668
rect 22568 33588 27856 33652
rect 27920 33588 27940 33652
rect 22568 33572 27940 33588
rect 22568 33508 27856 33572
rect 27920 33508 27940 33572
rect 22568 33492 27940 33508
rect 22568 33428 27856 33492
rect 27920 33428 27940 33492
rect 22568 33412 27940 33428
rect 22568 33348 27856 33412
rect 27920 33348 27940 33412
rect 22568 33332 27940 33348
rect 22568 33268 27856 33332
rect 27920 33268 27940 33332
rect 22568 33252 27940 33268
rect 22568 33188 27856 33252
rect 27920 33188 27940 33252
rect 22568 33172 27940 33188
rect 22568 33108 27856 33172
rect 27920 33108 27940 33172
rect 22568 33092 27940 33108
rect 22568 33028 27856 33092
rect 27920 33028 27940 33092
rect 22568 33012 27940 33028
rect 22568 32948 27856 33012
rect 27920 32948 27940 33012
rect 22568 32932 27940 32948
rect 22568 32868 27856 32932
rect 27920 32868 27940 32932
rect 22568 32852 27940 32868
rect 22568 32788 27856 32852
rect 27920 32788 27940 32852
rect 22568 32772 27940 32788
rect 22568 32708 27856 32772
rect 27920 32708 27940 32772
rect 22568 32692 27940 32708
rect 22568 32628 27856 32692
rect 27920 32628 27940 32692
rect 22568 32612 27940 32628
rect 22568 32548 27856 32612
rect 27920 32548 27940 32612
rect 22568 32532 27940 32548
rect 22568 32468 27856 32532
rect 27920 32468 27940 32532
rect 22568 32452 27940 32468
rect 22568 32388 27856 32452
rect 27920 32388 27940 32452
rect 22568 32372 27940 32388
rect 22568 32308 27856 32372
rect 27920 32308 27940 32372
rect 22568 32292 27940 32308
rect 22568 32228 27856 32292
rect 27920 32228 27940 32292
rect 22568 32212 27940 32228
rect 22568 32148 27856 32212
rect 27920 32148 27940 32212
rect 22568 32132 27940 32148
rect 22568 32068 27856 32132
rect 27920 32068 27940 32132
rect 22568 32040 27940 32068
rect 28180 37092 33552 37120
rect 28180 37028 33468 37092
rect 33532 37028 33552 37092
rect 28180 37012 33552 37028
rect 28180 36948 33468 37012
rect 33532 36948 33552 37012
rect 28180 36932 33552 36948
rect 28180 36868 33468 36932
rect 33532 36868 33552 36932
rect 28180 36852 33552 36868
rect 28180 36788 33468 36852
rect 33532 36788 33552 36852
rect 28180 36772 33552 36788
rect 28180 36708 33468 36772
rect 33532 36708 33552 36772
rect 28180 36692 33552 36708
rect 28180 36628 33468 36692
rect 33532 36628 33552 36692
rect 28180 36612 33552 36628
rect 28180 36548 33468 36612
rect 33532 36548 33552 36612
rect 28180 36532 33552 36548
rect 28180 36468 33468 36532
rect 33532 36468 33552 36532
rect 28180 36452 33552 36468
rect 28180 36388 33468 36452
rect 33532 36388 33552 36452
rect 28180 36372 33552 36388
rect 28180 36308 33468 36372
rect 33532 36308 33552 36372
rect 28180 36292 33552 36308
rect 28180 36228 33468 36292
rect 33532 36228 33552 36292
rect 28180 36212 33552 36228
rect 28180 36148 33468 36212
rect 33532 36148 33552 36212
rect 28180 36132 33552 36148
rect 28180 36068 33468 36132
rect 33532 36068 33552 36132
rect 28180 36052 33552 36068
rect 28180 35988 33468 36052
rect 33532 35988 33552 36052
rect 28180 35972 33552 35988
rect 28180 35908 33468 35972
rect 33532 35908 33552 35972
rect 28180 35892 33552 35908
rect 28180 35828 33468 35892
rect 33532 35828 33552 35892
rect 28180 35812 33552 35828
rect 28180 35748 33468 35812
rect 33532 35748 33552 35812
rect 28180 35732 33552 35748
rect 28180 35668 33468 35732
rect 33532 35668 33552 35732
rect 28180 35652 33552 35668
rect 28180 35588 33468 35652
rect 33532 35588 33552 35652
rect 28180 35572 33552 35588
rect 28180 35508 33468 35572
rect 33532 35508 33552 35572
rect 28180 35492 33552 35508
rect 28180 35428 33468 35492
rect 33532 35428 33552 35492
rect 28180 35412 33552 35428
rect 28180 35348 33468 35412
rect 33532 35348 33552 35412
rect 28180 35332 33552 35348
rect 28180 35268 33468 35332
rect 33532 35268 33552 35332
rect 28180 35252 33552 35268
rect 28180 35188 33468 35252
rect 33532 35188 33552 35252
rect 28180 35172 33552 35188
rect 28180 35108 33468 35172
rect 33532 35108 33552 35172
rect 28180 35092 33552 35108
rect 28180 35028 33468 35092
rect 33532 35028 33552 35092
rect 28180 35012 33552 35028
rect 28180 34948 33468 35012
rect 33532 34948 33552 35012
rect 28180 34932 33552 34948
rect 28180 34868 33468 34932
rect 33532 34868 33552 34932
rect 28180 34852 33552 34868
rect 28180 34788 33468 34852
rect 33532 34788 33552 34852
rect 28180 34772 33552 34788
rect 28180 34708 33468 34772
rect 33532 34708 33552 34772
rect 28180 34692 33552 34708
rect 28180 34628 33468 34692
rect 33532 34628 33552 34692
rect 28180 34612 33552 34628
rect 28180 34548 33468 34612
rect 33532 34548 33552 34612
rect 28180 34532 33552 34548
rect 28180 34468 33468 34532
rect 33532 34468 33552 34532
rect 28180 34452 33552 34468
rect 28180 34388 33468 34452
rect 33532 34388 33552 34452
rect 28180 34372 33552 34388
rect 28180 34308 33468 34372
rect 33532 34308 33552 34372
rect 28180 34292 33552 34308
rect 28180 34228 33468 34292
rect 33532 34228 33552 34292
rect 28180 34212 33552 34228
rect 28180 34148 33468 34212
rect 33532 34148 33552 34212
rect 28180 34132 33552 34148
rect 28180 34068 33468 34132
rect 33532 34068 33552 34132
rect 28180 34052 33552 34068
rect 28180 33988 33468 34052
rect 33532 33988 33552 34052
rect 28180 33972 33552 33988
rect 28180 33908 33468 33972
rect 33532 33908 33552 33972
rect 28180 33892 33552 33908
rect 28180 33828 33468 33892
rect 33532 33828 33552 33892
rect 28180 33812 33552 33828
rect 28180 33748 33468 33812
rect 33532 33748 33552 33812
rect 28180 33732 33552 33748
rect 28180 33668 33468 33732
rect 33532 33668 33552 33732
rect 28180 33652 33552 33668
rect 28180 33588 33468 33652
rect 33532 33588 33552 33652
rect 28180 33572 33552 33588
rect 28180 33508 33468 33572
rect 33532 33508 33552 33572
rect 28180 33492 33552 33508
rect 28180 33428 33468 33492
rect 33532 33428 33552 33492
rect 28180 33412 33552 33428
rect 28180 33348 33468 33412
rect 33532 33348 33552 33412
rect 28180 33332 33552 33348
rect 28180 33268 33468 33332
rect 33532 33268 33552 33332
rect 28180 33252 33552 33268
rect 28180 33188 33468 33252
rect 33532 33188 33552 33252
rect 28180 33172 33552 33188
rect 28180 33108 33468 33172
rect 33532 33108 33552 33172
rect 28180 33092 33552 33108
rect 28180 33028 33468 33092
rect 33532 33028 33552 33092
rect 28180 33012 33552 33028
rect 28180 32948 33468 33012
rect 33532 32948 33552 33012
rect 28180 32932 33552 32948
rect 28180 32868 33468 32932
rect 33532 32868 33552 32932
rect 28180 32852 33552 32868
rect 28180 32788 33468 32852
rect 33532 32788 33552 32852
rect 28180 32772 33552 32788
rect 28180 32708 33468 32772
rect 33532 32708 33552 32772
rect 28180 32692 33552 32708
rect 28180 32628 33468 32692
rect 33532 32628 33552 32692
rect 28180 32612 33552 32628
rect 28180 32548 33468 32612
rect 33532 32548 33552 32612
rect 28180 32532 33552 32548
rect 28180 32468 33468 32532
rect 33532 32468 33552 32532
rect 28180 32452 33552 32468
rect 28180 32388 33468 32452
rect 33532 32388 33552 32452
rect 28180 32372 33552 32388
rect 28180 32308 33468 32372
rect 33532 32308 33552 32372
rect 28180 32292 33552 32308
rect 28180 32228 33468 32292
rect 33532 32228 33552 32292
rect 28180 32212 33552 32228
rect 28180 32148 33468 32212
rect 33532 32148 33552 32212
rect 28180 32132 33552 32148
rect 28180 32068 33468 32132
rect 33532 32068 33552 32132
rect 28180 32040 33552 32068
rect 33792 37092 39164 37120
rect 33792 37028 39080 37092
rect 39144 37028 39164 37092
rect 33792 37012 39164 37028
rect 33792 36948 39080 37012
rect 39144 36948 39164 37012
rect 33792 36932 39164 36948
rect 33792 36868 39080 36932
rect 39144 36868 39164 36932
rect 33792 36852 39164 36868
rect 33792 36788 39080 36852
rect 39144 36788 39164 36852
rect 33792 36772 39164 36788
rect 33792 36708 39080 36772
rect 39144 36708 39164 36772
rect 33792 36692 39164 36708
rect 33792 36628 39080 36692
rect 39144 36628 39164 36692
rect 33792 36612 39164 36628
rect 33792 36548 39080 36612
rect 39144 36548 39164 36612
rect 33792 36532 39164 36548
rect 33792 36468 39080 36532
rect 39144 36468 39164 36532
rect 33792 36452 39164 36468
rect 33792 36388 39080 36452
rect 39144 36388 39164 36452
rect 33792 36372 39164 36388
rect 33792 36308 39080 36372
rect 39144 36308 39164 36372
rect 33792 36292 39164 36308
rect 33792 36228 39080 36292
rect 39144 36228 39164 36292
rect 33792 36212 39164 36228
rect 33792 36148 39080 36212
rect 39144 36148 39164 36212
rect 33792 36132 39164 36148
rect 33792 36068 39080 36132
rect 39144 36068 39164 36132
rect 33792 36052 39164 36068
rect 33792 35988 39080 36052
rect 39144 35988 39164 36052
rect 33792 35972 39164 35988
rect 33792 35908 39080 35972
rect 39144 35908 39164 35972
rect 33792 35892 39164 35908
rect 33792 35828 39080 35892
rect 39144 35828 39164 35892
rect 33792 35812 39164 35828
rect 33792 35748 39080 35812
rect 39144 35748 39164 35812
rect 33792 35732 39164 35748
rect 33792 35668 39080 35732
rect 39144 35668 39164 35732
rect 33792 35652 39164 35668
rect 33792 35588 39080 35652
rect 39144 35588 39164 35652
rect 33792 35572 39164 35588
rect 33792 35508 39080 35572
rect 39144 35508 39164 35572
rect 33792 35492 39164 35508
rect 33792 35428 39080 35492
rect 39144 35428 39164 35492
rect 33792 35412 39164 35428
rect 33792 35348 39080 35412
rect 39144 35348 39164 35412
rect 33792 35332 39164 35348
rect 33792 35268 39080 35332
rect 39144 35268 39164 35332
rect 33792 35252 39164 35268
rect 33792 35188 39080 35252
rect 39144 35188 39164 35252
rect 33792 35172 39164 35188
rect 33792 35108 39080 35172
rect 39144 35108 39164 35172
rect 33792 35092 39164 35108
rect 33792 35028 39080 35092
rect 39144 35028 39164 35092
rect 33792 35012 39164 35028
rect 33792 34948 39080 35012
rect 39144 34948 39164 35012
rect 33792 34932 39164 34948
rect 33792 34868 39080 34932
rect 39144 34868 39164 34932
rect 33792 34852 39164 34868
rect 33792 34788 39080 34852
rect 39144 34788 39164 34852
rect 33792 34772 39164 34788
rect 33792 34708 39080 34772
rect 39144 34708 39164 34772
rect 33792 34692 39164 34708
rect 33792 34628 39080 34692
rect 39144 34628 39164 34692
rect 33792 34612 39164 34628
rect 33792 34548 39080 34612
rect 39144 34548 39164 34612
rect 33792 34532 39164 34548
rect 33792 34468 39080 34532
rect 39144 34468 39164 34532
rect 33792 34452 39164 34468
rect 33792 34388 39080 34452
rect 39144 34388 39164 34452
rect 33792 34372 39164 34388
rect 33792 34308 39080 34372
rect 39144 34308 39164 34372
rect 33792 34292 39164 34308
rect 33792 34228 39080 34292
rect 39144 34228 39164 34292
rect 33792 34212 39164 34228
rect 33792 34148 39080 34212
rect 39144 34148 39164 34212
rect 33792 34132 39164 34148
rect 33792 34068 39080 34132
rect 39144 34068 39164 34132
rect 33792 34052 39164 34068
rect 33792 33988 39080 34052
rect 39144 33988 39164 34052
rect 33792 33972 39164 33988
rect 33792 33908 39080 33972
rect 39144 33908 39164 33972
rect 33792 33892 39164 33908
rect 33792 33828 39080 33892
rect 39144 33828 39164 33892
rect 33792 33812 39164 33828
rect 33792 33748 39080 33812
rect 39144 33748 39164 33812
rect 33792 33732 39164 33748
rect 33792 33668 39080 33732
rect 39144 33668 39164 33732
rect 33792 33652 39164 33668
rect 33792 33588 39080 33652
rect 39144 33588 39164 33652
rect 33792 33572 39164 33588
rect 33792 33508 39080 33572
rect 39144 33508 39164 33572
rect 33792 33492 39164 33508
rect 33792 33428 39080 33492
rect 39144 33428 39164 33492
rect 33792 33412 39164 33428
rect 33792 33348 39080 33412
rect 39144 33348 39164 33412
rect 33792 33332 39164 33348
rect 33792 33268 39080 33332
rect 39144 33268 39164 33332
rect 33792 33252 39164 33268
rect 33792 33188 39080 33252
rect 39144 33188 39164 33252
rect 33792 33172 39164 33188
rect 33792 33108 39080 33172
rect 39144 33108 39164 33172
rect 33792 33092 39164 33108
rect 33792 33028 39080 33092
rect 39144 33028 39164 33092
rect 33792 33012 39164 33028
rect 33792 32948 39080 33012
rect 39144 32948 39164 33012
rect 33792 32932 39164 32948
rect 33792 32868 39080 32932
rect 39144 32868 39164 32932
rect 33792 32852 39164 32868
rect 33792 32788 39080 32852
rect 39144 32788 39164 32852
rect 33792 32772 39164 32788
rect 33792 32708 39080 32772
rect 39144 32708 39164 32772
rect 33792 32692 39164 32708
rect 33792 32628 39080 32692
rect 39144 32628 39164 32692
rect 33792 32612 39164 32628
rect 33792 32548 39080 32612
rect 39144 32548 39164 32612
rect 33792 32532 39164 32548
rect 33792 32468 39080 32532
rect 39144 32468 39164 32532
rect 33792 32452 39164 32468
rect 33792 32388 39080 32452
rect 39144 32388 39164 32452
rect 33792 32372 39164 32388
rect 33792 32308 39080 32372
rect 39144 32308 39164 32372
rect 33792 32292 39164 32308
rect 33792 32228 39080 32292
rect 39144 32228 39164 32292
rect 33792 32212 39164 32228
rect 33792 32148 39080 32212
rect 39144 32148 39164 32212
rect 33792 32132 39164 32148
rect 33792 32068 39080 32132
rect 39144 32068 39164 32132
rect 33792 32040 39164 32068
rect -39164 31772 -33792 31800
rect -39164 31708 -33876 31772
rect -33812 31708 -33792 31772
rect -39164 31692 -33792 31708
rect -39164 31628 -33876 31692
rect -33812 31628 -33792 31692
rect -39164 31612 -33792 31628
rect -39164 31548 -33876 31612
rect -33812 31548 -33792 31612
rect -39164 31532 -33792 31548
rect -39164 31468 -33876 31532
rect -33812 31468 -33792 31532
rect -39164 31452 -33792 31468
rect -39164 31388 -33876 31452
rect -33812 31388 -33792 31452
rect -39164 31372 -33792 31388
rect -39164 31308 -33876 31372
rect -33812 31308 -33792 31372
rect -39164 31292 -33792 31308
rect -39164 31228 -33876 31292
rect -33812 31228 -33792 31292
rect -39164 31212 -33792 31228
rect -39164 31148 -33876 31212
rect -33812 31148 -33792 31212
rect -39164 31132 -33792 31148
rect -39164 31068 -33876 31132
rect -33812 31068 -33792 31132
rect -39164 31052 -33792 31068
rect -39164 30988 -33876 31052
rect -33812 30988 -33792 31052
rect -39164 30972 -33792 30988
rect -39164 30908 -33876 30972
rect -33812 30908 -33792 30972
rect -39164 30892 -33792 30908
rect -39164 30828 -33876 30892
rect -33812 30828 -33792 30892
rect -39164 30812 -33792 30828
rect -39164 30748 -33876 30812
rect -33812 30748 -33792 30812
rect -39164 30732 -33792 30748
rect -39164 30668 -33876 30732
rect -33812 30668 -33792 30732
rect -39164 30652 -33792 30668
rect -39164 30588 -33876 30652
rect -33812 30588 -33792 30652
rect -39164 30572 -33792 30588
rect -39164 30508 -33876 30572
rect -33812 30508 -33792 30572
rect -39164 30492 -33792 30508
rect -39164 30428 -33876 30492
rect -33812 30428 -33792 30492
rect -39164 30412 -33792 30428
rect -39164 30348 -33876 30412
rect -33812 30348 -33792 30412
rect -39164 30332 -33792 30348
rect -39164 30268 -33876 30332
rect -33812 30268 -33792 30332
rect -39164 30252 -33792 30268
rect -39164 30188 -33876 30252
rect -33812 30188 -33792 30252
rect -39164 30172 -33792 30188
rect -39164 30108 -33876 30172
rect -33812 30108 -33792 30172
rect -39164 30092 -33792 30108
rect -39164 30028 -33876 30092
rect -33812 30028 -33792 30092
rect -39164 30012 -33792 30028
rect -39164 29948 -33876 30012
rect -33812 29948 -33792 30012
rect -39164 29932 -33792 29948
rect -39164 29868 -33876 29932
rect -33812 29868 -33792 29932
rect -39164 29852 -33792 29868
rect -39164 29788 -33876 29852
rect -33812 29788 -33792 29852
rect -39164 29772 -33792 29788
rect -39164 29708 -33876 29772
rect -33812 29708 -33792 29772
rect -39164 29692 -33792 29708
rect -39164 29628 -33876 29692
rect -33812 29628 -33792 29692
rect -39164 29612 -33792 29628
rect -39164 29548 -33876 29612
rect -33812 29548 -33792 29612
rect -39164 29532 -33792 29548
rect -39164 29468 -33876 29532
rect -33812 29468 -33792 29532
rect -39164 29452 -33792 29468
rect -39164 29388 -33876 29452
rect -33812 29388 -33792 29452
rect -39164 29372 -33792 29388
rect -39164 29308 -33876 29372
rect -33812 29308 -33792 29372
rect -39164 29292 -33792 29308
rect -39164 29228 -33876 29292
rect -33812 29228 -33792 29292
rect -39164 29212 -33792 29228
rect -39164 29148 -33876 29212
rect -33812 29148 -33792 29212
rect -39164 29132 -33792 29148
rect -39164 29068 -33876 29132
rect -33812 29068 -33792 29132
rect -39164 29052 -33792 29068
rect -39164 28988 -33876 29052
rect -33812 28988 -33792 29052
rect -39164 28972 -33792 28988
rect -39164 28908 -33876 28972
rect -33812 28908 -33792 28972
rect -39164 28892 -33792 28908
rect -39164 28828 -33876 28892
rect -33812 28828 -33792 28892
rect -39164 28812 -33792 28828
rect -39164 28748 -33876 28812
rect -33812 28748 -33792 28812
rect -39164 28732 -33792 28748
rect -39164 28668 -33876 28732
rect -33812 28668 -33792 28732
rect -39164 28652 -33792 28668
rect -39164 28588 -33876 28652
rect -33812 28588 -33792 28652
rect -39164 28572 -33792 28588
rect -39164 28508 -33876 28572
rect -33812 28508 -33792 28572
rect -39164 28492 -33792 28508
rect -39164 28428 -33876 28492
rect -33812 28428 -33792 28492
rect -39164 28412 -33792 28428
rect -39164 28348 -33876 28412
rect -33812 28348 -33792 28412
rect -39164 28332 -33792 28348
rect -39164 28268 -33876 28332
rect -33812 28268 -33792 28332
rect -39164 28252 -33792 28268
rect -39164 28188 -33876 28252
rect -33812 28188 -33792 28252
rect -39164 28172 -33792 28188
rect -39164 28108 -33876 28172
rect -33812 28108 -33792 28172
rect -39164 28092 -33792 28108
rect -39164 28028 -33876 28092
rect -33812 28028 -33792 28092
rect -39164 28012 -33792 28028
rect -39164 27948 -33876 28012
rect -33812 27948 -33792 28012
rect -39164 27932 -33792 27948
rect -39164 27868 -33876 27932
rect -33812 27868 -33792 27932
rect -39164 27852 -33792 27868
rect -39164 27788 -33876 27852
rect -33812 27788 -33792 27852
rect -39164 27772 -33792 27788
rect -39164 27708 -33876 27772
rect -33812 27708 -33792 27772
rect -39164 27692 -33792 27708
rect -39164 27628 -33876 27692
rect -33812 27628 -33792 27692
rect -39164 27612 -33792 27628
rect -39164 27548 -33876 27612
rect -33812 27548 -33792 27612
rect -39164 27532 -33792 27548
rect -39164 27468 -33876 27532
rect -33812 27468 -33792 27532
rect -39164 27452 -33792 27468
rect -39164 27388 -33876 27452
rect -33812 27388 -33792 27452
rect -39164 27372 -33792 27388
rect -39164 27308 -33876 27372
rect -33812 27308 -33792 27372
rect -39164 27292 -33792 27308
rect -39164 27228 -33876 27292
rect -33812 27228 -33792 27292
rect -39164 27212 -33792 27228
rect -39164 27148 -33876 27212
rect -33812 27148 -33792 27212
rect -39164 27132 -33792 27148
rect -39164 27068 -33876 27132
rect -33812 27068 -33792 27132
rect -39164 27052 -33792 27068
rect -39164 26988 -33876 27052
rect -33812 26988 -33792 27052
rect -39164 26972 -33792 26988
rect -39164 26908 -33876 26972
rect -33812 26908 -33792 26972
rect -39164 26892 -33792 26908
rect -39164 26828 -33876 26892
rect -33812 26828 -33792 26892
rect -39164 26812 -33792 26828
rect -39164 26748 -33876 26812
rect -33812 26748 -33792 26812
rect -39164 26720 -33792 26748
rect -33552 31772 -28180 31800
rect -33552 31708 -28264 31772
rect -28200 31708 -28180 31772
rect -33552 31692 -28180 31708
rect -33552 31628 -28264 31692
rect -28200 31628 -28180 31692
rect -33552 31612 -28180 31628
rect -33552 31548 -28264 31612
rect -28200 31548 -28180 31612
rect -33552 31532 -28180 31548
rect -33552 31468 -28264 31532
rect -28200 31468 -28180 31532
rect -33552 31452 -28180 31468
rect -33552 31388 -28264 31452
rect -28200 31388 -28180 31452
rect -33552 31372 -28180 31388
rect -33552 31308 -28264 31372
rect -28200 31308 -28180 31372
rect -33552 31292 -28180 31308
rect -33552 31228 -28264 31292
rect -28200 31228 -28180 31292
rect -33552 31212 -28180 31228
rect -33552 31148 -28264 31212
rect -28200 31148 -28180 31212
rect -33552 31132 -28180 31148
rect -33552 31068 -28264 31132
rect -28200 31068 -28180 31132
rect -33552 31052 -28180 31068
rect -33552 30988 -28264 31052
rect -28200 30988 -28180 31052
rect -33552 30972 -28180 30988
rect -33552 30908 -28264 30972
rect -28200 30908 -28180 30972
rect -33552 30892 -28180 30908
rect -33552 30828 -28264 30892
rect -28200 30828 -28180 30892
rect -33552 30812 -28180 30828
rect -33552 30748 -28264 30812
rect -28200 30748 -28180 30812
rect -33552 30732 -28180 30748
rect -33552 30668 -28264 30732
rect -28200 30668 -28180 30732
rect -33552 30652 -28180 30668
rect -33552 30588 -28264 30652
rect -28200 30588 -28180 30652
rect -33552 30572 -28180 30588
rect -33552 30508 -28264 30572
rect -28200 30508 -28180 30572
rect -33552 30492 -28180 30508
rect -33552 30428 -28264 30492
rect -28200 30428 -28180 30492
rect -33552 30412 -28180 30428
rect -33552 30348 -28264 30412
rect -28200 30348 -28180 30412
rect -33552 30332 -28180 30348
rect -33552 30268 -28264 30332
rect -28200 30268 -28180 30332
rect -33552 30252 -28180 30268
rect -33552 30188 -28264 30252
rect -28200 30188 -28180 30252
rect -33552 30172 -28180 30188
rect -33552 30108 -28264 30172
rect -28200 30108 -28180 30172
rect -33552 30092 -28180 30108
rect -33552 30028 -28264 30092
rect -28200 30028 -28180 30092
rect -33552 30012 -28180 30028
rect -33552 29948 -28264 30012
rect -28200 29948 -28180 30012
rect -33552 29932 -28180 29948
rect -33552 29868 -28264 29932
rect -28200 29868 -28180 29932
rect -33552 29852 -28180 29868
rect -33552 29788 -28264 29852
rect -28200 29788 -28180 29852
rect -33552 29772 -28180 29788
rect -33552 29708 -28264 29772
rect -28200 29708 -28180 29772
rect -33552 29692 -28180 29708
rect -33552 29628 -28264 29692
rect -28200 29628 -28180 29692
rect -33552 29612 -28180 29628
rect -33552 29548 -28264 29612
rect -28200 29548 -28180 29612
rect -33552 29532 -28180 29548
rect -33552 29468 -28264 29532
rect -28200 29468 -28180 29532
rect -33552 29452 -28180 29468
rect -33552 29388 -28264 29452
rect -28200 29388 -28180 29452
rect -33552 29372 -28180 29388
rect -33552 29308 -28264 29372
rect -28200 29308 -28180 29372
rect -33552 29292 -28180 29308
rect -33552 29228 -28264 29292
rect -28200 29228 -28180 29292
rect -33552 29212 -28180 29228
rect -33552 29148 -28264 29212
rect -28200 29148 -28180 29212
rect -33552 29132 -28180 29148
rect -33552 29068 -28264 29132
rect -28200 29068 -28180 29132
rect -33552 29052 -28180 29068
rect -33552 28988 -28264 29052
rect -28200 28988 -28180 29052
rect -33552 28972 -28180 28988
rect -33552 28908 -28264 28972
rect -28200 28908 -28180 28972
rect -33552 28892 -28180 28908
rect -33552 28828 -28264 28892
rect -28200 28828 -28180 28892
rect -33552 28812 -28180 28828
rect -33552 28748 -28264 28812
rect -28200 28748 -28180 28812
rect -33552 28732 -28180 28748
rect -33552 28668 -28264 28732
rect -28200 28668 -28180 28732
rect -33552 28652 -28180 28668
rect -33552 28588 -28264 28652
rect -28200 28588 -28180 28652
rect -33552 28572 -28180 28588
rect -33552 28508 -28264 28572
rect -28200 28508 -28180 28572
rect -33552 28492 -28180 28508
rect -33552 28428 -28264 28492
rect -28200 28428 -28180 28492
rect -33552 28412 -28180 28428
rect -33552 28348 -28264 28412
rect -28200 28348 -28180 28412
rect -33552 28332 -28180 28348
rect -33552 28268 -28264 28332
rect -28200 28268 -28180 28332
rect -33552 28252 -28180 28268
rect -33552 28188 -28264 28252
rect -28200 28188 -28180 28252
rect -33552 28172 -28180 28188
rect -33552 28108 -28264 28172
rect -28200 28108 -28180 28172
rect -33552 28092 -28180 28108
rect -33552 28028 -28264 28092
rect -28200 28028 -28180 28092
rect -33552 28012 -28180 28028
rect -33552 27948 -28264 28012
rect -28200 27948 -28180 28012
rect -33552 27932 -28180 27948
rect -33552 27868 -28264 27932
rect -28200 27868 -28180 27932
rect -33552 27852 -28180 27868
rect -33552 27788 -28264 27852
rect -28200 27788 -28180 27852
rect -33552 27772 -28180 27788
rect -33552 27708 -28264 27772
rect -28200 27708 -28180 27772
rect -33552 27692 -28180 27708
rect -33552 27628 -28264 27692
rect -28200 27628 -28180 27692
rect -33552 27612 -28180 27628
rect -33552 27548 -28264 27612
rect -28200 27548 -28180 27612
rect -33552 27532 -28180 27548
rect -33552 27468 -28264 27532
rect -28200 27468 -28180 27532
rect -33552 27452 -28180 27468
rect -33552 27388 -28264 27452
rect -28200 27388 -28180 27452
rect -33552 27372 -28180 27388
rect -33552 27308 -28264 27372
rect -28200 27308 -28180 27372
rect -33552 27292 -28180 27308
rect -33552 27228 -28264 27292
rect -28200 27228 -28180 27292
rect -33552 27212 -28180 27228
rect -33552 27148 -28264 27212
rect -28200 27148 -28180 27212
rect -33552 27132 -28180 27148
rect -33552 27068 -28264 27132
rect -28200 27068 -28180 27132
rect -33552 27052 -28180 27068
rect -33552 26988 -28264 27052
rect -28200 26988 -28180 27052
rect -33552 26972 -28180 26988
rect -33552 26908 -28264 26972
rect -28200 26908 -28180 26972
rect -33552 26892 -28180 26908
rect -33552 26828 -28264 26892
rect -28200 26828 -28180 26892
rect -33552 26812 -28180 26828
rect -33552 26748 -28264 26812
rect -28200 26748 -28180 26812
rect -33552 26720 -28180 26748
rect -27940 31772 -22568 31800
rect -27940 31708 -22652 31772
rect -22588 31708 -22568 31772
rect -27940 31692 -22568 31708
rect -27940 31628 -22652 31692
rect -22588 31628 -22568 31692
rect -27940 31612 -22568 31628
rect -27940 31548 -22652 31612
rect -22588 31548 -22568 31612
rect -27940 31532 -22568 31548
rect -27940 31468 -22652 31532
rect -22588 31468 -22568 31532
rect -27940 31452 -22568 31468
rect -27940 31388 -22652 31452
rect -22588 31388 -22568 31452
rect -27940 31372 -22568 31388
rect -27940 31308 -22652 31372
rect -22588 31308 -22568 31372
rect -27940 31292 -22568 31308
rect -27940 31228 -22652 31292
rect -22588 31228 -22568 31292
rect -27940 31212 -22568 31228
rect -27940 31148 -22652 31212
rect -22588 31148 -22568 31212
rect -27940 31132 -22568 31148
rect -27940 31068 -22652 31132
rect -22588 31068 -22568 31132
rect -27940 31052 -22568 31068
rect -27940 30988 -22652 31052
rect -22588 30988 -22568 31052
rect -27940 30972 -22568 30988
rect -27940 30908 -22652 30972
rect -22588 30908 -22568 30972
rect -27940 30892 -22568 30908
rect -27940 30828 -22652 30892
rect -22588 30828 -22568 30892
rect -27940 30812 -22568 30828
rect -27940 30748 -22652 30812
rect -22588 30748 -22568 30812
rect -27940 30732 -22568 30748
rect -27940 30668 -22652 30732
rect -22588 30668 -22568 30732
rect -27940 30652 -22568 30668
rect -27940 30588 -22652 30652
rect -22588 30588 -22568 30652
rect -27940 30572 -22568 30588
rect -27940 30508 -22652 30572
rect -22588 30508 -22568 30572
rect -27940 30492 -22568 30508
rect -27940 30428 -22652 30492
rect -22588 30428 -22568 30492
rect -27940 30412 -22568 30428
rect -27940 30348 -22652 30412
rect -22588 30348 -22568 30412
rect -27940 30332 -22568 30348
rect -27940 30268 -22652 30332
rect -22588 30268 -22568 30332
rect -27940 30252 -22568 30268
rect -27940 30188 -22652 30252
rect -22588 30188 -22568 30252
rect -27940 30172 -22568 30188
rect -27940 30108 -22652 30172
rect -22588 30108 -22568 30172
rect -27940 30092 -22568 30108
rect -27940 30028 -22652 30092
rect -22588 30028 -22568 30092
rect -27940 30012 -22568 30028
rect -27940 29948 -22652 30012
rect -22588 29948 -22568 30012
rect -27940 29932 -22568 29948
rect -27940 29868 -22652 29932
rect -22588 29868 -22568 29932
rect -27940 29852 -22568 29868
rect -27940 29788 -22652 29852
rect -22588 29788 -22568 29852
rect -27940 29772 -22568 29788
rect -27940 29708 -22652 29772
rect -22588 29708 -22568 29772
rect -27940 29692 -22568 29708
rect -27940 29628 -22652 29692
rect -22588 29628 -22568 29692
rect -27940 29612 -22568 29628
rect -27940 29548 -22652 29612
rect -22588 29548 -22568 29612
rect -27940 29532 -22568 29548
rect -27940 29468 -22652 29532
rect -22588 29468 -22568 29532
rect -27940 29452 -22568 29468
rect -27940 29388 -22652 29452
rect -22588 29388 -22568 29452
rect -27940 29372 -22568 29388
rect -27940 29308 -22652 29372
rect -22588 29308 -22568 29372
rect -27940 29292 -22568 29308
rect -27940 29228 -22652 29292
rect -22588 29228 -22568 29292
rect -27940 29212 -22568 29228
rect -27940 29148 -22652 29212
rect -22588 29148 -22568 29212
rect -27940 29132 -22568 29148
rect -27940 29068 -22652 29132
rect -22588 29068 -22568 29132
rect -27940 29052 -22568 29068
rect -27940 28988 -22652 29052
rect -22588 28988 -22568 29052
rect -27940 28972 -22568 28988
rect -27940 28908 -22652 28972
rect -22588 28908 -22568 28972
rect -27940 28892 -22568 28908
rect -27940 28828 -22652 28892
rect -22588 28828 -22568 28892
rect -27940 28812 -22568 28828
rect -27940 28748 -22652 28812
rect -22588 28748 -22568 28812
rect -27940 28732 -22568 28748
rect -27940 28668 -22652 28732
rect -22588 28668 -22568 28732
rect -27940 28652 -22568 28668
rect -27940 28588 -22652 28652
rect -22588 28588 -22568 28652
rect -27940 28572 -22568 28588
rect -27940 28508 -22652 28572
rect -22588 28508 -22568 28572
rect -27940 28492 -22568 28508
rect -27940 28428 -22652 28492
rect -22588 28428 -22568 28492
rect -27940 28412 -22568 28428
rect -27940 28348 -22652 28412
rect -22588 28348 -22568 28412
rect -27940 28332 -22568 28348
rect -27940 28268 -22652 28332
rect -22588 28268 -22568 28332
rect -27940 28252 -22568 28268
rect -27940 28188 -22652 28252
rect -22588 28188 -22568 28252
rect -27940 28172 -22568 28188
rect -27940 28108 -22652 28172
rect -22588 28108 -22568 28172
rect -27940 28092 -22568 28108
rect -27940 28028 -22652 28092
rect -22588 28028 -22568 28092
rect -27940 28012 -22568 28028
rect -27940 27948 -22652 28012
rect -22588 27948 -22568 28012
rect -27940 27932 -22568 27948
rect -27940 27868 -22652 27932
rect -22588 27868 -22568 27932
rect -27940 27852 -22568 27868
rect -27940 27788 -22652 27852
rect -22588 27788 -22568 27852
rect -27940 27772 -22568 27788
rect -27940 27708 -22652 27772
rect -22588 27708 -22568 27772
rect -27940 27692 -22568 27708
rect -27940 27628 -22652 27692
rect -22588 27628 -22568 27692
rect -27940 27612 -22568 27628
rect -27940 27548 -22652 27612
rect -22588 27548 -22568 27612
rect -27940 27532 -22568 27548
rect -27940 27468 -22652 27532
rect -22588 27468 -22568 27532
rect -27940 27452 -22568 27468
rect -27940 27388 -22652 27452
rect -22588 27388 -22568 27452
rect -27940 27372 -22568 27388
rect -27940 27308 -22652 27372
rect -22588 27308 -22568 27372
rect -27940 27292 -22568 27308
rect -27940 27228 -22652 27292
rect -22588 27228 -22568 27292
rect -27940 27212 -22568 27228
rect -27940 27148 -22652 27212
rect -22588 27148 -22568 27212
rect -27940 27132 -22568 27148
rect -27940 27068 -22652 27132
rect -22588 27068 -22568 27132
rect -27940 27052 -22568 27068
rect -27940 26988 -22652 27052
rect -22588 26988 -22568 27052
rect -27940 26972 -22568 26988
rect -27940 26908 -22652 26972
rect -22588 26908 -22568 26972
rect -27940 26892 -22568 26908
rect -27940 26828 -22652 26892
rect -22588 26828 -22568 26892
rect -27940 26812 -22568 26828
rect -27940 26748 -22652 26812
rect -22588 26748 -22568 26812
rect -27940 26720 -22568 26748
rect -22328 31772 -16956 31800
rect -22328 31708 -17040 31772
rect -16976 31708 -16956 31772
rect -22328 31692 -16956 31708
rect -22328 31628 -17040 31692
rect -16976 31628 -16956 31692
rect -22328 31612 -16956 31628
rect -22328 31548 -17040 31612
rect -16976 31548 -16956 31612
rect -22328 31532 -16956 31548
rect -22328 31468 -17040 31532
rect -16976 31468 -16956 31532
rect -22328 31452 -16956 31468
rect -22328 31388 -17040 31452
rect -16976 31388 -16956 31452
rect -22328 31372 -16956 31388
rect -22328 31308 -17040 31372
rect -16976 31308 -16956 31372
rect -22328 31292 -16956 31308
rect -22328 31228 -17040 31292
rect -16976 31228 -16956 31292
rect -22328 31212 -16956 31228
rect -22328 31148 -17040 31212
rect -16976 31148 -16956 31212
rect -22328 31132 -16956 31148
rect -22328 31068 -17040 31132
rect -16976 31068 -16956 31132
rect -22328 31052 -16956 31068
rect -22328 30988 -17040 31052
rect -16976 30988 -16956 31052
rect -22328 30972 -16956 30988
rect -22328 30908 -17040 30972
rect -16976 30908 -16956 30972
rect -22328 30892 -16956 30908
rect -22328 30828 -17040 30892
rect -16976 30828 -16956 30892
rect -22328 30812 -16956 30828
rect -22328 30748 -17040 30812
rect -16976 30748 -16956 30812
rect -22328 30732 -16956 30748
rect -22328 30668 -17040 30732
rect -16976 30668 -16956 30732
rect -22328 30652 -16956 30668
rect -22328 30588 -17040 30652
rect -16976 30588 -16956 30652
rect -22328 30572 -16956 30588
rect -22328 30508 -17040 30572
rect -16976 30508 -16956 30572
rect -22328 30492 -16956 30508
rect -22328 30428 -17040 30492
rect -16976 30428 -16956 30492
rect -22328 30412 -16956 30428
rect -22328 30348 -17040 30412
rect -16976 30348 -16956 30412
rect -22328 30332 -16956 30348
rect -22328 30268 -17040 30332
rect -16976 30268 -16956 30332
rect -22328 30252 -16956 30268
rect -22328 30188 -17040 30252
rect -16976 30188 -16956 30252
rect -22328 30172 -16956 30188
rect -22328 30108 -17040 30172
rect -16976 30108 -16956 30172
rect -22328 30092 -16956 30108
rect -22328 30028 -17040 30092
rect -16976 30028 -16956 30092
rect -22328 30012 -16956 30028
rect -22328 29948 -17040 30012
rect -16976 29948 -16956 30012
rect -22328 29932 -16956 29948
rect -22328 29868 -17040 29932
rect -16976 29868 -16956 29932
rect -22328 29852 -16956 29868
rect -22328 29788 -17040 29852
rect -16976 29788 -16956 29852
rect -22328 29772 -16956 29788
rect -22328 29708 -17040 29772
rect -16976 29708 -16956 29772
rect -22328 29692 -16956 29708
rect -22328 29628 -17040 29692
rect -16976 29628 -16956 29692
rect -22328 29612 -16956 29628
rect -22328 29548 -17040 29612
rect -16976 29548 -16956 29612
rect -22328 29532 -16956 29548
rect -22328 29468 -17040 29532
rect -16976 29468 -16956 29532
rect -22328 29452 -16956 29468
rect -22328 29388 -17040 29452
rect -16976 29388 -16956 29452
rect -22328 29372 -16956 29388
rect -22328 29308 -17040 29372
rect -16976 29308 -16956 29372
rect -22328 29292 -16956 29308
rect -22328 29228 -17040 29292
rect -16976 29228 -16956 29292
rect -22328 29212 -16956 29228
rect -22328 29148 -17040 29212
rect -16976 29148 -16956 29212
rect -22328 29132 -16956 29148
rect -22328 29068 -17040 29132
rect -16976 29068 -16956 29132
rect -22328 29052 -16956 29068
rect -22328 28988 -17040 29052
rect -16976 28988 -16956 29052
rect -22328 28972 -16956 28988
rect -22328 28908 -17040 28972
rect -16976 28908 -16956 28972
rect -22328 28892 -16956 28908
rect -22328 28828 -17040 28892
rect -16976 28828 -16956 28892
rect -22328 28812 -16956 28828
rect -22328 28748 -17040 28812
rect -16976 28748 -16956 28812
rect -22328 28732 -16956 28748
rect -22328 28668 -17040 28732
rect -16976 28668 -16956 28732
rect -22328 28652 -16956 28668
rect -22328 28588 -17040 28652
rect -16976 28588 -16956 28652
rect -22328 28572 -16956 28588
rect -22328 28508 -17040 28572
rect -16976 28508 -16956 28572
rect -22328 28492 -16956 28508
rect -22328 28428 -17040 28492
rect -16976 28428 -16956 28492
rect -22328 28412 -16956 28428
rect -22328 28348 -17040 28412
rect -16976 28348 -16956 28412
rect -22328 28332 -16956 28348
rect -22328 28268 -17040 28332
rect -16976 28268 -16956 28332
rect -22328 28252 -16956 28268
rect -22328 28188 -17040 28252
rect -16976 28188 -16956 28252
rect -22328 28172 -16956 28188
rect -22328 28108 -17040 28172
rect -16976 28108 -16956 28172
rect -22328 28092 -16956 28108
rect -22328 28028 -17040 28092
rect -16976 28028 -16956 28092
rect -22328 28012 -16956 28028
rect -22328 27948 -17040 28012
rect -16976 27948 -16956 28012
rect -22328 27932 -16956 27948
rect -22328 27868 -17040 27932
rect -16976 27868 -16956 27932
rect -22328 27852 -16956 27868
rect -22328 27788 -17040 27852
rect -16976 27788 -16956 27852
rect -22328 27772 -16956 27788
rect -22328 27708 -17040 27772
rect -16976 27708 -16956 27772
rect -22328 27692 -16956 27708
rect -22328 27628 -17040 27692
rect -16976 27628 -16956 27692
rect -22328 27612 -16956 27628
rect -22328 27548 -17040 27612
rect -16976 27548 -16956 27612
rect -22328 27532 -16956 27548
rect -22328 27468 -17040 27532
rect -16976 27468 -16956 27532
rect -22328 27452 -16956 27468
rect -22328 27388 -17040 27452
rect -16976 27388 -16956 27452
rect -22328 27372 -16956 27388
rect -22328 27308 -17040 27372
rect -16976 27308 -16956 27372
rect -22328 27292 -16956 27308
rect -22328 27228 -17040 27292
rect -16976 27228 -16956 27292
rect -22328 27212 -16956 27228
rect -22328 27148 -17040 27212
rect -16976 27148 -16956 27212
rect -22328 27132 -16956 27148
rect -22328 27068 -17040 27132
rect -16976 27068 -16956 27132
rect -22328 27052 -16956 27068
rect -22328 26988 -17040 27052
rect -16976 26988 -16956 27052
rect -22328 26972 -16956 26988
rect -22328 26908 -17040 26972
rect -16976 26908 -16956 26972
rect -22328 26892 -16956 26908
rect -22328 26828 -17040 26892
rect -16976 26828 -16956 26892
rect -22328 26812 -16956 26828
rect -22328 26748 -17040 26812
rect -16976 26748 -16956 26812
rect -22328 26720 -16956 26748
rect -16716 31772 -11344 31800
rect -16716 31708 -11428 31772
rect -11364 31708 -11344 31772
rect -16716 31692 -11344 31708
rect -16716 31628 -11428 31692
rect -11364 31628 -11344 31692
rect -16716 31612 -11344 31628
rect -16716 31548 -11428 31612
rect -11364 31548 -11344 31612
rect -16716 31532 -11344 31548
rect -16716 31468 -11428 31532
rect -11364 31468 -11344 31532
rect -16716 31452 -11344 31468
rect -16716 31388 -11428 31452
rect -11364 31388 -11344 31452
rect -16716 31372 -11344 31388
rect -16716 31308 -11428 31372
rect -11364 31308 -11344 31372
rect -16716 31292 -11344 31308
rect -16716 31228 -11428 31292
rect -11364 31228 -11344 31292
rect -16716 31212 -11344 31228
rect -16716 31148 -11428 31212
rect -11364 31148 -11344 31212
rect -16716 31132 -11344 31148
rect -16716 31068 -11428 31132
rect -11364 31068 -11344 31132
rect -16716 31052 -11344 31068
rect -16716 30988 -11428 31052
rect -11364 30988 -11344 31052
rect -16716 30972 -11344 30988
rect -16716 30908 -11428 30972
rect -11364 30908 -11344 30972
rect -16716 30892 -11344 30908
rect -16716 30828 -11428 30892
rect -11364 30828 -11344 30892
rect -16716 30812 -11344 30828
rect -16716 30748 -11428 30812
rect -11364 30748 -11344 30812
rect -16716 30732 -11344 30748
rect -16716 30668 -11428 30732
rect -11364 30668 -11344 30732
rect -16716 30652 -11344 30668
rect -16716 30588 -11428 30652
rect -11364 30588 -11344 30652
rect -16716 30572 -11344 30588
rect -16716 30508 -11428 30572
rect -11364 30508 -11344 30572
rect -16716 30492 -11344 30508
rect -16716 30428 -11428 30492
rect -11364 30428 -11344 30492
rect -16716 30412 -11344 30428
rect -16716 30348 -11428 30412
rect -11364 30348 -11344 30412
rect -16716 30332 -11344 30348
rect -16716 30268 -11428 30332
rect -11364 30268 -11344 30332
rect -16716 30252 -11344 30268
rect -16716 30188 -11428 30252
rect -11364 30188 -11344 30252
rect -16716 30172 -11344 30188
rect -16716 30108 -11428 30172
rect -11364 30108 -11344 30172
rect -16716 30092 -11344 30108
rect -16716 30028 -11428 30092
rect -11364 30028 -11344 30092
rect -16716 30012 -11344 30028
rect -16716 29948 -11428 30012
rect -11364 29948 -11344 30012
rect -16716 29932 -11344 29948
rect -16716 29868 -11428 29932
rect -11364 29868 -11344 29932
rect -16716 29852 -11344 29868
rect -16716 29788 -11428 29852
rect -11364 29788 -11344 29852
rect -16716 29772 -11344 29788
rect -16716 29708 -11428 29772
rect -11364 29708 -11344 29772
rect -16716 29692 -11344 29708
rect -16716 29628 -11428 29692
rect -11364 29628 -11344 29692
rect -16716 29612 -11344 29628
rect -16716 29548 -11428 29612
rect -11364 29548 -11344 29612
rect -16716 29532 -11344 29548
rect -16716 29468 -11428 29532
rect -11364 29468 -11344 29532
rect -16716 29452 -11344 29468
rect -16716 29388 -11428 29452
rect -11364 29388 -11344 29452
rect -16716 29372 -11344 29388
rect -16716 29308 -11428 29372
rect -11364 29308 -11344 29372
rect -16716 29292 -11344 29308
rect -16716 29228 -11428 29292
rect -11364 29228 -11344 29292
rect -16716 29212 -11344 29228
rect -16716 29148 -11428 29212
rect -11364 29148 -11344 29212
rect -16716 29132 -11344 29148
rect -16716 29068 -11428 29132
rect -11364 29068 -11344 29132
rect -16716 29052 -11344 29068
rect -16716 28988 -11428 29052
rect -11364 28988 -11344 29052
rect -16716 28972 -11344 28988
rect -16716 28908 -11428 28972
rect -11364 28908 -11344 28972
rect -16716 28892 -11344 28908
rect -16716 28828 -11428 28892
rect -11364 28828 -11344 28892
rect -16716 28812 -11344 28828
rect -16716 28748 -11428 28812
rect -11364 28748 -11344 28812
rect -16716 28732 -11344 28748
rect -16716 28668 -11428 28732
rect -11364 28668 -11344 28732
rect -16716 28652 -11344 28668
rect -16716 28588 -11428 28652
rect -11364 28588 -11344 28652
rect -16716 28572 -11344 28588
rect -16716 28508 -11428 28572
rect -11364 28508 -11344 28572
rect -16716 28492 -11344 28508
rect -16716 28428 -11428 28492
rect -11364 28428 -11344 28492
rect -16716 28412 -11344 28428
rect -16716 28348 -11428 28412
rect -11364 28348 -11344 28412
rect -16716 28332 -11344 28348
rect -16716 28268 -11428 28332
rect -11364 28268 -11344 28332
rect -16716 28252 -11344 28268
rect -16716 28188 -11428 28252
rect -11364 28188 -11344 28252
rect -16716 28172 -11344 28188
rect -16716 28108 -11428 28172
rect -11364 28108 -11344 28172
rect -16716 28092 -11344 28108
rect -16716 28028 -11428 28092
rect -11364 28028 -11344 28092
rect -16716 28012 -11344 28028
rect -16716 27948 -11428 28012
rect -11364 27948 -11344 28012
rect -16716 27932 -11344 27948
rect -16716 27868 -11428 27932
rect -11364 27868 -11344 27932
rect -16716 27852 -11344 27868
rect -16716 27788 -11428 27852
rect -11364 27788 -11344 27852
rect -16716 27772 -11344 27788
rect -16716 27708 -11428 27772
rect -11364 27708 -11344 27772
rect -16716 27692 -11344 27708
rect -16716 27628 -11428 27692
rect -11364 27628 -11344 27692
rect -16716 27612 -11344 27628
rect -16716 27548 -11428 27612
rect -11364 27548 -11344 27612
rect -16716 27532 -11344 27548
rect -16716 27468 -11428 27532
rect -11364 27468 -11344 27532
rect -16716 27452 -11344 27468
rect -16716 27388 -11428 27452
rect -11364 27388 -11344 27452
rect -16716 27372 -11344 27388
rect -16716 27308 -11428 27372
rect -11364 27308 -11344 27372
rect -16716 27292 -11344 27308
rect -16716 27228 -11428 27292
rect -11364 27228 -11344 27292
rect -16716 27212 -11344 27228
rect -16716 27148 -11428 27212
rect -11364 27148 -11344 27212
rect -16716 27132 -11344 27148
rect -16716 27068 -11428 27132
rect -11364 27068 -11344 27132
rect -16716 27052 -11344 27068
rect -16716 26988 -11428 27052
rect -11364 26988 -11344 27052
rect -16716 26972 -11344 26988
rect -16716 26908 -11428 26972
rect -11364 26908 -11344 26972
rect -16716 26892 -11344 26908
rect -16716 26828 -11428 26892
rect -11364 26828 -11344 26892
rect -16716 26812 -11344 26828
rect -16716 26748 -11428 26812
rect -11364 26748 -11344 26812
rect -16716 26720 -11344 26748
rect -11104 31772 -5732 31800
rect -11104 31708 -5816 31772
rect -5752 31708 -5732 31772
rect -11104 31692 -5732 31708
rect -11104 31628 -5816 31692
rect -5752 31628 -5732 31692
rect -11104 31612 -5732 31628
rect -11104 31548 -5816 31612
rect -5752 31548 -5732 31612
rect -11104 31532 -5732 31548
rect -11104 31468 -5816 31532
rect -5752 31468 -5732 31532
rect -11104 31452 -5732 31468
rect -11104 31388 -5816 31452
rect -5752 31388 -5732 31452
rect -11104 31372 -5732 31388
rect -11104 31308 -5816 31372
rect -5752 31308 -5732 31372
rect -11104 31292 -5732 31308
rect -11104 31228 -5816 31292
rect -5752 31228 -5732 31292
rect -11104 31212 -5732 31228
rect -11104 31148 -5816 31212
rect -5752 31148 -5732 31212
rect -11104 31132 -5732 31148
rect -11104 31068 -5816 31132
rect -5752 31068 -5732 31132
rect -11104 31052 -5732 31068
rect -11104 30988 -5816 31052
rect -5752 30988 -5732 31052
rect -11104 30972 -5732 30988
rect -11104 30908 -5816 30972
rect -5752 30908 -5732 30972
rect -11104 30892 -5732 30908
rect -11104 30828 -5816 30892
rect -5752 30828 -5732 30892
rect -11104 30812 -5732 30828
rect -11104 30748 -5816 30812
rect -5752 30748 -5732 30812
rect -11104 30732 -5732 30748
rect -11104 30668 -5816 30732
rect -5752 30668 -5732 30732
rect -11104 30652 -5732 30668
rect -11104 30588 -5816 30652
rect -5752 30588 -5732 30652
rect -11104 30572 -5732 30588
rect -11104 30508 -5816 30572
rect -5752 30508 -5732 30572
rect -11104 30492 -5732 30508
rect -11104 30428 -5816 30492
rect -5752 30428 -5732 30492
rect -11104 30412 -5732 30428
rect -11104 30348 -5816 30412
rect -5752 30348 -5732 30412
rect -11104 30332 -5732 30348
rect -11104 30268 -5816 30332
rect -5752 30268 -5732 30332
rect -11104 30252 -5732 30268
rect -11104 30188 -5816 30252
rect -5752 30188 -5732 30252
rect -11104 30172 -5732 30188
rect -11104 30108 -5816 30172
rect -5752 30108 -5732 30172
rect -11104 30092 -5732 30108
rect -11104 30028 -5816 30092
rect -5752 30028 -5732 30092
rect -11104 30012 -5732 30028
rect -11104 29948 -5816 30012
rect -5752 29948 -5732 30012
rect -11104 29932 -5732 29948
rect -11104 29868 -5816 29932
rect -5752 29868 -5732 29932
rect -11104 29852 -5732 29868
rect -11104 29788 -5816 29852
rect -5752 29788 -5732 29852
rect -11104 29772 -5732 29788
rect -11104 29708 -5816 29772
rect -5752 29708 -5732 29772
rect -11104 29692 -5732 29708
rect -11104 29628 -5816 29692
rect -5752 29628 -5732 29692
rect -11104 29612 -5732 29628
rect -11104 29548 -5816 29612
rect -5752 29548 -5732 29612
rect -11104 29532 -5732 29548
rect -11104 29468 -5816 29532
rect -5752 29468 -5732 29532
rect -11104 29452 -5732 29468
rect -11104 29388 -5816 29452
rect -5752 29388 -5732 29452
rect -11104 29372 -5732 29388
rect -11104 29308 -5816 29372
rect -5752 29308 -5732 29372
rect -11104 29292 -5732 29308
rect -11104 29228 -5816 29292
rect -5752 29228 -5732 29292
rect -11104 29212 -5732 29228
rect -11104 29148 -5816 29212
rect -5752 29148 -5732 29212
rect -11104 29132 -5732 29148
rect -11104 29068 -5816 29132
rect -5752 29068 -5732 29132
rect -11104 29052 -5732 29068
rect -11104 28988 -5816 29052
rect -5752 28988 -5732 29052
rect -11104 28972 -5732 28988
rect -11104 28908 -5816 28972
rect -5752 28908 -5732 28972
rect -11104 28892 -5732 28908
rect -11104 28828 -5816 28892
rect -5752 28828 -5732 28892
rect -11104 28812 -5732 28828
rect -11104 28748 -5816 28812
rect -5752 28748 -5732 28812
rect -11104 28732 -5732 28748
rect -11104 28668 -5816 28732
rect -5752 28668 -5732 28732
rect -11104 28652 -5732 28668
rect -11104 28588 -5816 28652
rect -5752 28588 -5732 28652
rect -11104 28572 -5732 28588
rect -11104 28508 -5816 28572
rect -5752 28508 -5732 28572
rect -11104 28492 -5732 28508
rect -11104 28428 -5816 28492
rect -5752 28428 -5732 28492
rect -11104 28412 -5732 28428
rect -11104 28348 -5816 28412
rect -5752 28348 -5732 28412
rect -11104 28332 -5732 28348
rect -11104 28268 -5816 28332
rect -5752 28268 -5732 28332
rect -11104 28252 -5732 28268
rect -11104 28188 -5816 28252
rect -5752 28188 -5732 28252
rect -11104 28172 -5732 28188
rect -11104 28108 -5816 28172
rect -5752 28108 -5732 28172
rect -11104 28092 -5732 28108
rect -11104 28028 -5816 28092
rect -5752 28028 -5732 28092
rect -11104 28012 -5732 28028
rect -11104 27948 -5816 28012
rect -5752 27948 -5732 28012
rect -11104 27932 -5732 27948
rect -11104 27868 -5816 27932
rect -5752 27868 -5732 27932
rect -11104 27852 -5732 27868
rect -11104 27788 -5816 27852
rect -5752 27788 -5732 27852
rect -11104 27772 -5732 27788
rect -11104 27708 -5816 27772
rect -5752 27708 -5732 27772
rect -11104 27692 -5732 27708
rect -11104 27628 -5816 27692
rect -5752 27628 -5732 27692
rect -11104 27612 -5732 27628
rect -11104 27548 -5816 27612
rect -5752 27548 -5732 27612
rect -11104 27532 -5732 27548
rect -11104 27468 -5816 27532
rect -5752 27468 -5732 27532
rect -11104 27452 -5732 27468
rect -11104 27388 -5816 27452
rect -5752 27388 -5732 27452
rect -11104 27372 -5732 27388
rect -11104 27308 -5816 27372
rect -5752 27308 -5732 27372
rect -11104 27292 -5732 27308
rect -11104 27228 -5816 27292
rect -5752 27228 -5732 27292
rect -11104 27212 -5732 27228
rect -11104 27148 -5816 27212
rect -5752 27148 -5732 27212
rect -11104 27132 -5732 27148
rect -11104 27068 -5816 27132
rect -5752 27068 -5732 27132
rect -11104 27052 -5732 27068
rect -11104 26988 -5816 27052
rect -5752 26988 -5732 27052
rect -11104 26972 -5732 26988
rect -11104 26908 -5816 26972
rect -5752 26908 -5732 26972
rect -11104 26892 -5732 26908
rect -11104 26828 -5816 26892
rect -5752 26828 -5732 26892
rect -11104 26812 -5732 26828
rect -11104 26748 -5816 26812
rect -5752 26748 -5732 26812
rect -11104 26720 -5732 26748
rect -5492 31772 -120 31800
rect -5492 31708 -204 31772
rect -140 31708 -120 31772
rect -5492 31692 -120 31708
rect -5492 31628 -204 31692
rect -140 31628 -120 31692
rect -5492 31612 -120 31628
rect -5492 31548 -204 31612
rect -140 31548 -120 31612
rect -5492 31532 -120 31548
rect -5492 31468 -204 31532
rect -140 31468 -120 31532
rect -5492 31452 -120 31468
rect -5492 31388 -204 31452
rect -140 31388 -120 31452
rect -5492 31372 -120 31388
rect -5492 31308 -204 31372
rect -140 31308 -120 31372
rect -5492 31292 -120 31308
rect -5492 31228 -204 31292
rect -140 31228 -120 31292
rect -5492 31212 -120 31228
rect -5492 31148 -204 31212
rect -140 31148 -120 31212
rect -5492 31132 -120 31148
rect -5492 31068 -204 31132
rect -140 31068 -120 31132
rect -5492 31052 -120 31068
rect -5492 30988 -204 31052
rect -140 30988 -120 31052
rect -5492 30972 -120 30988
rect -5492 30908 -204 30972
rect -140 30908 -120 30972
rect -5492 30892 -120 30908
rect -5492 30828 -204 30892
rect -140 30828 -120 30892
rect -5492 30812 -120 30828
rect -5492 30748 -204 30812
rect -140 30748 -120 30812
rect -5492 30732 -120 30748
rect -5492 30668 -204 30732
rect -140 30668 -120 30732
rect -5492 30652 -120 30668
rect -5492 30588 -204 30652
rect -140 30588 -120 30652
rect -5492 30572 -120 30588
rect -5492 30508 -204 30572
rect -140 30508 -120 30572
rect -5492 30492 -120 30508
rect -5492 30428 -204 30492
rect -140 30428 -120 30492
rect -5492 30412 -120 30428
rect -5492 30348 -204 30412
rect -140 30348 -120 30412
rect -5492 30332 -120 30348
rect -5492 30268 -204 30332
rect -140 30268 -120 30332
rect -5492 30252 -120 30268
rect -5492 30188 -204 30252
rect -140 30188 -120 30252
rect -5492 30172 -120 30188
rect -5492 30108 -204 30172
rect -140 30108 -120 30172
rect -5492 30092 -120 30108
rect -5492 30028 -204 30092
rect -140 30028 -120 30092
rect -5492 30012 -120 30028
rect -5492 29948 -204 30012
rect -140 29948 -120 30012
rect -5492 29932 -120 29948
rect -5492 29868 -204 29932
rect -140 29868 -120 29932
rect -5492 29852 -120 29868
rect -5492 29788 -204 29852
rect -140 29788 -120 29852
rect -5492 29772 -120 29788
rect -5492 29708 -204 29772
rect -140 29708 -120 29772
rect -5492 29692 -120 29708
rect -5492 29628 -204 29692
rect -140 29628 -120 29692
rect -5492 29612 -120 29628
rect -5492 29548 -204 29612
rect -140 29548 -120 29612
rect -5492 29532 -120 29548
rect -5492 29468 -204 29532
rect -140 29468 -120 29532
rect -5492 29452 -120 29468
rect -5492 29388 -204 29452
rect -140 29388 -120 29452
rect -5492 29372 -120 29388
rect -5492 29308 -204 29372
rect -140 29308 -120 29372
rect -5492 29292 -120 29308
rect -5492 29228 -204 29292
rect -140 29228 -120 29292
rect -5492 29212 -120 29228
rect -5492 29148 -204 29212
rect -140 29148 -120 29212
rect -5492 29132 -120 29148
rect -5492 29068 -204 29132
rect -140 29068 -120 29132
rect -5492 29052 -120 29068
rect -5492 28988 -204 29052
rect -140 28988 -120 29052
rect -5492 28972 -120 28988
rect -5492 28908 -204 28972
rect -140 28908 -120 28972
rect -5492 28892 -120 28908
rect -5492 28828 -204 28892
rect -140 28828 -120 28892
rect -5492 28812 -120 28828
rect -5492 28748 -204 28812
rect -140 28748 -120 28812
rect -5492 28732 -120 28748
rect -5492 28668 -204 28732
rect -140 28668 -120 28732
rect -5492 28652 -120 28668
rect -5492 28588 -204 28652
rect -140 28588 -120 28652
rect -5492 28572 -120 28588
rect -5492 28508 -204 28572
rect -140 28508 -120 28572
rect -5492 28492 -120 28508
rect -5492 28428 -204 28492
rect -140 28428 -120 28492
rect -5492 28412 -120 28428
rect -5492 28348 -204 28412
rect -140 28348 -120 28412
rect -5492 28332 -120 28348
rect -5492 28268 -204 28332
rect -140 28268 -120 28332
rect -5492 28252 -120 28268
rect -5492 28188 -204 28252
rect -140 28188 -120 28252
rect -5492 28172 -120 28188
rect -5492 28108 -204 28172
rect -140 28108 -120 28172
rect -5492 28092 -120 28108
rect -5492 28028 -204 28092
rect -140 28028 -120 28092
rect -5492 28012 -120 28028
rect -5492 27948 -204 28012
rect -140 27948 -120 28012
rect -5492 27932 -120 27948
rect -5492 27868 -204 27932
rect -140 27868 -120 27932
rect -5492 27852 -120 27868
rect -5492 27788 -204 27852
rect -140 27788 -120 27852
rect -5492 27772 -120 27788
rect -5492 27708 -204 27772
rect -140 27708 -120 27772
rect -5492 27692 -120 27708
rect -5492 27628 -204 27692
rect -140 27628 -120 27692
rect -5492 27612 -120 27628
rect -5492 27548 -204 27612
rect -140 27548 -120 27612
rect -5492 27532 -120 27548
rect -5492 27468 -204 27532
rect -140 27468 -120 27532
rect -5492 27452 -120 27468
rect -5492 27388 -204 27452
rect -140 27388 -120 27452
rect -5492 27372 -120 27388
rect -5492 27308 -204 27372
rect -140 27308 -120 27372
rect -5492 27292 -120 27308
rect -5492 27228 -204 27292
rect -140 27228 -120 27292
rect -5492 27212 -120 27228
rect -5492 27148 -204 27212
rect -140 27148 -120 27212
rect -5492 27132 -120 27148
rect -5492 27068 -204 27132
rect -140 27068 -120 27132
rect -5492 27052 -120 27068
rect -5492 26988 -204 27052
rect -140 26988 -120 27052
rect -5492 26972 -120 26988
rect -5492 26908 -204 26972
rect -140 26908 -120 26972
rect -5492 26892 -120 26908
rect -5492 26828 -204 26892
rect -140 26828 -120 26892
rect -5492 26812 -120 26828
rect -5492 26748 -204 26812
rect -140 26748 -120 26812
rect -5492 26720 -120 26748
rect 120 31772 5492 31800
rect 120 31708 5408 31772
rect 5472 31708 5492 31772
rect 120 31692 5492 31708
rect 120 31628 5408 31692
rect 5472 31628 5492 31692
rect 120 31612 5492 31628
rect 120 31548 5408 31612
rect 5472 31548 5492 31612
rect 120 31532 5492 31548
rect 120 31468 5408 31532
rect 5472 31468 5492 31532
rect 120 31452 5492 31468
rect 120 31388 5408 31452
rect 5472 31388 5492 31452
rect 120 31372 5492 31388
rect 120 31308 5408 31372
rect 5472 31308 5492 31372
rect 120 31292 5492 31308
rect 120 31228 5408 31292
rect 5472 31228 5492 31292
rect 120 31212 5492 31228
rect 120 31148 5408 31212
rect 5472 31148 5492 31212
rect 120 31132 5492 31148
rect 120 31068 5408 31132
rect 5472 31068 5492 31132
rect 120 31052 5492 31068
rect 120 30988 5408 31052
rect 5472 30988 5492 31052
rect 120 30972 5492 30988
rect 120 30908 5408 30972
rect 5472 30908 5492 30972
rect 120 30892 5492 30908
rect 120 30828 5408 30892
rect 5472 30828 5492 30892
rect 120 30812 5492 30828
rect 120 30748 5408 30812
rect 5472 30748 5492 30812
rect 120 30732 5492 30748
rect 120 30668 5408 30732
rect 5472 30668 5492 30732
rect 120 30652 5492 30668
rect 120 30588 5408 30652
rect 5472 30588 5492 30652
rect 120 30572 5492 30588
rect 120 30508 5408 30572
rect 5472 30508 5492 30572
rect 120 30492 5492 30508
rect 120 30428 5408 30492
rect 5472 30428 5492 30492
rect 120 30412 5492 30428
rect 120 30348 5408 30412
rect 5472 30348 5492 30412
rect 120 30332 5492 30348
rect 120 30268 5408 30332
rect 5472 30268 5492 30332
rect 120 30252 5492 30268
rect 120 30188 5408 30252
rect 5472 30188 5492 30252
rect 120 30172 5492 30188
rect 120 30108 5408 30172
rect 5472 30108 5492 30172
rect 120 30092 5492 30108
rect 120 30028 5408 30092
rect 5472 30028 5492 30092
rect 120 30012 5492 30028
rect 120 29948 5408 30012
rect 5472 29948 5492 30012
rect 120 29932 5492 29948
rect 120 29868 5408 29932
rect 5472 29868 5492 29932
rect 120 29852 5492 29868
rect 120 29788 5408 29852
rect 5472 29788 5492 29852
rect 120 29772 5492 29788
rect 120 29708 5408 29772
rect 5472 29708 5492 29772
rect 120 29692 5492 29708
rect 120 29628 5408 29692
rect 5472 29628 5492 29692
rect 120 29612 5492 29628
rect 120 29548 5408 29612
rect 5472 29548 5492 29612
rect 120 29532 5492 29548
rect 120 29468 5408 29532
rect 5472 29468 5492 29532
rect 120 29452 5492 29468
rect 120 29388 5408 29452
rect 5472 29388 5492 29452
rect 120 29372 5492 29388
rect 120 29308 5408 29372
rect 5472 29308 5492 29372
rect 120 29292 5492 29308
rect 120 29228 5408 29292
rect 5472 29228 5492 29292
rect 120 29212 5492 29228
rect 120 29148 5408 29212
rect 5472 29148 5492 29212
rect 120 29132 5492 29148
rect 120 29068 5408 29132
rect 5472 29068 5492 29132
rect 120 29052 5492 29068
rect 120 28988 5408 29052
rect 5472 28988 5492 29052
rect 120 28972 5492 28988
rect 120 28908 5408 28972
rect 5472 28908 5492 28972
rect 120 28892 5492 28908
rect 120 28828 5408 28892
rect 5472 28828 5492 28892
rect 120 28812 5492 28828
rect 120 28748 5408 28812
rect 5472 28748 5492 28812
rect 120 28732 5492 28748
rect 120 28668 5408 28732
rect 5472 28668 5492 28732
rect 120 28652 5492 28668
rect 120 28588 5408 28652
rect 5472 28588 5492 28652
rect 120 28572 5492 28588
rect 120 28508 5408 28572
rect 5472 28508 5492 28572
rect 120 28492 5492 28508
rect 120 28428 5408 28492
rect 5472 28428 5492 28492
rect 120 28412 5492 28428
rect 120 28348 5408 28412
rect 5472 28348 5492 28412
rect 120 28332 5492 28348
rect 120 28268 5408 28332
rect 5472 28268 5492 28332
rect 120 28252 5492 28268
rect 120 28188 5408 28252
rect 5472 28188 5492 28252
rect 120 28172 5492 28188
rect 120 28108 5408 28172
rect 5472 28108 5492 28172
rect 120 28092 5492 28108
rect 120 28028 5408 28092
rect 5472 28028 5492 28092
rect 120 28012 5492 28028
rect 120 27948 5408 28012
rect 5472 27948 5492 28012
rect 120 27932 5492 27948
rect 120 27868 5408 27932
rect 5472 27868 5492 27932
rect 120 27852 5492 27868
rect 120 27788 5408 27852
rect 5472 27788 5492 27852
rect 120 27772 5492 27788
rect 120 27708 5408 27772
rect 5472 27708 5492 27772
rect 120 27692 5492 27708
rect 120 27628 5408 27692
rect 5472 27628 5492 27692
rect 120 27612 5492 27628
rect 120 27548 5408 27612
rect 5472 27548 5492 27612
rect 120 27532 5492 27548
rect 120 27468 5408 27532
rect 5472 27468 5492 27532
rect 120 27452 5492 27468
rect 120 27388 5408 27452
rect 5472 27388 5492 27452
rect 120 27372 5492 27388
rect 120 27308 5408 27372
rect 5472 27308 5492 27372
rect 120 27292 5492 27308
rect 120 27228 5408 27292
rect 5472 27228 5492 27292
rect 120 27212 5492 27228
rect 120 27148 5408 27212
rect 5472 27148 5492 27212
rect 120 27132 5492 27148
rect 120 27068 5408 27132
rect 5472 27068 5492 27132
rect 120 27052 5492 27068
rect 120 26988 5408 27052
rect 5472 26988 5492 27052
rect 120 26972 5492 26988
rect 120 26908 5408 26972
rect 5472 26908 5492 26972
rect 120 26892 5492 26908
rect 120 26828 5408 26892
rect 5472 26828 5492 26892
rect 120 26812 5492 26828
rect 120 26748 5408 26812
rect 5472 26748 5492 26812
rect 120 26720 5492 26748
rect 5732 31772 11104 31800
rect 5732 31708 11020 31772
rect 11084 31708 11104 31772
rect 5732 31692 11104 31708
rect 5732 31628 11020 31692
rect 11084 31628 11104 31692
rect 5732 31612 11104 31628
rect 5732 31548 11020 31612
rect 11084 31548 11104 31612
rect 5732 31532 11104 31548
rect 5732 31468 11020 31532
rect 11084 31468 11104 31532
rect 5732 31452 11104 31468
rect 5732 31388 11020 31452
rect 11084 31388 11104 31452
rect 5732 31372 11104 31388
rect 5732 31308 11020 31372
rect 11084 31308 11104 31372
rect 5732 31292 11104 31308
rect 5732 31228 11020 31292
rect 11084 31228 11104 31292
rect 5732 31212 11104 31228
rect 5732 31148 11020 31212
rect 11084 31148 11104 31212
rect 5732 31132 11104 31148
rect 5732 31068 11020 31132
rect 11084 31068 11104 31132
rect 5732 31052 11104 31068
rect 5732 30988 11020 31052
rect 11084 30988 11104 31052
rect 5732 30972 11104 30988
rect 5732 30908 11020 30972
rect 11084 30908 11104 30972
rect 5732 30892 11104 30908
rect 5732 30828 11020 30892
rect 11084 30828 11104 30892
rect 5732 30812 11104 30828
rect 5732 30748 11020 30812
rect 11084 30748 11104 30812
rect 5732 30732 11104 30748
rect 5732 30668 11020 30732
rect 11084 30668 11104 30732
rect 5732 30652 11104 30668
rect 5732 30588 11020 30652
rect 11084 30588 11104 30652
rect 5732 30572 11104 30588
rect 5732 30508 11020 30572
rect 11084 30508 11104 30572
rect 5732 30492 11104 30508
rect 5732 30428 11020 30492
rect 11084 30428 11104 30492
rect 5732 30412 11104 30428
rect 5732 30348 11020 30412
rect 11084 30348 11104 30412
rect 5732 30332 11104 30348
rect 5732 30268 11020 30332
rect 11084 30268 11104 30332
rect 5732 30252 11104 30268
rect 5732 30188 11020 30252
rect 11084 30188 11104 30252
rect 5732 30172 11104 30188
rect 5732 30108 11020 30172
rect 11084 30108 11104 30172
rect 5732 30092 11104 30108
rect 5732 30028 11020 30092
rect 11084 30028 11104 30092
rect 5732 30012 11104 30028
rect 5732 29948 11020 30012
rect 11084 29948 11104 30012
rect 5732 29932 11104 29948
rect 5732 29868 11020 29932
rect 11084 29868 11104 29932
rect 5732 29852 11104 29868
rect 5732 29788 11020 29852
rect 11084 29788 11104 29852
rect 5732 29772 11104 29788
rect 5732 29708 11020 29772
rect 11084 29708 11104 29772
rect 5732 29692 11104 29708
rect 5732 29628 11020 29692
rect 11084 29628 11104 29692
rect 5732 29612 11104 29628
rect 5732 29548 11020 29612
rect 11084 29548 11104 29612
rect 5732 29532 11104 29548
rect 5732 29468 11020 29532
rect 11084 29468 11104 29532
rect 5732 29452 11104 29468
rect 5732 29388 11020 29452
rect 11084 29388 11104 29452
rect 5732 29372 11104 29388
rect 5732 29308 11020 29372
rect 11084 29308 11104 29372
rect 5732 29292 11104 29308
rect 5732 29228 11020 29292
rect 11084 29228 11104 29292
rect 5732 29212 11104 29228
rect 5732 29148 11020 29212
rect 11084 29148 11104 29212
rect 5732 29132 11104 29148
rect 5732 29068 11020 29132
rect 11084 29068 11104 29132
rect 5732 29052 11104 29068
rect 5732 28988 11020 29052
rect 11084 28988 11104 29052
rect 5732 28972 11104 28988
rect 5732 28908 11020 28972
rect 11084 28908 11104 28972
rect 5732 28892 11104 28908
rect 5732 28828 11020 28892
rect 11084 28828 11104 28892
rect 5732 28812 11104 28828
rect 5732 28748 11020 28812
rect 11084 28748 11104 28812
rect 5732 28732 11104 28748
rect 5732 28668 11020 28732
rect 11084 28668 11104 28732
rect 5732 28652 11104 28668
rect 5732 28588 11020 28652
rect 11084 28588 11104 28652
rect 5732 28572 11104 28588
rect 5732 28508 11020 28572
rect 11084 28508 11104 28572
rect 5732 28492 11104 28508
rect 5732 28428 11020 28492
rect 11084 28428 11104 28492
rect 5732 28412 11104 28428
rect 5732 28348 11020 28412
rect 11084 28348 11104 28412
rect 5732 28332 11104 28348
rect 5732 28268 11020 28332
rect 11084 28268 11104 28332
rect 5732 28252 11104 28268
rect 5732 28188 11020 28252
rect 11084 28188 11104 28252
rect 5732 28172 11104 28188
rect 5732 28108 11020 28172
rect 11084 28108 11104 28172
rect 5732 28092 11104 28108
rect 5732 28028 11020 28092
rect 11084 28028 11104 28092
rect 5732 28012 11104 28028
rect 5732 27948 11020 28012
rect 11084 27948 11104 28012
rect 5732 27932 11104 27948
rect 5732 27868 11020 27932
rect 11084 27868 11104 27932
rect 5732 27852 11104 27868
rect 5732 27788 11020 27852
rect 11084 27788 11104 27852
rect 5732 27772 11104 27788
rect 5732 27708 11020 27772
rect 11084 27708 11104 27772
rect 5732 27692 11104 27708
rect 5732 27628 11020 27692
rect 11084 27628 11104 27692
rect 5732 27612 11104 27628
rect 5732 27548 11020 27612
rect 11084 27548 11104 27612
rect 5732 27532 11104 27548
rect 5732 27468 11020 27532
rect 11084 27468 11104 27532
rect 5732 27452 11104 27468
rect 5732 27388 11020 27452
rect 11084 27388 11104 27452
rect 5732 27372 11104 27388
rect 5732 27308 11020 27372
rect 11084 27308 11104 27372
rect 5732 27292 11104 27308
rect 5732 27228 11020 27292
rect 11084 27228 11104 27292
rect 5732 27212 11104 27228
rect 5732 27148 11020 27212
rect 11084 27148 11104 27212
rect 5732 27132 11104 27148
rect 5732 27068 11020 27132
rect 11084 27068 11104 27132
rect 5732 27052 11104 27068
rect 5732 26988 11020 27052
rect 11084 26988 11104 27052
rect 5732 26972 11104 26988
rect 5732 26908 11020 26972
rect 11084 26908 11104 26972
rect 5732 26892 11104 26908
rect 5732 26828 11020 26892
rect 11084 26828 11104 26892
rect 5732 26812 11104 26828
rect 5732 26748 11020 26812
rect 11084 26748 11104 26812
rect 5732 26720 11104 26748
rect 11344 31772 16716 31800
rect 11344 31708 16632 31772
rect 16696 31708 16716 31772
rect 11344 31692 16716 31708
rect 11344 31628 16632 31692
rect 16696 31628 16716 31692
rect 11344 31612 16716 31628
rect 11344 31548 16632 31612
rect 16696 31548 16716 31612
rect 11344 31532 16716 31548
rect 11344 31468 16632 31532
rect 16696 31468 16716 31532
rect 11344 31452 16716 31468
rect 11344 31388 16632 31452
rect 16696 31388 16716 31452
rect 11344 31372 16716 31388
rect 11344 31308 16632 31372
rect 16696 31308 16716 31372
rect 11344 31292 16716 31308
rect 11344 31228 16632 31292
rect 16696 31228 16716 31292
rect 11344 31212 16716 31228
rect 11344 31148 16632 31212
rect 16696 31148 16716 31212
rect 11344 31132 16716 31148
rect 11344 31068 16632 31132
rect 16696 31068 16716 31132
rect 11344 31052 16716 31068
rect 11344 30988 16632 31052
rect 16696 30988 16716 31052
rect 11344 30972 16716 30988
rect 11344 30908 16632 30972
rect 16696 30908 16716 30972
rect 11344 30892 16716 30908
rect 11344 30828 16632 30892
rect 16696 30828 16716 30892
rect 11344 30812 16716 30828
rect 11344 30748 16632 30812
rect 16696 30748 16716 30812
rect 11344 30732 16716 30748
rect 11344 30668 16632 30732
rect 16696 30668 16716 30732
rect 11344 30652 16716 30668
rect 11344 30588 16632 30652
rect 16696 30588 16716 30652
rect 11344 30572 16716 30588
rect 11344 30508 16632 30572
rect 16696 30508 16716 30572
rect 11344 30492 16716 30508
rect 11344 30428 16632 30492
rect 16696 30428 16716 30492
rect 11344 30412 16716 30428
rect 11344 30348 16632 30412
rect 16696 30348 16716 30412
rect 11344 30332 16716 30348
rect 11344 30268 16632 30332
rect 16696 30268 16716 30332
rect 11344 30252 16716 30268
rect 11344 30188 16632 30252
rect 16696 30188 16716 30252
rect 11344 30172 16716 30188
rect 11344 30108 16632 30172
rect 16696 30108 16716 30172
rect 11344 30092 16716 30108
rect 11344 30028 16632 30092
rect 16696 30028 16716 30092
rect 11344 30012 16716 30028
rect 11344 29948 16632 30012
rect 16696 29948 16716 30012
rect 11344 29932 16716 29948
rect 11344 29868 16632 29932
rect 16696 29868 16716 29932
rect 11344 29852 16716 29868
rect 11344 29788 16632 29852
rect 16696 29788 16716 29852
rect 11344 29772 16716 29788
rect 11344 29708 16632 29772
rect 16696 29708 16716 29772
rect 11344 29692 16716 29708
rect 11344 29628 16632 29692
rect 16696 29628 16716 29692
rect 11344 29612 16716 29628
rect 11344 29548 16632 29612
rect 16696 29548 16716 29612
rect 11344 29532 16716 29548
rect 11344 29468 16632 29532
rect 16696 29468 16716 29532
rect 11344 29452 16716 29468
rect 11344 29388 16632 29452
rect 16696 29388 16716 29452
rect 11344 29372 16716 29388
rect 11344 29308 16632 29372
rect 16696 29308 16716 29372
rect 11344 29292 16716 29308
rect 11344 29228 16632 29292
rect 16696 29228 16716 29292
rect 11344 29212 16716 29228
rect 11344 29148 16632 29212
rect 16696 29148 16716 29212
rect 11344 29132 16716 29148
rect 11344 29068 16632 29132
rect 16696 29068 16716 29132
rect 11344 29052 16716 29068
rect 11344 28988 16632 29052
rect 16696 28988 16716 29052
rect 11344 28972 16716 28988
rect 11344 28908 16632 28972
rect 16696 28908 16716 28972
rect 11344 28892 16716 28908
rect 11344 28828 16632 28892
rect 16696 28828 16716 28892
rect 11344 28812 16716 28828
rect 11344 28748 16632 28812
rect 16696 28748 16716 28812
rect 11344 28732 16716 28748
rect 11344 28668 16632 28732
rect 16696 28668 16716 28732
rect 11344 28652 16716 28668
rect 11344 28588 16632 28652
rect 16696 28588 16716 28652
rect 11344 28572 16716 28588
rect 11344 28508 16632 28572
rect 16696 28508 16716 28572
rect 11344 28492 16716 28508
rect 11344 28428 16632 28492
rect 16696 28428 16716 28492
rect 11344 28412 16716 28428
rect 11344 28348 16632 28412
rect 16696 28348 16716 28412
rect 11344 28332 16716 28348
rect 11344 28268 16632 28332
rect 16696 28268 16716 28332
rect 11344 28252 16716 28268
rect 11344 28188 16632 28252
rect 16696 28188 16716 28252
rect 11344 28172 16716 28188
rect 11344 28108 16632 28172
rect 16696 28108 16716 28172
rect 11344 28092 16716 28108
rect 11344 28028 16632 28092
rect 16696 28028 16716 28092
rect 11344 28012 16716 28028
rect 11344 27948 16632 28012
rect 16696 27948 16716 28012
rect 11344 27932 16716 27948
rect 11344 27868 16632 27932
rect 16696 27868 16716 27932
rect 11344 27852 16716 27868
rect 11344 27788 16632 27852
rect 16696 27788 16716 27852
rect 11344 27772 16716 27788
rect 11344 27708 16632 27772
rect 16696 27708 16716 27772
rect 11344 27692 16716 27708
rect 11344 27628 16632 27692
rect 16696 27628 16716 27692
rect 11344 27612 16716 27628
rect 11344 27548 16632 27612
rect 16696 27548 16716 27612
rect 11344 27532 16716 27548
rect 11344 27468 16632 27532
rect 16696 27468 16716 27532
rect 11344 27452 16716 27468
rect 11344 27388 16632 27452
rect 16696 27388 16716 27452
rect 11344 27372 16716 27388
rect 11344 27308 16632 27372
rect 16696 27308 16716 27372
rect 11344 27292 16716 27308
rect 11344 27228 16632 27292
rect 16696 27228 16716 27292
rect 11344 27212 16716 27228
rect 11344 27148 16632 27212
rect 16696 27148 16716 27212
rect 11344 27132 16716 27148
rect 11344 27068 16632 27132
rect 16696 27068 16716 27132
rect 11344 27052 16716 27068
rect 11344 26988 16632 27052
rect 16696 26988 16716 27052
rect 11344 26972 16716 26988
rect 11344 26908 16632 26972
rect 16696 26908 16716 26972
rect 11344 26892 16716 26908
rect 11344 26828 16632 26892
rect 16696 26828 16716 26892
rect 11344 26812 16716 26828
rect 11344 26748 16632 26812
rect 16696 26748 16716 26812
rect 11344 26720 16716 26748
rect 16956 31772 22328 31800
rect 16956 31708 22244 31772
rect 22308 31708 22328 31772
rect 16956 31692 22328 31708
rect 16956 31628 22244 31692
rect 22308 31628 22328 31692
rect 16956 31612 22328 31628
rect 16956 31548 22244 31612
rect 22308 31548 22328 31612
rect 16956 31532 22328 31548
rect 16956 31468 22244 31532
rect 22308 31468 22328 31532
rect 16956 31452 22328 31468
rect 16956 31388 22244 31452
rect 22308 31388 22328 31452
rect 16956 31372 22328 31388
rect 16956 31308 22244 31372
rect 22308 31308 22328 31372
rect 16956 31292 22328 31308
rect 16956 31228 22244 31292
rect 22308 31228 22328 31292
rect 16956 31212 22328 31228
rect 16956 31148 22244 31212
rect 22308 31148 22328 31212
rect 16956 31132 22328 31148
rect 16956 31068 22244 31132
rect 22308 31068 22328 31132
rect 16956 31052 22328 31068
rect 16956 30988 22244 31052
rect 22308 30988 22328 31052
rect 16956 30972 22328 30988
rect 16956 30908 22244 30972
rect 22308 30908 22328 30972
rect 16956 30892 22328 30908
rect 16956 30828 22244 30892
rect 22308 30828 22328 30892
rect 16956 30812 22328 30828
rect 16956 30748 22244 30812
rect 22308 30748 22328 30812
rect 16956 30732 22328 30748
rect 16956 30668 22244 30732
rect 22308 30668 22328 30732
rect 16956 30652 22328 30668
rect 16956 30588 22244 30652
rect 22308 30588 22328 30652
rect 16956 30572 22328 30588
rect 16956 30508 22244 30572
rect 22308 30508 22328 30572
rect 16956 30492 22328 30508
rect 16956 30428 22244 30492
rect 22308 30428 22328 30492
rect 16956 30412 22328 30428
rect 16956 30348 22244 30412
rect 22308 30348 22328 30412
rect 16956 30332 22328 30348
rect 16956 30268 22244 30332
rect 22308 30268 22328 30332
rect 16956 30252 22328 30268
rect 16956 30188 22244 30252
rect 22308 30188 22328 30252
rect 16956 30172 22328 30188
rect 16956 30108 22244 30172
rect 22308 30108 22328 30172
rect 16956 30092 22328 30108
rect 16956 30028 22244 30092
rect 22308 30028 22328 30092
rect 16956 30012 22328 30028
rect 16956 29948 22244 30012
rect 22308 29948 22328 30012
rect 16956 29932 22328 29948
rect 16956 29868 22244 29932
rect 22308 29868 22328 29932
rect 16956 29852 22328 29868
rect 16956 29788 22244 29852
rect 22308 29788 22328 29852
rect 16956 29772 22328 29788
rect 16956 29708 22244 29772
rect 22308 29708 22328 29772
rect 16956 29692 22328 29708
rect 16956 29628 22244 29692
rect 22308 29628 22328 29692
rect 16956 29612 22328 29628
rect 16956 29548 22244 29612
rect 22308 29548 22328 29612
rect 16956 29532 22328 29548
rect 16956 29468 22244 29532
rect 22308 29468 22328 29532
rect 16956 29452 22328 29468
rect 16956 29388 22244 29452
rect 22308 29388 22328 29452
rect 16956 29372 22328 29388
rect 16956 29308 22244 29372
rect 22308 29308 22328 29372
rect 16956 29292 22328 29308
rect 16956 29228 22244 29292
rect 22308 29228 22328 29292
rect 16956 29212 22328 29228
rect 16956 29148 22244 29212
rect 22308 29148 22328 29212
rect 16956 29132 22328 29148
rect 16956 29068 22244 29132
rect 22308 29068 22328 29132
rect 16956 29052 22328 29068
rect 16956 28988 22244 29052
rect 22308 28988 22328 29052
rect 16956 28972 22328 28988
rect 16956 28908 22244 28972
rect 22308 28908 22328 28972
rect 16956 28892 22328 28908
rect 16956 28828 22244 28892
rect 22308 28828 22328 28892
rect 16956 28812 22328 28828
rect 16956 28748 22244 28812
rect 22308 28748 22328 28812
rect 16956 28732 22328 28748
rect 16956 28668 22244 28732
rect 22308 28668 22328 28732
rect 16956 28652 22328 28668
rect 16956 28588 22244 28652
rect 22308 28588 22328 28652
rect 16956 28572 22328 28588
rect 16956 28508 22244 28572
rect 22308 28508 22328 28572
rect 16956 28492 22328 28508
rect 16956 28428 22244 28492
rect 22308 28428 22328 28492
rect 16956 28412 22328 28428
rect 16956 28348 22244 28412
rect 22308 28348 22328 28412
rect 16956 28332 22328 28348
rect 16956 28268 22244 28332
rect 22308 28268 22328 28332
rect 16956 28252 22328 28268
rect 16956 28188 22244 28252
rect 22308 28188 22328 28252
rect 16956 28172 22328 28188
rect 16956 28108 22244 28172
rect 22308 28108 22328 28172
rect 16956 28092 22328 28108
rect 16956 28028 22244 28092
rect 22308 28028 22328 28092
rect 16956 28012 22328 28028
rect 16956 27948 22244 28012
rect 22308 27948 22328 28012
rect 16956 27932 22328 27948
rect 16956 27868 22244 27932
rect 22308 27868 22328 27932
rect 16956 27852 22328 27868
rect 16956 27788 22244 27852
rect 22308 27788 22328 27852
rect 16956 27772 22328 27788
rect 16956 27708 22244 27772
rect 22308 27708 22328 27772
rect 16956 27692 22328 27708
rect 16956 27628 22244 27692
rect 22308 27628 22328 27692
rect 16956 27612 22328 27628
rect 16956 27548 22244 27612
rect 22308 27548 22328 27612
rect 16956 27532 22328 27548
rect 16956 27468 22244 27532
rect 22308 27468 22328 27532
rect 16956 27452 22328 27468
rect 16956 27388 22244 27452
rect 22308 27388 22328 27452
rect 16956 27372 22328 27388
rect 16956 27308 22244 27372
rect 22308 27308 22328 27372
rect 16956 27292 22328 27308
rect 16956 27228 22244 27292
rect 22308 27228 22328 27292
rect 16956 27212 22328 27228
rect 16956 27148 22244 27212
rect 22308 27148 22328 27212
rect 16956 27132 22328 27148
rect 16956 27068 22244 27132
rect 22308 27068 22328 27132
rect 16956 27052 22328 27068
rect 16956 26988 22244 27052
rect 22308 26988 22328 27052
rect 16956 26972 22328 26988
rect 16956 26908 22244 26972
rect 22308 26908 22328 26972
rect 16956 26892 22328 26908
rect 16956 26828 22244 26892
rect 22308 26828 22328 26892
rect 16956 26812 22328 26828
rect 16956 26748 22244 26812
rect 22308 26748 22328 26812
rect 16956 26720 22328 26748
rect 22568 31772 27940 31800
rect 22568 31708 27856 31772
rect 27920 31708 27940 31772
rect 22568 31692 27940 31708
rect 22568 31628 27856 31692
rect 27920 31628 27940 31692
rect 22568 31612 27940 31628
rect 22568 31548 27856 31612
rect 27920 31548 27940 31612
rect 22568 31532 27940 31548
rect 22568 31468 27856 31532
rect 27920 31468 27940 31532
rect 22568 31452 27940 31468
rect 22568 31388 27856 31452
rect 27920 31388 27940 31452
rect 22568 31372 27940 31388
rect 22568 31308 27856 31372
rect 27920 31308 27940 31372
rect 22568 31292 27940 31308
rect 22568 31228 27856 31292
rect 27920 31228 27940 31292
rect 22568 31212 27940 31228
rect 22568 31148 27856 31212
rect 27920 31148 27940 31212
rect 22568 31132 27940 31148
rect 22568 31068 27856 31132
rect 27920 31068 27940 31132
rect 22568 31052 27940 31068
rect 22568 30988 27856 31052
rect 27920 30988 27940 31052
rect 22568 30972 27940 30988
rect 22568 30908 27856 30972
rect 27920 30908 27940 30972
rect 22568 30892 27940 30908
rect 22568 30828 27856 30892
rect 27920 30828 27940 30892
rect 22568 30812 27940 30828
rect 22568 30748 27856 30812
rect 27920 30748 27940 30812
rect 22568 30732 27940 30748
rect 22568 30668 27856 30732
rect 27920 30668 27940 30732
rect 22568 30652 27940 30668
rect 22568 30588 27856 30652
rect 27920 30588 27940 30652
rect 22568 30572 27940 30588
rect 22568 30508 27856 30572
rect 27920 30508 27940 30572
rect 22568 30492 27940 30508
rect 22568 30428 27856 30492
rect 27920 30428 27940 30492
rect 22568 30412 27940 30428
rect 22568 30348 27856 30412
rect 27920 30348 27940 30412
rect 22568 30332 27940 30348
rect 22568 30268 27856 30332
rect 27920 30268 27940 30332
rect 22568 30252 27940 30268
rect 22568 30188 27856 30252
rect 27920 30188 27940 30252
rect 22568 30172 27940 30188
rect 22568 30108 27856 30172
rect 27920 30108 27940 30172
rect 22568 30092 27940 30108
rect 22568 30028 27856 30092
rect 27920 30028 27940 30092
rect 22568 30012 27940 30028
rect 22568 29948 27856 30012
rect 27920 29948 27940 30012
rect 22568 29932 27940 29948
rect 22568 29868 27856 29932
rect 27920 29868 27940 29932
rect 22568 29852 27940 29868
rect 22568 29788 27856 29852
rect 27920 29788 27940 29852
rect 22568 29772 27940 29788
rect 22568 29708 27856 29772
rect 27920 29708 27940 29772
rect 22568 29692 27940 29708
rect 22568 29628 27856 29692
rect 27920 29628 27940 29692
rect 22568 29612 27940 29628
rect 22568 29548 27856 29612
rect 27920 29548 27940 29612
rect 22568 29532 27940 29548
rect 22568 29468 27856 29532
rect 27920 29468 27940 29532
rect 22568 29452 27940 29468
rect 22568 29388 27856 29452
rect 27920 29388 27940 29452
rect 22568 29372 27940 29388
rect 22568 29308 27856 29372
rect 27920 29308 27940 29372
rect 22568 29292 27940 29308
rect 22568 29228 27856 29292
rect 27920 29228 27940 29292
rect 22568 29212 27940 29228
rect 22568 29148 27856 29212
rect 27920 29148 27940 29212
rect 22568 29132 27940 29148
rect 22568 29068 27856 29132
rect 27920 29068 27940 29132
rect 22568 29052 27940 29068
rect 22568 28988 27856 29052
rect 27920 28988 27940 29052
rect 22568 28972 27940 28988
rect 22568 28908 27856 28972
rect 27920 28908 27940 28972
rect 22568 28892 27940 28908
rect 22568 28828 27856 28892
rect 27920 28828 27940 28892
rect 22568 28812 27940 28828
rect 22568 28748 27856 28812
rect 27920 28748 27940 28812
rect 22568 28732 27940 28748
rect 22568 28668 27856 28732
rect 27920 28668 27940 28732
rect 22568 28652 27940 28668
rect 22568 28588 27856 28652
rect 27920 28588 27940 28652
rect 22568 28572 27940 28588
rect 22568 28508 27856 28572
rect 27920 28508 27940 28572
rect 22568 28492 27940 28508
rect 22568 28428 27856 28492
rect 27920 28428 27940 28492
rect 22568 28412 27940 28428
rect 22568 28348 27856 28412
rect 27920 28348 27940 28412
rect 22568 28332 27940 28348
rect 22568 28268 27856 28332
rect 27920 28268 27940 28332
rect 22568 28252 27940 28268
rect 22568 28188 27856 28252
rect 27920 28188 27940 28252
rect 22568 28172 27940 28188
rect 22568 28108 27856 28172
rect 27920 28108 27940 28172
rect 22568 28092 27940 28108
rect 22568 28028 27856 28092
rect 27920 28028 27940 28092
rect 22568 28012 27940 28028
rect 22568 27948 27856 28012
rect 27920 27948 27940 28012
rect 22568 27932 27940 27948
rect 22568 27868 27856 27932
rect 27920 27868 27940 27932
rect 22568 27852 27940 27868
rect 22568 27788 27856 27852
rect 27920 27788 27940 27852
rect 22568 27772 27940 27788
rect 22568 27708 27856 27772
rect 27920 27708 27940 27772
rect 22568 27692 27940 27708
rect 22568 27628 27856 27692
rect 27920 27628 27940 27692
rect 22568 27612 27940 27628
rect 22568 27548 27856 27612
rect 27920 27548 27940 27612
rect 22568 27532 27940 27548
rect 22568 27468 27856 27532
rect 27920 27468 27940 27532
rect 22568 27452 27940 27468
rect 22568 27388 27856 27452
rect 27920 27388 27940 27452
rect 22568 27372 27940 27388
rect 22568 27308 27856 27372
rect 27920 27308 27940 27372
rect 22568 27292 27940 27308
rect 22568 27228 27856 27292
rect 27920 27228 27940 27292
rect 22568 27212 27940 27228
rect 22568 27148 27856 27212
rect 27920 27148 27940 27212
rect 22568 27132 27940 27148
rect 22568 27068 27856 27132
rect 27920 27068 27940 27132
rect 22568 27052 27940 27068
rect 22568 26988 27856 27052
rect 27920 26988 27940 27052
rect 22568 26972 27940 26988
rect 22568 26908 27856 26972
rect 27920 26908 27940 26972
rect 22568 26892 27940 26908
rect 22568 26828 27856 26892
rect 27920 26828 27940 26892
rect 22568 26812 27940 26828
rect 22568 26748 27856 26812
rect 27920 26748 27940 26812
rect 22568 26720 27940 26748
rect 28180 31772 33552 31800
rect 28180 31708 33468 31772
rect 33532 31708 33552 31772
rect 28180 31692 33552 31708
rect 28180 31628 33468 31692
rect 33532 31628 33552 31692
rect 28180 31612 33552 31628
rect 28180 31548 33468 31612
rect 33532 31548 33552 31612
rect 28180 31532 33552 31548
rect 28180 31468 33468 31532
rect 33532 31468 33552 31532
rect 28180 31452 33552 31468
rect 28180 31388 33468 31452
rect 33532 31388 33552 31452
rect 28180 31372 33552 31388
rect 28180 31308 33468 31372
rect 33532 31308 33552 31372
rect 28180 31292 33552 31308
rect 28180 31228 33468 31292
rect 33532 31228 33552 31292
rect 28180 31212 33552 31228
rect 28180 31148 33468 31212
rect 33532 31148 33552 31212
rect 28180 31132 33552 31148
rect 28180 31068 33468 31132
rect 33532 31068 33552 31132
rect 28180 31052 33552 31068
rect 28180 30988 33468 31052
rect 33532 30988 33552 31052
rect 28180 30972 33552 30988
rect 28180 30908 33468 30972
rect 33532 30908 33552 30972
rect 28180 30892 33552 30908
rect 28180 30828 33468 30892
rect 33532 30828 33552 30892
rect 28180 30812 33552 30828
rect 28180 30748 33468 30812
rect 33532 30748 33552 30812
rect 28180 30732 33552 30748
rect 28180 30668 33468 30732
rect 33532 30668 33552 30732
rect 28180 30652 33552 30668
rect 28180 30588 33468 30652
rect 33532 30588 33552 30652
rect 28180 30572 33552 30588
rect 28180 30508 33468 30572
rect 33532 30508 33552 30572
rect 28180 30492 33552 30508
rect 28180 30428 33468 30492
rect 33532 30428 33552 30492
rect 28180 30412 33552 30428
rect 28180 30348 33468 30412
rect 33532 30348 33552 30412
rect 28180 30332 33552 30348
rect 28180 30268 33468 30332
rect 33532 30268 33552 30332
rect 28180 30252 33552 30268
rect 28180 30188 33468 30252
rect 33532 30188 33552 30252
rect 28180 30172 33552 30188
rect 28180 30108 33468 30172
rect 33532 30108 33552 30172
rect 28180 30092 33552 30108
rect 28180 30028 33468 30092
rect 33532 30028 33552 30092
rect 28180 30012 33552 30028
rect 28180 29948 33468 30012
rect 33532 29948 33552 30012
rect 28180 29932 33552 29948
rect 28180 29868 33468 29932
rect 33532 29868 33552 29932
rect 28180 29852 33552 29868
rect 28180 29788 33468 29852
rect 33532 29788 33552 29852
rect 28180 29772 33552 29788
rect 28180 29708 33468 29772
rect 33532 29708 33552 29772
rect 28180 29692 33552 29708
rect 28180 29628 33468 29692
rect 33532 29628 33552 29692
rect 28180 29612 33552 29628
rect 28180 29548 33468 29612
rect 33532 29548 33552 29612
rect 28180 29532 33552 29548
rect 28180 29468 33468 29532
rect 33532 29468 33552 29532
rect 28180 29452 33552 29468
rect 28180 29388 33468 29452
rect 33532 29388 33552 29452
rect 28180 29372 33552 29388
rect 28180 29308 33468 29372
rect 33532 29308 33552 29372
rect 28180 29292 33552 29308
rect 28180 29228 33468 29292
rect 33532 29228 33552 29292
rect 28180 29212 33552 29228
rect 28180 29148 33468 29212
rect 33532 29148 33552 29212
rect 28180 29132 33552 29148
rect 28180 29068 33468 29132
rect 33532 29068 33552 29132
rect 28180 29052 33552 29068
rect 28180 28988 33468 29052
rect 33532 28988 33552 29052
rect 28180 28972 33552 28988
rect 28180 28908 33468 28972
rect 33532 28908 33552 28972
rect 28180 28892 33552 28908
rect 28180 28828 33468 28892
rect 33532 28828 33552 28892
rect 28180 28812 33552 28828
rect 28180 28748 33468 28812
rect 33532 28748 33552 28812
rect 28180 28732 33552 28748
rect 28180 28668 33468 28732
rect 33532 28668 33552 28732
rect 28180 28652 33552 28668
rect 28180 28588 33468 28652
rect 33532 28588 33552 28652
rect 28180 28572 33552 28588
rect 28180 28508 33468 28572
rect 33532 28508 33552 28572
rect 28180 28492 33552 28508
rect 28180 28428 33468 28492
rect 33532 28428 33552 28492
rect 28180 28412 33552 28428
rect 28180 28348 33468 28412
rect 33532 28348 33552 28412
rect 28180 28332 33552 28348
rect 28180 28268 33468 28332
rect 33532 28268 33552 28332
rect 28180 28252 33552 28268
rect 28180 28188 33468 28252
rect 33532 28188 33552 28252
rect 28180 28172 33552 28188
rect 28180 28108 33468 28172
rect 33532 28108 33552 28172
rect 28180 28092 33552 28108
rect 28180 28028 33468 28092
rect 33532 28028 33552 28092
rect 28180 28012 33552 28028
rect 28180 27948 33468 28012
rect 33532 27948 33552 28012
rect 28180 27932 33552 27948
rect 28180 27868 33468 27932
rect 33532 27868 33552 27932
rect 28180 27852 33552 27868
rect 28180 27788 33468 27852
rect 33532 27788 33552 27852
rect 28180 27772 33552 27788
rect 28180 27708 33468 27772
rect 33532 27708 33552 27772
rect 28180 27692 33552 27708
rect 28180 27628 33468 27692
rect 33532 27628 33552 27692
rect 28180 27612 33552 27628
rect 28180 27548 33468 27612
rect 33532 27548 33552 27612
rect 28180 27532 33552 27548
rect 28180 27468 33468 27532
rect 33532 27468 33552 27532
rect 28180 27452 33552 27468
rect 28180 27388 33468 27452
rect 33532 27388 33552 27452
rect 28180 27372 33552 27388
rect 28180 27308 33468 27372
rect 33532 27308 33552 27372
rect 28180 27292 33552 27308
rect 28180 27228 33468 27292
rect 33532 27228 33552 27292
rect 28180 27212 33552 27228
rect 28180 27148 33468 27212
rect 33532 27148 33552 27212
rect 28180 27132 33552 27148
rect 28180 27068 33468 27132
rect 33532 27068 33552 27132
rect 28180 27052 33552 27068
rect 28180 26988 33468 27052
rect 33532 26988 33552 27052
rect 28180 26972 33552 26988
rect 28180 26908 33468 26972
rect 33532 26908 33552 26972
rect 28180 26892 33552 26908
rect 28180 26828 33468 26892
rect 33532 26828 33552 26892
rect 28180 26812 33552 26828
rect 28180 26748 33468 26812
rect 33532 26748 33552 26812
rect 28180 26720 33552 26748
rect 33792 31772 39164 31800
rect 33792 31708 39080 31772
rect 39144 31708 39164 31772
rect 33792 31692 39164 31708
rect 33792 31628 39080 31692
rect 39144 31628 39164 31692
rect 33792 31612 39164 31628
rect 33792 31548 39080 31612
rect 39144 31548 39164 31612
rect 33792 31532 39164 31548
rect 33792 31468 39080 31532
rect 39144 31468 39164 31532
rect 33792 31452 39164 31468
rect 33792 31388 39080 31452
rect 39144 31388 39164 31452
rect 33792 31372 39164 31388
rect 33792 31308 39080 31372
rect 39144 31308 39164 31372
rect 33792 31292 39164 31308
rect 33792 31228 39080 31292
rect 39144 31228 39164 31292
rect 33792 31212 39164 31228
rect 33792 31148 39080 31212
rect 39144 31148 39164 31212
rect 33792 31132 39164 31148
rect 33792 31068 39080 31132
rect 39144 31068 39164 31132
rect 33792 31052 39164 31068
rect 33792 30988 39080 31052
rect 39144 30988 39164 31052
rect 33792 30972 39164 30988
rect 33792 30908 39080 30972
rect 39144 30908 39164 30972
rect 33792 30892 39164 30908
rect 33792 30828 39080 30892
rect 39144 30828 39164 30892
rect 33792 30812 39164 30828
rect 33792 30748 39080 30812
rect 39144 30748 39164 30812
rect 33792 30732 39164 30748
rect 33792 30668 39080 30732
rect 39144 30668 39164 30732
rect 33792 30652 39164 30668
rect 33792 30588 39080 30652
rect 39144 30588 39164 30652
rect 33792 30572 39164 30588
rect 33792 30508 39080 30572
rect 39144 30508 39164 30572
rect 33792 30492 39164 30508
rect 33792 30428 39080 30492
rect 39144 30428 39164 30492
rect 33792 30412 39164 30428
rect 33792 30348 39080 30412
rect 39144 30348 39164 30412
rect 33792 30332 39164 30348
rect 33792 30268 39080 30332
rect 39144 30268 39164 30332
rect 33792 30252 39164 30268
rect 33792 30188 39080 30252
rect 39144 30188 39164 30252
rect 33792 30172 39164 30188
rect 33792 30108 39080 30172
rect 39144 30108 39164 30172
rect 33792 30092 39164 30108
rect 33792 30028 39080 30092
rect 39144 30028 39164 30092
rect 33792 30012 39164 30028
rect 33792 29948 39080 30012
rect 39144 29948 39164 30012
rect 33792 29932 39164 29948
rect 33792 29868 39080 29932
rect 39144 29868 39164 29932
rect 33792 29852 39164 29868
rect 33792 29788 39080 29852
rect 39144 29788 39164 29852
rect 33792 29772 39164 29788
rect 33792 29708 39080 29772
rect 39144 29708 39164 29772
rect 33792 29692 39164 29708
rect 33792 29628 39080 29692
rect 39144 29628 39164 29692
rect 33792 29612 39164 29628
rect 33792 29548 39080 29612
rect 39144 29548 39164 29612
rect 33792 29532 39164 29548
rect 33792 29468 39080 29532
rect 39144 29468 39164 29532
rect 33792 29452 39164 29468
rect 33792 29388 39080 29452
rect 39144 29388 39164 29452
rect 33792 29372 39164 29388
rect 33792 29308 39080 29372
rect 39144 29308 39164 29372
rect 33792 29292 39164 29308
rect 33792 29228 39080 29292
rect 39144 29228 39164 29292
rect 33792 29212 39164 29228
rect 33792 29148 39080 29212
rect 39144 29148 39164 29212
rect 33792 29132 39164 29148
rect 33792 29068 39080 29132
rect 39144 29068 39164 29132
rect 33792 29052 39164 29068
rect 33792 28988 39080 29052
rect 39144 28988 39164 29052
rect 33792 28972 39164 28988
rect 33792 28908 39080 28972
rect 39144 28908 39164 28972
rect 33792 28892 39164 28908
rect 33792 28828 39080 28892
rect 39144 28828 39164 28892
rect 33792 28812 39164 28828
rect 33792 28748 39080 28812
rect 39144 28748 39164 28812
rect 33792 28732 39164 28748
rect 33792 28668 39080 28732
rect 39144 28668 39164 28732
rect 33792 28652 39164 28668
rect 33792 28588 39080 28652
rect 39144 28588 39164 28652
rect 33792 28572 39164 28588
rect 33792 28508 39080 28572
rect 39144 28508 39164 28572
rect 33792 28492 39164 28508
rect 33792 28428 39080 28492
rect 39144 28428 39164 28492
rect 33792 28412 39164 28428
rect 33792 28348 39080 28412
rect 39144 28348 39164 28412
rect 33792 28332 39164 28348
rect 33792 28268 39080 28332
rect 39144 28268 39164 28332
rect 33792 28252 39164 28268
rect 33792 28188 39080 28252
rect 39144 28188 39164 28252
rect 33792 28172 39164 28188
rect 33792 28108 39080 28172
rect 39144 28108 39164 28172
rect 33792 28092 39164 28108
rect 33792 28028 39080 28092
rect 39144 28028 39164 28092
rect 33792 28012 39164 28028
rect 33792 27948 39080 28012
rect 39144 27948 39164 28012
rect 33792 27932 39164 27948
rect 33792 27868 39080 27932
rect 39144 27868 39164 27932
rect 33792 27852 39164 27868
rect 33792 27788 39080 27852
rect 39144 27788 39164 27852
rect 33792 27772 39164 27788
rect 33792 27708 39080 27772
rect 39144 27708 39164 27772
rect 33792 27692 39164 27708
rect 33792 27628 39080 27692
rect 39144 27628 39164 27692
rect 33792 27612 39164 27628
rect 33792 27548 39080 27612
rect 39144 27548 39164 27612
rect 33792 27532 39164 27548
rect 33792 27468 39080 27532
rect 39144 27468 39164 27532
rect 33792 27452 39164 27468
rect 33792 27388 39080 27452
rect 39144 27388 39164 27452
rect 33792 27372 39164 27388
rect 33792 27308 39080 27372
rect 39144 27308 39164 27372
rect 33792 27292 39164 27308
rect 33792 27228 39080 27292
rect 39144 27228 39164 27292
rect 33792 27212 39164 27228
rect 33792 27148 39080 27212
rect 39144 27148 39164 27212
rect 33792 27132 39164 27148
rect 33792 27068 39080 27132
rect 39144 27068 39164 27132
rect 33792 27052 39164 27068
rect 33792 26988 39080 27052
rect 39144 26988 39164 27052
rect 33792 26972 39164 26988
rect 33792 26908 39080 26972
rect 39144 26908 39164 26972
rect 33792 26892 39164 26908
rect 33792 26828 39080 26892
rect 39144 26828 39164 26892
rect 33792 26812 39164 26828
rect 33792 26748 39080 26812
rect 39144 26748 39164 26812
rect 33792 26720 39164 26748
rect -39164 26452 -33792 26480
rect -39164 26388 -33876 26452
rect -33812 26388 -33792 26452
rect -39164 26372 -33792 26388
rect -39164 26308 -33876 26372
rect -33812 26308 -33792 26372
rect -39164 26292 -33792 26308
rect -39164 26228 -33876 26292
rect -33812 26228 -33792 26292
rect -39164 26212 -33792 26228
rect -39164 26148 -33876 26212
rect -33812 26148 -33792 26212
rect -39164 26132 -33792 26148
rect -39164 26068 -33876 26132
rect -33812 26068 -33792 26132
rect -39164 26052 -33792 26068
rect -39164 25988 -33876 26052
rect -33812 25988 -33792 26052
rect -39164 25972 -33792 25988
rect -39164 25908 -33876 25972
rect -33812 25908 -33792 25972
rect -39164 25892 -33792 25908
rect -39164 25828 -33876 25892
rect -33812 25828 -33792 25892
rect -39164 25812 -33792 25828
rect -39164 25748 -33876 25812
rect -33812 25748 -33792 25812
rect -39164 25732 -33792 25748
rect -39164 25668 -33876 25732
rect -33812 25668 -33792 25732
rect -39164 25652 -33792 25668
rect -39164 25588 -33876 25652
rect -33812 25588 -33792 25652
rect -39164 25572 -33792 25588
rect -39164 25508 -33876 25572
rect -33812 25508 -33792 25572
rect -39164 25492 -33792 25508
rect -39164 25428 -33876 25492
rect -33812 25428 -33792 25492
rect -39164 25412 -33792 25428
rect -39164 25348 -33876 25412
rect -33812 25348 -33792 25412
rect -39164 25332 -33792 25348
rect -39164 25268 -33876 25332
rect -33812 25268 -33792 25332
rect -39164 25252 -33792 25268
rect -39164 25188 -33876 25252
rect -33812 25188 -33792 25252
rect -39164 25172 -33792 25188
rect -39164 25108 -33876 25172
rect -33812 25108 -33792 25172
rect -39164 25092 -33792 25108
rect -39164 25028 -33876 25092
rect -33812 25028 -33792 25092
rect -39164 25012 -33792 25028
rect -39164 24948 -33876 25012
rect -33812 24948 -33792 25012
rect -39164 24932 -33792 24948
rect -39164 24868 -33876 24932
rect -33812 24868 -33792 24932
rect -39164 24852 -33792 24868
rect -39164 24788 -33876 24852
rect -33812 24788 -33792 24852
rect -39164 24772 -33792 24788
rect -39164 24708 -33876 24772
rect -33812 24708 -33792 24772
rect -39164 24692 -33792 24708
rect -39164 24628 -33876 24692
rect -33812 24628 -33792 24692
rect -39164 24612 -33792 24628
rect -39164 24548 -33876 24612
rect -33812 24548 -33792 24612
rect -39164 24532 -33792 24548
rect -39164 24468 -33876 24532
rect -33812 24468 -33792 24532
rect -39164 24452 -33792 24468
rect -39164 24388 -33876 24452
rect -33812 24388 -33792 24452
rect -39164 24372 -33792 24388
rect -39164 24308 -33876 24372
rect -33812 24308 -33792 24372
rect -39164 24292 -33792 24308
rect -39164 24228 -33876 24292
rect -33812 24228 -33792 24292
rect -39164 24212 -33792 24228
rect -39164 24148 -33876 24212
rect -33812 24148 -33792 24212
rect -39164 24132 -33792 24148
rect -39164 24068 -33876 24132
rect -33812 24068 -33792 24132
rect -39164 24052 -33792 24068
rect -39164 23988 -33876 24052
rect -33812 23988 -33792 24052
rect -39164 23972 -33792 23988
rect -39164 23908 -33876 23972
rect -33812 23908 -33792 23972
rect -39164 23892 -33792 23908
rect -39164 23828 -33876 23892
rect -33812 23828 -33792 23892
rect -39164 23812 -33792 23828
rect -39164 23748 -33876 23812
rect -33812 23748 -33792 23812
rect -39164 23732 -33792 23748
rect -39164 23668 -33876 23732
rect -33812 23668 -33792 23732
rect -39164 23652 -33792 23668
rect -39164 23588 -33876 23652
rect -33812 23588 -33792 23652
rect -39164 23572 -33792 23588
rect -39164 23508 -33876 23572
rect -33812 23508 -33792 23572
rect -39164 23492 -33792 23508
rect -39164 23428 -33876 23492
rect -33812 23428 -33792 23492
rect -39164 23412 -33792 23428
rect -39164 23348 -33876 23412
rect -33812 23348 -33792 23412
rect -39164 23332 -33792 23348
rect -39164 23268 -33876 23332
rect -33812 23268 -33792 23332
rect -39164 23252 -33792 23268
rect -39164 23188 -33876 23252
rect -33812 23188 -33792 23252
rect -39164 23172 -33792 23188
rect -39164 23108 -33876 23172
rect -33812 23108 -33792 23172
rect -39164 23092 -33792 23108
rect -39164 23028 -33876 23092
rect -33812 23028 -33792 23092
rect -39164 23012 -33792 23028
rect -39164 22948 -33876 23012
rect -33812 22948 -33792 23012
rect -39164 22932 -33792 22948
rect -39164 22868 -33876 22932
rect -33812 22868 -33792 22932
rect -39164 22852 -33792 22868
rect -39164 22788 -33876 22852
rect -33812 22788 -33792 22852
rect -39164 22772 -33792 22788
rect -39164 22708 -33876 22772
rect -33812 22708 -33792 22772
rect -39164 22692 -33792 22708
rect -39164 22628 -33876 22692
rect -33812 22628 -33792 22692
rect -39164 22612 -33792 22628
rect -39164 22548 -33876 22612
rect -33812 22548 -33792 22612
rect -39164 22532 -33792 22548
rect -39164 22468 -33876 22532
rect -33812 22468 -33792 22532
rect -39164 22452 -33792 22468
rect -39164 22388 -33876 22452
rect -33812 22388 -33792 22452
rect -39164 22372 -33792 22388
rect -39164 22308 -33876 22372
rect -33812 22308 -33792 22372
rect -39164 22292 -33792 22308
rect -39164 22228 -33876 22292
rect -33812 22228 -33792 22292
rect -39164 22212 -33792 22228
rect -39164 22148 -33876 22212
rect -33812 22148 -33792 22212
rect -39164 22132 -33792 22148
rect -39164 22068 -33876 22132
rect -33812 22068 -33792 22132
rect -39164 22052 -33792 22068
rect -39164 21988 -33876 22052
rect -33812 21988 -33792 22052
rect -39164 21972 -33792 21988
rect -39164 21908 -33876 21972
rect -33812 21908 -33792 21972
rect -39164 21892 -33792 21908
rect -39164 21828 -33876 21892
rect -33812 21828 -33792 21892
rect -39164 21812 -33792 21828
rect -39164 21748 -33876 21812
rect -33812 21748 -33792 21812
rect -39164 21732 -33792 21748
rect -39164 21668 -33876 21732
rect -33812 21668 -33792 21732
rect -39164 21652 -33792 21668
rect -39164 21588 -33876 21652
rect -33812 21588 -33792 21652
rect -39164 21572 -33792 21588
rect -39164 21508 -33876 21572
rect -33812 21508 -33792 21572
rect -39164 21492 -33792 21508
rect -39164 21428 -33876 21492
rect -33812 21428 -33792 21492
rect -39164 21400 -33792 21428
rect -33552 26452 -28180 26480
rect -33552 26388 -28264 26452
rect -28200 26388 -28180 26452
rect -33552 26372 -28180 26388
rect -33552 26308 -28264 26372
rect -28200 26308 -28180 26372
rect -33552 26292 -28180 26308
rect -33552 26228 -28264 26292
rect -28200 26228 -28180 26292
rect -33552 26212 -28180 26228
rect -33552 26148 -28264 26212
rect -28200 26148 -28180 26212
rect -33552 26132 -28180 26148
rect -33552 26068 -28264 26132
rect -28200 26068 -28180 26132
rect -33552 26052 -28180 26068
rect -33552 25988 -28264 26052
rect -28200 25988 -28180 26052
rect -33552 25972 -28180 25988
rect -33552 25908 -28264 25972
rect -28200 25908 -28180 25972
rect -33552 25892 -28180 25908
rect -33552 25828 -28264 25892
rect -28200 25828 -28180 25892
rect -33552 25812 -28180 25828
rect -33552 25748 -28264 25812
rect -28200 25748 -28180 25812
rect -33552 25732 -28180 25748
rect -33552 25668 -28264 25732
rect -28200 25668 -28180 25732
rect -33552 25652 -28180 25668
rect -33552 25588 -28264 25652
rect -28200 25588 -28180 25652
rect -33552 25572 -28180 25588
rect -33552 25508 -28264 25572
rect -28200 25508 -28180 25572
rect -33552 25492 -28180 25508
rect -33552 25428 -28264 25492
rect -28200 25428 -28180 25492
rect -33552 25412 -28180 25428
rect -33552 25348 -28264 25412
rect -28200 25348 -28180 25412
rect -33552 25332 -28180 25348
rect -33552 25268 -28264 25332
rect -28200 25268 -28180 25332
rect -33552 25252 -28180 25268
rect -33552 25188 -28264 25252
rect -28200 25188 -28180 25252
rect -33552 25172 -28180 25188
rect -33552 25108 -28264 25172
rect -28200 25108 -28180 25172
rect -33552 25092 -28180 25108
rect -33552 25028 -28264 25092
rect -28200 25028 -28180 25092
rect -33552 25012 -28180 25028
rect -33552 24948 -28264 25012
rect -28200 24948 -28180 25012
rect -33552 24932 -28180 24948
rect -33552 24868 -28264 24932
rect -28200 24868 -28180 24932
rect -33552 24852 -28180 24868
rect -33552 24788 -28264 24852
rect -28200 24788 -28180 24852
rect -33552 24772 -28180 24788
rect -33552 24708 -28264 24772
rect -28200 24708 -28180 24772
rect -33552 24692 -28180 24708
rect -33552 24628 -28264 24692
rect -28200 24628 -28180 24692
rect -33552 24612 -28180 24628
rect -33552 24548 -28264 24612
rect -28200 24548 -28180 24612
rect -33552 24532 -28180 24548
rect -33552 24468 -28264 24532
rect -28200 24468 -28180 24532
rect -33552 24452 -28180 24468
rect -33552 24388 -28264 24452
rect -28200 24388 -28180 24452
rect -33552 24372 -28180 24388
rect -33552 24308 -28264 24372
rect -28200 24308 -28180 24372
rect -33552 24292 -28180 24308
rect -33552 24228 -28264 24292
rect -28200 24228 -28180 24292
rect -33552 24212 -28180 24228
rect -33552 24148 -28264 24212
rect -28200 24148 -28180 24212
rect -33552 24132 -28180 24148
rect -33552 24068 -28264 24132
rect -28200 24068 -28180 24132
rect -33552 24052 -28180 24068
rect -33552 23988 -28264 24052
rect -28200 23988 -28180 24052
rect -33552 23972 -28180 23988
rect -33552 23908 -28264 23972
rect -28200 23908 -28180 23972
rect -33552 23892 -28180 23908
rect -33552 23828 -28264 23892
rect -28200 23828 -28180 23892
rect -33552 23812 -28180 23828
rect -33552 23748 -28264 23812
rect -28200 23748 -28180 23812
rect -33552 23732 -28180 23748
rect -33552 23668 -28264 23732
rect -28200 23668 -28180 23732
rect -33552 23652 -28180 23668
rect -33552 23588 -28264 23652
rect -28200 23588 -28180 23652
rect -33552 23572 -28180 23588
rect -33552 23508 -28264 23572
rect -28200 23508 -28180 23572
rect -33552 23492 -28180 23508
rect -33552 23428 -28264 23492
rect -28200 23428 -28180 23492
rect -33552 23412 -28180 23428
rect -33552 23348 -28264 23412
rect -28200 23348 -28180 23412
rect -33552 23332 -28180 23348
rect -33552 23268 -28264 23332
rect -28200 23268 -28180 23332
rect -33552 23252 -28180 23268
rect -33552 23188 -28264 23252
rect -28200 23188 -28180 23252
rect -33552 23172 -28180 23188
rect -33552 23108 -28264 23172
rect -28200 23108 -28180 23172
rect -33552 23092 -28180 23108
rect -33552 23028 -28264 23092
rect -28200 23028 -28180 23092
rect -33552 23012 -28180 23028
rect -33552 22948 -28264 23012
rect -28200 22948 -28180 23012
rect -33552 22932 -28180 22948
rect -33552 22868 -28264 22932
rect -28200 22868 -28180 22932
rect -33552 22852 -28180 22868
rect -33552 22788 -28264 22852
rect -28200 22788 -28180 22852
rect -33552 22772 -28180 22788
rect -33552 22708 -28264 22772
rect -28200 22708 -28180 22772
rect -33552 22692 -28180 22708
rect -33552 22628 -28264 22692
rect -28200 22628 -28180 22692
rect -33552 22612 -28180 22628
rect -33552 22548 -28264 22612
rect -28200 22548 -28180 22612
rect -33552 22532 -28180 22548
rect -33552 22468 -28264 22532
rect -28200 22468 -28180 22532
rect -33552 22452 -28180 22468
rect -33552 22388 -28264 22452
rect -28200 22388 -28180 22452
rect -33552 22372 -28180 22388
rect -33552 22308 -28264 22372
rect -28200 22308 -28180 22372
rect -33552 22292 -28180 22308
rect -33552 22228 -28264 22292
rect -28200 22228 -28180 22292
rect -33552 22212 -28180 22228
rect -33552 22148 -28264 22212
rect -28200 22148 -28180 22212
rect -33552 22132 -28180 22148
rect -33552 22068 -28264 22132
rect -28200 22068 -28180 22132
rect -33552 22052 -28180 22068
rect -33552 21988 -28264 22052
rect -28200 21988 -28180 22052
rect -33552 21972 -28180 21988
rect -33552 21908 -28264 21972
rect -28200 21908 -28180 21972
rect -33552 21892 -28180 21908
rect -33552 21828 -28264 21892
rect -28200 21828 -28180 21892
rect -33552 21812 -28180 21828
rect -33552 21748 -28264 21812
rect -28200 21748 -28180 21812
rect -33552 21732 -28180 21748
rect -33552 21668 -28264 21732
rect -28200 21668 -28180 21732
rect -33552 21652 -28180 21668
rect -33552 21588 -28264 21652
rect -28200 21588 -28180 21652
rect -33552 21572 -28180 21588
rect -33552 21508 -28264 21572
rect -28200 21508 -28180 21572
rect -33552 21492 -28180 21508
rect -33552 21428 -28264 21492
rect -28200 21428 -28180 21492
rect -33552 21400 -28180 21428
rect -27940 26452 -22568 26480
rect -27940 26388 -22652 26452
rect -22588 26388 -22568 26452
rect -27940 26372 -22568 26388
rect -27940 26308 -22652 26372
rect -22588 26308 -22568 26372
rect -27940 26292 -22568 26308
rect -27940 26228 -22652 26292
rect -22588 26228 -22568 26292
rect -27940 26212 -22568 26228
rect -27940 26148 -22652 26212
rect -22588 26148 -22568 26212
rect -27940 26132 -22568 26148
rect -27940 26068 -22652 26132
rect -22588 26068 -22568 26132
rect -27940 26052 -22568 26068
rect -27940 25988 -22652 26052
rect -22588 25988 -22568 26052
rect -27940 25972 -22568 25988
rect -27940 25908 -22652 25972
rect -22588 25908 -22568 25972
rect -27940 25892 -22568 25908
rect -27940 25828 -22652 25892
rect -22588 25828 -22568 25892
rect -27940 25812 -22568 25828
rect -27940 25748 -22652 25812
rect -22588 25748 -22568 25812
rect -27940 25732 -22568 25748
rect -27940 25668 -22652 25732
rect -22588 25668 -22568 25732
rect -27940 25652 -22568 25668
rect -27940 25588 -22652 25652
rect -22588 25588 -22568 25652
rect -27940 25572 -22568 25588
rect -27940 25508 -22652 25572
rect -22588 25508 -22568 25572
rect -27940 25492 -22568 25508
rect -27940 25428 -22652 25492
rect -22588 25428 -22568 25492
rect -27940 25412 -22568 25428
rect -27940 25348 -22652 25412
rect -22588 25348 -22568 25412
rect -27940 25332 -22568 25348
rect -27940 25268 -22652 25332
rect -22588 25268 -22568 25332
rect -27940 25252 -22568 25268
rect -27940 25188 -22652 25252
rect -22588 25188 -22568 25252
rect -27940 25172 -22568 25188
rect -27940 25108 -22652 25172
rect -22588 25108 -22568 25172
rect -27940 25092 -22568 25108
rect -27940 25028 -22652 25092
rect -22588 25028 -22568 25092
rect -27940 25012 -22568 25028
rect -27940 24948 -22652 25012
rect -22588 24948 -22568 25012
rect -27940 24932 -22568 24948
rect -27940 24868 -22652 24932
rect -22588 24868 -22568 24932
rect -27940 24852 -22568 24868
rect -27940 24788 -22652 24852
rect -22588 24788 -22568 24852
rect -27940 24772 -22568 24788
rect -27940 24708 -22652 24772
rect -22588 24708 -22568 24772
rect -27940 24692 -22568 24708
rect -27940 24628 -22652 24692
rect -22588 24628 -22568 24692
rect -27940 24612 -22568 24628
rect -27940 24548 -22652 24612
rect -22588 24548 -22568 24612
rect -27940 24532 -22568 24548
rect -27940 24468 -22652 24532
rect -22588 24468 -22568 24532
rect -27940 24452 -22568 24468
rect -27940 24388 -22652 24452
rect -22588 24388 -22568 24452
rect -27940 24372 -22568 24388
rect -27940 24308 -22652 24372
rect -22588 24308 -22568 24372
rect -27940 24292 -22568 24308
rect -27940 24228 -22652 24292
rect -22588 24228 -22568 24292
rect -27940 24212 -22568 24228
rect -27940 24148 -22652 24212
rect -22588 24148 -22568 24212
rect -27940 24132 -22568 24148
rect -27940 24068 -22652 24132
rect -22588 24068 -22568 24132
rect -27940 24052 -22568 24068
rect -27940 23988 -22652 24052
rect -22588 23988 -22568 24052
rect -27940 23972 -22568 23988
rect -27940 23908 -22652 23972
rect -22588 23908 -22568 23972
rect -27940 23892 -22568 23908
rect -27940 23828 -22652 23892
rect -22588 23828 -22568 23892
rect -27940 23812 -22568 23828
rect -27940 23748 -22652 23812
rect -22588 23748 -22568 23812
rect -27940 23732 -22568 23748
rect -27940 23668 -22652 23732
rect -22588 23668 -22568 23732
rect -27940 23652 -22568 23668
rect -27940 23588 -22652 23652
rect -22588 23588 -22568 23652
rect -27940 23572 -22568 23588
rect -27940 23508 -22652 23572
rect -22588 23508 -22568 23572
rect -27940 23492 -22568 23508
rect -27940 23428 -22652 23492
rect -22588 23428 -22568 23492
rect -27940 23412 -22568 23428
rect -27940 23348 -22652 23412
rect -22588 23348 -22568 23412
rect -27940 23332 -22568 23348
rect -27940 23268 -22652 23332
rect -22588 23268 -22568 23332
rect -27940 23252 -22568 23268
rect -27940 23188 -22652 23252
rect -22588 23188 -22568 23252
rect -27940 23172 -22568 23188
rect -27940 23108 -22652 23172
rect -22588 23108 -22568 23172
rect -27940 23092 -22568 23108
rect -27940 23028 -22652 23092
rect -22588 23028 -22568 23092
rect -27940 23012 -22568 23028
rect -27940 22948 -22652 23012
rect -22588 22948 -22568 23012
rect -27940 22932 -22568 22948
rect -27940 22868 -22652 22932
rect -22588 22868 -22568 22932
rect -27940 22852 -22568 22868
rect -27940 22788 -22652 22852
rect -22588 22788 -22568 22852
rect -27940 22772 -22568 22788
rect -27940 22708 -22652 22772
rect -22588 22708 -22568 22772
rect -27940 22692 -22568 22708
rect -27940 22628 -22652 22692
rect -22588 22628 -22568 22692
rect -27940 22612 -22568 22628
rect -27940 22548 -22652 22612
rect -22588 22548 -22568 22612
rect -27940 22532 -22568 22548
rect -27940 22468 -22652 22532
rect -22588 22468 -22568 22532
rect -27940 22452 -22568 22468
rect -27940 22388 -22652 22452
rect -22588 22388 -22568 22452
rect -27940 22372 -22568 22388
rect -27940 22308 -22652 22372
rect -22588 22308 -22568 22372
rect -27940 22292 -22568 22308
rect -27940 22228 -22652 22292
rect -22588 22228 -22568 22292
rect -27940 22212 -22568 22228
rect -27940 22148 -22652 22212
rect -22588 22148 -22568 22212
rect -27940 22132 -22568 22148
rect -27940 22068 -22652 22132
rect -22588 22068 -22568 22132
rect -27940 22052 -22568 22068
rect -27940 21988 -22652 22052
rect -22588 21988 -22568 22052
rect -27940 21972 -22568 21988
rect -27940 21908 -22652 21972
rect -22588 21908 -22568 21972
rect -27940 21892 -22568 21908
rect -27940 21828 -22652 21892
rect -22588 21828 -22568 21892
rect -27940 21812 -22568 21828
rect -27940 21748 -22652 21812
rect -22588 21748 -22568 21812
rect -27940 21732 -22568 21748
rect -27940 21668 -22652 21732
rect -22588 21668 -22568 21732
rect -27940 21652 -22568 21668
rect -27940 21588 -22652 21652
rect -22588 21588 -22568 21652
rect -27940 21572 -22568 21588
rect -27940 21508 -22652 21572
rect -22588 21508 -22568 21572
rect -27940 21492 -22568 21508
rect -27940 21428 -22652 21492
rect -22588 21428 -22568 21492
rect -27940 21400 -22568 21428
rect -22328 26452 -16956 26480
rect -22328 26388 -17040 26452
rect -16976 26388 -16956 26452
rect -22328 26372 -16956 26388
rect -22328 26308 -17040 26372
rect -16976 26308 -16956 26372
rect -22328 26292 -16956 26308
rect -22328 26228 -17040 26292
rect -16976 26228 -16956 26292
rect -22328 26212 -16956 26228
rect -22328 26148 -17040 26212
rect -16976 26148 -16956 26212
rect -22328 26132 -16956 26148
rect -22328 26068 -17040 26132
rect -16976 26068 -16956 26132
rect -22328 26052 -16956 26068
rect -22328 25988 -17040 26052
rect -16976 25988 -16956 26052
rect -22328 25972 -16956 25988
rect -22328 25908 -17040 25972
rect -16976 25908 -16956 25972
rect -22328 25892 -16956 25908
rect -22328 25828 -17040 25892
rect -16976 25828 -16956 25892
rect -22328 25812 -16956 25828
rect -22328 25748 -17040 25812
rect -16976 25748 -16956 25812
rect -22328 25732 -16956 25748
rect -22328 25668 -17040 25732
rect -16976 25668 -16956 25732
rect -22328 25652 -16956 25668
rect -22328 25588 -17040 25652
rect -16976 25588 -16956 25652
rect -22328 25572 -16956 25588
rect -22328 25508 -17040 25572
rect -16976 25508 -16956 25572
rect -22328 25492 -16956 25508
rect -22328 25428 -17040 25492
rect -16976 25428 -16956 25492
rect -22328 25412 -16956 25428
rect -22328 25348 -17040 25412
rect -16976 25348 -16956 25412
rect -22328 25332 -16956 25348
rect -22328 25268 -17040 25332
rect -16976 25268 -16956 25332
rect -22328 25252 -16956 25268
rect -22328 25188 -17040 25252
rect -16976 25188 -16956 25252
rect -22328 25172 -16956 25188
rect -22328 25108 -17040 25172
rect -16976 25108 -16956 25172
rect -22328 25092 -16956 25108
rect -22328 25028 -17040 25092
rect -16976 25028 -16956 25092
rect -22328 25012 -16956 25028
rect -22328 24948 -17040 25012
rect -16976 24948 -16956 25012
rect -22328 24932 -16956 24948
rect -22328 24868 -17040 24932
rect -16976 24868 -16956 24932
rect -22328 24852 -16956 24868
rect -22328 24788 -17040 24852
rect -16976 24788 -16956 24852
rect -22328 24772 -16956 24788
rect -22328 24708 -17040 24772
rect -16976 24708 -16956 24772
rect -22328 24692 -16956 24708
rect -22328 24628 -17040 24692
rect -16976 24628 -16956 24692
rect -22328 24612 -16956 24628
rect -22328 24548 -17040 24612
rect -16976 24548 -16956 24612
rect -22328 24532 -16956 24548
rect -22328 24468 -17040 24532
rect -16976 24468 -16956 24532
rect -22328 24452 -16956 24468
rect -22328 24388 -17040 24452
rect -16976 24388 -16956 24452
rect -22328 24372 -16956 24388
rect -22328 24308 -17040 24372
rect -16976 24308 -16956 24372
rect -22328 24292 -16956 24308
rect -22328 24228 -17040 24292
rect -16976 24228 -16956 24292
rect -22328 24212 -16956 24228
rect -22328 24148 -17040 24212
rect -16976 24148 -16956 24212
rect -22328 24132 -16956 24148
rect -22328 24068 -17040 24132
rect -16976 24068 -16956 24132
rect -22328 24052 -16956 24068
rect -22328 23988 -17040 24052
rect -16976 23988 -16956 24052
rect -22328 23972 -16956 23988
rect -22328 23908 -17040 23972
rect -16976 23908 -16956 23972
rect -22328 23892 -16956 23908
rect -22328 23828 -17040 23892
rect -16976 23828 -16956 23892
rect -22328 23812 -16956 23828
rect -22328 23748 -17040 23812
rect -16976 23748 -16956 23812
rect -22328 23732 -16956 23748
rect -22328 23668 -17040 23732
rect -16976 23668 -16956 23732
rect -22328 23652 -16956 23668
rect -22328 23588 -17040 23652
rect -16976 23588 -16956 23652
rect -22328 23572 -16956 23588
rect -22328 23508 -17040 23572
rect -16976 23508 -16956 23572
rect -22328 23492 -16956 23508
rect -22328 23428 -17040 23492
rect -16976 23428 -16956 23492
rect -22328 23412 -16956 23428
rect -22328 23348 -17040 23412
rect -16976 23348 -16956 23412
rect -22328 23332 -16956 23348
rect -22328 23268 -17040 23332
rect -16976 23268 -16956 23332
rect -22328 23252 -16956 23268
rect -22328 23188 -17040 23252
rect -16976 23188 -16956 23252
rect -22328 23172 -16956 23188
rect -22328 23108 -17040 23172
rect -16976 23108 -16956 23172
rect -22328 23092 -16956 23108
rect -22328 23028 -17040 23092
rect -16976 23028 -16956 23092
rect -22328 23012 -16956 23028
rect -22328 22948 -17040 23012
rect -16976 22948 -16956 23012
rect -22328 22932 -16956 22948
rect -22328 22868 -17040 22932
rect -16976 22868 -16956 22932
rect -22328 22852 -16956 22868
rect -22328 22788 -17040 22852
rect -16976 22788 -16956 22852
rect -22328 22772 -16956 22788
rect -22328 22708 -17040 22772
rect -16976 22708 -16956 22772
rect -22328 22692 -16956 22708
rect -22328 22628 -17040 22692
rect -16976 22628 -16956 22692
rect -22328 22612 -16956 22628
rect -22328 22548 -17040 22612
rect -16976 22548 -16956 22612
rect -22328 22532 -16956 22548
rect -22328 22468 -17040 22532
rect -16976 22468 -16956 22532
rect -22328 22452 -16956 22468
rect -22328 22388 -17040 22452
rect -16976 22388 -16956 22452
rect -22328 22372 -16956 22388
rect -22328 22308 -17040 22372
rect -16976 22308 -16956 22372
rect -22328 22292 -16956 22308
rect -22328 22228 -17040 22292
rect -16976 22228 -16956 22292
rect -22328 22212 -16956 22228
rect -22328 22148 -17040 22212
rect -16976 22148 -16956 22212
rect -22328 22132 -16956 22148
rect -22328 22068 -17040 22132
rect -16976 22068 -16956 22132
rect -22328 22052 -16956 22068
rect -22328 21988 -17040 22052
rect -16976 21988 -16956 22052
rect -22328 21972 -16956 21988
rect -22328 21908 -17040 21972
rect -16976 21908 -16956 21972
rect -22328 21892 -16956 21908
rect -22328 21828 -17040 21892
rect -16976 21828 -16956 21892
rect -22328 21812 -16956 21828
rect -22328 21748 -17040 21812
rect -16976 21748 -16956 21812
rect -22328 21732 -16956 21748
rect -22328 21668 -17040 21732
rect -16976 21668 -16956 21732
rect -22328 21652 -16956 21668
rect -22328 21588 -17040 21652
rect -16976 21588 -16956 21652
rect -22328 21572 -16956 21588
rect -22328 21508 -17040 21572
rect -16976 21508 -16956 21572
rect -22328 21492 -16956 21508
rect -22328 21428 -17040 21492
rect -16976 21428 -16956 21492
rect -22328 21400 -16956 21428
rect -16716 26452 -11344 26480
rect -16716 26388 -11428 26452
rect -11364 26388 -11344 26452
rect -16716 26372 -11344 26388
rect -16716 26308 -11428 26372
rect -11364 26308 -11344 26372
rect -16716 26292 -11344 26308
rect -16716 26228 -11428 26292
rect -11364 26228 -11344 26292
rect -16716 26212 -11344 26228
rect -16716 26148 -11428 26212
rect -11364 26148 -11344 26212
rect -16716 26132 -11344 26148
rect -16716 26068 -11428 26132
rect -11364 26068 -11344 26132
rect -16716 26052 -11344 26068
rect -16716 25988 -11428 26052
rect -11364 25988 -11344 26052
rect -16716 25972 -11344 25988
rect -16716 25908 -11428 25972
rect -11364 25908 -11344 25972
rect -16716 25892 -11344 25908
rect -16716 25828 -11428 25892
rect -11364 25828 -11344 25892
rect -16716 25812 -11344 25828
rect -16716 25748 -11428 25812
rect -11364 25748 -11344 25812
rect -16716 25732 -11344 25748
rect -16716 25668 -11428 25732
rect -11364 25668 -11344 25732
rect -16716 25652 -11344 25668
rect -16716 25588 -11428 25652
rect -11364 25588 -11344 25652
rect -16716 25572 -11344 25588
rect -16716 25508 -11428 25572
rect -11364 25508 -11344 25572
rect -16716 25492 -11344 25508
rect -16716 25428 -11428 25492
rect -11364 25428 -11344 25492
rect -16716 25412 -11344 25428
rect -16716 25348 -11428 25412
rect -11364 25348 -11344 25412
rect -16716 25332 -11344 25348
rect -16716 25268 -11428 25332
rect -11364 25268 -11344 25332
rect -16716 25252 -11344 25268
rect -16716 25188 -11428 25252
rect -11364 25188 -11344 25252
rect -16716 25172 -11344 25188
rect -16716 25108 -11428 25172
rect -11364 25108 -11344 25172
rect -16716 25092 -11344 25108
rect -16716 25028 -11428 25092
rect -11364 25028 -11344 25092
rect -16716 25012 -11344 25028
rect -16716 24948 -11428 25012
rect -11364 24948 -11344 25012
rect -16716 24932 -11344 24948
rect -16716 24868 -11428 24932
rect -11364 24868 -11344 24932
rect -16716 24852 -11344 24868
rect -16716 24788 -11428 24852
rect -11364 24788 -11344 24852
rect -16716 24772 -11344 24788
rect -16716 24708 -11428 24772
rect -11364 24708 -11344 24772
rect -16716 24692 -11344 24708
rect -16716 24628 -11428 24692
rect -11364 24628 -11344 24692
rect -16716 24612 -11344 24628
rect -16716 24548 -11428 24612
rect -11364 24548 -11344 24612
rect -16716 24532 -11344 24548
rect -16716 24468 -11428 24532
rect -11364 24468 -11344 24532
rect -16716 24452 -11344 24468
rect -16716 24388 -11428 24452
rect -11364 24388 -11344 24452
rect -16716 24372 -11344 24388
rect -16716 24308 -11428 24372
rect -11364 24308 -11344 24372
rect -16716 24292 -11344 24308
rect -16716 24228 -11428 24292
rect -11364 24228 -11344 24292
rect -16716 24212 -11344 24228
rect -16716 24148 -11428 24212
rect -11364 24148 -11344 24212
rect -16716 24132 -11344 24148
rect -16716 24068 -11428 24132
rect -11364 24068 -11344 24132
rect -16716 24052 -11344 24068
rect -16716 23988 -11428 24052
rect -11364 23988 -11344 24052
rect -16716 23972 -11344 23988
rect -16716 23908 -11428 23972
rect -11364 23908 -11344 23972
rect -16716 23892 -11344 23908
rect -16716 23828 -11428 23892
rect -11364 23828 -11344 23892
rect -16716 23812 -11344 23828
rect -16716 23748 -11428 23812
rect -11364 23748 -11344 23812
rect -16716 23732 -11344 23748
rect -16716 23668 -11428 23732
rect -11364 23668 -11344 23732
rect -16716 23652 -11344 23668
rect -16716 23588 -11428 23652
rect -11364 23588 -11344 23652
rect -16716 23572 -11344 23588
rect -16716 23508 -11428 23572
rect -11364 23508 -11344 23572
rect -16716 23492 -11344 23508
rect -16716 23428 -11428 23492
rect -11364 23428 -11344 23492
rect -16716 23412 -11344 23428
rect -16716 23348 -11428 23412
rect -11364 23348 -11344 23412
rect -16716 23332 -11344 23348
rect -16716 23268 -11428 23332
rect -11364 23268 -11344 23332
rect -16716 23252 -11344 23268
rect -16716 23188 -11428 23252
rect -11364 23188 -11344 23252
rect -16716 23172 -11344 23188
rect -16716 23108 -11428 23172
rect -11364 23108 -11344 23172
rect -16716 23092 -11344 23108
rect -16716 23028 -11428 23092
rect -11364 23028 -11344 23092
rect -16716 23012 -11344 23028
rect -16716 22948 -11428 23012
rect -11364 22948 -11344 23012
rect -16716 22932 -11344 22948
rect -16716 22868 -11428 22932
rect -11364 22868 -11344 22932
rect -16716 22852 -11344 22868
rect -16716 22788 -11428 22852
rect -11364 22788 -11344 22852
rect -16716 22772 -11344 22788
rect -16716 22708 -11428 22772
rect -11364 22708 -11344 22772
rect -16716 22692 -11344 22708
rect -16716 22628 -11428 22692
rect -11364 22628 -11344 22692
rect -16716 22612 -11344 22628
rect -16716 22548 -11428 22612
rect -11364 22548 -11344 22612
rect -16716 22532 -11344 22548
rect -16716 22468 -11428 22532
rect -11364 22468 -11344 22532
rect -16716 22452 -11344 22468
rect -16716 22388 -11428 22452
rect -11364 22388 -11344 22452
rect -16716 22372 -11344 22388
rect -16716 22308 -11428 22372
rect -11364 22308 -11344 22372
rect -16716 22292 -11344 22308
rect -16716 22228 -11428 22292
rect -11364 22228 -11344 22292
rect -16716 22212 -11344 22228
rect -16716 22148 -11428 22212
rect -11364 22148 -11344 22212
rect -16716 22132 -11344 22148
rect -16716 22068 -11428 22132
rect -11364 22068 -11344 22132
rect -16716 22052 -11344 22068
rect -16716 21988 -11428 22052
rect -11364 21988 -11344 22052
rect -16716 21972 -11344 21988
rect -16716 21908 -11428 21972
rect -11364 21908 -11344 21972
rect -16716 21892 -11344 21908
rect -16716 21828 -11428 21892
rect -11364 21828 -11344 21892
rect -16716 21812 -11344 21828
rect -16716 21748 -11428 21812
rect -11364 21748 -11344 21812
rect -16716 21732 -11344 21748
rect -16716 21668 -11428 21732
rect -11364 21668 -11344 21732
rect -16716 21652 -11344 21668
rect -16716 21588 -11428 21652
rect -11364 21588 -11344 21652
rect -16716 21572 -11344 21588
rect -16716 21508 -11428 21572
rect -11364 21508 -11344 21572
rect -16716 21492 -11344 21508
rect -16716 21428 -11428 21492
rect -11364 21428 -11344 21492
rect -16716 21400 -11344 21428
rect -11104 26452 -5732 26480
rect -11104 26388 -5816 26452
rect -5752 26388 -5732 26452
rect -11104 26372 -5732 26388
rect -11104 26308 -5816 26372
rect -5752 26308 -5732 26372
rect -11104 26292 -5732 26308
rect -11104 26228 -5816 26292
rect -5752 26228 -5732 26292
rect -11104 26212 -5732 26228
rect -11104 26148 -5816 26212
rect -5752 26148 -5732 26212
rect -11104 26132 -5732 26148
rect -11104 26068 -5816 26132
rect -5752 26068 -5732 26132
rect -11104 26052 -5732 26068
rect -11104 25988 -5816 26052
rect -5752 25988 -5732 26052
rect -11104 25972 -5732 25988
rect -11104 25908 -5816 25972
rect -5752 25908 -5732 25972
rect -11104 25892 -5732 25908
rect -11104 25828 -5816 25892
rect -5752 25828 -5732 25892
rect -11104 25812 -5732 25828
rect -11104 25748 -5816 25812
rect -5752 25748 -5732 25812
rect -11104 25732 -5732 25748
rect -11104 25668 -5816 25732
rect -5752 25668 -5732 25732
rect -11104 25652 -5732 25668
rect -11104 25588 -5816 25652
rect -5752 25588 -5732 25652
rect -11104 25572 -5732 25588
rect -11104 25508 -5816 25572
rect -5752 25508 -5732 25572
rect -11104 25492 -5732 25508
rect -11104 25428 -5816 25492
rect -5752 25428 -5732 25492
rect -11104 25412 -5732 25428
rect -11104 25348 -5816 25412
rect -5752 25348 -5732 25412
rect -11104 25332 -5732 25348
rect -11104 25268 -5816 25332
rect -5752 25268 -5732 25332
rect -11104 25252 -5732 25268
rect -11104 25188 -5816 25252
rect -5752 25188 -5732 25252
rect -11104 25172 -5732 25188
rect -11104 25108 -5816 25172
rect -5752 25108 -5732 25172
rect -11104 25092 -5732 25108
rect -11104 25028 -5816 25092
rect -5752 25028 -5732 25092
rect -11104 25012 -5732 25028
rect -11104 24948 -5816 25012
rect -5752 24948 -5732 25012
rect -11104 24932 -5732 24948
rect -11104 24868 -5816 24932
rect -5752 24868 -5732 24932
rect -11104 24852 -5732 24868
rect -11104 24788 -5816 24852
rect -5752 24788 -5732 24852
rect -11104 24772 -5732 24788
rect -11104 24708 -5816 24772
rect -5752 24708 -5732 24772
rect -11104 24692 -5732 24708
rect -11104 24628 -5816 24692
rect -5752 24628 -5732 24692
rect -11104 24612 -5732 24628
rect -11104 24548 -5816 24612
rect -5752 24548 -5732 24612
rect -11104 24532 -5732 24548
rect -11104 24468 -5816 24532
rect -5752 24468 -5732 24532
rect -11104 24452 -5732 24468
rect -11104 24388 -5816 24452
rect -5752 24388 -5732 24452
rect -11104 24372 -5732 24388
rect -11104 24308 -5816 24372
rect -5752 24308 -5732 24372
rect -11104 24292 -5732 24308
rect -11104 24228 -5816 24292
rect -5752 24228 -5732 24292
rect -11104 24212 -5732 24228
rect -11104 24148 -5816 24212
rect -5752 24148 -5732 24212
rect -11104 24132 -5732 24148
rect -11104 24068 -5816 24132
rect -5752 24068 -5732 24132
rect -11104 24052 -5732 24068
rect -11104 23988 -5816 24052
rect -5752 23988 -5732 24052
rect -11104 23972 -5732 23988
rect -11104 23908 -5816 23972
rect -5752 23908 -5732 23972
rect -11104 23892 -5732 23908
rect -11104 23828 -5816 23892
rect -5752 23828 -5732 23892
rect -11104 23812 -5732 23828
rect -11104 23748 -5816 23812
rect -5752 23748 -5732 23812
rect -11104 23732 -5732 23748
rect -11104 23668 -5816 23732
rect -5752 23668 -5732 23732
rect -11104 23652 -5732 23668
rect -11104 23588 -5816 23652
rect -5752 23588 -5732 23652
rect -11104 23572 -5732 23588
rect -11104 23508 -5816 23572
rect -5752 23508 -5732 23572
rect -11104 23492 -5732 23508
rect -11104 23428 -5816 23492
rect -5752 23428 -5732 23492
rect -11104 23412 -5732 23428
rect -11104 23348 -5816 23412
rect -5752 23348 -5732 23412
rect -11104 23332 -5732 23348
rect -11104 23268 -5816 23332
rect -5752 23268 -5732 23332
rect -11104 23252 -5732 23268
rect -11104 23188 -5816 23252
rect -5752 23188 -5732 23252
rect -11104 23172 -5732 23188
rect -11104 23108 -5816 23172
rect -5752 23108 -5732 23172
rect -11104 23092 -5732 23108
rect -11104 23028 -5816 23092
rect -5752 23028 -5732 23092
rect -11104 23012 -5732 23028
rect -11104 22948 -5816 23012
rect -5752 22948 -5732 23012
rect -11104 22932 -5732 22948
rect -11104 22868 -5816 22932
rect -5752 22868 -5732 22932
rect -11104 22852 -5732 22868
rect -11104 22788 -5816 22852
rect -5752 22788 -5732 22852
rect -11104 22772 -5732 22788
rect -11104 22708 -5816 22772
rect -5752 22708 -5732 22772
rect -11104 22692 -5732 22708
rect -11104 22628 -5816 22692
rect -5752 22628 -5732 22692
rect -11104 22612 -5732 22628
rect -11104 22548 -5816 22612
rect -5752 22548 -5732 22612
rect -11104 22532 -5732 22548
rect -11104 22468 -5816 22532
rect -5752 22468 -5732 22532
rect -11104 22452 -5732 22468
rect -11104 22388 -5816 22452
rect -5752 22388 -5732 22452
rect -11104 22372 -5732 22388
rect -11104 22308 -5816 22372
rect -5752 22308 -5732 22372
rect -11104 22292 -5732 22308
rect -11104 22228 -5816 22292
rect -5752 22228 -5732 22292
rect -11104 22212 -5732 22228
rect -11104 22148 -5816 22212
rect -5752 22148 -5732 22212
rect -11104 22132 -5732 22148
rect -11104 22068 -5816 22132
rect -5752 22068 -5732 22132
rect -11104 22052 -5732 22068
rect -11104 21988 -5816 22052
rect -5752 21988 -5732 22052
rect -11104 21972 -5732 21988
rect -11104 21908 -5816 21972
rect -5752 21908 -5732 21972
rect -11104 21892 -5732 21908
rect -11104 21828 -5816 21892
rect -5752 21828 -5732 21892
rect -11104 21812 -5732 21828
rect -11104 21748 -5816 21812
rect -5752 21748 -5732 21812
rect -11104 21732 -5732 21748
rect -11104 21668 -5816 21732
rect -5752 21668 -5732 21732
rect -11104 21652 -5732 21668
rect -11104 21588 -5816 21652
rect -5752 21588 -5732 21652
rect -11104 21572 -5732 21588
rect -11104 21508 -5816 21572
rect -5752 21508 -5732 21572
rect -11104 21492 -5732 21508
rect -11104 21428 -5816 21492
rect -5752 21428 -5732 21492
rect -11104 21400 -5732 21428
rect -5492 26452 -120 26480
rect -5492 26388 -204 26452
rect -140 26388 -120 26452
rect -5492 26372 -120 26388
rect -5492 26308 -204 26372
rect -140 26308 -120 26372
rect -5492 26292 -120 26308
rect -5492 26228 -204 26292
rect -140 26228 -120 26292
rect -5492 26212 -120 26228
rect -5492 26148 -204 26212
rect -140 26148 -120 26212
rect -5492 26132 -120 26148
rect -5492 26068 -204 26132
rect -140 26068 -120 26132
rect -5492 26052 -120 26068
rect -5492 25988 -204 26052
rect -140 25988 -120 26052
rect -5492 25972 -120 25988
rect -5492 25908 -204 25972
rect -140 25908 -120 25972
rect -5492 25892 -120 25908
rect -5492 25828 -204 25892
rect -140 25828 -120 25892
rect -5492 25812 -120 25828
rect -5492 25748 -204 25812
rect -140 25748 -120 25812
rect -5492 25732 -120 25748
rect -5492 25668 -204 25732
rect -140 25668 -120 25732
rect -5492 25652 -120 25668
rect -5492 25588 -204 25652
rect -140 25588 -120 25652
rect -5492 25572 -120 25588
rect -5492 25508 -204 25572
rect -140 25508 -120 25572
rect -5492 25492 -120 25508
rect -5492 25428 -204 25492
rect -140 25428 -120 25492
rect -5492 25412 -120 25428
rect -5492 25348 -204 25412
rect -140 25348 -120 25412
rect -5492 25332 -120 25348
rect -5492 25268 -204 25332
rect -140 25268 -120 25332
rect -5492 25252 -120 25268
rect -5492 25188 -204 25252
rect -140 25188 -120 25252
rect -5492 25172 -120 25188
rect -5492 25108 -204 25172
rect -140 25108 -120 25172
rect -5492 25092 -120 25108
rect -5492 25028 -204 25092
rect -140 25028 -120 25092
rect -5492 25012 -120 25028
rect -5492 24948 -204 25012
rect -140 24948 -120 25012
rect -5492 24932 -120 24948
rect -5492 24868 -204 24932
rect -140 24868 -120 24932
rect -5492 24852 -120 24868
rect -5492 24788 -204 24852
rect -140 24788 -120 24852
rect -5492 24772 -120 24788
rect -5492 24708 -204 24772
rect -140 24708 -120 24772
rect -5492 24692 -120 24708
rect -5492 24628 -204 24692
rect -140 24628 -120 24692
rect -5492 24612 -120 24628
rect -5492 24548 -204 24612
rect -140 24548 -120 24612
rect -5492 24532 -120 24548
rect -5492 24468 -204 24532
rect -140 24468 -120 24532
rect -5492 24452 -120 24468
rect -5492 24388 -204 24452
rect -140 24388 -120 24452
rect -5492 24372 -120 24388
rect -5492 24308 -204 24372
rect -140 24308 -120 24372
rect -5492 24292 -120 24308
rect -5492 24228 -204 24292
rect -140 24228 -120 24292
rect -5492 24212 -120 24228
rect -5492 24148 -204 24212
rect -140 24148 -120 24212
rect -5492 24132 -120 24148
rect -5492 24068 -204 24132
rect -140 24068 -120 24132
rect -5492 24052 -120 24068
rect -5492 23988 -204 24052
rect -140 23988 -120 24052
rect -5492 23972 -120 23988
rect -5492 23908 -204 23972
rect -140 23908 -120 23972
rect -5492 23892 -120 23908
rect -5492 23828 -204 23892
rect -140 23828 -120 23892
rect -5492 23812 -120 23828
rect -5492 23748 -204 23812
rect -140 23748 -120 23812
rect -5492 23732 -120 23748
rect -5492 23668 -204 23732
rect -140 23668 -120 23732
rect -5492 23652 -120 23668
rect -5492 23588 -204 23652
rect -140 23588 -120 23652
rect -5492 23572 -120 23588
rect -5492 23508 -204 23572
rect -140 23508 -120 23572
rect -5492 23492 -120 23508
rect -5492 23428 -204 23492
rect -140 23428 -120 23492
rect -5492 23412 -120 23428
rect -5492 23348 -204 23412
rect -140 23348 -120 23412
rect -5492 23332 -120 23348
rect -5492 23268 -204 23332
rect -140 23268 -120 23332
rect -5492 23252 -120 23268
rect -5492 23188 -204 23252
rect -140 23188 -120 23252
rect -5492 23172 -120 23188
rect -5492 23108 -204 23172
rect -140 23108 -120 23172
rect -5492 23092 -120 23108
rect -5492 23028 -204 23092
rect -140 23028 -120 23092
rect -5492 23012 -120 23028
rect -5492 22948 -204 23012
rect -140 22948 -120 23012
rect -5492 22932 -120 22948
rect -5492 22868 -204 22932
rect -140 22868 -120 22932
rect -5492 22852 -120 22868
rect -5492 22788 -204 22852
rect -140 22788 -120 22852
rect -5492 22772 -120 22788
rect -5492 22708 -204 22772
rect -140 22708 -120 22772
rect -5492 22692 -120 22708
rect -5492 22628 -204 22692
rect -140 22628 -120 22692
rect -5492 22612 -120 22628
rect -5492 22548 -204 22612
rect -140 22548 -120 22612
rect -5492 22532 -120 22548
rect -5492 22468 -204 22532
rect -140 22468 -120 22532
rect -5492 22452 -120 22468
rect -5492 22388 -204 22452
rect -140 22388 -120 22452
rect -5492 22372 -120 22388
rect -5492 22308 -204 22372
rect -140 22308 -120 22372
rect -5492 22292 -120 22308
rect -5492 22228 -204 22292
rect -140 22228 -120 22292
rect -5492 22212 -120 22228
rect -5492 22148 -204 22212
rect -140 22148 -120 22212
rect -5492 22132 -120 22148
rect -5492 22068 -204 22132
rect -140 22068 -120 22132
rect -5492 22052 -120 22068
rect -5492 21988 -204 22052
rect -140 21988 -120 22052
rect -5492 21972 -120 21988
rect -5492 21908 -204 21972
rect -140 21908 -120 21972
rect -5492 21892 -120 21908
rect -5492 21828 -204 21892
rect -140 21828 -120 21892
rect -5492 21812 -120 21828
rect -5492 21748 -204 21812
rect -140 21748 -120 21812
rect -5492 21732 -120 21748
rect -5492 21668 -204 21732
rect -140 21668 -120 21732
rect -5492 21652 -120 21668
rect -5492 21588 -204 21652
rect -140 21588 -120 21652
rect -5492 21572 -120 21588
rect -5492 21508 -204 21572
rect -140 21508 -120 21572
rect -5492 21492 -120 21508
rect -5492 21428 -204 21492
rect -140 21428 -120 21492
rect -5492 21400 -120 21428
rect 120 26452 5492 26480
rect 120 26388 5408 26452
rect 5472 26388 5492 26452
rect 120 26372 5492 26388
rect 120 26308 5408 26372
rect 5472 26308 5492 26372
rect 120 26292 5492 26308
rect 120 26228 5408 26292
rect 5472 26228 5492 26292
rect 120 26212 5492 26228
rect 120 26148 5408 26212
rect 5472 26148 5492 26212
rect 120 26132 5492 26148
rect 120 26068 5408 26132
rect 5472 26068 5492 26132
rect 120 26052 5492 26068
rect 120 25988 5408 26052
rect 5472 25988 5492 26052
rect 120 25972 5492 25988
rect 120 25908 5408 25972
rect 5472 25908 5492 25972
rect 120 25892 5492 25908
rect 120 25828 5408 25892
rect 5472 25828 5492 25892
rect 120 25812 5492 25828
rect 120 25748 5408 25812
rect 5472 25748 5492 25812
rect 120 25732 5492 25748
rect 120 25668 5408 25732
rect 5472 25668 5492 25732
rect 120 25652 5492 25668
rect 120 25588 5408 25652
rect 5472 25588 5492 25652
rect 120 25572 5492 25588
rect 120 25508 5408 25572
rect 5472 25508 5492 25572
rect 120 25492 5492 25508
rect 120 25428 5408 25492
rect 5472 25428 5492 25492
rect 120 25412 5492 25428
rect 120 25348 5408 25412
rect 5472 25348 5492 25412
rect 120 25332 5492 25348
rect 120 25268 5408 25332
rect 5472 25268 5492 25332
rect 120 25252 5492 25268
rect 120 25188 5408 25252
rect 5472 25188 5492 25252
rect 120 25172 5492 25188
rect 120 25108 5408 25172
rect 5472 25108 5492 25172
rect 120 25092 5492 25108
rect 120 25028 5408 25092
rect 5472 25028 5492 25092
rect 120 25012 5492 25028
rect 120 24948 5408 25012
rect 5472 24948 5492 25012
rect 120 24932 5492 24948
rect 120 24868 5408 24932
rect 5472 24868 5492 24932
rect 120 24852 5492 24868
rect 120 24788 5408 24852
rect 5472 24788 5492 24852
rect 120 24772 5492 24788
rect 120 24708 5408 24772
rect 5472 24708 5492 24772
rect 120 24692 5492 24708
rect 120 24628 5408 24692
rect 5472 24628 5492 24692
rect 120 24612 5492 24628
rect 120 24548 5408 24612
rect 5472 24548 5492 24612
rect 120 24532 5492 24548
rect 120 24468 5408 24532
rect 5472 24468 5492 24532
rect 120 24452 5492 24468
rect 120 24388 5408 24452
rect 5472 24388 5492 24452
rect 120 24372 5492 24388
rect 120 24308 5408 24372
rect 5472 24308 5492 24372
rect 120 24292 5492 24308
rect 120 24228 5408 24292
rect 5472 24228 5492 24292
rect 120 24212 5492 24228
rect 120 24148 5408 24212
rect 5472 24148 5492 24212
rect 120 24132 5492 24148
rect 120 24068 5408 24132
rect 5472 24068 5492 24132
rect 120 24052 5492 24068
rect 120 23988 5408 24052
rect 5472 23988 5492 24052
rect 120 23972 5492 23988
rect 120 23908 5408 23972
rect 5472 23908 5492 23972
rect 120 23892 5492 23908
rect 120 23828 5408 23892
rect 5472 23828 5492 23892
rect 120 23812 5492 23828
rect 120 23748 5408 23812
rect 5472 23748 5492 23812
rect 120 23732 5492 23748
rect 120 23668 5408 23732
rect 5472 23668 5492 23732
rect 120 23652 5492 23668
rect 120 23588 5408 23652
rect 5472 23588 5492 23652
rect 120 23572 5492 23588
rect 120 23508 5408 23572
rect 5472 23508 5492 23572
rect 120 23492 5492 23508
rect 120 23428 5408 23492
rect 5472 23428 5492 23492
rect 120 23412 5492 23428
rect 120 23348 5408 23412
rect 5472 23348 5492 23412
rect 120 23332 5492 23348
rect 120 23268 5408 23332
rect 5472 23268 5492 23332
rect 120 23252 5492 23268
rect 120 23188 5408 23252
rect 5472 23188 5492 23252
rect 120 23172 5492 23188
rect 120 23108 5408 23172
rect 5472 23108 5492 23172
rect 120 23092 5492 23108
rect 120 23028 5408 23092
rect 5472 23028 5492 23092
rect 120 23012 5492 23028
rect 120 22948 5408 23012
rect 5472 22948 5492 23012
rect 120 22932 5492 22948
rect 120 22868 5408 22932
rect 5472 22868 5492 22932
rect 120 22852 5492 22868
rect 120 22788 5408 22852
rect 5472 22788 5492 22852
rect 120 22772 5492 22788
rect 120 22708 5408 22772
rect 5472 22708 5492 22772
rect 120 22692 5492 22708
rect 120 22628 5408 22692
rect 5472 22628 5492 22692
rect 120 22612 5492 22628
rect 120 22548 5408 22612
rect 5472 22548 5492 22612
rect 120 22532 5492 22548
rect 120 22468 5408 22532
rect 5472 22468 5492 22532
rect 120 22452 5492 22468
rect 120 22388 5408 22452
rect 5472 22388 5492 22452
rect 120 22372 5492 22388
rect 120 22308 5408 22372
rect 5472 22308 5492 22372
rect 120 22292 5492 22308
rect 120 22228 5408 22292
rect 5472 22228 5492 22292
rect 120 22212 5492 22228
rect 120 22148 5408 22212
rect 5472 22148 5492 22212
rect 120 22132 5492 22148
rect 120 22068 5408 22132
rect 5472 22068 5492 22132
rect 120 22052 5492 22068
rect 120 21988 5408 22052
rect 5472 21988 5492 22052
rect 120 21972 5492 21988
rect 120 21908 5408 21972
rect 5472 21908 5492 21972
rect 120 21892 5492 21908
rect 120 21828 5408 21892
rect 5472 21828 5492 21892
rect 120 21812 5492 21828
rect 120 21748 5408 21812
rect 5472 21748 5492 21812
rect 120 21732 5492 21748
rect 120 21668 5408 21732
rect 5472 21668 5492 21732
rect 120 21652 5492 21668
rect 120 21588 5408 21652
rect 5472 21588 5492 21652
rect 120 21572 5492 21588
rect 120 21508 5408 21572
rect 5472 21508 5492 21572
rect 120 21492 5492 21508
rect 120 21428 5408 21492
rect 5472 21428 5492 21492
rect 120 21400 5492 21428
rect 5732 26452 11104 26480
rect 5732 26388 11020 26452
rect 11084 26388 11104 26452
rect 5732 26372 11104 26388
rect 5732 26308 11020 26372
rect 11084 26308 11104 26372
rect 5732 26292 11104 26308
rect 5732 26228 11020 26292
rect 11084 26228 11104 26292
rect 5732 26212 11104 26228
rect 5732 26148 11020 26212
rect 11084 26148 11104 26212
rect 5732 26132 11104 26148
rect 5732 26068 11020 26132
rect 11084 26068 11104 26132
rect 5732 26052 11104 26068
rect 5732 25988 11020 26052
rect 11084 25988 11104 26052
rect 5732 25972 11104 25988
rect 5732 25908 11020 25972
rect 11084 25908 11104 25972
rect 5732 25892 11104 25908
rect 5732 25828 11020 25892
rect 11084 25828 11104 25892
rect 5732 25812 11104 25828
rect 5732 25748 11020 25812
rect 11084 25748 11104 25812
rect 5732 25732 11104 25748
rect 5732 25668 11020 25732
rect 11084 25668 11104 25732
rect 5732 25652 11104 25668
rect 5732 25588 11020 25652
rect 11084 25588 11104 25652
rect 5732 25572 11104 25588
rect 5732 25508 11020 25572
rect 11084 25508 11104 25572
rect 5732 25492 11104 25508
rect 5732 25428 11020 25492
rect 11084 25428 11104 25492
rect 5732 25412 11104 25428
rect 5732 25348 11020 25412
rect 11084 25348 11104 25412
rect 5732 25332 11104 25348
rect 5732 25268 11020 25332
rect 11084 25268 11104 25332
rect 5732 25252 11104 25268
rect 5732 25188 11020 25252
rect 11084 25188 11104 25252
rect 5732 25172 11104 25188
rect 5732 25108 11020 25172
rect 11084 25108 11104 25172
rect 5732 25092 11104 25108
rect 5732 25028 11020 25092
rect 11084 25028 11104 25092
rect 5732 25012 11104 25028
rect 5732 24948 11020 25012
rect 11084 24948 11104 25012
rect 5732 24932 11104 24948
rect 5732 24868 11020 24932
rect 11084 24868 11104 24932
rect 5732 24852 11104 24868
rect 5732 24788 11020 24852
rect 11084 24788 11104 24852
rect 5732 24772 11104 24788
rect 5732 24708 11020 24772
rect 11084 24708 11104 24772
rect 5732 24692 11104 24708
rect 5732 24628 11020 24692
rect 11084 24628 11104 24692
rect 5732 24612 11104 24628
rect 5732 24548 11020 24612
rect 11084 24548 11104 24612
rect 5732 24532 11104 24548
rect 5732 24468 11020 24532
rect 11084 24468 11104 24532
rect 5732 24452 11104 24468
rect 5732 24388 11020 24452
rect 11084 24388 11104 24452
rect 5732 24372 11104 24388
rect 5732 24308 11020 24372
rect 11084 24308 11104 24372
rect 5732 24292 11104 24308
rect 5732 24228 11020 24292
rect 11084 24228 11104 24292
rect 5732 24212 11104 24228
rect 5732 24148 11020 24212
rect 11084 24148 11104 24212
rect 5732 24132 11104 24148
rect 5732 24068 11020 24132
rect 11084 24068 11104 24132
rect 5732 24052 11104 24068
rect 5732 23988 11020 24052
rect 11084 23988 11104 24052
rect 5732 23972 11104 23988
rect 5732 23908 11020 23972
rect 11084 23908 11104 23972
rect 5732 23892 11104 23908
rect 5732 23828 11020 23892
rect 11084 23828 11104 23892
rect 5732 23812 11104 23828
rect 5732 23748 11020 23812
rect 11084 23748 11104 23812
rect 5732 23732 11104 23748
rect 5732 23668 11020 23732
rect 11084 23668 11104 23732
rect 5732 23652 11104 23668
rect 5732 23588 11020 23652
rect 11084 23588 11104 23652
rect 5732 23572 11104 23588
rect 5732 23508 11020 23572
rect 11084 23508 11104 23572
rect 5732 23492 11104 23508
rect 5732 23428 11020 23492
rect 11084 23428 11104 23492
rect 5732 23412 11104 23428
rect 5732 23348 11020 23412
rect 11084 23348 11104 23412
rect 5732 23332 11104 23348
rect 5732 23268 11020 23332
rect 11084 23268 11104 23332
rect 5732 23252 11104 23268
rect 5732 23188 11020 23252
rect 11084 23188 11104 23252
rect 5732 23172 11104 23188
rect 5732 23108 11020 23172
rect 11084 23108 11104 23172
rect 5732 23092 11104 23108
rect 5732 23028 11020 23092
rect 11084 23028 11104 23092
rect 5732 23012 11104 23028
rect 5732 22948 11020 23012
rect 11084 22948 11104 23012
rect 5732 22932 11104 22948
rect 5732 22868 11020 22932
rect 11084 22868 11104 22932
rect 5732 22852 11104 22868
rect 5732 22788 11020 22852
rect 11084 22788 11104 22852
rect 5732 22772 11104 22788
rect 5732 22708 11020 22772
rect 11084 22708 11104 22772
rect 5732 22692 11104 22708
rect 5732 22628 11020 22692
rect 11084 22628 11104 22692
rect 5732 22612 11104 22628
rect 5732 22548 11020 22612
rect 11084 22548 11104 22612
rect 5732 22532 11104 22548
rect 5732 22468 11020 22532
rect 11084 22468 11104 22532
rect 5732 22452 11104 22468
rect 5732 22388 11020 22452
rect 11084 22388 11104 22452
rect 5732 22372 11104 22388
rect 5732 22308 11020 22372
rect 11084 22308 11104 22372
rect 5732 22292 11104 22308
rect 5732 22228 11020 22292
rect 11084 22228 11104 22292
rect 5732 22212 11104 22228
rect 5732 22148 11020 22212
rect 11084 22148 11104 22212
rect 5732 22132 11104 22148
rect 5732 22068 11020 22132
rect 11084 22068 11104 22132
rect 5732 22052 11104 22068
rect 5732 21988 11020 22052
rect 11084 21988 11104 22052
rect 5732 21972 11104 21988
rect 5732 21908 11020 21972
rect 11084 21908 11104 21972
rect 5732 21892 11104 21908
rect 5732 21828 11020 21892
rect 11084 21828 11104 21892
rect 5732 21812 11104 21828
rect 5732 21748 11020 21812
rect 11084 21748 11104 21812
rect 5732 21732 11104 21748
rect 5732 21668 11020 21732
rect 11084 21668 11104 21732
rect 5732 21652 11104 21668
rect 5732 21588 11020 21652
rect 11084 21588 11104 21652
rect 5732 21572 11104 21588
rect 5732 21508 11020 21572
rect 11084 21508 11104 21572
rect 5732 21492 11104 21508
rect 5732 21428 11020 21492
rect 11084 21428 11104 21492
rect 5732 21400 11104 21428
rect 11344 26452 16716 26480
rect 11344 26388 16632 26452
rect 16696 26388 16716 26452
rect 11344 26372 16716 26388
rect 11344 26308 16632 26372
rect 16696 26308 16716 26372
rect 11344 26292 16716 26308
rect 11344 26228 16632 26292
rect 16696 26228 16716 26292
rect 11344 26212 16716 26228
rect 11344 26148 16632 26212
rect 16696 26148 16716 26212
rect 11344 26132 16716 26148
rect 11344 26068 16632 26132
rect 16696 26068 16716 26132
rect 11344 26052 16716 26068
rect 11344 25988 16632 26052
rect 16696 25988 16716 26052
rect 11344 25972 16716 25988
rect 11344 25908 16632 25972
rect 16696 25908 16716 25972
rect 11344 25892 16716 25908
rect 11344 25828 16632 25892
rect 16696 25828 16716 25892
rect 11344 25812 16716 25828
rect 11344 25748 16632 25812
rect 16696 25748 16716 25812
rect 11344 25732 16716 25748
rect 11344 25668 16632 25732
rect 16696 25668 16716 25732
rect 11344 25652 16716 25668
rect 11344 25588 16632 25652
rect 16696 25588 16716 25652
rect 11344 25572 16716 25588
rect 11344 25508 16632 25572
rect 16696 25508 16716 25572
rect 11344 25492 16716 25508
rect 11344 25428 16632 25492
rect 16696 25428 16716 25492
rect 11344 25412 16716 25428
rect 11344 25348 16632 25412
rect 16696 25348 16716 25412
rect 11344 25332 16716 25348
rect 11344 25268 16632 25332
rect 16696 25268 16716 25332
rect 11344 25252 16716 25268
rect 11344 25188 16632 25252
rect 16696 25188 16716 25252
rect 11344 25172 16716 25188
rect 11344 25108 16632 25172
rect 16696 25108 16716 25172
rect 11344 25092 16716 25108
rect 11344 25028 16632 25092
rect 16696 25028 16716 25092
rect 11344 25012 16716 25028
rect 11344 24948 16632 25012
rect 16696 24948 16716 25012
rect 11344 24932 16716 24948
rect 11344 24868 16632 24932
rect 16696 24868 16716 24932
rect 11344 24852 16716 24868
rect 11344 24788 16632 24852
rect 16696 24788 16716 24852
rect 11344 24772 16716 24788
rect 11344 24708 16632 24772
rect 16696 24708 16716 24772
rect 11344 24692 16716 24708
rect 11344 24628 16632 24692
rect 16696 24628 16716 24692
rect 11344 24612 16716 24628
rect 11344 24548 16632 24612
rect 16696 24548 16716 24612
rect 11344 24532 16716 24548
rect 11344 24468 16632 24532
rect 16696 24468 16716 24532
rect 11344 24452 16716 24468
rect 11344 24388 16632 24452
rect 16696 24388 16716 24452
rect 11344 24372 16716 24388
rect 11344 24308 16632 24372
rect 16696 24308 16716 24372
rect 11344 24292 16716 24308
rect 11344 24228 16632 24292
rect 16696 24228 16716 24292
rect 11344 24212 16716 24228
rect 11344 24148 16632 24212
rect 16696 24148 16716 24212
rect 11344 24132 16716 24148
rect 11344 24068 16632 24132
rect 16696 24068 16716 24132
rect 11344 24052 16716 24068
rect 11344 23988 16632 24052
rect 16696 23988 16716 24052
rect 11344 23972 16716 23988
rect 11344 23908 16632 23972
rect 16696 23908 16716 23972
rect 11344 23892 16716 23908
rect 11344 23828 16632 23892
rect 16696 23828 16716 23892
rect 11344 23812 16716 23828
rect 11344 23748 16632 23812
rect 16696 23748 16716 23812
rect 11344 23732 16716 23748
rect 11344 23668 16632 23732
rect 16696 23668 16716 23732
rect 11344 23652 16716 23668
rect 11344 23588 16632 23652
rect 16696 23588 16716 23652
rect 11344 23572 16716 23588
rect 11344 23508 16632 23572
rect 16696 23508 16716 23572
rect 11344 23492 16716 23508
rect 11344 23428 16632 23492
rect 16696 23428 16716 23492
rect 11344 23412 16716 23428
rect 11344 23348 16632 23412
rect 16696 23348 16716 23412
rect 11344 23332 16716 23348
rect 11344 23268 16632 23332
rect 16696 23268 16716 23332
rect 11344 23252 16716 23268
rect 11344 23188 16632 23252
rect 16696 23188 16716 23252
rect 11344 23172 16716 23188
rect 11344 23108 16632 23172
rect 16696 23108 16716 23172
rect 11344 23092 16716 23108
rect 11344 23028 16632 23092
rect 16696 23028 16716 23092
rect 11344 23012 16716 23028
rect 11344 22948 16632 23012
rect 16696 22948 16716 23012
rect 11344 22932 16716 22948
rect 11344 22868 16632 22932
rect 16696 22868 16716 22932
rect 11344 22852 16716 22868
rect 11344 22788 16632 22852
rect 16696 22788 16716 22852
rect 11344 22772 16716 22788
rect 11344 22708 16632 22772
rect 16696 22708 16716 22772
rect 11344 22692 16716 22708
rect 11344 22628 16632 22692
rect 16696 22628 16716 22692
rect 11344 22612 16716 22628
rect 11344 22548 16632 22612
rect 16696 22548 16716 22612
rect 11344 22532 16716 22548
rect 11344 22468 16632 22532
rect 16696 22468 16716 22532
rect 11344 22452 16716 22468
rect 11344 22388 16632 22452
rect 16696 22388 16716 22452
rect 11344 22372 16716 22388
rect 11344 22308 16632 22372
rect 16696 22308 16716 22372
rect 11344 22292 16716 22308
rect 11344 22228 16632 22292
rect 16696 22228 16716 22292
rect 11344 22212 16716 22228
rect 11344 22148 16632 22212
rect 16696 22148 16716 22212
rect 11344 22132 16716 22148
rect 11344 22068 16632 22132
rect 16696 22068 16716 22132
rect 11344 22052 16716 22068
rect 11344 21988 16632 22052
rect 16696 21988 16716 22052
rect 11344 21972 16716 21988
rect 11344 21908 16632 21972
rect 16696 21908 16716 21972
rect 11344 21892 16716 21908
rect 11344 21828 16632 21892
rect 16696 21828 16716 21892
rect 11344 21812 16716 21828
rect 11344 21748 16632 21812
rect 16696 21748 16716 21812
rect 11344 21732 16716 21748
rect 11344 21668 16632 21732
rect 16696 21668 16716 21732
rect 11344 21652 16716 21668
rect 11344 21588 16632 21652
rect 16696 21588 16716 21652
rect 11344 21572 16716 21588
rect 11344 21508 16632 21572
rect 16696 21508 16716 21572
rect 11344 21492 16716 21508
rect 11344 21428 16632 21492
rect 16696 21428 16716 21492
rect 11344 21400 16716 21428
rect 16956 26452 22328 26480
rect 16956 26388 22244 26452
rect 22308 26388 22328 26452
rect 16956 26372 22328 26388
rect 16956 26308 22244 26372
rect 22308 26308 22328 26372
rect 16956 26292 22328 26308
rect 16956 26228 22244 26292
rect 22308 26228 22328 26292
rect 16956 26212 22328 26228
rect 16956 26148 22244 26212
rect 22308 26148 22328 26212
rect 16956 26132 22328 26148
rect 16956 26068 22244 26132
rect 22308 26068 22328 26132
rect 16956 26052 22328 26068
rect 16956 25988 22244 26052
rect 22308 25988 22328 26052
rect 16956 25972 22328 25988
rect 16956 25908 22244 25972
rect 22308 25908 22328 25972
rect 16956 25892 22328 25908
rect 16956 25828 22244 25892
rect 22308 25828 22328 25892
rect 16956 25812 22328 25828
rect 16956 25748 22244 25812
rect 22308 25748 22328 25812
rect 16956 25732 22328 25748
rect 16956 25668 22244 25732
rect 22308 25668 22328 25732
rect 16956 25652 22328 25668
rect 16956 25588 22244 25652
rect 22308 25588 22328 25652
rect 16956 25572 22328 25588
rect 16956 25508 22244 25572
rect 22308 25508 22328 25572
rect 16956 25492 22328 25508
rect 16956 25428 22244 25492
rect 22308 25428 22328 25492
rect 16956 25412 22328 25428
rect 16956 25348 22244 25412
rect 22308 25348 22328 25412
rect 16956 25332 22328 25348
rect 16956 25268 22244 25332
rect 22308 25268 22328 25332
rect 16956 25252 22328 25268
rect 16956 25188 22244 25252
rect 22308 25188 22328 25252
rect 16956 25172 22328 25188
rect 16956 25108 22244 25172
rect 22308 25108 22328 25172
rect 16956 25092 22328 25108
rect 16956 25028 22244 25092
rect 22308 25028 22328 25092
rect 16956 25012 22328 25028
rect 16956 24948 22244 25012
rect 22308 24948 22328 25012
rect 16956 24932 22328 24948
rect 16956 24868 22244 24932
rect 22308 24868 22328 24932
rect 16956 24852 22328 24868
rect 16956 24788 22244 24852
rect 22308 24788 22328 24852
rect 16956 24772 22328 24788
rect 16956 24708 22244 24772
rect 22308 24708 22328 24772
rect 16956 24692 22328 24708
rect 16956 24628 22244 24692
rect 22308 24628 22328 24692
rect 16956 24612 22328 24628
rect 16956 24548 22244 24612
rect 22308 24548 22328 24612
rect 16956 24532 22328 24548
rect 16956 24468 22244 24532
rect 22308 24468 22328 24532
rect 16956 24452 22328 24468
rect 16956 24388 22244 24452
rect 22308 24388 22328 24452
rect 16956 24372 22328 24388
rect 16956 24308 22244 24372
rect 22308 24308 22328 24372
rect 16956 24292 22328 24308
rect 16956 24228 22244 24292
rect 22308 24228 22328 24292
rect 16956 24212 22328 24228
rect 16956 24148 22244 24212
rect 22308 24148 22328 24212
rect 16956 24132 22328 24148
rect 16956 24068 22244 24132
rect 22308 24068 22328 24132
rect 16956 24052 22328 24068
rect 16956 23988 22244 24052
rect 22308 23988 22328 24052
rect 16956 23972 22328 23988
rect 16956 23908 22244 23972
rect 22308 23908 22328 23972
rect 16956 23892 22328 23908
rect 16956 23828 22244 23892
rect 22308 23828 22328 23892
rect 16956 23812 22328 23828
rect 16956 23748 22244 23812
rect 22308 23748 22328 23812
rect 16956 23732 22328 23748
rect 16956 23668 22244 23732
rect 22308 23668 22328 23732
rect 16956 23652 22328 23668
rect 16956 23588 22244 23652
rect 22308 23588 22328 23652
rect 16956 23572 22328 23588
rect 16956 23508 22244 23572
rect 22308 23508 22328 23572
rect 16956 23492 22328 23508
rect 16956 23428 22244 23492
rect 22308 23428 22328 23492
rect 16956 23412 22328 23428
rect 16956 23348 22244 23412
rect 22308 23348 22328 23412
rect 16956 23332 22328 23348
rect 16956 23268 22244 23332
rect 22308 23268 22328 23332
rect 16956 23252 22328 23268
rect 16956 23188 22244 23252
rect 22308 23188 22328 23252
rect 16956 23172 22328 23188
rect 16956 23108 22244 23172
rect 22308 23108 22328 23172
rect 16956 23092 22328 23108
rect 16956 23028 22244 23092
rect 22308 23028 22328 23092
rect 16956 23012 22328 23028
rect 16956 22948 22244 23012
rect 22308 22948 22328 23012
rect 16956 22932 22328 22948
rect 16956 22868 22244 22932
rect 22308 22868 22328 22932
rect 16956 22852 22328 22868
rect 16956 22788 22244 22852
rect 22308 22788 22328 22852
rect 16956 22772 22328 22788
rect 16956 22708 22244 22772
rect 22308 22708 22328 22772
rect 16956 22692 22328 22708
rect 16956 22628 22244 22692
rect 22308 22628 22328 22692
rect 16956 22612 22328 22628
rect 16956 22548 22244 22612
rect 22308 22548 22328 22612
rect 16956 22532 22328 22548
rect 16956 22468 22244 22532
rect 22308 22468 22328 22532
rect 16956 22452 22328 22468
rect 16956 22388 22244 22452
rect 22308 22388 22328 22452
rect 16956 22372 22328 22388
rect 16956 22308 22244 22372
rect 22308 22308 22328 22372
rect 16956 22292 22328 22308
rect 16956 22228 22244 22292
rect 22308 22228 22328 22292
rect 16956 22212 22328 22228
rect 16956 22148 22244 22212
rect 22308 22148 22328 22212
rect 16956 22132 22328 22148
rect 16956 22068 22244 22132
rect 22308 22068 22328 22132
rect 16956 22052 22328 22068
rect 16956 21988 22244 22052
rect 22308 21988 22328 22052
rect 16956 21972 22328 21988
rect 16956 21908 22244 21972
rect 22308 21908 22328 21972
rect 16956 21892 22328 21908
rect 16956 21828 22244 21892
rect 22308 21828 22328 21892
rect 16956 21812 22328 21828
rect 16956 21748 22244 21812
rect 22308 21748 22328 21812
rect 16956 21732 22328 21748
rect 16956 21668 22244 21732
rect 22308 21668 22328 21732
rect 16956 21652 22328 21668
rect 16956 21588 22244 21652
rect 22308 21588 22328 21652
rect 16956 21572 22328 21588
rect 16956 21508 22244 21572
rect 22308 21508 22328 21572
rect 16956 21492 22328 21508
rect 16956 21428 22244 21492
rect 22308 21428 22328 21492
rect 16956 21400 22328 21428
rect 22568 26452 27940 26480
rect 22568 26388 27856 26452
rect 27920 26388 27940 26452
rect 22568 26372 27940 26388
rect 22568 26308 27856 26372
rect 27920 26308 27940 26372
rect 22568 26292 27940 26308
rect 22568 26228 27856 26292
rect 27920 26228 27940 26292
rect 22568 26212 27940 26228
rect 22568 26148 27856 26212
rect 27920 26148 27940 26212
rect 22568 26132 27940 26148
rect 22568 26068 27856 26132
rect 27920 26068 27940 26132
rect 22568 26052 27940 26068
rect 22568 25988 27856 26052
rect 27920 25988 27940 26052
rect 22568 25972 27940 25988
rect 22568 25908 27856 25972
rect 27920 25908 27940 25972
rect 22568 25892 27940 25908
rect 22568 25828 27856 25892
rect 27920 25828 27940 25892
rect 22568 25812 27940 25828
rect 22568 25748 27856 25812
rect 27920 25748 27940 25812
rect 22568 25732 27940 25748
rect 22568 25668 27856 25732
rect 27920 25668 27940 25732
rect 22568 25652 27940 25668
rect 22568 25588 27856 25652
rect 27920 25588 27940 25652
rect 22568 25572 27940 25588
rect 22568 25508 27856 25572
rect 27920 25508 27940 25572
rect 22568 25492 27940 25508
rect 22568 25428 27856 25492
rect 27920 25428 27940 25492
rect 22568 25412 27940 25428
rect 22568 25348 27856 25412
rect 27920 25348 27940 25412
rect 22568 25332 27940 25348
rect 22568 25268 27856 25332
rect 27920 25268 27940 25332
rect 22568 25252 27940 25268
rect 22568 25188 27856 25252
rect 27920 25188 27940 25252
rect 22568 25172 27940 25188
rect 22568 25108 27856 25172
rect 27920 25108 27940 25172
rect 22568 25092 27940 25108
rect 22568 25028 27856 25092
rect 27920 25028 27940 25092
rect 22568 25012 27940 25028
rect 22568 24948 27856 25012
rect 27920 24948 27940 25012
rect 22568 24932 27940 24948
rect 22568 24868 27856 24932
rect 27920 24868 27940 24932
rect 22568 24852 27940 24868
rect 22568 24788 27856 24852
rect 27920 24788 27940 24852
rect 22568 24772 27940 24788
rect 22568 24708 27856 24772
rect 27920 24708 27940 24772
rect 22568 24692 27940 24708
rect 22568 24628 27856 24692
rect 27920 24628 27940 24692
rect 22568 24612 27940 24628
rect 22568 24548 27856 24612
rect 27920 24548 27940 24612
rect 22568 24532 27940 24548
rect 22568 24468 27856 24532
rect 27920 24468 27940 24532
rect 22568 24452 27940 24468
rect 22568 24388 27856 24452
rect 27920 24388 27940 24452
rect 22568 24372 27940 24388
rect 22568 24308 27856 24372
rect 27920 24308 27940 24372
rect 22568 24292 27940 24308
rect 22568 24228 27856 24292
rect 27920 24228 27940 24292
rect 22568 24212 27940 24228
rect 22568 24148 27856 24212
rect 27920 24148 27940 24212
rect 22568 24132 27940 24148
rect 22568 24068 27856 24132
rect 27920 24068 27940 24132
rect 22568 24052 27940 24068
rect 22568 23988 27856 24052
rect 27920 23988 27940 24052
rect 22568 23972 27940 23988
rect 22568 23908 27856 23972
rect 27920 23908 27940 23972
rect 22568 23892 27940 23908
rect 22568 23828 27856 23892
rect 27920 23828 27940 23892
rect 22568 23812 27940 23828
rect 22568 23748 27856 23812
rect 27920 23748 27940 23812
rect 22568 23732 27940 23748
rect 22568 23668 27856 23732
rect 27920 23668 27940 23732
rect 22568 23652 27940 23668
rect 22568 23588 27856 23652
rect 27920 23588 27940 23652
rect 22568 23572 27940 23588
rect 22568 23508 27856 23572
rect 27920 23508 27940 23572
rect 22568 23492 27940 23508
rect 22568 23428 27856 23492
rect 27920 23428 27940 23492
rect 22568 23412 27940 23428
rect 22568 23348 27856 23412
rect 27920 23348 27940 23412
rect 22568 23332 27940 23348
rect 22568 23268 27856 23332
rect 27920 23268 27940 23332
rect 22568 23252 27940 23268
rect 22568 23188 27856 23252
rect 27920 23188 27940 23252
rect 22568 23172 27940 23188
rect 22568 23108 27856 23172
rect 27920 23108 27940 23172
rect 22568 23092 27940 23108
rect 22568 23028 27856 23092
rect 27920 23028 27940 23092
rect 22568 23012 27940 23028
rect 22568 22948 27856 23012
rect 27920 22948 27940 23012
rect 22568 22932 27940 22948
rect 22568 22868 27856 22932
rect 27920 22868 27940 22932
rect 22568 22852 27940 22868
rect 22568 22788 27856 22852
rect 27920 22788 27940 22852
rect 22568 22772 27940 22788
rect 22568 22708 27856 22772
rect 27920 22708 27940 22772
rect 22568 22692 27940 22708
rect 22568 22628 27856 22692
rect 27920 22628 27940 22692
rect 22568 22612 27940 22628
rect 22568 22548 27856 22612
rect 27920 22548 27940 22612
rect 22568 22532 27940 22548
rect 22568 22468 27856 22532
rect 27920 22468 27940 22532
rect 22568 22452 27940 22468
rect 22568 22388 27856 22452
rect 27920 22388 27940 22452
rect 22568 22372 27940 22388
rect 22568 22308 27856 22372
rect 27920 22308 27940 22372
rect 22568 22292 27940 22308
rect 22568 22228 27856 22292
rect 27920 22228 27940 22292
rect 22568 22212 27940 22228
rect 22568 22148 27856 22212
rect 27920 22148 27940 22212
rect 22568 22132 27940 22148
rect 22568 22068 27856 22132
rect 27920 22068 27940 22132
rect 22568 22052 27940 22068
rect 22568 21988 27856 22052
rect 27920 21988 27940 22052
rect 22568 21972 27940 21988
rect 22568 21908 27856 21972
rect 27920 21908 27940 21972
rect 22568 21892 27940 21908
rect 22568 21828 27856 21892
rect 27920 21828 27940 21892
rect 22568 21812 27940 21828
rect 22568 21748 27856 21812
rect 27920 21748 27940 21812
rect 22568 21732 27940 21748
rect 22568 21668 27856 21732
rect 27920 21668 27940 21732
rect 22568 21652 27940 21668
rect 22568 21588 27856 21652
rect 27920 21588 27940 21652
rect 22568 21572 27940 21588
rect 22568 21508 27856 21572
rect 27920 21508 27940 21572
rect 22568 21492 27940 21508
rect 22568 21428 27856 21492
rect 27920 21428 27940 21492
rect 22568 21400 27940 21428
rect 28180 26452 33552 26480
rect 28180 26388 33468 26452
rect 33532 26388 33552 26452
rect 28180 26372 33552 26388
rect 28180 26308 33468 26372
rect 33532 26308 33552 26372
rect 28180 26292 33552 26308
rect 28180 26228 33468 26292
rect 33532 26228 33552 26292
rect 28180 26212 33552 26228
rect 28180 26148 33468 26212
rect 33532 26148 33552 26212
rect 28180 26132 33552 26148
rect 28180 26068 33468 26132
rect 33532 26068 33552 26132
rect 28180 26052 33552 26068
rect 28180 25988 33468 26052
rect 33532 25988 33552 26052
rect 28180 25972 33552 25988
rect 28180 25908 33468 25972
rect 33532 25908 33552 25972
rect 28180 25892 33552 25908
rect 28180 25828 33468 25892
rect 33532 25828 33552 25892
rect 28180 25812 33552 25828
rect 28180 25748 33468 25812
rect 33532 25748 33552 25812
rect 28180 25732 33552 25748
rect 28180 25668 33468 25732
rect 33532 25668 33552 25732
rect 28180 25652 33552 25668
rect 28180 25588 33468 25652
rect 33532 25588 33552 25652
rect 28180 25572 33552 25588
rect 28180 25508 33468 25572
rect 33532 25508 33552 25572
rect 28180 25492 33552 25508
rect 28180 25428 33468 25492
rect 33532 25428 33552 25492
rect 28180 25412 33552 25428
rect 28180 25348 33468 25412
rect 33532 25348 33552 25412
rect 28180 25332 33552 25348
rect 28180 25268 33468 25332
rect 33532 25268 33552 25332
rect 28180 25252 33552 25268
rect 28180 25188 33468 25252
rect 33532 25188 33552 25252
rect 28180 25172 33552 25188
rect 28180 25108 33468 25172
rect 33532 25108 33552 25172
rect 28180 25092 33552 25108
rect 28180 25028 33468 25092
rect 33532 25028 33552 25092
rect 28180 25012 33552 25028
rect 28180 24948 33468 25012
rect 33532 24948 33552 25012
rect 28180 24932 33552 24948
rect 28180 24868 33468 24932
rect 33532 24868 33552 24932
rect 28180 24852 33552 24868
rect 28180 24788 33468 24852
rect 33532 24788 33552 24852
rect 28180 24772 33552 24788
rect 28180 24708 33468 24772
rect 33532 24708 33552 24772
rect 28180 24692 33552 24708
rect 28180 24628 33468 24692
rect 33532 24628 33552 24692
rect 28180 24612 33552 24628
rect 28180 24548 33468 24612
rect 33532 24548 33552 24612
rect 28180 24532 33552 24548
rect 28180 24468 33468 24532
rect 33532 24468 33552 24532
rect 28180 24452 33552 24468
rect 28180 24388 33468 24452
rect 33532 24388 33552 24452
rect 28180 24372 33552 24388
rect 28180 24308 33468 24372
rect 33532 24308 33552 24372
rect 28180 24292 33552 24308
rect 28180 24228 33468 24292
rect 33532 24228 33552 24292
rect 28180 24212 33552 24228
rect 28180 24148 33468 24212
rect 33532 24148 33552 24212
rect 28180 24132 33552 24148
rect 28180 24068 33468 24132
rect 33532 24068 33552 24132
rect 28180 24052 33552 24068
rect 28180 23988 33468 24052
rect 33532 23988 33552 24052
rect 28180 23972 33552 23988
rect 28180 23908 33468 23972
rect 33532 23908 33552 23972
rect 28180 23892 33552 23908
rect 28180 23828 33468 23892
rect 33532 23828 33552 23892
rect 28180 23812 33552 23828
rect 28180 23748 33468 23812
rect 33532 23748 33552 23812
rect 28180 23732 33552 23748
rect 28180 23668 33468 23732
rect 33532 23668 33552 23732
rect 28180 23652 33552 23668
rect 28180 23588 33468 23652
rect 33532 23588 33552 23652
rect 28180 23572 33552 23588
rect 28180 23508 33468 23572
rect 33532 23508 33552 23572
rect 28180 23492 33552 23508
rect 28180 23428 33468 23492
rect 33532 23428 33552 23492
rect 28180 23412 33552 23428
rect 28180 23348 33468 23412
rect 33532 23348 33552 23412
rect 28180 23332 33552 23348
rect 28180 23268 33468 23332
rect 33532 23268 33552 23332
rect 28180 23252 33552 23268
rect 28180 23188 33468 23252
rect 33532 23188 33552 23252
rect 28180 23172 33552 23188
rect 28180 23108 33468 23172
rect 33532 23108 33552 23172
rect 28180 23092 33552 23108
rect 28180 23028 33468 23092
rect 33532 23028 33552 23092
rect 28180 23012 33552 23028
rect 28180 22948 33468 23012
rect 33532 22948 33552 23012
rect 28180 22932 33552 22948
rect 28180 22868 33468 22932
rect 33532 22868 33552 22932
rect 28180 22852 33552 22868
rect 28180 22788 33468 22852
rect 33532 22788 33552 22852
rect 28180 22772 33552 22788
rect 28180 22708 33468 22772
rect 33532 22708 33552 22772
rect 28180 22692 33552 22708
rect 28180 22628 33468 22692
rect 33532 22628 33552 22692
rect 28180 22612 33552 22628
rect 28180 22548 33468 22612
rect 33532 22548 33552 22612
rect 28180 22532 33552 22548
rect 28180 22468 33468 22532
rect 33532 22468 33552 22532
rect 28180 22452 33552 22468
rect 28180 22388 33468 22452
rect 33532 22388 33552 22452
rect 28180 22372 33552 22388
rect 28180 22308 33468 22372
rect 33532 22308 33552 22372
rect 28180 22292 33552 22308
rect 28180 22228 33468 22292
rect 33532 22228 33552 22292
rect 28180 22212 33552 22228
rect 28180 22148 33468 22212
rect 33532 22148 33552 22212
rect 28180 22132 33552 22148
rect 28180 22068 33468 22132
rect 33532 22068 33552 22132
rect 28180 22052 33552 22068
rect 28180 21988 33468 22052
rect 33532 21988 33552 22052
rect 28180 21972 33552 21988
rect 28180 21908 33468 21972
rect 33532 21908 33552 21972
rect 28180 21892 33552 21908
rect 28180 21828 33468 21892
rect 33532 21828 33552 21892
rect 28180 21812 33552 21828
rect 28180 21748 33468 21812
rect 33532 21748 33552 21812
rect 28180 21732 33552 21748
rect 28180 21668 33468 21732
rect 33532 21668 33552 21732
rect 28180 21652 33552 21668
rect 28180 21588 33468 21652
rect 33532 21588 33552 21652
rect 28180 21572 33552 21588
rect 28180 21508 33468 21572
rect 33532 21508 33552 21572
rect 28180 21492 33552 21508
rect 28180 21428 33468 21492
rect 33532 21428 33552 21492
rect 28180 21400 33552 21428
rect 33792 26452 39164 26480
rect 33792 26388 39080 26452
rect 39144 26388 39164 26452
rect 33792 26372 39164 26388
rect 33792 26308 39080 26372
rect 39144 26308 39164 26372
rect 33792 26292 39164 26308
rect 33792 26228 39080 26292
rect 39144 26228 39164 26292
rect 33792 26212 39164 26228
rect 33792 26148 39080 26212
rect 39144 26148 39164 26212
rect 33792 26132 39164 26148
rect 33792 26068 39080 26132
rect 39144 26068 39164 26132
rect 33792 26052 39164 26068
rect 33792 25988 39080 26052
rect 39144 25988 39164 26052
rect 33792 25972 39164 25988
rect 33792 25908 39080 25972
rect 39144 25908 39164 25972
rect 33792 25892 39164 25908
rect 33792 25828 39080 25892
rect 39144 25828 39164 25892
rect 33792 25812 39164 25828
rect 33792 25748 39080 25812
rect 39144 25748 39164 25812
rect 33792 25732 39164 25748
rect 33792 25668 39080 25732
rect 39144 25668 39164 25732
rect 33792 25652 39164 25668
rect 33792 25588 39080 25652
rect 39144 25588 39164 25652
rect 33792 25572 39164 25588
rect 33792 25508 39080 25572
rect 39144 25508 39164 25572
rect 33792 25492 39164 25508
rect 33792 25428 39080 25492
rect 39144 25428 39164 25492
rect 33792 25412 39164 25428
rect 33792 25348 39080 25412
rect 39144 25348 39164 25412
rect 33792 25332 39164 25348
rect 33792 25268 39080 25332
rect 39144 25268 39164 25332
rect 33792 25252 39164 25268
rect 33792 25188 39080 25252
rect 39144 25188 39164 25252
rect 33792 25172 39164 25188
rect 33792 25108 39080 25172
rect 39144 25108 39164 25172
rect 33792 25092 39164 25108
rect 33792 25028 39080 25092
rect 39144 25028 39164 25092
rect 33792 25012 39164 25028
rect 33792 24948 39080 25012
rect 39144 24948 39164 25012
rect 33792 24932 39164 24948
rect 33792 24868 39080 24932
rect 39144 24868 39164 24932
rect 33792 24852 39164 24868
rect 33792 24788 39080 24852
rect 39144 24788 39164 24852
rect 33792 24772 39164 24788
rect 33792 24708 39080 24772
rect 39144 24708 39164 24772
rect 33792 24692 39164 24708
rect 33792 24628 39080 24692
rect 39144 24628 39164 24692
rect 33792 24612 39164 24628
rect 33792 24548 39080 24612
rect 39144 24548 39164 24612
rect 33792 24532 39164 24548
rect 33792 24468 39080 24532
rect 39144 24468 39164 24532
rect 33792 24452 39164 24468
rect 33792 24388 39080 24452
rect 39144 24388 39164 24452
rect 33792 24372 39164 24388
rect 33792 24308 39080 24372
rect 39144 24308 39164 24372
rect 33792 24292 39164 24308
rect 33792 24228 39080 24292
rect 39144 24228 39164 24292
rect 33792 24212 39164 24228
rect 33792 24148 39080 24212
rect 39144 24148 39164 24212
rect 33792 24132 39164 24148
rect 33792 24068 39080 24132
rect 39144 24068 39164 24132
rect 33792 24052 39164 24068
rect 33792 23988 39080 24052
rect 39144 23988 39164 24052
rect 33792 23972 39164 23988
rect 33792 23908 39080 23972
rect 39144 23908 39164 23972
rect 33792 23892 39164 23908
rect 33792 23828 39080 23892
rect 39144 23828 39164 23892
rect 33792 23812 39164 23828
rect 33792 23748 39080 23812
rect 39144 23748 39164 23812
rect 33792 23732 39164 23748
rect 33792 23668 39080 23732
rect 39144 23668 39164 23732
rect 33792 23652 39164 23668
rect 33792 23588 39080 23652
rect 39144 23588 39164 23652
rect 33792 23572 39164 23588
rect 33792 23508 39080 23572
rect 39144 23508 39164 23572
rect 33792 23492 39164 23508
rect 33792 23428 39080 23492
rect 39144 23428 39164 23492
rect 33792 23412 39164 23428
rect 33792 23348 39080 23412
rect 39144 23348 39164 23412
rect 33792 23332 39164 23348
rect 33792 23268 39080 23332
rect 39144 23268 39164 23332
rect 33792 23252 39164 23268
rect 33792 23188 39080 23252
rect 39144 23188 39164 23252
rect 33792 23172 39164 23188
rect 33792 23108 39080 23172
rect 39144 23108 39164 23172
rect 33792 23092 39164 23108
rect 33792 23028 39080 23092
rect 39144 23028 39164 23092
rect 33792 23012 39164 23028
rect 33792 22948 39080 23012
rect 39144 22948 39164 23012
rect 33792 22932 39164 22948
rect 33792 22868 39080 22932
rect 39144 22868 39164 22932
rect 33792 22852 39164 22868
rect 33792 22788 39080 22852
rect 39144 22788 39164 22852
rect 33792 22772 39164 22788
rect 33792 22708 39080 22772
rect 39144 22708 39164 22772
rect 33792 22692 39164 22708
rect 33792 22628 39080 22692
rect 39144 22628 39164 22692
rect 33792 22612 39164 22628
rect 33792 22548 39080 22612
rect 39144 22548 39164 22612
rect 33792 22532 39164 22548
rect 33792 22468 39080 22532
rect 39144 22468 39164 22532
rect 33792 22452 39164 22468
rect 33792 22388 39080 22452
rect 39144 22388 39164 22452
rect 33792 22372 39164 22388
rect 33792 22308 39080 22372
rect 39144 22308 39164 22372
rect 33792 22292 39164 22308
rect 33792 22228 39080 22292
rect 39144 22228 39164 22292
rect 33792 22212 39164 22228
rect 33792 22148 39080 22212
rect 39144 22148 39164 22212
rect 33792 22132 39164 22148
rect 33792 22068 39080 22132
rect 39144 22068 39164 22132
rect 33792 22052 39164 22068
rect 33792 21988 39080 22052
rect 39144 21988 39164 22052
rect 33792 21972 39164 21988
rect 33792 21908 39080 21972
rect 39144 21908 39164 21972
rect 33792 21892 39164 21908
rect 33792 21828 39080 21892
rect 39144 21828 39164 21892
rect 33792 21812 39164 21828
rect 33792 21748 39080 21812
rect 39144 21748 39164 21812
rect 33792 21732 39164 21748
rect 33792 21668 39080 21732
rect 39144 21668 39164 21732
rect 33792 21652 39164 21668
rect 33792 21588 39080 21652
rect 39144 21588 39164 21652
rect 33792 21572 39164 21588
rect 33792 21508 39080 21572
rect 39144 21508 39164 21572
rect 33792 21492 39164 21508
rect 33792 21428 39080 21492
rect 39144 21428 39164 21492
rect 33792 21400 39164 21428
rect -39164 21132 -33792 21160
rect -39164 21068 -33876 21132
rect -33812 21068 -33792 21132
rect -39164 21052 -33792 21068
rect -39164 20988 -33876 21052
rect -33812 20988 -33792 21052
rect -39164 20972 -33792 20988
rect -39164 20908 -33876 20972
rect -33812 20908 -33792 20972
rect -39164 20892 -33792 20908
rect -39164 20828 -33876 20892
rect -33812 20828 -33792 20892
rect -39164 20812 -33792 20828
rect -39164 20748 -33876 20812
rect -33812 20748 -33792 20812
rect -39164 20732 -33792 20748
rect -39164 20668 -33876 20732
rect -33812 20668 -33792 20732
rect -39164 20652 -33792 20668
rect -39164 20588 -33876 20652
rect -33812 20588 -33792 20652
rect -39164 20572 -33792 20588
rect -39164 20508 -33876 20572
rect -33812 20508 -33792 20572
rect -39164 20492 -33792 20508
rect -39164 20428 -33876 20492
rect -33812 20428 -33792 20492
rect -39164 20412 -33792 20428
rect -39164 20348 -33876 20412
rect -33812 20348 -33792 20412
rect -39164 20332 -33792 20348
rect -39164 20268 -33876 20332
rect -33812 20268 -33792 20332
rect -39164 20252 -33792 20268
rect -39164 20188 -33876 20252
rect -33812 20188 -33792 20252
rect -39164 20172 -33792 20188
rect -39164 20108 -33876 20172
rect -33812 20108 -33792 20172
rect -39164 20092 -33792 20108
rect -39164 20028 -33876 20092
rect -33812 20028 -33792 20092
rect -39164 20012 -33792 20028
rect -39164 19948 -33876 20012
rect -33812 19948 -33792 20012
rect -39164 19932 -33792 19948
rect -39164 19868 -33876 19932
rect -33812 19868 -33792 19932
rect -39164 19852 -33792 19868
rect -39164 19788 -33876 19852
rect -33812 19788 -33792 19852
rect -39164 19772 -33792 19788
rect -39164 19708 -33876 19772
rect -33812 19708 -33792 19772
rect -39164 19692 -33792 19708
rect -39164 19628 -33876 19692
rect -33812 19628 -33792 19692
rect -39164 19612 -33792 19628
rect -39164 19548 -33876 19612
rect -33812 19548 -33792 19612
rect -39164 19532 -33792 19548
rect -39164 19468 -33876 19532
rect -33812 19468 -33792 19532
rect -39164 19452 -33792 19468
rect -39164 19388 -33876 19452
rect -33812 19388 -33792 19452
rect -39164 19372 -33792 19388
rect -39164 19308 -33876 19372
rect -33812 19308 -33792 19372
rect -39164 19292 -33792 19308
rect -39164 19228 -33876 19292
rect -33812 19228 -33792 19292
rect -39164 19212 -33792 19228
rect -39164 19148 -33876 19212
rect -33812 19148 -33792 19212
rect -39164 19132 -33792 19148
rect -39164 19068 -33876 19132
rect -33812 19068 -33792 19132
rect -39164 19052 -33792 19068
rect -39164 18988 -33876 19052
rect -33812 18988 -33792 19052
rect -39164 18972 -33792 18988
rect -39164 18908 -33876 18972
rect -33812 18908 -33792 18972
rect -39164 18892 -33792 18908
rect -39164 18828 -33876 18892
rect -33812 18828 -33792 18892
rect -39164 18812 -33792 18828
rect -39164 18748 -33876 18812
rect -33812 18748 -33792 18812
rect -39164 18732 -33792 18748
rect -39164 18668 -33876 18732
rect -33812 18668 -33792 18732
rect -39164 18652 -33792 18668
rect -39164 18588 -33876 18652
rect -33812 18588 -33792 18652
rect -39164 18572 -33792 18588
rect -39164 18508 -33876 18572
rect -33812 18508 -33792 18572
rect -39164 18492 -33792 18508
rect -39164 18428 -33876 18492
rect -33812 18428 -33792 18492
rect -39164 18412 -33792 18428
rect -39164 18348 -33876 18412
rect -33812 18348 -33792 18412
rect -39164 18332 -33792 18348
rect -39164 18268 -33876 18332
rect -33812 18268 -33792 18332
rect -39164 18252 -33792 18268
rect -39164 18188 -33876 18252
rect -33812 18188 -33792 18252
rect -39164 18172 -33792 18188
rect -39164 18108 -33876 18172
rect -33812 18108 -33792 18172
rect -39164 18092 -33792 18108
rect -39164 18028 -33876 18092
rect -33812 18028 -33792 18092
rect -39164 18012 -33792 18028
rect -39164 17948 -33876 18012
rect -33812 17948 -33792 18012
rect -39164 17932 -33792 17948
rect -39164 17868 -33876 17932
rect -33812 17868 -33792 17932
rect -39164 17852 -33792 17868
rect -39164 17788 -33876 17852
rect -33812 17788 -33792 17852
rect -39164 17772 -33792 17788
rect -39164 17708 -33876 17772
rect -33812 17708 -33792 17772
rect -39164 17692 -33792 17708
rect -39164 17628 -33876 17692
rect -33812 17628 -33792 17692
rect -39164 17612 -33792 17628
rect -39164 17548 -33876 17612
rect -33812 17548 -33792 17612
rect -39164 17532 -33792 17548
rect -39164 17468 -33876 17532
rect -33812 17468 -33792 17532
rect -39164 17452 -33792 17468
rect -39164 17388 -33876 17452
rect -33812 17388 -33792 17452
rect -39164 17372 -33792 17388
rect -39164 17308 -33876 17372
rect -33812 17308 -33792 17372
rect -39164 17292 -33792 17308
rect -39164 17228 -33876 17292
rect -33812 17228 -33792 17292
rect -39164 17212 -33792 17228
rect -39164 17148 -33876 17212
rect -33812 17148 -33792 17212
rect -39164 17132 -33792 17148
rect -39164 17068 -33876 17132
rect -33812 17068 -33792 17132
rect -39164 17052 -33792 17068
rect -39164 16988 -33876 17052
rect -33812 16988 -33792 17052
rect -39164 16972 -33792 16988
rect -39164 16908 -33876 16972
rect -33812 16908 -33792 16972
rect -39164 16892 -33792 16908
rect -39164 16828 -33876 16892
rect -33812 16828 -33792 16892
rect -39164 16812 -33792 16828
rect -39164 16748 -33876 16812
rect -33812 16748 -33792 16812
rect -39164 16732 -33792 16748
rect -39164 16668 -33876 16732
rect -33812 16668 -33792 16732
rect -39164 16652 -33792 16668
rect -39164 16588 -33876 16652
rect -33812 16588 -33792 16652
rect -39164 16572 -33792 16588
rect -39164 16508 -33876 16572
rect -33812 16508 -33792 16572
rect -39164 16492 -33792 16508
rect -39164 16428 -33876 16492
rect -33812 16428 -33792 16492
rect -39164 16412 -33792 16428
rect -39164 16348 -33876 16412
rect -33812 16348 -33792 16412
rect -39164 16332 -33792 16348
rect -39164 16268 -33876 16332
rect -33812 16268 -33792 16332
rect -39164 16252 -33792 16268
rect -39164 16188 -33876 16252
rect -33812 16188 -33792 16252
rect -39164 16172 -33792 16188
rect -39164 16108 -33876 16172
rect -33812 16108 -33792 16172
rect -39164 16080 -33792 16108
rect -33552 21132 -28180 21160
rect -33552 21068 -28264 21132
rect -28200 21068 -28180 21132
rect -33552 21052 -28180 21068
rect -33552 20988 -28264 21052
rect -28200 20988 -28180 21052
rect -33552 20972 -28180 20988
rect -33552 20908 -28264 20972
rect -28200 20908 -28180 20972
rect -33552 20892 -28180 20908
rect -33552 20828 -28264 20892
rect -28200 20828 -28180 20892
rect -33552 20812 -28180 20828
rect -33552 20748 -28264 20812
rect -28200 20748 -28180 20812
rect -33552 20732 -28180 20748
rect -33552 20668 -28264 20732
rect -28200 20668 -28180 20732
rect -33552 20652 -28180 20668
rect -33552 20588 -28264 20652
rect -28200 20588 -28180 20652
rect -33552 20572 -28180 20588
rect -33552 20508 -28264 20572
rect -28200 20508 -28180 20572
rect -33552 20492 -28180 20508
rect -33552 20428 -28264 20492
rect -28200 20428 -28180 20492
rect -33552 20412 -28180 20428
rect -33552 20348 -28264 20412
rect -28200 20348 -28180 20412
rect -33552 20332 -28180 20348
rect -33552 20268 -28264 20332
rect -28200 20268 -28180 20332
rect -33552 20252 -28180 20268
rect -33552 20188 -28264 20252
rect -28200 20188 -28180 20252
rect -33552 20172 -28180 20188
rect -33552 20108 -28264 20172
rect -28200 20108 -28180 20172
rect -33552 20092 -28180 20108
rect -33552 20028 -28264 20092
rect -28200 20028 -28180 20092
rect -33552 20012 -28180 20028
rect -33552 19948 -28264 20012
rect -28200 19948 -28180 20012
rect -33552 19932 -28180 19948
rect -33552 19868 -28264 19932
rect -28200 19868 -28180 19932
rect -33552 19852 -28180 19868
rect -33552 19788 -28264 19852
rect -28200 19788 -28180 19852
rect -33552 19772 -28180 19788
rect -33552 19708 -28264 19772
rect -28200 19708 -28180 19772
rect -33552 19692 -28180 19708
rect -33552 19628 -28264 19692
rect -28200 19628 -28180 19692
rect -33552 19612 -28180 19628
rect -33552 19548 -28264 19612
rect -28200 19548 -28180 19612
rect -33552 19532 -28180 19548
rect -33552 19468 -28264 19532
rect -28200 19468 -28180 19532
rect -33552 19452 -28180 19468
rect -33552 19388 -28264 19452
rect -28200 19388 -28180 19452
rect -33552 19372 -28180 19388
rect -33552 19308 -28264 19372
rect -28200 19308 -28180 19372
rect -33552 19292 -28180 19308
rect -33552 19228 -28264 19292
rect -28200 19228 -28180 19292
rect -33552 19212 -28180 19228
rect -33552 19148 -28264 19212
rect -28200 19148 -28180 19212
rect -33552 19132 -28180 19148
rect -33552 19068 -28264 19132
rect -28200 19068 -28180 19132
rect -33552 19052 -28180 19068
rect -33552 18988 -28264 19052
rect -28200 18988 -28180 19052
rect -33552 18972 -28180 18988
rect -33552 18908 -28264 18972
rect -28200 18908 -28180 18972
rect -33552 18892 -28180 18908
rect -33552 18828 -28264 18892
rect -28200 18828 -28180 18892
rect -33552 18812 -28180 18828
rect -33552 18748 -28264 18812
rect -28200 18748 -28180 18812
rect -33552 18732 -28180 18748
rect -33552 18668 -28264 18732
rect -28200 18668 -28180 18732
rect -33552 18652 -28180 18668
rect -33552 18588 -28264 18652
rect -28200 18588 -28180 18652
rect -33552 18572 -28180 18588
rect -33552 18508 -28264 18572
rect -28200 18508 -28180 18572
rect -33552 18492 -28180 18508
rect -33552 18428 -28264 18492
rect -28200 18428 -28180 18492
rect -33552 18412 -28180 18428
rect -33552 18348 -28264 18412
rect -28200 18348 -28180 18412
rect -33552 18332 -28180 18348
rect -33552 18268 -28264 18332
rect -28200 18268 -28180 18332
rect -33552 18252 -28180 18268
rect -33552 18188 -28264 18252
rect -28200 18188 -28180 18252
rect -33552 18172 -28180 18188
rect -33552 18108 -28264 18172
rect -28200 18108 -28180 18172
rect -33552 18092 -28180 18108
rect -33552 18028 -28264 18092
rect -28200 18028 -28180 18092
rect -33552 18012 -28180 18028
rect -33552 17948 -28264 18012
rect -28200 17948 -28180 18012
rect -33552 17932 -28180 17948
rect -33552 17868 -28264 17932
rect -28200 17868 -28180 17932
rect -33552 17852 -28180 17868
rect -33552 17788 -28264 17852
rect -28200 17788 -28180 17852
rect -33552 17772 -28180 17788
rect -33552 17708 -28264 17772
rect -28200 17708 -28180 17772
rect -33552 17692 -28180 17708
rect -33552 17628 -28264 17692
rect -28200 17628 -28180 17692
rect -33552 17612 -28180 17628
rect -33552 17548 -28264 17612
rect -28200 17548 -28180 17612
rect -33552 17532 -28180 17548
rect -33552 17468 -28264 17532
rect -28200 17468 -28180 17532
rect -33552 17452 -28180 17468
rect -33552 17388 -28264 17452
rect -28200 17388 -28180 17452
rect -33552 17372 -28180 17388
rect -33552 17308 -28264 17372
rect -28200 17308 -28180 17372
rect -33552 17292 -28180 17308
rect -33552 17228 -28264 17292
rect -28200 17228 -28180 17292
rect -33552 17212 -28180 17228
rect -33552 17148 -28264 17212
rect -28200 17148 -28180 17212
rect -33552 17132 -28180 17148
rect -33552 17068 -28264 17132
rect -28200 17068 -28180 17132
rect -33552 17052 -28180 17068
rect -33552 16988 -28264 17052
rect -28200 16988 -28180 17052
rect -33552 16972 -28180 16988
rect -33552 16908 -28264 16972
rect -28200 16908 -28180 16972
rect -33552 16892 -28180 16908
rect -33552 16828 -28264 16892
rect -28200 16828 -28180 16892
rect -33552 16812 -28180 16828
rect -33552 16748 -28264 16812
rect -28200 16748 -28180 16812
rect -33552 16732 -28180 16748
rect -33552 16668 -28264 16732
rect -28200 16668 -28180 16732
rect -33552 16652 -28180 16668
rect -33552 16588 -28264 16652
rect -28200 16588 -28180 16652
rect -33552 16572 -28180 16588
rect -33552 16508 -28264 16572
rect -28200 16508 -28180 16572
rect -33552 16492 -28180 16508
rect -33552 16428 -28264 16492
rect -28200 16428 -28180 16492
rect -33552 16412 -28180 16428
rect -33552 16348 -28264 16412
rect -28200 16348 -28180 16412
rect -33552 16332 -28180 16348
rect -33552 16268 -28264 16332
rect -28200 16268 -28180 16332
rect -33552 16252 -28180 16268
rect -33552 16188 -28264 16252
rect -28200 16188 -28180 16252
rect -33552 16172 -28180 16188
rect -33552 16108 -28264 16172
rect -28200 16108 -28180 16172
rect -33552 16080 -28180 16108
rect -27940 21132 -22568 21160
rect -27940 21068 -22652 21132
rect -22588 21068 -22568 21132
rect -27940 21052 -22568 21068
rect -27940 20988 -22652 21052
rect -22588 20988 -22568 21052
rect -27940 20972 -22568 20988
rect -27940 20908 -22652 20972
rect -22588 20908 -22568 20972
rect -27940 20892 -22568 20908
rect -27940 20828 -22652 20892
rect -22588 20828 -22568 20892
rect -27940 20812 -22568 20828
rect -27940 20748 -22652 20812
rect -22588 20748 -22568 20812
rect -27940 20732 -22568 20748
rect -27940 20668 -22652 20732
rect -22588 20668 -22568 20732
rect -27940 20652 -22568 20668
rect -27940 20588 -22652 20652
rect -22588 20588 -22568 20652
rect -27940 20572 -22568 20588
rect -27940 20508 -22652 20572
rect -22588 20508 -22568 20572
rect -27940 20492 -22568 20508
rect -27940 20428 -22652 20492
rect -22588 20428 -22568 20492
rect -27940 20412 -22568 20428
rect -27940 20348 -22652 20412
rect -22588 20348 -22568 20412
rect -27940 20332 -22568 20348
rect -27940 20268 -22652 20332
rect -22588 20268 -22568 20332
rect -27940 20252 -22568 20268
rect -27940 20188 -22652 20252
rect -22588 20188 -22568 20252
rect -27940 20172 -22568 20188
rect -27940 20108 -22652 20172
rect -22588 20108 -22568 20172
rect -27940 20092 -22568 20108
rect -27940 20028 -22652 20092
rect -22588 20028 -22568 20092
rect -27940 20012 -22568 20028
rect -27940 19948 -22652 20012
rect -22588 19948 -22568 20012
rect -27940 19932 -22568 19948
rect -27940 19868 -22652 19932
rect -22588 19868 -22568 19932
rect -27940 19852 -22568 19868
rect -27940 19788 -22652 19852
rect -22588 19788 -22568 19852
rect -27940 19772 -22568 19788
rect -27940 19708 -22652 19772
rect -22588 19708 -22568 19772
rect -27940 19692 -22568 19708
rect -27940 19628 -22652 19692
rect -22588 19628 -22568 19692
rect -27940 19612 -22568 19628
rect -27940 19548 -22652 19612
rect -22588 19548 -22568 19612
rect -27940 19532 -22568 19548
rect -27940 19468 -22652 19532
rect -22588 19468 -22568 19532
rect -27940 19452 -22568 19468
rect -27940 19388 -22652 19452
rect -22588 19388 -22568 19452
rect -27940 19372 -22568 19388
rect -27940 19308 -22652 19372
rect -22588 19308 -22568 19372
rect -27940 19292 -22568 19308
rect -27940 19228 -22652 19292
rect -22588 19228 -22568 19292
rect -27940 19212 -22568 19228
rect -27940 19148 -22652 19212
rect -22588 19148 -22568 19212
rect -27940 19132 -22568 19148
rect -27940 19068 -22652 19132
rect -22588 19068 -22568 19132
rect -27940 19052 -22568 19068
rect -27940 18988 -22652 19052
rect -22588 18988 -22568 19052
rect -27940 18972 -22568 18988
rect -27940 18908 -22652 18972
rect -22588 18908 -22568 18972
rect -27940 18892 -22568 18908
rect -27940 18828 -22652 18892
rect -22588 18828 -22568 18892
rect -27940 18812 -22568 18828
rect -27940 18748 -22652 18812
rect -22588 18748 -22568 18812
rect -27940 18732 -22568 18748
rect -27940 18668 -22652 18732
rect -22588 18668 -22568 18732
rect -27940 18652 -22568 18668
rect -27940 18588 -22652 18652
rect -22588 18588 -22568 18652
rect -27940 18572 -22568 18588
rect -27940 18508 -22652 18572
rect -22588 18508 -22568 18572
rect -27940 18492 -22568 18508
rect -27940 18428 -22652 18492
rect -22588 18428 -22568 18492
rect -27940 18412 -22568 18428
rect -27940 18348 -22652 18412
rect -22588 18348 -22568 18412
rect -27940 18332 -22568 18348
rect -27940 18268 -22652 18332
rect -22588 18268 -22568 18332
rect -27940 18252 -22568 18268
rect -27940 18188 -22652 18252
rect -22588 18188 -22568 18252
rect -27940 18172 -22568 18188
rect -27940 18108 -22652 18172
rect -22588 18108 -22568 18172
rect -27940 18092 -22568 18108
rect -27940 18028 -22652 18092
rect -22588 18028 -22568 18092
rect -27940 18012 -22568 18028
rect -27940 17948 -22652 18012
rect -22588 17948 -22568 18012
rect -27940 17932 -22568 17948
rect -27940 17868 -22652 17932
rect -22588 17868 -22568 17932
rect -27940 17852 -22568 17868
rect -27940 17788 -22652 17852
rect -22588 17788 -22568 17852
rect -27940 17772 -22568 17788
rect -27940 17708 -22652 17772
rect -22588 17708 -22568 17772
rect -27940 17692 -22568 17708
rect -27940 17628 -22652 17692
rect -22588 17628 -22568 17692
rect -27940 17612 -22568 17628
rect -27940 17548 -22652 17612
rect -22588 17548 -22568 17612
rect -27940 17532 -22568 17548
rect -27940 17468 -22652 17532
rect -22588 17468 -22568 17532
rect -27940 17452 -22568 17468
rect -27940 17388 -22652 17452
rect -22588 17388 -22568 17452
rect -27940 17372 -22568 17388
rect -27940 17308 -22652 17372
rect -22588 17308 -22568 17372
rect -27940 17292 -22568 17308
rect -27940 17228 -22652 17292
rect -22588 17228 -22568 17292
rect -27940 17212 -22568 17228
rect -27940 17148 -22652 17212
rect -22588 17148 -22568 17212
rect -27940 17132 -22568 17148
rect -27940 17068 -22652 17132
rect -22588 17068 -22568 17132
rect -27940 17052 -22568 17068
rect -27940 16988 -22652 17052
rect -22588 16988 -22568 17052
rect -27940 16972 -22568 16988
rect -27940 16908 -22652 16972
rect -22588 16908 -22568 16972
rect -27940 16892 -22568 16908
rect -27940 16828 -22652 16892
rect -22588 16828 -22568 16892
rect -27940 16812 -22568 16828
rect -27940 16748 -22652 16812
rect -22588 16748 -22568 16812
rect -27940 16732 -22568 16748
rect -27940 16668 -22652 16732
rect -22588 16668 -22568 16732
rect -27940 16652 -22568 16668
rect -27940 16588 -22652 16652
rect -22588 16588 -22568 16652
rect -27940 16572 -22568 16588
rect -27940 16508 -22652 16572
rect -22588 16508 -22568 16572
rect -27940 16492 -22568 16508
rect -27940 16428 -22652 16492
rect -22588 16428 -22568 16492
rect -27940 16412 -22568 16428
rect -27940 16348 -22652 16412
rect -22588 16348 -22568 16412
rect -27940 16332 -22568 16348
rect -27940 16268 -22652 16332
rect -22588 16268 -22568 16332
rect -27940 16252 -22568 16268
rect -27940 16188 -22652 16252
rect -22588 16188 -22568 16252
rect -27940 16172 -22568 16188
rect -27940 16108 -22652 16172
rect -22588 16108 -22568 16172
rect -27940 16080 -22568 16108
rect -22328 21132 -16956 21160
rect -22328 21068 -17040 21132
rect -16976 21068 -16956 21132
rect -22328 21052 -16956 21068
rect -22328 20988 -17040 21052
rect -16976 20988 -16956 21052
rect -22328 20972 -16956 20988
rect -22328 20908 -17040 20972
rect -16976 20908 -16956 20972
rect -22328 20892 -16956 20908
rect -22328 20828 -17040 20892
rect -16976 20828 -16956 20892
rect -22328 20812 -16956 20828
rect -22328 20748 -17040 20812
rect -16976 20748 -16956 20812
rect -22328 20732 -16956 20748
rect -22328 20668 -17040 20732
rect -16976 20668 -16956 20732
rect -22328 20652 -16956 20668
rect -22328 20588 -17040 20652
rect -16976 20588 -16956 20652
rect -22328 20572 -16956 20588
rect -22328 20508 -17040 20572
rect -16976 20508 -16956 20572
rect -22328 20492 -16956 20508
rect -22328 20428 -17040 20492
rect -16976 20428 -16956 20492
rect -22328 20412 -16956 20428
rect -22328 20348 -17040 20412
rect -16976 20348 -16956 20412
rect -22328 20332 -16956 20348
rect -22328 20268 -17040 20332
rect -16976 20268 -16956 20332
rect -22328 20252 -16956 20268
rect -22328 20188 -17040 20252
rect -16976 20188 -16956 20252
rect -22328 20172 -16956 20188
rect -22328 20108 -17040 20172
rect -16976 20108 -16956 20172
rect -22328 20092 -16956 20108
rect -22328 20028 -17040 20092
rect -16976 20028 -16956 20092
rect -22328 20012 -16956 20028
rect -22328 19948 -17040 20012
rect -16976 19948 -16956 20012
rect -22328 19932 -16956 19948
rect -22328 19868 -17040 19932
rect -16976 19868 -16956 19932
rect -22328 19852 -16956 19868
rect -22328 19788 -17040 19852
rect -16976 19788 -16956 19852
rect -22328 19772 -16956 19788
rect -22328 19708 -17040 19772
rect -16976 19708 -16956 19772
rect -22328 19692 -16956 19708
rect -22328 19628 -17040 19692
rect -16976 19628 -16956 19692
rect -22328 19612 -16956 19628
rect -22328 19548 -17040 19612
rect -16976 19548 -16956 19612
rect -22328 19532 -16956 19548
rect -22328 19468 -17040 19532
rect -16976 19468 -16956 19532
rect -22328 19452 -16956 19468
rect -22328 19388 -17040 19452
rect -16976 19388 -16956 19452
rect -22328 19372 -16956 19388
rect -22328 19308 -17040 19372
rect -16976 19308 -16956 19372
rect -22328 19292 -16956 19308
rect -22328 19228 -17040 19292
rect -16976 19228 -16956 19292
rect -22328 19212 -16956 19228
rect -22328 19148 -17040 19212
rect -16976 19148 -16956 19212
rect -22328 19132 -16956 19148
rect -22328 19068 -17040 19132
rect -16976 19068 -16956 19132
rect -22328 19052 -16956 19068
rect -22328 18988 -17040 19052
rect -16976 18988 -16956 19052
rect -22328 18972 -16956 18988
rect -22328 18908 -17040 18972
rect -16976 18908 -16956 18972
rect -22328 18892 -16956 18908
rect -22328 18828 -17040 18892
rect -16976 18828 -16956 18892
rect -22328 18812 -16956 18828
rect -22328 18748 -17040 18812
rect -16976 18748 -16956 18812
rect -22328 18732 -16956 18748
rect -22328 18668 -17040 18732
rect -16976 18668 -16956 18732
rect -22328 18652 -16956 18668
rect -22328 18588 -17040 18652
rect -16976 18588 -16956 18652
rect -22328 18572 -16956 18588
rect -22328 18508 -17040 18572
rect -16976 18508 -16956 18572
rect -22328 18492 -16956 18508
rect -22328 18428 -17040 18492
rect -16976 18428 -16956 18492
rect -22328 18412 -16956 18428
rect -22328 18348 -17040 18412
rect -16976 18348 -16956 18412
rect -22328 18332 -16956 18348
rect -22328 18268 -17040 18332
rect -16976 18268 -16956 18332
rect -22328 18252 -16956 18268
rect -22328 18188 -17040 18252
rect -16976 18188 -16956 18252
rect -22328 18172 -16956 18188
rect -22328 18108 -17040 18172
rect -16976 18108 -16956 18172
rect -22328 18092 -16956 18108
rect -22328 18028 -17040 18092
rect -16976 18028 -16956 18092
rect -22328 18012 -16956 18028
rect -22328 17948 -17040 18012
rect -16976 17948 -16956 18012
rect -22328 17932 -16956 17948
rect -22328 17868 -17040 17932
rect -16976 17868 -16956 17932
rect -22328 17852 -16956 17868
rect -22328 17788 -17040 17852
rect -16976 17788 -16956 17852
rect -22328 17772 -16956 17788
rect -22328 17708 -17040 17772
rect -16976 17708 -16956 17772
rect -22328 17692 -16956 17708
rect -22328 17628 -17040 17692
rect -16976 17628 -16956 17692
rect -22328 17612 -16956 17628
rect -22328 17548 -17040 17612
rect -16976 17548 -16956 17612
rect -22328 17532 -16956 17548
rect -22328 17468 -17040 17532
rect -16976 17468 -16956 17532
rect -22328 17452 -16956 17468
rect -22328 17388 -17040 17452
rect -16976 17388 -16956 17452
rect -22328 17372 -16956 17388
rect -22328 17308 -17040 17372
rect -16976 17308 -16956 17372
rect -22328 17292 -16956 17308
rect -22328 17228 -17040 17292
rect -16976 17228 -16956 17292
rect -22328 17212 -16956 17228
rect -22328 17148 -17040 17212
rect -16976 17148 -16956 17212
rect -22328 17132 -16956 17148
rect -22328 17068 -17040 17132
rect -16976 17068 -16956 17132
rect -22328 17052 -16956 17068
rect -22328 16988 -17040 17052
rect -16976 16988 -16956 17052
rect -22328 16972 -16956 16988
rect -22328 16908 -17040 16972
rect -16976 16908 -16956 16972
rect -22328 16892 -16956 16908
rect -22328 16828 -17040 16892
rect -16976 16828 -16956 16892
rect -22328 16812 -16956 16828
rect -22328 16748 -17040 16812
rect -16976 16748 -16956 16812
rect -22328 16732 -16956 16748
rect -22328 16668 -17040 16732
rect -16976 16668 -16956 16732
rect -22328 16652 -16956 16668
rect -22328 16588 -17040 16652
rect -16976 16588 -16956 16652
rect -22328 16572 -16956 16588
rect -22328 16508 -17040 16572
rect -16976 16508 -16956 16572
rect -22328 16492 -16956 16508
rect -22328 16428 -17040 16492
rect -16976 16428 -16956 16492
rect -22328 16412 -16956 16428
rect -22328 16348 -17040 16412
rect -16976 16348 -16956 16412
rect -22328 16332 -16956 16348
rect -22328 16268 -17040 16332
rect -16976 16268 -16956 16332
rect -22328 16252 -16956 16268
rect -22328 16188 -17040 16252
rect -16976 16188 -16956 16252
rect -22328 16172 -16956 16188
rect -22328 16108 -17040 16172
rect -16976 16108 -16956 16172
rect -22328 16080 -16956 16108
rect -16716 21132 -11344 21160
rect -16716 21068 -11428 21132
rect -11364 21068 -11344 21132
rect -16716 21052 -11344 21068
rect -16716 20988 -11428 21052
rect -11364 20988 -11344 21052
rect -16716 20972 -11344 20988
rect -16716 20908 -11428 20972
rect -11364 20908 -11344 20972
rect -16716 20892 -11344 20908
rect -16716 20828 -11428 20892
rect -11364 20828 -11344 20892
rect -16716 20812 -11344 20828
rect -16716 20748 -11428 20812
rect -11364 20748 -11344 20812
rect -16716 20732 -11344 20748
rect -16716 20668 -11428 20732
rect -11364 20668 -11344 20732
rect -16716 20652 -11344 20668
rect -16716 20588 -11428 20652
rect -11364 20588 -11344 20652
rect -16716 20572 -11344 20588
rect -16716 20508 -11428 20572
rect -11364 20508 -11344 20572
rect -16716 20492 -11344 20508
rect -16716 20428 -11428 20492
rect -11364 20428 -11344 20492
rect -16716 20412 -11344 20428
rect -16716 20348 -11428 20412
rect -11364 20348 -11344 20412
rect -16716 20332 -11344 20348
rect -16716 20268 -11428 20332
rect -11364 20268 -11344 20332
rect -16716 20252 -11344 20268
rect -16716 20188 -11428 20252
rect -11364 20188 -11344 20252
rect -16716 20172 -11344 20188
rect -16716 20108 -11428 20172
rect -11364 20108 -11344 20172
rect -16716 20092 -11344 20108
rect -16716 20028 -11428 20092
rect -11364 20028 -11344 20092
rect -16716 20012 -11344 20028
rect -16716 19948 -11428 20012
rect -11364 19948 -11344 20012
rect -16716 19932 -11344 19948
rect -16716 19868 -11428 19932
rect -11364 19868 -11344 19932
rect -16716 19852 -11344 19868
rect -16716 19788 -11428 19852
rect -11364 19788 -11344 19852
rect -16716 19772 -11344 19788
rect -16716 19708 -11428 19772
rect -11364 19708 -11344 19772
rect -16716 19692 -11344 19708
rect -16716 19628 -11428 19692
rect -11364 19628 -11344 19692
rect -16716 19612 -11344 19628
rect -16716 19548 -11428 19612
rect -11364 19548 -11344 19612
rect -16716 19532 -11344 19548
rect -16716 19468 -11428 19532
rect -11364 19468 -11344 19532
rect -16716 19452 -11344 19468
rect -16716 19388 -11428 19452
rect -11364 19388 -11344 19452
rect -16716 19372 -11344 19388
rect -16716 19308 -11428 19372
rect -11364 19308 -11344 19372
rect -16716 19292 -11344 19308
rect -16716 19228 -11428 19292
rect -11364 19228 -11344 19292
rect -16716 19212 -11344 19228
rect -16716 19148 -11428 19212
rect -11364 19148 -11344 19212
rect -16716 19132 -11344 19148
rect -16716 19068 -11428 19132
rect -11364 19068 -11344 19132
rect -16716 19052 -11344 19068
rect -16716 18988 -11428 19052
rect -11364 18988 -11344 19052
rect -16716 18972 -11344 18988
rect -16716 18908 -11428 18972
rect -11364 18908 -11344 18972
rect -16716 18892 -11344 18908
rect -16716 18828 -11428 18892
rect -11364 18828 -11344 18892
rect -16716 18812 -11344 18828
rect -16716 18748 -11428 18812
rect -11364 18748 -11344 18812
rect -16716 18732 -11344 18748
rect -16716 18668 -11428 18732
rect -11364 18668 -11344 18732
rect -16716 18652 -11344 18668
rect -16716 18588 -11428 18652
rect -11364 18588 -11344 18652
rect -16716 18572 -11344 18588
rect -16716 18508 -11428 18572
rect -11364 18508 -11344 18572
rect -16716 18492 -11344 18508
rect -16716 18428 -11428 18492
rect -11364 18428 -11344 18492
rect -16716 18412 -11344 18428
rect -16716 18348 -11428 18412
rect -11364 18348 -11344 18412
rect -16716 18332 -11344 18348
rect -16716 18268 -11428 18332
rect -11364 18268 -11344 18332
rect -16716 18252 -11344 18268
rect -16716 18188 -11428 18252
rect -11364 18188 -11344 18252
rect -16716 18172 -11344 18188
rect -16716 18108 -11428 18172
rect -11364 18108 -11344 18172
rect -16716 18092 -11344 18108
rect -16716 18028 -11428 18092
rect -11364 18028 -11344 18092
rect -16716 18012 -11344 18028
rect -16716 17948 -11428 18012
rect -11364 17948 -11344 18012
rect -16716 17932 -11344 17948
rect -16716 17868 -11428 17932
rect -11364 17868 -11344 17932
rect -16716 17852 -11344 17868
rect -16716 17788 -11428 17852
rect -11364 17788 -11344 17852
rect -16716 17772 -11344 17788
rect -16716 17708 -11428 17772
rect -11364 17708 -11344 17772
rect -16716 17692 -11344 17708
rect -16716 17628 -11428 17692
rect -11364 17628 -11344 17692
rect -16716 17612 -11344 17628
rect -16716 17548 -11428 17612
rect -11364 17548 -11344 17612
rect -16716 17532 -11344 17548
rect -16716 17468 -11428 17532
rect -11364 17468 -11344 17532
rect -16716 17452 -11344 17468
rect -16716 17388 -11428 17452
rect -11364 17388 -11344 17452
rect -16716 17372 -11344 17388
rect -16716 17308 -11428 17372
rect -11364 17308 -11344 17372
rect -16716 17292 -11344 17308
rect -16716 17228 -11428 17292
rect -11364 17228 -11344 17292
rect -16716 17212 -11344 17228
rect -16716 17148 -11428 17212
rect -11364 17148 -11344 17212
rect -16716 17132 -11344 17148
rect -16716 17068 -11428 17132
rect -11364 17068 -11344 17132
rect -16716 17052 -11344 17068
rect -16716 16988 -11428 17052
rect -11364 16988 -11344 17052
rect -16716 16972 -11344 16988
rect -16716 16908 -11428 16972
rect -11364 16908 -11344 16972
rect -16716 16892 -11344 16908
rect -16716 16828 -11428 16892
rect -11364 16828 -11344 16892
rect -16716 16812 -11344 16828
rect -16716 16748 -11428 16812
rect -11364 16748 -11344 16812
rect -16716 16732 -11344 16748
rect -16716 16668 -11428 16732
rect -11364 16668 -11344 16732
rect -16716 16652 -11344 16668
rect -16716 16588 -11428 16652
rect -11364 16588 -11344 16652
rect -16716 16572 -11344 16588
rect -16716 16508 -11428 16572
rect -11364 16508 -11344 16572
rect -16716 16492 -11344 16508
rect -16716 16428 -11428 16492
rect -11364 16428 -11344 16492
rect -16716 16412 -11344 16428
rect -16716 16348 -11428 16412
rect -11364 16348 -11344 16412
rect -16716 16332 -11344 16348
rect -16716 16268 -11428 16332
rect -11364 16268 -11344 16332
rect -16716 16252 -11344 16268
rect -16716 16188 -11428 16252
rect -11364 16188 -11344 16252
rect -16716 16172 -11344 16188
rect -16716 16108 -11428 16172
rect -11364 16108 -11344 16172
rect -16716 16080 -11344 16108
rect -11104 21132 -5732 21160
rect -11104 21068 -5816 21132
rect -5752 21068 -5732 21132
rect -11104 21052 -5732 21068
rect -11104 20988 -5816 21052
rect -5752 20988 -5732 21052
rect -11104 20972 -5732 20988
rect -11104 20908 -5816 20972
rect -5752 20908 -5732 20972
rect -11104 20892 -5732 20908
rect -11104 20828 -5816 20892
rect -5752 20828 -5732 20892
rect -11104 20812 -5732 20828
rect -11104 20748 -5816 20812
rect -5752 20748 -5732 20812
rect -11104 20732 -5732 20748
rect -11104 20668 -5816 20732
rect -5752 20668 -5732 20732
rect -11104 20652 -5732 20668
rect -11104 20588 -5816 20652
rect -5752 20588 -5732 20652
rect -11104 20572 -5732 20588
rect -11104 20508 -5816 20572
rect -5752 20508 -5732 20572
rect -11104 20492 -5732 20508
rect -11104 20428 -5816 20492
rect -5752 20428 -5732 20492
rect -11104 20412 -5732 20428
rect -11104 20348 -5816 20412
rect -5752 20348 -5732 20412
rect -11104 20332 -5732 20348
rect -11104 20268 -5816 20332
rect -5752 20268 -5732 20332
rect -11104 20252 -5732 20268
rect -11104 20188 -5816 20252
rect -5752 20188 -5732 20252
rect -11104 20172 -5732 20188
rect -11104 20108 -5816 20172
rect -5752 20108 -5732 20172
rect -11104 20092 -5732 20108
rect -11104 20028 -5816 20092
rect -5752 20028 -5732 20092
rect -11104 20012 -5732 20028
rect -11104 19948 -5816 20012
rect -5752 19948 -5732 20012
rect -11104 19932 -5732 19948
rect -11104 19868 -5816 19932
rect -5752 19868 -5732 19932
rect -11104 19852 -5732 19868
rect -11104 19788 -5816 19852
rect -5752 19788 -5732 19852
rect -11104 19772 -5732 19788
rect -11104 19708 -5816 19772
rect -5752 19708 -5732 19772
rect -11104 19692 -5732 19708
rect -11104 19628 -5816 19692
rect -5752 19628 -5732 19692
rect -11104 19612 -5732 19628
rect -11104 19548 -5816 19612
rect -5752 19548 -5732 19612
rect -11104 19532 -5732 19548
rect -11104 19468 -5816 19532
rect -5752 19468 -5732 19532
rect -11104 19452 -5732 19468
rect -11104 19388 -5816 19452
rect -5752 19388 -5732 19452
rect -11104 19372 -5732 19388
rect -11104 19308 -5816 19372
rect -5752 19308 -5732 19372
rect -11104 19292 -5732 19308
rect -11104 19228 -5816 19292
rect -5752 19228 -5732 19292
rect -11104 19212 -5732 19228
rect -11104 19148 -5816 19212
rect -5752 19148 -5732 19212
rect -11104 19132 -5732 19148
rect -11104 19068 -5816 19132
rect -5752 19068 -5732 19132
rect -11104 19052 -5732 19068
rect -11104 18988 -5816 19052
rect -5752 18988 -5732 19052
rect -11104 18972 -5732 18988
rect -11104 18908 -5816 18972
rect -5752 18908 -5732 18972
rect -11104 18892 -5732 18908
rect -11104 18828 -5816 18892
rect -5752 18828 -5732 18892
rect -11104 18812 -5732 18828
rect -11104 18748 -5816 18812
rect -5752 18748 -5732 18812
rect -11104 18732 -5732 18748
rect -11104 18668 -5816 18732
rect -5752 18668 -5732 18732
rect -11104 18652 -5732 18668
rect -11104 18588 -5816 18652
rect -5752 18588 -5732 18652
rect -11104 18572 -5732 18588
rect -11104 18508 -5816 18572
rect -5752 18508 -5732 18572
rect -11104 18492 -5732 18508
rect -11104 18428 -5816 18492
rect -5752 18428 -5732 18492
rect -11104 18412 -5732 18428
rect -11104 18348 -5816 18412
rect -5752 18348 -5732 18412
rect -11104 18332 -5732 18348
rect -11104 18268 -5816 18332
rect -5752 18268 -5732 18332
rect -11104 18252 -5732 18268
rect -11104 18188 -5816 18252
rect -5752 18188 -5732 18252
rect -11104 18172 -5732 18188
rect -11104 18108 -5816 18172
rect -5752 18108 -5732 18172
rect -11104 18092 -5732 18108
rect -11104 18028 -5816 18092
rect -5752 18028 -5732 18092
rect -11104 18012 -5732 18028
rect -11104 17948 -5816 18012
rect -5752 17948 -5732 18012
rect -11104 17932 -5732 17948
rect -11104 17868 -5816 17932
rect -5752 17868 -5732 17932
rect -11104 17852 -5732 17868
rect -11104 17788 -5816 17852
rect -5752 17788 -5732 17852
rect -11104 17772 -5732 17788
rect -11104 17708 -5816 17772
rect -5752 17708 -5732 17772
rect -11104 17692 -5732 17708
rect -11104 17628 -5816 17692
rect -5752 17628 -5732 17692
rect -11104 17612 -5732 17628
rect -11104 17548 -5816 17612
rect -5752 17548 -5732 17612
rect -11104 17532 -5732 17548
rect -11104 17468 -5816 17532
rect -5752 17468 -5732 17532
rect -11104 17452 -5732 17468
rect -11104 17388 -5816 17452
rect -5752 17388 -5732 17452
rect -11104 17372 -5732 17388
rect -11104 17308 -5816 17372
rect -5752 17308 -5732 17372
rect -11104 17292 -5732 17308
rect -11104 17228 -5816 17292
rect -5752 17228 -5732 17292
rect -11104 17212 -5732 17228
rect -11104 17148 -5816 17212
rect -5752 17148 -5732 17212
rect -11104 17132 -5732 17148
rect -11104 17068 -5816 17132
rect -5752 17068 -5732 17132
rect -11104 17052 -5732 17068
rect -11104 16988 -5816 17052
rect -5752 16988 -5732 17052
rect -11104 16972 -5732 16988
rect -11104 16908 -5816 16972
rect -5752 16908 -5732 16972
rect -11104 16892 -5732 16908
rect -11104 16828 -5816 16892
rect -5752 16828 -5732 16892
rect -11104 16812 -5732 16828
rect -11104 16748 -5816 16812
rect -5752 16748 -5732 16812
rect -11104 16732 -5732 16748
rect -11104 16668 -5816 16732
rect -5752 16668 -5732 16732
rect -11104 16652 -5732 16668
rect -11104 16588 -5816 16652
rect -5752 16588 -5732 16652
rect -11104 16572 -5732 16588
rect -11104 16508 -5816 16572
rect -5752 16508 -5732 16572
rect -11104 16492 -5732 16508
rect -11104 16428 -5816 16492
rect -5752 16428 -5732 16492
rect -11104 16412 -5732 16428
rect -11104 16348 -5816 16412
rect -5752 16348 -5732 16412
rect -11104 16332 -5732 16348
rect -11104 16268 -5816 16332
rect -5752 16268 -5732 16332
rect -11104 16252 -5732 16268
rect -11104 16188 -5816 16252
rect -5752 16188 -5732 16252
rect -11104 16172 -5732 16188
rect -11104 16108 -5816 16172
rect -5752 16108 -5732 16172
rect -11104 16080 -5732 16108
rect -5492 21132 -120 21160
rect -5492 21068 -204 21132
rect -140 21068 -120 21132
rect -5492 21052 -120 21068
rect -5492 20988 -204 21052
rect -140 20988 -120 21052
rect -5492 20972 -120 20988
rect -5492 20908 -204 20972
rect -140 20908 -120 20972
rect -5492 20892 -120 20908
rect -5492 20828 -204 20892
rect -140 20828 -120 20892
rect -5492 20812 -120 20828
rect -5492 20748 -204 20812
rect -140 20748 -120 20812
rect -5492 20732 -120 20748
rect -5492 20668 -204 20732
rect -140 20668 -120 20732
rect -5492 20652 -120 20668
rect -5492 20588 -204 20652
rect -140 20588 -120 20652
rect -5492 20572 -120 20588
rect -5492 20508 -204 20572
rect -140 20508 -120 20572
rect -5492 20492 -120 20508
rect -5492 20428 -204 20492
rect -140 20428 -120 20492
rect -5492 20412 -120 20428
rect -5492 20348 -204 20412
rect -140 20348 -120 20412
rect -5492 20332 -120 20348
rect -5492 20268 -204 20332
rect -140 20268 -120 20332
rect -5492 20252 -120 20268
rect -5492 20188 -204 20252
rect -140 20188 -120 20252
rect -5492 20172 -120 20188
rect -5492 20108 -204 20172
rect -140 20108 -120 20172
rect -5492 20092 -120 20108
rect -5492 20028 -204 20092
rect -140 20028 -120 20092
rect -5492 20012 -120 20028
rect -5492 19948 -204 20012
rect -140 19948 -120 20012
rect -5492 19932 -120 19948
rect -5492 19868 -204 19932
rect -140 19868 -120 19932
rect -5492 19852 -120 19868
rect -5492 19788 -204 19852
rect -140 19788 -120 19852
rect -5492 19772 -120 19788
rect -5492 19708 -204 19772
rect -140 19708 -120 19772
rect -5492 19692 -120 19708
rect -5492 19628 -204 19692
rect -140 19628 -120 19692
rect -5492 19612 -120 19628
rect -5492 19548 -204 19612
rect -140 19548 -120 19612
rect -5492 19532 -120 19548
rect -5492 19468 -204 19532
rect -140 19468 -120 19532
rect -5492 19452 -120 19468
rect -5492 19388 -204 19452
rect -140 19388 -120 19452
rect -5492 19372 -120 19388
rect -5492 19308 -204 19372
rect -140 19308 -120 19372
rect -5492 19292 -120 19308
rect -5492 19228 -204 19292
rect -140 19228 -120 19292
rect -5492 19212 -120 19228
rect -5492 19148 -204 19212
rect -140 19148 -120 19212
rect -5492 19132 -120 19148
rect -5492 19068 -204 19132
rect -140 19068 -120 19132
rect -5492 19052 -120 19068
rect -5492 18988 -204 19052
rect -140 18988 -120 19052
rect -5492 18972 -120 18988
rect -5492 18908 -204 18972
rect -140 18908 -120 18972
rect -5492 18892 -120 18908
rect -5492 18828 -204 18892
rect -140 18828 -120 18892
rect -5492 18812 -120 18828
rect -5492 18748 -204 18812
rect -140 18748 -120 18812
rect -5492 18732 -120 18748
rect -5492 18668 -204 18732
rect -140 18668 -120 18732
rect -5492 18652 -120 18668
rect -5492 18588 -204 18652
rect -140 18588 -120 18652
rect -5492 18572 -120 18588
rect -5492 18508 -204 18572
rect -140 18508 -120 18572
rect -5492 18492 -120 18508
rect -5492 18428 -204 18492
rect -140 18428 -120 18492
rect -5492 18412 -120 18428
rect -5492 18348 -204 18412
rect -140 18348 -120 18412
rect -5492 18332 -120 18348
rect -5492 18268 -204 18332
rect -140 18268 -120 18332
rect -5492 18252 -120 18268
rect -5492 18188 -204 18252
rect -140 18188 -120 18252
rect -5492 18172 -120 18188
rect -5492 18108 -204 18172
rect -140 18108 -120 18172
rect -5492 18092 -120 18108
rect -5492 18028 -204 18092
rect -140 18028 -120 18092
rect -5492 18012 -120 18028
rect -5492 17948 -204 18012
rect -140 17948 -120 18012
rect -5492 17932 -120 17948
rect -5492 17868 -204 17932
rect -140 17868 -120 17932
rect -5492 17852 -120 17868
rect -5492 17788 -204 17852
rect -140 17788 -120 17852
rect -5492 17772 -120 17788
rect -5492 17708 -204 17772
rect -140 17708 -120 17772
rect -5492 17692 -120 17708
rect -5492 17628 -204 17692
rect -140 17628 -120 17692
rect -5492 17612 -120 17628
rect -5492 17548 -204 17612
rect -140 17548 -120 17612
rect -5492 17532 -120 17548
rect -5492 17468 -204 17532
rect -140 17468 -120 17532
rect -5492 17452 -120 17468
rect -5492 17388 -204 17452
rect -140 17388 -120 17452
rect -5492 17372 -120 17388
rect -5492 17308 -204 17372
rect -140 17308 -120 17372
rect -5492 17292 -120 17308
rect -5492 17228 -204 17292
rect -140 17228 -120 17292
rect -5492 17212 -120 17228
rect -5492 17148 -204 17212
rect -140 17148 -120 17212
rect -5492 17132 -120 17148
rect -5492 17068 -204 17132
rect -140 17068 -120 17132
rect -5492 17052 -120 17068
rect -5492 16988 -204 17052
rect -140 16988 -120 17052
rect -5492 16972 -120 16988
rect -5492 16908 -204 16972
rect -140 16908 -120 16972
rect -5492 16892 -120 16908
rect -5492 16828 -204 16892
rect -140 16828 -120 16892
rect -5492 16812 -120 16828
rect -5492 16748 -204 16812
rect -140 16748 -120 16812
rect -5492 16732 -120 16748
rect -5492 16668 -204 16732
rect -140 16668 -120 16732
rect -5492 16652 -120 16668
rect -5492 16588 -204 16652
rect -140 16588 -120 16652
rect -5492 16572 -120 16588
rect -5492 16508 -204 16572
rect -140 16508 -120 16572
rect -5492 16492 -120 16508
rect -5492 16428 -204 16492
rect -140 16428 -120 16492
rect -5492 16412 -120 16428
rect -5492 16348 -204 16412
rect -140 16348 -120 16412
rect -5492 16332 -120 16348
rect -5492 16268 -204 16332
rect -140 16268 -120 16332
rect -5492 16252 -120 16268
rect -5492 16188 -204 16252
rect -140 16188 -120 16252
rect -5492 16172 -120 16188
rect -5492 16108 -204 16172
rect -140 16108 -120 16172
rect -5492 16080 -120 16108
rect 120 21132 5492 21160
rect 120 21068 5408 21132
rect 5472 21068 5492 21132
rect 120 21052 5492 21068
rect 120 20988 5408 21052
rect 5472 20988 5492 21052
rect 120 20972 5492 20988
rect 120 20908 5408 20972
rect 5472 20908 5492 20972
rect 120 20892 5492 20908
rect 120 20828 5408 20892
rect 5472 20828 5492 20892
rect 120 20812 5492 20828
rect 120 20748 5408 20812
rect 5472 20748 5492 20812
rect 120 20732 5492 20748
rect 120 20668 5408 20732
rect 5472 20668 5492 20732
rect 120 20652 5492 20668
rect 120 20588 5408 20652
rect 5472 20588 5492 20652
rect 120 20572 5492 20588
rect 120 20508 5408 20572
rect 5472 20508 5492 20572
rect 120 20492 5492 20508
rect 120 20428 5408 20492
rect 5472 20428 5492 20492
rect 120 20412 5492 20428
rect 120 20348 5408 20412
rect 5472 20348 5492 20412
rect 120 20332 5492 20348
rect 120 20268 5408 20332
rect 5472 20268 5492 20332
rect 120 20252 5492 20268
rect 120 20188 5408 20252
rect 5472 20188 5492 20252
rect 120 20172 5492 20188
rect 120 20108 5408 20172
rect 5472 20108 5492 20172
rect 120 20092 5492 20108
rect 120 20028 5408 20092
rect 5472 20028 5492 20092
rect 120 20012 5492 20028
rect 120 19948 5408 20012
rect 5472 19948 5492 20012
rect 120 19932 5492 19948
rect 120 19868 5408 19932
rect 5472 19868 5492 19932
rect 120 19852 5492 19868
rect 120 19788 5408 19852
rect 5472 19788 5492 19852
rect 120 19772 5492 19788
rect 120 19708 5408 19772
rect 5472 19708 5492 19772
rect 120 19692 5492 19708
rect 120 19628 5408 19692
rect 5472 19628 5492 19692
rect 120 19612 5492 19628
rect 120 19548 5408 19612
rect 5472 19548 5492 19612
rect 120 19532 5492 19548
rect 120 19468 5408 19532
rect 5472 19468 5492 19532
rect 120 19452 5492 19468
rect 120 19388 5408 19452
rect 5472 19388 5492 19452
rect 120 19372 5492 19388
rect 120 19308 5408 19372
rect 5472 19308 5492 19372
rect 120 19292 5492 19308
rect 120 19228 5408 19292
rect 5472 19228 5492 19292
rect 120 19212 5492 19228
rect 120 19148 5408 19212
rect 5472 19148 5492 19212
rect 120 19132 5492 19148
rect 120 19068 5408 19132
rect 5472 19068 5492 19132
rect 120 19052 5492 19068
rect 120 18988 5408 19052
rect 5472 18988 5492 19052
rect 120 18972 5492 18988
rect 120 18908 5408 18972
rect 5472 18908 5492 18972
rect 120 18892 5492 18908
rect 120 18828 5408 18892
rect 5472 18828 5492 18892
rect 120 18812 5492 18828
rect 120 18748 5408 18812
rect 5472 18748 5492 18812
rect 120 18732 5492 18748
rect 120 18668 5408 18732
rect 5472 18668 5492 18732
rect 120 18652 5492 18668
rect 120 18588 5408 18652
rect 5472 18588 5492 18652
rect 120 18572 5492 18588
rect 120 18508 5408 18572
rect 5472 18508 5492 18572
rect 120 18492 5492 18508
rect 120 18428 5408 18492
rect 5472 18428 5492 18492
rect 120 18412 5492 18428
rect 120 18348 5408 18412
rect 5472 18348 5492 18412
rect 120 18332 5492 18348
rect 120 18268 5408 18332
rect 5472 18268 5492 18332
rect 120 18252 5492 18268
rect 120 18188 5408 18252
rect 5472 18188 5492 18252
rect 120 18172 5492 18188
rect 120 18108 5408 18172
rect 5472 18108 5492 18172
rect 120 18092 5492 18108
rect 120 18028 5408 18092
rect 5472 18028 5492 18092
rect 120 18012 5492 18028
rect 120 17948 5408 18012
rect 5472 17948 5492 18012
rect 120 17932 5492 17948
rect 120 17868 5408 17932
rect 5472 17868 5492 17932
rect 120 17852 5492 17868
rect 120 17788 5408 17852
rect 5472 17788 5492 17852
rect 120 17772 5492 17788
rect 120 17708 5408 17772
rect 5472 17708 5492 17772
rect 120 17692 5492 17708
rect 120 17628 5408 17692
rect 5472 17628 5492 17692
rect 120 17612 5492 17628
rect 120 17548 5408 17612
rect 5472 17548 5492 17612
rect 120 17532 5492 17548
rect 120 17468 5408 17532
rect 5472 17468 5492 17532
rect 120 17452 5492 17468
rect 120 17388 5408 17452
rect 5472 17388 5492 17452
rect 120 17372 5492 17388
rect 120 17308 5408 17372
rect 5472 17308 5492 17372
rect 120 17292 5492 17308
rect 120 17228 5408 17292
rect 5472 17228 5492 17292
rect 120 17212 5492 17228
rect 120 17148 5408 17212
rect 5472 17148 5492 17212
rect 120 17132 5492 17148
rect 120 17068 5408 17132
rect 5472 17068 5492 17132
rect 120 17052 5492 17068
rect 120 16988 5408 17052
rect 5472 16988 5492 17052
rect 120 16972 5492 16988
rect 120 16908 5408 16972
rect 5472 16908 5492 16972
rect 120 16892 5492 16908
rect 120 16828 5408 16892
rect 5472 16828 5492 16892
rect 120 16812 5492 16828
rect 120 16748 5408 16812
rect 5472 16748 5492 16812
rect 120 16732 5492 16748
rect 120 16668 5408 16732
rect 5472 16668 5492 16732
rect 120 16652 5492 16668
rect 120 16588 5408 16652
rect 5472 16588 5492 16652
rect 120 16572 5492 16588
rect 120 16508 5408 16572
rect 5472 16508 5492 16572
rect 120 16492 5492 16508
rect 120 16428 5408 16492
rect 5472 16428 5492 16492
rect 120 16412 5492 16428
rect 120 16348 5408 16412
rect 5472 16348 5492 16412
rect 120 16332 5492 16348
rect 120 16268 5408 16332
rect 5472 16268 5492 16332
rect 120 16252 5492 16268
rect 120 16188 5408 16252
rect 5472 16188 5492 16252
rect 120 16172 5492 16188
rect 120 16108 5408 16172
rect 5472 16108 5492 16172
rect 120 16080 5492 16108
rect 5732 21132 11104 21160
rect 5732 21068 11020 21132
rect 11084 21068 11104 21132
rect 5732 21052 11104 21068
rect 5732 20988 11020 21052
rect 11084 20988 11104 21052
rect 5732 20972 11104 20988
rect 5732 20908 11020 20972
rect 11084 20908 11104 20972
rect 5732 20892 11104 20908
rect 5732 20828 11020 20892
rect 11084 20828 11104 20892
rect 5732 20812 11104 20828
rect 5732 20748 11020 20812
rect 11084 20748 11104 20812
rect 5732 20732 11104 20748
rect 5732 20668 11020 20732
rect 11084 20668 11104 20732
rect 5732 20652 11104 20668
rect 5732 20588 11020 20652
rect 11084 20588 11104 20652
rect 5732 20572 11104 20588
rect 5732 20508 11020 20572
rect 11084 20508 11104 20572
rect 5732 20492 11104 20508
rect 5732 20428 11020 20492
rect 11084 20428 11104 20492
rect 5732 20412 11104 20428
rect 5732 20348 11020 20412
rect 11084 20348 11104 20412
rect 5732 20332 11104 20348
rect 5732 20268 11020 20332
rect 11084 20268 11104 20332
rect 5732 20252 11104 20268
rect 5732 20188 11020 20252
rect 11084 20188 11104 20252
rect 5732 20172 11104 20188
rect 5732 20108 11020 20172
rect 11084 20108 11104 20172
rect 5732 20092 11104 20108
rect 5732 20028 11020 20092
rect 11084 20028 11104 20092
rect 5732 20012 11104 20028
rect 5732 19948 11020 20012
rect 11084 19948 11104 20012
rect 5732 19932 11104 19948
rect 5732 19868 11020 19932
rect 11084 19868 11104 19932
rect 5732 19852 11104 19868
rect 5732 19788 11020 19852
rect 11084 19788 11104 19852
rect 5732 19772 11104 19788
rect 5732 19708 11020 19772
rect 11084 19708 11104 19772
rect 5732 19692 11104 19708
rect 5732 19628 11020 19692
rect 11084 19628 11104 19692
rect 5732 19612 11104 19628
rect 5732 19548 11020 19612
rect 11084 19548 11104 19612
rect 5732 19532 11104 19548
rect 5732 19468 11020 19532
rect 11084 19468 11104 19532
rect 5732 19452 11104 19468
rect 5732 19388 11020 19452
rect 11084 19388 11104 19452
rect 5732 19372 11104 19388
rect 5732 19308 11020 19372
rect 11084 19308 11104 19372
rect 5732 19292 11104 19308
rect 5732 19228 11020 19292
rect 11084 19228 11104 19292
rect 5732 19212 11104 19228
rect 5732 19148 11020 19212
rect 11084 19148 11104 19212
rect 5732 19132 11104 19148
rect 5732 19068 11020 19132
rect 11084 19068 11104 19132
rect 5732 19052 11104 19068
rect 5732 18988 11020 19052
rect 11084 18988 11104 19052
rect 5732 18972 11104 18988
rect 5732 18908 11020 18972
rect 11084 18908 11104 18972
rect 5732 18892 11104 18908
rect 5732 18828 11020 18892
rect 11084 18828 11104 18892
rect 5732 18812 11104 18828
rect 5732 18748 11020 18812
rect 11084 18748 11104 18812
rect 5732 18732 11104 18748
rect 5732 18668 11020 18732
rect 11084 18668 11104 18732
rect 5732 18652 11104 18668
rect 5732 18588 11020 18652
rect 11084 18588 11104 18652
rect 5732 18572 11104 18588
rect 5732 18508 11020 18572
rect 11084 18508 11104 18572
rect 5732 18492 11104 18508
rect 5732 18428 11020 18492
rect 11084 18428 11104 18492
rect 5732 18412 11104 18428
rect 5732 18348 11020 18412
rect 11084 18348 11104 18412
rect 5732 18332 11104 18348
rect 5732 18268 11020 18332
rect 11084 18268 11104 18332
rect 5732 18252 11104 18268
rect 5732 18188 11020 18252
rect 11084 18188 11104 18252
rect 5732 18172 11104 18188
rect 5732 18108 11020 18172
rect 11084 18108 11104 18172
rect 5732 18092 11104 18108
rect 5732 18028 11020 18092
rect 11084 18028 11104 18092
rect 5732 18012 11104 18028
rect 5732 17948 11020 18012
rect 11084 17948 11104 18012
rect 5732 17932 11104 17948
rect 5732 17868 11020 17932
rect 11084 17868 11104 17932
rect 5732 17852 11104 17868
rect 5732 17788 11020 17852
rect 11084 17788 11104 17852
rect 5732 17772 11104 17788
rect 5732 17708 11020 17772
rect 11084 17708 11104 17772
rect 5732 17692 11104 17708
rect 5732 17628 11020 17692
rect 11084 17628 11104 17692
rect 5732 17612 11104 17628
rect 5732 17548 11020 17612
rect 11084 17548 11104 17612
rect 5732 17532 11104 17548
rect 5732 17468 11020 17532
rect 11084 17468 11104 17532
rect 5732 17452 11104 17468
rect 5732 17388 11020 17452
rect 11084 17388 11104 17452
rect 5732 17372 11104 17388
rect 5732 17308 11020 17372
rect 11084 17308 11104 17372
rect 5732 17292 11104 17308
rect 5732 17228 11020 17292
rect 11084 17228 11104 17292
rect 5732 17212 11104 17228
rect 5732 17148 11020 17212
rect 11084 17148 11104 17212
rect 5732 17132 11104 17148
rect 5732 17068 11020 17132
rect 11084 17068 11104 17132
rect 5732 17052 11104 17068
rect 5732 16988 11020 17052
rect 11084 16988 11104 17052
rect 5732 16972 11104 16988
rect 5732 16908 11020 16972
rect 11084 16908 11104 16972
rect 5732 16892 11104 16908
rect 5732 16828 11020 16892
rect 11084 16828 11104 16892
rect 5732 16812 11104 16828
rect 5732 16748 11020 16812
rect 11084 16748 11104 16812
rect 5732 16732 11104 16748
rect 5732 16668 11020 16732
rect 11084 16668 11104 16732
rect 5732 16652 11104 16668
rect 5732 16588 11020 16652
rect 11084 16588 11104 16652
rect 5732 16572 11104 16588
rect 5732 16508 11020 16572
rect 11084 16508 11104 16572
rect 5732 16492 11104 16508
rect 5732 16428 11020 16492
rect 11084 16428 11104 16492
rect 5732 16412 11104 16428
rect 5732 16348 11020 16412
rect 11084 16348 11104 16412
rect 5732 16332 11104 16348
rect 5732 16268 11020 16332
rect 11084 16268 11104 16332
rect 5732 16252 11104 16268
rect 5732 16188 11020 16252
rect 11084 16188 11104 16252
rect 5732 16172 11104 16188
rect 5732 16108 11020 16172
rect 11084 16108 11104 16172
rect 5732 16080 11104 16108
rect 11344 21132 16716 21160
rect 11344 21068 16632 21132
rect 16696 21068 16716 21132
rect 11344 21052 16716 21068
rect 11344 20988 16632 21052
rect 16696 20988 16716 21052
rect 11344 20972 16716 20988
rect 11344 20908 16632 20972
rect 16696 20908 16716 20972
rect 11344 20892 16716 20908
rect 11344 20828 16632 20892
rect 16696 20828 16716 20892
rect 11344 20812 16716 20828
rect 11344 20748 16632 20812
rect 16696 20748 16716 20812
rect 11344 20732 16716 20748
rect 11344 20668 16632 20732
rect 16696 20668 16716 20732
rect 11344 20652 16716 20668
rect 11344 20588 16632 20652
rect 16696 20588 16716 20652
rect 11344 20572 16716 20588
rect 11344 20508 16632 20572
rect 16696 20508 16716 20572
rect 11344 20492 16716 20508
rect 11344 20428 16632 20492
rect 16696 20428 16716 20492
rect 11344 20412 16716 20428
rect 11344 20348 16632 20412
rect 16696 20348 16716 20412
rect 11344 20332 16716 20348
rect 11344 20268 16632 20332
rect 16696 20268 16716 20332
rect 11344 20252 16716 20268
rect 11344 20188 16632 20252
rect 16696 20188 16716 20252
rect 11344 20172 16716 20188
rect 11344 20108 16632 20172
rect 16696 20108 16716 20172
rect 11344 20092 16716 20108
rect 11344 20028 16632 20092
rect 16696 20028 16716 20092
rect 11344 20012 16716 20028
rect 11344 19948 16632 20012
rect 16696 19948 16716 20012
rect 11344 19932 16716 19948
rect 11344 19868 16632 19932
rect 16696 19868 16716 19932
rect 11344 19852 16716 19868
rect 11344 19788 16632 19852
rect 16696 19788 16716 19852
rect 11344 19772 16716 19788
rect 11344 19708 16632 19772
rect 16696 19708 16716 19772
rect 11344 19692 16716 19708
rect 11344 19628 16632 19692
rect 16696 19628 16716 19692
rect 11344 19612 16716 19628
rect 11344 19548 16632 19612
rect 16696 19548 16716 19612
rect 11344 19532 16716 19548
rect 11344 19468 16632 19532
rect 16696 19468 16716 19532
rect 11344 19452 16716 19468
rect 11344 19388 16632 19452
rect 16696 19388 16716 19452
rect 11344 19372 16716 19388
rect 11344 19308 16632 19372
rect 16696 19308 16716 19372
rect 11344 19292 16716 19308
rect 11344 19228 16632 19292
rect 16696 19228 16716 19292
rect 11344 19212 16716 19228
rect 11344 19148 16632 19212
rect 16696 19148 16716 19212
rect 11344 19132 16716 19148
rect 11344 19068 16632 19132
rect 16696 19068 16716 19132
rect 11344 19052 16716 19068
rect 11344 18988 16632 19052
rect 16696 18988 16716 19052
rect 11344 18972 16716 18988
rect 11344 18908 16632 18972
rect 16696 18908 16716 18972
rect 11344 18892 16716 18908
rect 11344 18828 16632 18892
rect 16696 18828 16716 18892
rect 11344 18812 16716 18828
rect 11344 18748 16632 18812
rect 16696 18748 16716 18812
rect 11344 18732 16716 18748
rect 11344 18668 16632 18732
rect 16696 18668 16716 18732
rect 11344 18652 16716 18668
rect 11344 18588 16632 18652
rect 16696 18588 16716 18652
rect 11344 18572 16716 18588
rect 11344 18508 16632 18572
rect 16696 18508 16716 18572
rect 11344 18492 16716 18508
rect 11344 18428 16632 18492
rect 16696 18428 16716 18492
rect 11344 18412 16716 18428
rect 11344 18348 16632 18412
rect 16696 18348 16716 18412
rect 11344 18332 16716 18348
rect 11344 18268 16632 18332
rect 16696 18268 16716 18332
rect 11344 18252 16716 18268
rect 11344 18188 16632 18252
rect 16696 18188 16716 18252
rect 11344 18172 16716 18188
rect 11344 18108 16632 18172
rect 16696 18108 16716 18172
rect 11344 18092 16716 18108
rect 11344 18028 16632 18092
rect 16696 18028 16716 18092
rect 11344 18012 16716 18028
rect 11344 17948 16632 18012
rect 16696 17948 16716 18012
rect 11344 17932 16716 17948
rect 11344 17868 16632 17932
rect 16696 17868 16716 17932
rect 11344 17852 16716 17868
rect 11344 17788 16632 17852
rect 16696 17788 16716 17852
rect 11344 17772 16716 17788
rect 11344 17708 16632 17772
rect 16696 17708 16716 17772
rect 11344 17692 16716 17708
rect 11344 17628 16632 17692
rect 16696 17628 16716 17692
rect 11344 17612 16716 17628
rect 11344 17548 16632 17612
rect 16696 17548 16716 17612
rect 11344 17532 16716 17548
rect 11344 17468 16632 17532
rect 16696 17468 16716 17532
rect 11344 17452 16716 17468
rect 11344 17388 16632 17452
rect 16696 17388 16716 17452
rect 11344 17372 16716 17388
rect 11344 17308 16632 17372
rect 16696 17308 16716 17372
rect 11344 17292 16716 17308
rect 11344 17228 16632 17292
rect 16696 17228 16716 17292
rect 11344 17212 16716 17228
rect 11344 17148 16632 17212
rect 16696 17148 16716 17212
rect 11344 17132 16716 17148
rect 11344 17068 16632 17132
rect 16696 17068 16716 17132
rect 11344 17052 16716 17068
rect 11344 16988 16632 17052
rect 16696 16988 16716 17052
rect 11344 16972 16716 16988
rect 11344 16908 16632 16972
rect 16696 16908 16716 16972
rect 11344 16892 16716 16908
rect 11344 16828 16632 16892
rect 16696 16828 16716 16892
rect 11344 16812 16716 16828
rect 11344 16748 16632 16812
rect 16696 16748 16716 16812
rect 11344 16732 16716 16748
rect 11344 16668 16632 16732
rect 16696 16668 16716 16732
rect 11344 16652 16716 16668
rect 11344 16588 16632 16652
rect 16696 16588 16716 16652
rect 11344 16572 16716 16588
rect 11344 16508 16632 16572
rect 16696 16508 16716 16572
rect 11344 16492 16716 16508
rect 11344 16428 16632 16492
rect 16696 16428 16716 16492
rect 11344 16412 16716 16428
rect 11344 16348 16632 16412
rect 16696 16348 16716 16412
rect 11344 16332 16716 16348
rect 11344 16268 16632 16332
rect 16696 16268 16716 16332
rect 11344 16252 16716 16268
rect 11344 16188 16632 16252
rect 16696 16188 16716 16252
rect 11344 16172 16716 16188
rect 11344 16108 16632 16172
rect 16696 16108 16716 16172
rect 11344 16080 16716 16108
rect 16956 21132 22328 21160
rect 16956 21068 22244 21132
rect 22308 21068 22328 21132
rect 16956 21052 22328 21068
rect 16956 20988 22244 21052
rect 22308 20988 22328 21052
rect 16956 20972 22328 20988
rect 16956 20908 22244 20972
rect 22308 20908 22328 20972
rect 16956 20892 22328 20908
rect 16956 20828 22244 20892
rect 22308 20828 22328 20892
rect 16956 20812 22328 20828
rect 16956 20748 22244 20812
rect 22308 20748 22328 20812
rect 16956 20732 22328 20748
rect 16956 20668 22244 20732
rect 22308 20668 22328 20732
rect 16956 20652 22328 20668
rect 16956 20588 22244 20652
rect 22308 20588 22328 20652
rect 16956 20572 22328 20588
rect 16956 20508 22244 20572
rect 22308 20508 22328 20572
rect 16956 20492 22328 20508
rect 16956 20428 22244 20492
rect 22308 20428 22328 20492
rect 16956 20412 22328 20428
rect 16956 20348 22244 20412
rect 22308 20348 22328 20412
rect 16956 20332 22328 20348
rect 16956 20268 22244 20332
rect 22308 20268 22328 20332
rect 16956 20252 22328 20268
rect 16956 20188 22244 20252
rect 22308 20188 22328 20252
rect 16956 20172 22328 20188
rect 16956 20108 22244 20172
rect 22308 20108 22328 20172
rect 16956 20092 22328 20108
rect 16956 20028 22244 20092
rect 22308 20028 22328 20092
rect 16956 20012 22328 20028
rect 16956 19948 22244 20012
rect 22308 19948 22328 20012
rect 16956 19932 22328 19948
rect 16956 19868 22244 19932
rect 22308 19868 22328 19932
rect 16956 19852 22328 19868
rect 16956 19788 22244 19852
rect 22308 19788 22328 19852
rect 16956 19772 22328 19788
rect 16956 19708 22244 19772
rect 22308 19708 22328 19772
rect 16956 19692 22328 19708
rect 16956 19628 22244 19692
rect 22308 19628 22328 19692
rect 16956 19612 22328 19628
rect 16956 19548 22244 19612
rect 22308 19548 22328 19612
rect 16956 19532 22328 19548
rect 16956 19468 22244 19532
rect 22308 19468 22328 19532
rect 16956 19452 22328 19468
rect 16956 19388 22244 19452
rect 22308 19388 22328 19452
rect 16956 19372 22328 19388
rect 16956 19308 22244 19372
rect 22308 19308 22328 19372
rect 16956 19292 22328 19308
rect 16956 19228 22244 19292
rect 22308 19228 22328 19292
rect 16956 19212 22328 19228
rect 16956 19148 22244 19212
rect 22308 19148 22328 19212
rect 16956 19132 22328 19148
rect 16956 19068 22244 19132
rect 22308 19068 22328 19132
rect 16956 19052 22328 19068
rect 16956 18988 22244 19052
rect 22308 18988 22328 19052
rect 16956 18972 22328 18988
rect 16956 18908 22244 18972
rect 22308 18908 22328 18972
rect 16956 18892 22328 18908
rect 16956 18828 22244 18892
rect 22308 18828 22328 18892
rect 16956 18812 22328 18828
rect 16956 18748 22244 18812
rect 22308 18748 22328 18812
rect 16956 18732 22328 18748
rect 16956 18668 22244 18732
rect 22308 18668 22328 18732
rect 16956 18652 22328 18668
rect 16956 18588 22244 18652
rect 22308 18588 22328 18652
rect 16956 18572 22328 18588
rect 16956 18508 22244 18572
rect 22308 18508 22328 18572
rect 16956 18492 22328 18508
rect 16956 18428 22244 18492
rect 22308 18428 22328 18492
rect 16956 18412 22328 18428
rect 16956 18348 22244 18412
rect 22308 18348 22328 18412
rect 16956 18332 22328 18348
rect 16956 18268 22244 18332
rect 22308 18268 22328 18332
rect 16956 18252 22328 18268
rect 16956 18188 22244 18252
rect 22308 18188 22328 18252
rect 16956 18172 22328 18188
rect 16956 18108 22244 18172
rect 22308 18108 22328 18172
rect 16956 18092 22328 18108
rect 16956 18028 22244 18092
rect 22308 18028 22328 18092
rect 16956 18012 22328 18028
rect 16956 17948 22244 18012
rect 22308 17948 22328 18012
rect 16956 17932 22328 17948
rect 16956 17868 22244 17932
rect 22308 17868 22328 17932
rect 16956 17852 22328 17868
rect 16956 17788 22244 17852
rect 22308 17788 22328 17852
rect 16956 17772 22328 17788
rect 16956 17708 22244 17772
rect 22308 17708 22328 17772
rect 16956 17692 22328 17708
rect 16956 17628 22244 17692
rect 22308 17628 22328 17692
rect 16956 17612 22328 17628
rect 16956 17548 22244 17612
rect 22308 17548 22328 17612
rect 16956 17532 22328 17548
rect 16956 17468 22244 17532
rect 22308 17468 22328 17532
rect 16956 17452 22328 17468
rect 16956 17388 22244 17452
rect 22308 17388 22328 17452
rect 16956 17372 22328 17388
rect 16956 17308 22244 17372
rect 22308 17308 22328 17372
rect 16956 17292 22328 17308
rect 16956 17228 22244 17292
rect 22308 17228 22328 17292
rect 16956 17212 22328 17228
rect 16956 17148 22244 17212
rect 22308 17148 22328 17212
rect 16956 17132 22328 17148
rect 16956 17068 22244 17132
rect 22308 17068 22328 17132
rect 16956 17052 22328 17068
rect 16956 16988 22244 17052
rect 22308 16988 22328 17052
rect 16956 16972 22328 16988
rect 16956 16908 22244 16972
rect 22308 16908 22328 16972
rect 16956 16892 22328 16908
rect 16956 16828 22244 16892
rect 22308 16828 22328 16892
rect 16956 16812 22328 16828
rect 16956 16748 22244 16812
rect 22308 16748 22328 16812
rect 16956 16732 22328 16748
rect 16956 16668 22244 16732
rect 22308 16668 22328 16732
rect 16956 16652 22328 16668
rect 16956 16588 22244 16652
rect 22308 16588 22328 16652
rect 16956 16572 22328 16588
rect 16956 16508 22244 16572
rect 22308 16508 22328 16572
rect 16956 16492 22328 16508
rect 16956 16428 22244 16492
rect 22308 16428 22328 16492
rect 16956 16412 22328 16428
rect 16956 16348 22244 16412
rect 22308 16348 22328 16412
rect 16956 16332 22328 16348
rect 16956 16268 22244 16332
rect 22308 16268 22328 16332
rect 16956 16252 22328 16268
rect 16956 16188 22244 16252
rect 22308 16188 22328 16252
rect 16956 16172 22328 16188
rect 16956 16108 22244 16172
rect 22308 16108 22328 16172
rect 16956 16080 22328 16108
rect 22568 21132 27940 21160
rect 22568 21068 27856 21132
rect 27920 21068 27940 21132
rect 22568 21052 27940 21068
rect 22568 20988 27856 21052
rect 27920 20988 27940 21052
rect 22568 20972 27940 20988
rect 22568 20908 27856 20972
rect 27920 20908 27940 20972
rect 22568 20892 27940 20908
rect 22568 20828 27856 20892
rect 27920 20828 27940 20892
rect 22568 20812 27940 20828
rect 22568 20748 27856 20812
rect 27920 20748 27940 20812
rect 22568 20732 27940 20748
rect 22568 20668 27856 20732
rect 27920 20668 27940 20732
rect 22568 20652 27940 20668
rect 22568 20588 27856 20652
rect 27920 20588 27940 20652
rect 22568 20572 27940 20588
rect 22568 20508 27856 20572
rect 27920 20508 27940 20572
rect 22568 20492 27940 20508
rect 22568 20428 27856 20492
rect 27920 20428 27940 20492
rect 22568 20412 27940 20428
rect 22568 20348 27856 20412
rect 27920 20348 27940 20412
rect 22568 20332 27940 20348
rect 22568 20268 27856 20332
rect 27920 20268 27940 20332
rect 22568 20252 27940 20268
rect 22568 20188 27856 20252
rect 27920 20188 27940 20252
rect 22568 20172 27940 20188
rect 22568 20108 27856 20172
rect 27920 20108 27940 20172
rect 22568 20092 27940 20108
rect 22568 20028 27856 20092
rect 27920 20028 27940 20092
rect 22568 20012 27940 20028
rect 22568 19948 27856 20012
rect 27920 19948 27940 20012
rect 22568 19932 27940 19948
rect 22568 19868 27856 19932
rect 27920 19868 27940 19932
rect 22568 19852 27940 19868
rect 22568 19788 27856 19852
rect 27920 19788 27940 19852
rect 22568 19772 27940 19788
rect 22568 19708 27856 19772
rect 27920 19708 27940 19772
rect 22568 19692 27940 19708
rect 22568 19628 27856 19692
rect 27920 19628 27940 19692
rect 22568 19612 27940 19628
rect 22568 19548 27856 19612
rect 27920 19548 27940 19612
rect 22568 19532 27940 19548
rect 22568 19468 27856 19532
rect 27920 19468 27940 19532
rect 22568 19452 27940 19468
rect 22568 19388 27856 19452
rect 27920 19388 27940 19452
rect 22568 19372 27940 19388
rect 22568 19308 27856 19372
rect 27920 19308 27940 19372
rect 22568 19292 27940 19308
rect 22568 19228 27856 19292
rect 27920 19228 27940 19292
rect 22568 19212 27940 19228
rect 22568 19148 27856 19212
rect 27920 19148 27940 19212
rect 22568 19132 27940 19148
rect 22568 19068 27856 19132
rect 27920 19068 27940 19132
rect 22568 19052 27940 19068
rect 22568 18988 27856 19052
rect 27920 18988 27940 19052
rect 22568 18972 27940 18988
rect 22568 18908 27856 18972
rect 27920 18908 27940 18972
rect 22568 18892 27940 18908
rect 22568 18828 27856 18892
rect 27920 18828 27940 18892
rect 22568 18812 27940 18828
rect 22568 18748 27856 18812
rect 27920 18748 27940 18812
rect 22568 18732 27940 18748
rect 22568 18668 27856 18732
rect 27920 18668 27940 18732
rect 22568 18652 27940 18668
rect 22568 18588 27856 18652
rect 27920 18588 27940 18652
rect 22568 18572 27940 18588
rect 22568 18508 27856 18572
rect 27920 18508 27940 18572
rect 22568 18492 27940 18508
rect 22568 18428 27856 18492
rect 27920 18428 27940 18492
rect 22568 18412 27940 18428
rect 22568 18348 27856 18412
rect 27920 18348 27940 18412
rect 22568 18332 27940 18348
rect 22568 18268 27856 18332
rect 27920 18268 27940 18332
rect 22568 18252 27940 18268
rect 22568 18188 27856 18252
rect 27920 18188 27940 18252
rect 22568 18172 27940 18188
rect 22568 18108 27856 18172
rect 27920 18108 27940 18172
rect 22568 18092 27940 18108
rect 22568 18028 27856 18092
rect 27920 18028 27940 18092
rect 22568 18012 27940 18028
rect 22568 17948 27856 18012
rect 27920 17948 27940 18012
rect 22568 17932 27940 17948
rect 22568 17868 27856 17932
rect 27920 17868 27940 17932
rect 22568 17852 27940 17868
rect 22568 17788 27856 17852
rect 27920 17788 27940 17852
rect 22568 17772 27940 17788
rect 22568 17708 27856 17772
rect 27920 17708 27940 17772
rect 22568 17692 27940 17708
rect 22568 17628 27856 17692
rect 27920 17628 27940 17692
rect 22568 17612 27940 17628
rect 22568 17548 27856 17612
rect 27920 17548 27940 17612
rect 22568 17532 27940 17548
rect 22568 17468 27856 17532
rect 27920 17468 27940 17532
rect 22568 17452 27940 17468
rect 22568 17388 27856 17452
rect 27920 17388 27940 17452
rect 22568 17372 27940 17388
rect 22568 17308 27856 17372
rect 27920 17308 27940 17372
rect 22568 17292 27940 17308
rect 22568 17228 27856 17292
rect 27920 17228 27940 17292
rect 22568 17212 27940 17228
rect 22568 17148 27856 17212
rect 27920 17148 27940 17212
rect 22568 17132 27940 17148
rect 22568 17068 27856 17132
rect 27920 17068 27940 17132
rect 22568 17052 27940 17068
rect 22568 16988 27856 17052
rect 27920 16988 27940 17052
rect 22568 16972 27940 16988
rect 22568 16908 27856 16972
rect 27920 16908 27940 16972
rect 22568 16892 27940 16908
rect 22568 16828 27856 16892
rect 27920 16828 27940 16892
rect 22568 16812 27940 16828
rect 22568 16748 27856 16812
rect 27920 16748 27940 16812
rect 22568 16732 27940 16748
rect 22568 16668 27856 16732
rect 27920 16668 27940 16732
rect 22568 16652 27940 16668
rect 22568 16588 27856 16652
rect 27920 16588 27940 16652
rect 22568 16572 27940 16588
rect 22568 16508 27856 16572
rect 27920 16508 27940 16572
rect 22568 16492 27940 16508
rect 22568 16428 27856 16492
rect 27920 16428 27940 16492
rect 22568 16412 27940 16428
rect 22568 16348 27856 16412
rect 27920 16348 27940 16412
rect 22568 16332 27940 16348
rect 22568 16268 27856 16332
rect 27920 16268 27940 16332
rect 22568 16252 27940 16268
rect 22568 16188 27856 16252
rect 27920 16188 27940 16252
rect 22568 16172 27940 16188
rect 22568 16108 27856 16172
rect 27920 16108 27940 16172
rect 22568 16080 27940 16108
rect 28180 21132 33552 21160
rect 28180 21068 33468 21132
rect 33532 21068 33552 21132
rect 28180 21052 33552 21068
rect 28180 20988 33468 21052
rect 33532 20988 33552 21052
rect 28180 20972 33552 20988
rect 28180 20908 33468 20972
rect 33532 20908 33552 20972
rect 28180 20892 33552 20908
rect 28180 20828 33468 20892
rect 33532 20828 33552 20892
rect 28180 20812 33552 20828
rect 28180 20748 33468 20812
rect 33532 20748 33552 20812
rect 28180 20732 33552 20748
rect 28180 20668 33468 20732
rect 33532 20668 33552 20732
rect 28180 20652 33552 20668
rect 28180 20588 33468 20652
rect 33532 20588 33552 20652
rect 28180 20572 33552 20588
rect 28180 20508 33468 20572
rect 33532 20508 33552 20572
rect 28180 20492 33552 20508
rect 28180 20428 33468 20492
rect 33532 20428 33552 20492
rect 28180 20412 33552 20428
rect 28180 20348 33468 20412
rect 33532 20348 33552 20412
rect 28180 20332 33552 20348
rect 28180 20268 33468 20332
rect 33532 20268 33552 20332
rect 28180 20252 33552 20268
rect 28180 20188 33468 20252
rect 33532 20188 33552 20252
rect 28180 20172 33552 20188
rect 28180 20108 33468 20172
rect 33532 20108 33552 20172
rect 28180 20092 33552 20108
rect 28180 20028 33468 20092
rect 33532 20028 33552 20092
rect 28180 20012 33552 20028
rect 28180 19948 33468 20012
rect 33532 19948 33552 20012
rect 28180 19932 33552 19948
rect 28180 19868 33468 19932
rect 33532 19868 33552 19932
rect 28180 19852 33552 19868
rect 28180 19788 33468 19852
rect 33532 19788 33552 19852
rect 28180 19772 33552 19788
rect 28180 19708 33468 19772
rect 33532 19708 33552 19772
rect 28180 19692 33552 19708
rect 28180 19628 33468 19692
rect 33532 19628 33552 19692
rect 28180 19612 33552 19628
rect 28180 19548 33468 19612
rect 33532 19548 33552 19612
rect 28180 19532 33552 19548
rect 28180 19468 33468 19532
rect 33532 19468 33552 19532
rect 28180 19452 33552 19468
rect 28180 19388 33468 19452
rect 33532 19388 33552 19452
rect 28180 19372 33552 19388
rect 28180 19308 33468 19372
rect 33532 19308 33552 19372
rect 28180 19292 33552 19308
rect 28180 19228 33468 19292
rect 33532 19228 33552 19292
rect 28180 19212 33552 19228
rect 28180 19148 33468 19212
rect 33532 19148 33552 19212
rect 28180 19132 33552 19148
rect 28180 19068 33468 19132
rect 33532 19068 33552 19132
rect 28180 19052 33552 19068
rect 28180 18988 33468 19052
rect 33532 18988 33552 19052
rect 28180 18972 33552 18988
rect 28180 18908 33468 18972
rect 33532 18908 33552 18972
rect 28180 18892 33552 18908
rect 28180 18828 33468 18892
rect 33532 18828 33552 18892
rect 28180 18812 33552 18828
rect 28180 18748 33468 18812
rect 33532 18748 33552 18812
rect 28180 18732 33552 18748
rect 28180 18668 33468 18732
rect 33532 18668 33552 18732
rect 28180 18652 33552 18668
rect 28180 18588 33468 18652
rect 33532 18588 33552 18652
rect 28180 18572 33552 18588
rect 28180 18508 33468 18572
rect 33532 18508 33552 18572
rect 28180 18492 33552 18508
rect 28180 18428 33468 18492
rect 33532 18428 33552 18492
rect 28180 18412 33552 18428
rect 28180 18348 33468 18412
rect 33532 18348 33552 18412
rect 28180 18332 33552 18348
rect 28180 18268 33468 18332
rect 33532 18268 33552 18332
rect 28180 18252 33552 18268
rect 28180 18188 33468 18252
rect 33532 18188 33552 18252
rect 28180 18172 33552 18188
rect 28180 18108 33468 18172
rect 33532 18108 33552 18172
rect 28180 18092 33552 18108
rect 28180 18028 33468 18092
rect 33532 18028 33552 18092
rect 28180 18012 33552 18028
rect 28180 17948 33468 18012
rect 33532 17948 33552 18012
rect 28180 17932 33552 17948
rect 28180 17868 33468 17932
rect 33532 17868 33552 17932
rect 28180 17852 33552 17868
rect 28180 17788 33468 17852
rect 33532 17788 33552 17852
rect 28180 17772 33552 17788
rect 28180 17708 33468 17772
rect 33532 17708 33552 17772
rect 28180 17692 33552 17708
rect 28180 17628 33468 17692
rect 33532 17628 33552 17692
rect 28180 17612 33552 17628
rect 28180 17548 33468 17612
rect 33532 17548 33552 17612
rect 28180 17532 33552 17548
rect 28180 17468 33468 17532
rect 33532 17468 33552 17532
rect 28180 17452 33552 17468
rect 28180 17388 33468 17452
rect 33532 17388 33552 17452
rect 28180 17372 33552 17388
rect 28180 17308 33468 17372
rect 33532 17308 33552 17372
rect 28180 17292 33552 17308
rect 28180 17228 33468 17292
rect 33532 17228 33552 17292
rect 28180 17212 33552 17228
rect 28180 17148 33468 17212
rect 33532 17148 33552 17212
rect 28180 17132 33552 17148
rect 28180 17068 33468 17132
rect 33532 17068 33552 17132
rect 28180 17052 33552 17068
rect 28180 16988 33468 17052
rect 33532 16988 33552 17052
rect 28180 16972 33552 16988
rect 28180 16908 33468 16972
rect 33532 16908 33552 16972
rect 28180 16892 33552 16908
rect 28180 16828 33468 16892
rect 33532 16828 33552 16892
rect 28180 16812 33552 16828
rect 28180 16748 33468 16812
rect 33532 16748 33552 16812
rect 28180 16732 33552 16748
rect 28180 16668 33468 16732
rect 33532 16668 33552 16732
rect 28180 16652 33552 16668
rect 28180 16588 33468 16652
rect 33532 16588 33552 16652
rect 28180 16572 33552 16588
rect 28180 16508 33468 16572
rect 33532 16508 33552 16572
rect 28180 16492 33552 16508
rect 28180 16428 33468 16492
rect 33532 16428 33552 16492
rect 28180 16412 33552 16428
rect 28180 16348 33468 16412
rect 33532 16348 33552 16412
rect 28180 16332 33552 16348
rect 28180 16268 33468 16332
rect 33532 16268 33552 16332
rect 28180 16252 33552 16268
rect 28180 16188 33468 16252
rect 33532 16188 33552 16252
rect 28180 16172 33552 16188
rect 28180 16108 33468 16172
rect 33532 16108 33552 16172
rect 28180 16080 33552 16108
rect 33792 21132 39164 21160
rect 33792 21068 39080 21132
rect 39144 21068 39164 21132
rect 33792 21052 39164 21068
rect 33792 20988 39080 21052
rect 39144 20988 39164 21052
rect 33792 20972 39164 20988
rect 33792 20908 39080 20972
rect 39144 20908 39164 20972
rect 33792 20892 39164 20908
rect 33792 20828 39080 20892
rect 39144 20828 39164 20892
rect 33792 20812 39164 20828
rect 33792 20748 39080 20812
rect 39144 20748 39164 20812
rect 33792 20732 39164 20748
rect 33792 20668 39080 20732
rect 39144 20668 39164 20732
rect 33792 20652 39164 20668
rect 33792 20588 39080 20652
rect 39144 20588 39164 20652
rect 33792 20572 39164 20588
rect 33792 20508 39080 20572
rect 39144 20508 39164 20572
rect 33792 20492 39164 20508
rect 33792 20428 39080 20492
rect 39144 20428 39164 20492
rect 33792 20412 39164 20428
rect 33792 20348 39080 20412
rect 39144 20348 39164 20412
rect 33792 20332 39164 20348
rect 33792 20268 39080 20332
rect 39144 20268 39164 20332
rect 33792 20252 39164 20268
rect 33792 20188 39080 20252
rect 39144 20188 39164 20252
rect 33792 20172 39164 20188
rect 33792 20108 39080 20172
rect 39144 20108 39164 20172
rect 33792 20092 39164 20108
rect 33792 20028 39080 20092
rect 39144 20028 39164 20092
rect 33792 20012 39164 20028
rect 33792 19948 39080 20012
rect 39144 19948 39164 20012
rect 33792 19932 39164 19948
rect 33792 19868 39080 19932
rect 39144 19868 39164 19932
rect 33792 19852 39164 19868
rect 33792 19788 39080 19852
rect 39144 19788 39164 19852
rect 33792 19772 39164 19788
rect 33792 19708 39080 19772
rect 39144 19708 39164 19772
rect 33792 19692 39164 19708
rect 33792 19628 39080 19692
rect 39144 19628 39164 19692
rect 33792 19612 39164 19628
rect 33792 19548 39080 19612
rect 39144 19548 39164 19612
rect 33792 19532 39164 19548
rect 33792 19468 39080 19532
rect 39144 19468 39164 19532
rect 33792 19452 39164 19468
rect 33792 19388 39080 19452
rect 39144 19388 39164 19452
rect 33792 19372 39164 19388
rect 33792 19308 39080 19372
rect 39144 19308 39164 19372
rect 33792 19292 39164 19308
rect 33792 19228 39080 19292
rect 39144 19228 39164 19292
rect 33792 19212 39164 19228
rect 33792 19148 39080 19212
rect 39144 19148 39164 19212
rect 33792 19132 39164 19148
rect 33792 19068 39080 19132
rect 39144 19068 39164 19132
rect 33792 19052 39164 19068
rect 33792 18988 39080 19052
rect 39144 18988 39164 19052
rect 33792 18972 39164 18988
rect 33792 18908 39080 18972
rect 39144 18908 39164 18972
rect 33792 18892 39164 18908
rect 33792 18828 39080 18892
rect 39144 18828 39164 18892
rect 33792 18812 39164 18828
rect 33792 18748 39080 18812
rect 39144 18748 39164 18812
rect 33792 18732 39164 18748
rect 33792 18668 39080 18732
rect 39144 18668 39164 18732
rect 33792 18652 39164 18668
rect 33792 18588 39080 18652
rect 39144 18588 39164 18652
rect 33792 18572 39164 18588
rect 33792 18508 39080 18572
rect 39144 18508 39164 18572
rect 33792 18492 39164 18508
rect 33792 18428 39080 18492
rect 39144 18428 39164 18492
rect 33792 18412 39164 18428
rect 33792 18348 39080 18412
rect 39144 18348 39164 18412
rect 33792 18332 39164 18348
rect 33792 18268 39080 18332
rect 39144 18268 39164 18332
rect 33792 18252 39164 18268
rect 33792 18188 39080 18252
rect 39144 18188 39164 18252
rect 33792 18172 39164 18188
rect 33792 18108 39080 18172
rect 39144 18108 39164 18172
rect 33792 18092 39164 18108
rect 33792 18028 39080 18092
rect 39144 18028 39164 18092
rect 33792 18012 39164 18028
rect 33792 17948 39080 18012
rect 39144 17948 39164 18012
rect 33792 17932 39164 17948
rect 33792 17868 39080 17932
rect 39144 17868 39164 17932
rect 33792 17852 39164 17868
rect 33792 17788 39080 17852
rect 39144 17788 39164 17852
rect 33792 17772 39164 17788
rect 33792 17708 39080 17772
rect 39144 17708 39164 17772
rect 33792 17692 39164 17708
rect 33792 17628 39080 17692
rect 39144 17628 39164 17692
rect 33792 17612 39164 17628
rect 33792 17548 39080 17612
rect 39144 17548 39164 17612
rect 33792 17532 39164 17548
rect 33792 17468 39080 17532
rect 39144 17468 39164 17532
rect 33792 17452 39164 17468
rect 33792 17388 39080 17452
rect 39144 17388 39164 17452
rect 33792 17372 39164 17388
rect 33792 17308 39080 17372
rect 39144 17308 39164 17372
rect 33792 17292 39164 17308
rect 33792 17228 39080 17292
rect 39144 17228 39164 17292
rect 33792 17212 39164 17228
rect 33792 17148 39080 17212
rect 39144 17148 39164 17212
rect 33792 17132 39164 17148
rect 33792 17068 39080 17132
rect 39144 17068 39164 17132
rect 33792 17052 39164 17068
rect 33792 16988 39080 17052
rect 39144 16988 39164 17052
rect 33792 16972 39164 16988
rect 33792 16908 39080 16972
rect 39144 16908 39164 16972
rect 33792 16892 39164 16908
rect 33792 16828 39080 16892
rect 39144 16828 39164 16892
rect 33792 16812 39164 16828
rect 33792 16748 39080 16812
rect 39144 16748 39164 16812
rect 33792 16732 39164 16748
rect 33792 16668 39080 16732
rect 39144 16668 39164 16732
rect 33792 16652 39164 16668
rect 33792 16588 39080 16652
rect 39144 16588 39164 16652
rect 33792 16572 39164 16588
rect 33792 16508 39080 16572
rect 39144 16508 39164 16572
rect 33792 16492 39164 16508
rect 33792 16428 39080 16492
rect 39144 16428 39164 16492
rect 33792 16412 39164 16428
rect 33792 16348 39080 16412
rect 39144 16348 39164 16412
rect 33792 16332 39164 16348
rect 33792 16268 39080 16332
rect 39144 16268 39164 16332
rect 33792 16252 39164 16268
rect 33792 16188 39080 16252
rect 39144 16188 39164 16252
rect 33792 16172 39164 16188
rect 33792 16108 39080 16172
rect 39144 16108 39164 16172
rect 33792 16080 39164 16108
rect -39164 15812 -33792 15840
rect -39164 15748 -33876 15812
rect -33812 15748 -33792 15812
rect -39164 15732 -33792 15748
rect -39164 15668 -33876 15732
rect -33812 15668 -33792 15732
rect -39164 15652 -33792 15668
rect -39164 15588 -33876 15652
rect -33812 15588 -33792 15652
rect -39164 15572 -33792 15588
rect -39164 15508 -33876 15572
rect -33812 15508 -33792 15572
rect -39164 15492 -33792 15508
rect -39164 15428 -33876 15492
rect -33812 15428 -33792 15492
rect -39164 15412 -33792 15428
rect -39164 15348 -33876 15412
rect -33812 15348 -33792 15412
rect -39164 15332 -33792 15348
rect -39164 15268 -33876 15332
rect -33812 15268 -33792 15332
rect -39164 15252 -33792 15268
rect -39164 15188 -33876 15252
rect -33812 15188 -33792 15252
rect -39164 15172 -33792 15188
rect -39164 15108 -33876 15172
rect -33812 15108 -33792 15172
rect -39164 15092 -33792 15108
rect -39164 15028 -33876 15092
rect -33812 15028 -33792 15092
rect -39164 15012 -33792 15028
rect -39164 14948 -33876 15012
rect -33812 14948 -33792 15012
rect -39164 14932 -33792 14948
rect -39164 14868 -33876 14932
rect -33812 14868 -33792 14932
rect -39164 14852 -33792 14868
rect -39164 14788 -33876 14852
rect -33812 14788 -33792 14852
rect -39164 14772 -33792 14788
rect -39164 14708 -33876 14772
rect -33812 14708 -33792 14772
rect -39164 14692 -33792 14708
rect -39164 14628 -33876 14692
rect -33812 14628 -33792 14692
rect -39164 14612 -33792 14628
rect -39164 14548 -33876 14612
rect -33812 14548 -33792 14612
rect -39164 14532 -33792 14548
rect -39164 14468 -33876 14532
rect -33812 14468 -33792 14532
rect -39164 14452 -33792 14468
rect -39164 14388 -33876 14452
rect -33812 14388 -33792 14452
rect -39164 14372 -33792 14388
rect -39164 14308 -33876 14372
rect -33812 14308 -33792 14372
rect -39164 14292 -33792 14308
rect -39164 14228 -33876 14292
rect -33812 14228 -33792 14292
rect -39164 14212 -33792 14228
rect -39164 14148 -33876 14212
rect -33812 14148 -33792 14212
rect -39164 14132 -33792 14148
rect -39164 14068 -33876 14132
rect -33812 14068 -33792 14132
rect -39164 14052 -33792 14068
rect -39164 13988 -33876 14052
rect -33812 13988 -33792 14052
rect -39164 13972 -33792 13988
rect -39164 13908 -33876 13972
rect -33812 13908 -33792 13972
rect -39164 13892 -33792 13908
rect -39164 13828 -33876 13892
rect -33812 13828 -33792 13892
rect -39164 13812 -33792 13828
rect -39164 13748 -33876 13812
rect -33812 13748 -33792 13812
rect -39164 13732 -33792 13748
rect -39164 13668 -33876 13732
rect -33812 13668 -33792 13732
rect -39164 13652 -33792 13668
rect -39164 13588 -33876 13652
rect -33812 13588 -33792 13652
rect -39164 13572 -33792 13588
rect -39164 13508 -33876 13572
rect -33812 13508 -33792 13572
rect -39164 13492 -33792 13508
rect -39164 13428 -33876 13492
rect -33812 13428 -33792 13492
rect -39164 13412 -33792 13428
rect -39164 13348 -33876 13412
rect -33812 13348 -33792 13412
rect -39164 13332 -33792 13348
rect -39164 13268 -33876 13332
rect -33812 13268 -33792 13332
rect -39164 13252 -33792 13268
rect -39164 13188 -33876 13252
rect -33812 13188 -33792 13252
rect -39164 13172 -33792 13188
rect -39164 13108 -33876 13172
rect -33812 13108 -33792 13172
rect -39164 13092 -33792 13108
rect -39164 13028 -33876 13092
rect -33812 13028 -33792 13092
rect -39164 13012 -33792 13028
rect -39164 12948 -33876 13012
rect -33812 12948 -33792 13012
rect -39164 12932 -33792 12948
rect -39164 12868 -33876 12932
rect -33812 12868 -33792 12932
rect -39164 12852 -33792 12868
rect -39164 12788 -33876 12852
rect -33812 12788 -33792 12852
rect -39164 12772 -33792 12788
rect -39164 12708 -33876 12772
rect -33812 12708 -33792 12772
rect -39164 12692 -33792 12708
rect -39164 12628 -33876 12692
rect -33812 12628 -33792 12692
rect -39164 12612 -33792 12628
rect -39164 12548 -33876 12612
rect -33812 12548 -33792 12612
rect -39164 12532 -33792 12548
rect -39164 12468 -33876 12532
rect -33812 12468 -33792 12532
rect -39164 12452 -33792 12468
rect -39164 12388 -33876 12452
rect -33812 12388 -33792 12452
rect -39164 12372 -33792 12388
rect -39164 12308 -33876 12372
rect -33812 12308 -33792 12372
rect -39164 12292 -33792 12308
rect -39164 12228 -33876 12292
rect -33812 12228 -33792 12292
rect -39164 12212 -33792 12228
rect -39164 12148 -33876 12212
rect -33812 12148 -33792 12212
rect -39164 12132 -33792 12148
rect -39164 12068 -33876 12132
rect -33812 12068 -33792 12132
rect -39164 12052 -33792 12068
rect -39164 11988 -33876 12052
rect -33812 11988 -33792 12052
rect -39164 11972 -33792 11988
rect -39164 11908 -33876 11972
rect -33812 11908 -33792 11972
rect -39164 11892 -33792 11908
rect -39164 11828 -33876 11892
rect -33812 11828 -33792 11892
rect -39164 11812 -33792 11828
rect -39164 11748 -33876 11812
rect -33812 11748 -33792 11812
rect -39164 11732 -33792 11748
rect -39164 11668 -33876 11732
rect -33812 11668 -33792 11732
rect -39164 11652 -33792 11668
rect -39164 11588 -33876 11652
rect -33812 11588 -33792 11652
rect -39164 11572 -33792 11588
rect -39164 11508 -33876 11572
rect -33812 11508 -33792 11572
rect -39164 11492 -33792 11508
rect -39164 11428 -33876 11492
rect -33812 11428 -33792 11492
rect -39164 11412 -33792 11428
rect -39164 11348 -33876 11412
rect -33812 11348 -33792 11412
rect -39164 11332 -33792 11348
rect -39164 11268 -33876 11332
rect -33812 11268 -33792 11332
rect -39164 11252 -33792 11268
rect -39164 11188 -33876 11252
rect -33812 11188 -33792 11252
rect -39164 11172 -33792 11188
rect -39164 11108 -33876 11172
rect -33812 11108 -33792 11172
rect -39164 11092 -33792 11108
rect -39164 11028 -33876 11092
rect -33812 11028 -33792 11092
rect -39164 11012 -33792 11028
rect -39164 10948 -33876 11012
rect -33812 10948 -33792 11012
rect -39164 10932 -33792 10948
rect -39164 10868 -33876 10932
rect -33812 10868 -33792 10932
rect -39164 10852 -33792 10868
rect -39164 10788 -33876 10852
rect -33812 10788 -33792 10852
rect -39164 10760 -33792 10788
rect -33552 15812 -28180 15840
rect -33552 15748 -28264 15812
rect -28200 15748 -28180 15812
rect -33552 15732 -28180 15748
rect -33552 15668 -28264 15732
rect -28200 15668 -28180 15732
rect -33552 15652 -28180 15668
rect -33552 15588 -28264 15652
rect -28200 15588 -28180 15652
rect -33552 15572 -28180 15588
rect -33552 15508 -28264 15572
rect -28200 15508 -28180 15572
rect -33552 15492 -28180 15508
rect -33552 15428 -28264 15492
rect -28200 15428 -28180 15492
rect -33552 15412 -28180 15428
rect -33552 15348 -28264 15412
rect -28200 15348 -28180 15412
rect -33552 15332 -28180 15348
rect -33552 15268 -28264 15332
rect -28200 15268 -28180 15332
rect -33552 15252 -28180 15268
rect -33552 15188 -28264 15252
rect -28200 15188 -28180 15252
rect -33552 15172 -28180 15188
rect -33552 15108 -28264 15172
rect -28200 15108 -28180 15172
rect -33552 15092 -28180 15108
rect -33552 15028 -28264 15092
rect -28200 15028 -28180 15092
rect -33552 15012 -28180 15028
rect -33552 14948 -28264 15012
rect -28200 14948 -28180 15012
rect -33552 14932 -28180 14948
rect -33552 14868 -28264 14932
rect -28200 14868 -28180 14932
rect -33552 14852 -28180 14868
rect -33552 14788 -28264 14852
rect -28200 14788 -28180 14852
rect -33552 14772 -28180 14788
rect -33552 14708 -28264 14772
rect -28200 14708 -28180 14772
rect -33552 14692 -28180 14708
rect -33552 14628 -28264 14692
rect -28200 14628 -28180 14692
rect -33552 14612 -28180 14628
rect -33552 14548 -28264 14612
rect -28200 14548 -28180 14612
rect -33552 14532 -28180 14548
rect -33552 14468 -28264 14532
rect -28200 14468 -28180 14532
rect -33552 14452 -28180 14468
rect -33552 14388 -28264 14452
rect -28200 14388 -28180 14452
rect -33552 14372 -28180 14388
rect -33552 14308 -28264 14372
rect -28200 14308 -28180 14372
rect -33552 14292 -28180 14308
rect -33552 14228 -28264 14292
rect -28200 14228 -28180 14292
rect -33552 14212 -28180 14228
rect -33552 14148 -28264 14212
rect -28200 14148 -28180 14212
rect -33552 14132 -28180 14148
rect -33552 14068 -28264 14132
rect -28200 14068 -28180 14132
rect -33552 14052 -28180 14068
rect -33552 13988 -28264 14052
rect -28200 13988 -28180 14052
rect -33552 13972 -28180 13988
rect -33552 13908 -28264 13972
rect -28200 13908 -28180 13972
rect -33552 13892 -28180 13908
rect -33552 13828 -28264 13892
rect -28200 13828 -28180 13892
rect -33552 13812 -28180 13828
rect -33552 13748 -28264 13812
rect -28200 13748 -28180 13812
rect -33552 13732 -28180 13748
rect -33552 13668 -28264 13732
rect -28200 13668 -28180 13732
rect -33552 13652 -28180 13668
rect -33552 13588 -28264 13652
rect -28200 13588 -28180 13652
rect -33552 13572 -28180 13588
rect -33552 13508 -28264 13572
rect -28200 13508 -28180 13572
rect -33552 13492 -28180 13508
rect -33552 13428 -28264 13492
rect -28200 13428 -28180 13492
rect -33552 13412 -28180 13428
rect -33552 13348 -28264 13412
rect -28200 13348 -28180 13412
rect -33552 13332 -28180 13348
rect -33552 13268 -28264 13332
rect -28200 13268 -28180 13332
rect -33552 13252 -28180 13268
rect -33552 13188 -28264 13252
rect -28200 13188 -28180 13252
rect -33552 13172 -28180 13188
rect -33552 13108 -28264 13172
rect -28200 13108 -28180 13172
rect -33552 13092 -28180 13108
rect -33552 13028 -28264 13092
rect -28200 13028 -28180 13092
rect -33552 13012 -28180 13028
rect -33552 12948 -28264 13012
rect -28200 12948 -28180 13012
rect -33552 12932 -28180 12948
rect -33552 12868 -28264 12932
rect -28200 12868 -28180 12932
rect -33552 12852 -28180 12868
rect -33552 12788 -28264 12852
rect -28200 12788 -28180 12852
rect -33552 12772 -28180 12788
rect -33552 12708 -28264 12772
rect -28200 12708 -28180 12772
rect -33552 12692 -28180 12708
rect -33552 12628 -28264 12692
rect -28200 12628 -28180 12692
rect -33552 12612 -28180 12628
rect -33552 12548 -28264 12612
rect -28200 12548 -28180 12612
rect -33552 12532 -28180 12548
rect -33552 12468 -28264 12532
rect -28200 12468 -28180 12532
rect -33552 12452 -28180 12468
rect -33552 12388 -28264 12452
rect -28200 12388 -28180 12452
rect -33552 12372 -28180 12388
rect -33552 12308 -28264 12372
rect -28200 12308 -28180 12372
rect -33552 12292 -28180 12308
rect -33552 12228 -28264 12292
rect -28200 12228 -28180 12292
rect -33552 12212 -28180 12228
rect -33552 12148 -28264 12212
rect -28200 12148 -28180 12212
rect -33552 12132 -28180 12148
rect -33552 12068 -28264 12132
rect -28200 12068 -28180 12132
rect -33552 12052 -28180 12068
rect -33552 11988 -28264 12052
rect -28200 11988 -28180 12052
rect -33552 11972 -28180 11988
rect -33552 11908 -28264 11972
rect -28200 11908 -28180 11972
rect -33552 11892 -28180 11908
rect -33552 11828 -28264 11892
rect -28200 11828 -28180 11892
rect -33552 11812 -28180 11828
rect -33552 11748 -28264 11812
rect -28200 11748 -28180 11812
rect -33552 11732 -28180 11748
rect -33552 11668 -28264 11732
rect -28200 11668 -28180 11732
rect -33552 11652 -28180 11668
rect -33552 11588 -28264 11652
rect -28200 11588 -28180 11652
rect -33552 11572 -28180 11588
rect -33552 11508 -28264 11572
rect -28200 11508 -28180 11572
rect -33552 11492 -28180 11508
rect -33552 11428 -28264 11492
rect -28200 11428 -28180 11492
rect -33552 11412 -28180 11428
rect -33552 11348 -28264 11412
rect -28200 11348 -28180 11412
rect -33552 11332 -28180 11348
rect -33552 11268 -28264 11332
rect -28200 11268 -28180 11332
rect -33552 11252 -28180 11268
rect -33552 11188 -28264 11252
rect -28200 11188 -28180 11252
rect -33552 11172 -28180 11188
rect -33552 11108 -28264 11172
rect -28200 11108 -28180 11172
rect -33552 11092 -28180 11108
rect -33552 11028 -28264 11092
rect -28200 11028 -28180 11092
rect -33552 11012 -28180 11028
rect -33552 10948 -28264 11012
rect -28200 10948 -28180 11012
rect -33552 10932 -28180 10948
rect -33552 10868 -28264 10932
rect -28200 10868 -28180 10932
rect -33552 10852 -28180 10868
rect -33552 10788 -28264 10852
rect -28200 10788 -28180 10852
rect -33552 10760 -28180 10788
rect -27940 15812 -22568 15840
rect -27940 15748 -22652 15812
rect -22588 15748 -22568 15812
rect -27940 15732 -22568 15748
rect -27940 15668 -22652 15732
rect -22588 15668 -22568 15732
rect -27940 15652 -22568 15668
rect -27940 15588 -22652 15652
rect -22588 15588 -22568 15652
rect -27940 15572 -22568 15588
rect -27940 15508 -22652 15572
rect -22588 15508 -22568 15572
rect -27940 15492 -22568 15508
rect -27940 15428 -22652 15492
rect -22588 15428 -22568 15492
rect -27940 15412 -22568 15428
rect -27940 15348 -22652 15412
rect -22588 15348 -22568 15412
rect -27940 15332 -22568 15348
rect -27940 15268 -22652 15332
rect -22588 15268 -22568 15332
rect -27940 15252 -22568 15268
rect -27940 15188 -22652 15252
rect -22588 15188 -22568 15252
rect -27940 15172 -22568 15188
rect -27940 15108 -22652 15172
rect -22588 15108 -22568 15172
rect -27940 15092 -22568 15108
rect -27940 15028 -22652 15092
rect -22588 15028 -22568 15092
rect -27940 15012 -22568 15028
rect -27940 14948 -22652 15012
rect -22588 14948 -22568 15012
rect -27940 14932 -22568 14948
rect -27940 14868 -22652 14932
rect -22588 14868 -22568 14932
rect -27940 14852 -22568 14868
rect -27940 14788 -22652 14852
rect -22588 14788 -22568 14852
rect -27940 14772 -22568 14788
rect -27940 14708 -22652 14772
rect -22588 14708 -22568 14772
rect -27940 14692 -22568 14708
rect -27940 14628 -22652 14692
rect -22588 14628 -22568 14692
rect -27940 14612 -22568 14628
rect -27940 14548 -22652 14612
rect -22588 14548 -22568 14612
rect -27940 14532 -22568 14548
rect -27940 14468 -22652 14532
rect -22588 14468 -22568 14532
rect -27940 14452 -22568 14468
rect -27940 14388 -22652 14452
rect -22588 14388 -22568 14452
rect -27940 14372 -22568 14388
rect -27940 14308 -22652 14372
rect -22588 14308 -22568 14372
rect -27940 14292 -22568 14308
rect -27940 14228 -22652 14292
rect -22588 14228 -22568 14292
rect -27940 14212 -22568 14228
rect -27940 14148 -22652 14212
rect -22588 14148 -22568 14212
rect -27940 14132 -22568 14148
rect -27940 14068 -22652 14132
rect -22588 14068 -22568 14132
rect -27940 14052 -22568 14068
rect -27940 13988 -22652 14052
rect -22588 13988 -22568 14052
rect -27940 13972 -22568 13988
rect -27940 13908 -22652 13972
rect -22588 13908 -22568 13972
rect -27940 13892 -22568 13908
rect -27940 13828 -22652 13892
rect -22588 13828 -22568 13892
rect -27940 13812 -22568 13828
rect -27940 13748 -22652 13812
rect -22588 13748 -22568 13812
rect -27940 13732 -22568 13748
rect -27940 13668 -22652 13732
rect -22588 13668 -22568 13732
rect -27940 13652 -22568 13668
rect -27940 13588 -22652 13652
rect -22588 13588 -22568 13652
rect -27940 13572 -22568 13588
rect -27940 13508 -22652 13572
rect -22588 13508 -22568 13572
rect -27940 13492 -22568 13508
rect -27940 13428 -22652 13492
rect -22588 13428 -22568 13492
rect -27940 13412 -22568 13428
rect -27940 13348 -22652 13412
rect -22588 13348 -22568 13412
rect -27940 13332 -22568 13348
rect -27940 13268 -22652 13332
rect -22588 13268 -22568 13332
rect -27940 13252 -22568 13268
rect -27940 13188 -22652 13252
rect -22588 13188 -22568 13252
rect -27940 13172 -22568 13188
rect -27940 13108 -22652 13172
rect -22588 13108 -22568 13172
rect -27940 13092 -22568 13108
rect -27940 13028 -22652 13092
rect -22588 13028 -22568 13092
rect -27940 13012 -22568 13028
rect -27940 12948 -22652 13012
rect -22588 12948 -22568 13012
rect -27940 12932 -22568 12948
rect -27940 12868 -22652 12932
rect -22588 12868 -22568 12932
rect -27940 12852 -22568 12868
rect -27940 12788 -22652 12852
rect -22588 12788 -22568 12852
rect -27940 12772 -22568 12788
rect -27940 12708 -22652 12772
rect -22588 12708 -22568 12772
rect -27940 12692 -22568 12708
rect -27940 12628 -22652 12692
rect -22588 12628 -22568 12692
rect -27940 12612 -22568 12628
rect -27940 12548 -22652 12612
rect -22588 12548 -22568 12612
rect -27940 12532 -22568 12548
rect -27940 12468 -22652 12532
rect -22588 12468 -22568 12532
rect -27940 12452 -22568 12468
rect -27940 12388 -22652 12452
rect -22588 12388 -22568 12452
rect -27940 12372 -22568 12388
rect -27940 12308 -22652 12372
rect -22588 12308 -22568 12372
rect -27940 12292 -22568 12308
rect -27940 12228 -22652 12292
rect -22588 12228 -22568 12292
rect -27940 12212 -22568 12228
rect -27940 12148 -22652 12212
rect -22588 12148 -22568 12212
rect -27940 12132 -22568 12148
rect -27940 12068 -22652 12132
rect -22588 12068 -22568 12132
rect -27940 12052 -22568 12068
rect -27940 11988 -22652 12052
rect -22588 11988 -22568 12052
rect -27940 11972 -22568 11988
rect -27940 11908 -22652 11972
rect -22588 11908 -22568 11972
rect -27940 11892 -22568 11908
rect -27940 11828 -22652 11892
rect -22588 11828 -22568 11892
rect -27940 11812 -22568 11828
rect -27940 11748 -22652 11812
rect -22588 11748 -22568 11812
rect -27940 11732 -22568 11748
rect -27940 11668 -22652 11732
rect -22588 11668 -22568 11732
rect -27940 11652 -22568 11668
rect -27940 11588 -22652 11652
rect -22588 11588 -22568 11652
rect -27940 11572 -22568 11588
rect -27940 11508 -22652 11572
rect -22588 11508 -22568 11572
rect -27940 11492 -22568 11508
rect -27940 11428 -22652 11492
rect -22588 11428 -22568 11492
rect -27940 11412 -22568 11428
rect -27940 11348 -22652 11412
rect -22588 11348 -22568 11412
rect -27940 11332 -22568 11348
rect -27940 11268 -22652 11332
rect -22588 11268 -22568 11332
rect -27940 11252 -22568 11268
rect -27940 11188 -22652 11252
rect -22588 11188 -22568 11252
rect -27940 11172 -22568 11188
rect -27940 11108 -22652 11172
rect -22588 11108 -22568 11172
rect -27940 11092 -22568 11108
rect -27940 11028 -22652 11092
rect -22588 11028 -22568 11092
rect -27940 11012 -22568 11028
rect -27940 10948 -22652 11012
rect -22588 10948 -22568 11012
rect -27940 10932 -22568 10948
rect -27940 10868 -22652 10932
rect -22588 10868 -22568 10932
rect -27940 10852 -22568 10868
rect -27940 10788 -22652 10852
rect -22588 10788 -22568 10852
rect -27940 10760 -22568 10788
rect -22328 15812 -16956 15840
rect -22328 15748 -17040 15812
rect -16976 15748 -16956 15812
rect -22328 15732 -16956 15748
rect -22328 15668 -17040 15732
rect -16976 15668 -16956 15732
rect -22328 15652 -16956 15668
rect -22328 15588 -17040 15652
rect -16976 15588 -16956 15652
rect -22328 15572 -16956 15588
rect -22328 15508 -17040 15572
rect -16976 15508 -16956 15572
rect -22328 15492 -16956 15508
rect -22328 15428 -17040 15492
rect -16976 15428 -16956 15492
rect -22328 15412 -16956 15428
rect -22328 15348 -17040 15412
rect -16976 15348 -16956 15412
rect -22328 15332 -16956 15348
rect -22328 15268 -17040 15332
rect -16976 15268 -16956 15332
rect -22328 15252 -16956 15268
rect -22328 15188 -17040 15252
rect -16976 15188 -16956 15252
rect -22328 15172 -16956 15188
rect -22328 15108 -17040 15172
rect -16976 15108 -16956 15172
rect -22328 15092 -16956 15108
rect -22328 15028 -17040 15092
rect -16976 15028 -16956 15092
rect -22328 15012 -16956 15028
rect -22328 14948 -17040 15012
rect -16976 14948 -16956 15012
rect -22328 14932 -16956 14948
rect -22328 14868 -17040 14932
rect -16976 14868 -16956 14932
rect -22328 14852 -16956 14868
rect -22328 14788 -17040 14852
rect -16976 14788 -16956 14852
rect -22328 14772 -16956 14788
rect -22328 14708 -17040 14772
rect -16976 14708 -16956 14772
rect -22328 14692 -16956 14708
rect -22328 14628 -17040 14692
rect -16976 14628 -16956 14692
rect -22328 14612 -16956 14628
rect -22328 14548 -17040 14612
rect -16976 14548 -16956 14612
rect -22328 14532 -16956 14548
rect -22328 14468 -17040 14532
rect -16976 14468 -16956 14532
rect -22328 14452 -16956 14468
rect -22328 14388 -17040 14452
rect -16976 14388 -16956 14452
rect -22328 14372 -16956 14388
rect -22328 14308 -17040 14372
rect -16976 14308 -16956 14372
rect -22328 14292 -16956 14308
rect -22328 14228 -17040 14292
rect -16976 14228 -16956 14292
rect -22328 14212 -16956 14228
rect -22328 14148 -17040 14212
rect -16976 14148 -16956 14212
rect -22328 14132 -16956 14148
rect -22328 14068 -17040 14132
rect -16976 14068 -16956 14132
rect -22328 14052 -16956 14068
rect -22328 13988 -17040 14052
rect -16976 13988 -16956 14052
rect -22328 13972 -16956 13988
rect -22328 13908 -17040 13972
rect -16976 13908 -16956 13972
rect -22328 13892 -16956 13908
rect -22328 13828 -17040 13892
rect -16976 13828 -16956 13892
rect -22328 13812 -16956 13828
rect -22328 13748 -17040 13812
rect -16976 13748 -16956 13812
rect -22328 13732 -16956 13748
rect -22328 13668 -17040 13732
rect -16976 13668 -16956 13732
rect -22328 13652 -16956 13668
rect -22328 13588 -17040 13652
rect -16976 13588 -16956 13652
rect -22328 13572 -16956 13588
rect -22328 13508 -17040 13572
rect -16976 13508 -16956 13572
rect -22328 13492 -16956 13508
rect -22328 13428 -17040 13492
rect -16976 13428 -16956 13492
rect -22328 13412 -16956 13428
rect -22328 13348 -17040 13412
rect -16976 13348 -16956 13412
rect -22328 13332 -16956 13348
rect -22328 13268 -17040 13332
rect -16976 13268 -16956 13332
rect -22328 13252 -16956 13268
rect -22328 13188 -17040 13252
rect -16976 13188 -16956 13252
rect -22328 13172 -16956 13188
rect -22328 13108 -17040 13172
rect -16976 13108 -16956 13172
rect -22328 13092 -16956 13108
rect -22328 13028 -17040 13092
rect -16976 13028 -16956 13092
rect -22328 13012 -16956 13028
rect -22328 12948 -17040 13012
rect -16976 12948 -16956 13012
rect -22328 12932 -16956 12948
rect -22328 12868 -17040 12932
rect -16976 12868 -16956 12932
rect -22328 12852 -16956 12868
rect -22328 12788 -17040 12852
rect -16976 12788 -16956 12852
rect -22328 12772 -16956 12788
rect -22328 12708 -17040 12772
rect -16976 12708 -16956 12772
rect -22328 12692 -16956 12708
rect -22328 12628 -17040 12692
rect -16976 12628 -16956 12692
rect -22328 12612 -16956 12628
rect -22328 12548 -17040 12612
rect -16976 12548 -16956 12612
rect -22328 12532 -16956 12548
rect -22328 12468 -17040 12532
rect -16976 12468 -16956 12532
rect -22328 12452 -16956 12468
rect -22328 12388 -17040 12452
rect -16976 12388 -16956 12452
rect -22328 12372 -16956 12388
rect -22328 12308 -17040 12372
rect -16976 12308 -16956 12372
rect -22328 12292 -16956 12308
rect -22328 12228 -17040 12292
rect -16976 12228 -16956 12292
rect -22328 12212 -16956 12228
rect -22328 12148 -17040 12212
rect -16976 12148 -16956 12212
rect -22328 12132 -16956 12148
rect -22328 12068 -17040 12132
rect -16976 12068 -16956 12132
rect -22328 12052 -16956 12068
rect -22328 11988 -17040 12052
rect -16976 11988 -16956 12052
rect -22328 11972 -16956 11988
rect -22328 11908 -17040 11972
rect -16976 11908 -16956 11972
rect -22328 11892 -16956 11908
rect -22328 11828 -17040 11892
rect -16976 11828 -16956 11892
rect -22328 11812 -16956 11828
rect -22328 11748 -17040 11812
rect -16976 11748 -16956 11812
rect -22328 11732 -16956 11748
rect -22328 11668 -17040 11732
rect -16976 11668 -16956 11732
rect -22328 11652 -16956 11668
rect -22328 11588 -17040 11652
rect -16976 11588 -16956 11652
rect -22328 11572 -16956 11588
rect -22328 11508 -17040 11572
rect -16976 11508 -16956 11572
rect -22328 11492 -16956 11508
rect -22328 11428 -17040 11492
rect -16976 11428 -16956 11492
rect -22328 11412 -16956 11428
rect -22328 11348 -17040 11412
rect -16976 11348 -16956 11412
rect -22328 11332 -16956 11348
rect -22328 11268 -17040 11332
rect -16976 11268 -16956 11332
rect -22328 11252 -16956 11268
rect -22328 11188 -17040 11252
rect -16976 11188 -16956 11252
rect -22328 11172 -16956 11188
rect -22328 11108 -17040 11172
rect -16976 11108 -16956 11172
rect -22328 11092 -16956 11108
rect -22328 11028 -17040 11092
rect -16976 11028 -16956 11092
rect -22328 11012 -16956 11028
rect -22328 10948 -17040 11012
rect -16976 10948 -16956 11012
rect -22328 10932 -16956 10948
rect -22328 10868 -17040 10932
rect -16976 10868 -16956 10932
rect -22328 10852 -16956 10868
rect -22328 10788 -17040 10852
rect -16976 10788 -16956 10852
rect -22328 10760 -16956 10788
rect -16716 15812 -11344 15840
rect -16716 15748 -11428 15812
rect -11364 15748 -11344 15812
rect -16716 15732 -11344 15748
rect -16716 15668 -11428 15732
rect -11364 15668 -11344 15732
rect -16716 15652 -11344 15668
rect -16716 15588 -11428 15652
rect -11364 15588 -11344 15652
rect -16716 15572 -11344 15588
rect -16716 15508 -11428 15572
rect -11364 15508 -11344 15572
rect -16716 15492 -11344 15508
rect -16716 15428 -11428 15492
rect -11364 15428 -11344 15492
rect -16716 15412 -11344 15428
rect -16716 15348 -11428 15412
rect -11364 15348 -11344 15412
rect -16716 15332 -11344 15348
rect -16716 15268 -11428 15332
rect -11364 15268 -11344 15332
rect -16716 15252 -11344 15268
rect -16716 15188 -11428 15252
rect -11364 15188 -11344 15252
rect -16716 15172 -11344 15188
rect -16716 15108 -11428 15172
rect -11364 15108 -11344 15172
rect -16716 15092 -11344 15108
rect -16716 15028 -11428 15092
rect -11364 15028 -11344 15092
rect -16716 15012 -11344 15028
rect -16716 14948 -11428 15012
rect -11364 14948 -11344 15012
rect -16716 14932 -11344 14948
rect -16716 14868 -11428 14932
rect -11364 14868 -11344 14932
rect -16716 14852 -11344 14868
rect -16716 14788 -11428 14852
rect -11364 14788 -11344 14852
rect -16716 14772 -11344 14788
rect -16716 14708 -11428 14772
rect -11364 14708 -11344 14772
rect -16716 14692 -11344 14708
rect -16716 14628 -11428 14692
rect -11364 14628 -11344 14692
rect -16716 14612 -11344 14628
rect -16716 14548 -11428 14612
rect -11364 14548 -11344 14612
rect -16716 14532 -11344 14548
rect -16716 14468 -11428 14532
rect -11364 14468 -11344 14532
rect -16716 14452 -11344 14468
rect -16716 14388 -11428 14452
rect -11364 14388 -11344 14452
rect -16716 14372 -11344 14388
rect -16716 14308 -11428 14372
rect -11364 14308 -11344 14372
rect -16716 14292 -11344 14308
rect -16716 14228 -11428 14292
rect -11364 14228 -11344 14292
rect -16716 14212 -11344 14228
rect -16716 14148 -11428 14212
rect -11364 14148 -11344 14212
rect -16716 14132 -11344 14148
rect -16716 14068 -11428 14132
rect -11364 14068 -11344 14132
rect -16716 14052 -11344 14068
rect -16716 13988 -11428 14052
rect -11364 13988 -11344 14052
rect -16716 13972 -11344 13988
rect -16716 13908 -11428 13972
rect -11364 13908 -11344 13972
rect -16716 13892 -11344 13908
rect -16716 13828 -11428 13892
rect -11364 13828 -11344 13892
rect -16716 13812 -11344 13828
rect -16716 13748 -11428 13812
rect -11364 13748 -11344 13812
rect -16716 13732 -11344 13748
rect -16716 13668 -11428 13732
rect -11364 13668 -11344 13732
rect -16716 13652 -11344 13668
rect -16716 13588 -11428 13652
rect -11364 13588 -11344 13652
rect -16716 13572 -11344 13588
rect -16716 13508 -11428 13572
rect -11364 13508 -11344 13572
rect -16716 13492 -11344 13508
rect -16716 13428 -11428 13492
rect -11364 13428 -11344 13492
rect -16716 13412 -11344 13428
rect -16716 13348 -11428 13412
rect -11364 13348 -11344 13412
rect -16716 13332 -11344 13348
rect -16716 13268 -11428 13332
rect -11364 13268 -11344 13332
rect -16716 13252 -11344 13268
rect -16716 13188 -11428 13252
rect -11364 13188 -11344 13252
rect -16716 13172 -11344 13188
rect -16716 13108 -11428 13172
rect -11364 13108 -11344 13172
rect -16716 13092 -11344 13108
rect -16716 13028 -11428 13092
rect -11364 13028 -11344 13092
rect -16716 13012 -11344 13028
rect -16716 12948 -11428 13012
rect -11364 12948 -11344 13012
rect -16716 12932 -11344 12948
rect -16716 12868 -11428 12932
rect -11364 12868 -11344 12932
rect -16716 12852 -11344 12868
rect -16716 12788 -11428 12852
rect -11364 12788 -11344 12852
rect -16716 12772 -11344 12788
rect -16716 12708 -11428 12772
rect -11364 12708 -11344 12772
rect -16716 12692 -11344 12708
rect -16716 12628 -11428 12692
rect -11364 12628 -11344 12692
rect -16716 12612 -11344 12628
rect -16716 12548 -11428 12612
rect -11364 12548 -11344 12612
rect -16716 12532 -11344 12548
rect -16716 12468 -11428 12532
rect -11364 12468 -11344 12532
rect -16716 12452 -11344 12468
rect -16716 12388 -11428 12452
rect -11364 12388 -11344 12452
rect -16716 12372 -11344 12388
rect -16716 12308 -11428 12372
rect -11364 12308 -11344 12372
rect -16716 12292 -11344 12308
rect -16716 12228 -11428 12292
rect -11364 12228 -11344 12292
rect -16716 12212 -11344 12228
rect -16716 12148 -11428 12212
rect -11364 12148 -11344 12212
rect -16716 12132 -11344 12148
rect -16716 12068 -11428 12132
rect -11364 12068 -11344 12132
rect -16716 12052 -11344 12068
rect -16716 11988 -11428 12052
rect -11364 11988 -11344 12052
rect -16716 11972 -11344 11988
rect -16716 11908 -11428 11972
rect -11364 11908 -11344 11972
rect -16716 11892 -11344 11908
rect -16716 11828 -11428 11892
rect -11364 11828 -11344 11892
rect -16716 11812 -11344 11828
rect -16716 11748 -11428 11812
rect -11364 11748 -11344 11812
rect -16716 11732 -11344 11748
rect -16716 11668 -11428 11732
rect -11364 11668 -11344 11732
rect -16716 11652 -11344 11668
rect -16716 11588 -11428 11652
rect -11364 11588 -11344 11652
rect -16716 11572 -11344 11588
rect -16716 11508 -11428 11572
rect -11364 11508 -11344 11572
rect -16716 11492 -11344 11508
rect -16716 11428 -11428 11492
rect -11364 11428 -11344 11492
rect -16716 11412 -11344 11428
rect -16716 11348 -11428 11412
rect -11364 11348 -11344 11412
rect -16716 11332 -11344 11348
rect -16716 11268 -11428 11332
rect -11364 11268 -11344 11332
rect -16716 11252 -11344 11268
rect -16716 11188 -11428 11252
rect -11364 11188 -11344 11252
rect -16716 11172 -11344 11188
rect -16716 11108 -11428 11172
rect -11364 11108 -11344 11172
rect -16716 11092 -11344 11108
rect -16716 11028 -11428 11092
rect -11364 11028 -11344 11092
rect -16716 11012 -11344 11028
rect -16716 10948 -11428 11012
rect -11364 10948 -11344 11012
rect -16716 10932 -11344 10948
rect -16716 10868 -11428 10932
rect -11364 10868 -11344 10932
rect -16716 10852 -11344 10868
rect -16716 10788 -11428 10852
rect -11364 10788 -11344 10852
rect -16716 10760 -11344 10788
rect -11104 15812 -5732 15840
rect -11104 15748 -5816 15812
rect -5752 15748 -5732 15812
rect -11104 15732 -5732 15748
rect -11104 15668 -5816 15732
rect -5752 15668 -5732 15732
rect -11104 15652 -5732 15668
rect -11104 15588 -5816 15652
rect -5752 15588 -5732 15652
rect -11104 15572 -5732 15588
rect -11104 15508 -5816 15572
rect -5752 15508 -5732 15572
rect -11104 15492 -5732 15508
rect -11104 15428 -5816 15492
rect -5752 15428 -5732 15492
rect -11104 15412 -5732 15428
rect -11104 15348 -5816 15412
rect -5752 15348 -5732 15412
rect -11104 15332 -5732 15348
rect -11104 15268 -5816 15332
rect -5752 15268 -5732 15332
rect -11104 15252 -5732 15268
rect -11104 15188 -5816 15252
rect -5752 15188 -5732 15252
rect -11104 15172 -5732 15188
rect -11104 15108 -5816 15172
rect -5752 15108 -5732 15172
rect -11104 15092 -5732 15108
rect -11104 15028 -5816 15092
rect -5752 15028 -5732 15092
rect -11104 15012 -5732 15028
rect -11104 14948 -5816 15012
rect -5752 14948 -5732 15012
rect -11104 14932 -5732 14948
rect -11104 14868 -5816 14932
rect -5752 14868 -5732 14932
rect -11104 14852 -5732 14868
rect -11104 14788 -5816 14852
rect -5752 14788 -5732 14852
rect -11104 14772 -5732 14788
rect -11104 14708 -5816 14772
rect -5752 14708 -5732 14772
rect -11104 14692 -5732 14708
rect -11104 14628 -5816 14692
rect -5752 14628 -5732 14692
rect -11104 14612 -5732 14628
rect -11104 14548 -5816 14612
rect -5752 14548 -5732 14612
rect -11104 14532 -5732 14548
rect -11104 14468 -5816 14532
rect -5752 14468 -5732 14532
rect -11104 14452 -5732 14468
rect -11104 14388 -5816 14452
rect -5752 14388 -5732 14452
rect -11104 14372 -5732 14388
rect -11104 14308 -5816 14372
rect -5752 14308 -5732 14372
rect -11104 14292 -5732 14308
rect -11104 14228 -5816 14292
rect -5752 14228 -5732 14292
rect -11104 14212 -5732 14228
rect -11104 14148 -5816 14212
rect -5752 14148 -5732 14212
rect -11104 14132 -5732 14148
rect -11104 14068 -5816 14132
rect -5752 14068 -5732 14132
rect -11104 14052 -5732 14068
rect -11104 13988 -5816 14052
rect -5752 13988 -5732 14052
rect -11104 13972 -5732 13988
rect -11104 13908 -5816 13972
rect -5752 13908 -5732 13972
rect -11104 13892 -5732 13908
rect -11104 13828 -5816 13892
rect -5752 13828 -5732 13892
rect -11104 13812 -5732 13828
rect -11104 13748 -5816 13812
rect -5752 13748 -5732 13812
rect -11104 13732 -5732 13748
rect -11104 13668 -5816 13732
rect -5752 13668 -5732 13732
rect -11104 13652 -5732 13668
rect -11104 13588 -5816 13652
rect -5752 13588 -5732 13652
rect -11104 13572 -5732 13588
rect -11104 13508 -5816 13572
rect -5752 13508 -5732 13572
rect -11104 13492 -5732 13508
rect -11104 13428 -5816 13492
rect -5752 13428 -5732 13492
rect -11104 13412 -5732 13428
rect -11104 13348 -5816 13412
rect -5752 13348 -5732 13412
rect -11104 13332 -5732 13348
rect -11104 13268 -5816 13332
rect -5752 13268 -5732 13332
rect -11104 13252 -5732 13268
rect -11104 13188 -5816 13252
rect -5752 13188 -5732 13252
rect -11104 13172 -5732 13188
rect -11104 13108 -5816 13172
rect -5752 13108 -5732 13172
rect -11104 13092 -5732 13108
rect -11104 13028 -5816 13092
rect -5752 13028 -5732 13092
rect -11104 13012 -5732 13028
rect -11104 12948 -5816 13012
rect -5752 12948 -5732 13012
rect -11104 12932 -5732 12948
rect -11104 12868 -5816 12932
rect -5752 12868 -5732 12932
rect -11104 12852 -5732 12868
rect -11104 12788 -5816 12852
rect -5752 12788 -5732 12852
rect -11104 12772 -5732 12788
rect -11104 12708 -5816 12772
rect -5752 12708 -5732 12772
rect -11104 12692 -5732 12708
rect -11104 12628 -5816 12692
rect -5752 12628 -5732 12692
rect -11104 12612 -5732 12628
rect -11104 12548 -5816 12612
rect -5752 12548 -5732 12612
rect -11104 12532 -5732 12548
rect -11104 12468 -5816 12532
rect -5752 12468 -5732 12532
rect -11104 12452 -5732 12468
rect -11104 12388 -5816 12452
rect -5752 12388 -5732 12452
rect -11104 12372 -5732 12388
rect -11104 12308 -5816 12372
rect -5752 12308 -5732 12372
rect -11104 12292 -5732 12308
rect -11104 12228 -5816 12292
rect -5752 12228 -5732 12292
rect -11104 12212 -5732 12228
rect -11104 12148 -5816 12212
rect -5752 12148 -5732 12212
rect -11104 12132 -5732 12148
rect -11104 12068 -5816 12132
rect -5752 12068 -5732 12132
rect -11104 12052 -5732 12068
rect -11104 11988 -5816 12052
rect -5752 11988 -5732 12052
rect -11104 11972 -5732 11988
rect -11104 11908 -5816 11972
rect -5752 11908 -5732 11972
rect -11104 11892 -5732 11908
rect -11104 11828 -5816 11892
rect -5752 11828 -5732 11892
rect -11104 11812 -5732 11828
rect -11104 11748 -5816 11812
rect -5752 11748 -5732 11812
rect -11104 11732 -5732 11748
rect -11104 11668 -5816 11732
rect -5752 11668 -5732 11732
rect -11104 11652 -5732 11668
rect -11104 11588 -5816 11652
rect -5752 11588 -5732 11652
rect -11104 11572 -5732 11588
rect -11104 11508 -5816 11572
rect -5752 11508 -5732 11572
rect -11104 11492 -5732 11508
rect -11104 11428 -5816 11492
rect -5752 11428 -5732 11492
rect -11104 11412 -5732 11428
rect -11104 11348 -5816 11412
rect -5752 11348 -5732 11412
rect -11104 11332 -5732 11348
rect -11104 11268 -5816 11332
rect -5752 11268 -5732 11332
rect -11104 11252 -5732 11268
rect -11104 11188 -5816 11252
rect -5752 11188 -5732 11252
rect -11104 11172 -5732 11188
rect -11104 11108 -5816 11172
rect -5752 11108 -5732 11172
rect -11104 11092 -5732 11108
rect -11104 11028 -5816 11092
rect -5752 11028 -5732 11092
rect -11104 11012 -5732 11028
rect -11104 10948 -5816 11012
rect -5752 10948 -5732 11012
rect -11104 10932 -5732 10948
rect -11104 10868 -5816 10932
rect -5752 10868 -5732 10932
rect -11104 10852 -5732 10868
rect -11104 10788 -5816 10852
rect -5752 10788 -5732 10852
rect -11104 10760 -5732 10788
rect -5492 15812 -120 15840
rect -5492 15748 -204 15812
rect -140 15748 -120 15812
rect -5492 15732 -120 15748
rect -5492 15668 -204 15732
rect -140 15668 -120 15732
rect -5492 15652 -120 15668
rect -5492 15588 -204 15652
rect -140 15588 -120 15652
rect -5492 15572 -120 15588
rect -5492 15508 -204 15572
rect -140 15508 -120 15572
rect -5492 15492 -120 15508
rect -5492 15428 -204 15492
rect -140 15428 -120 15492
rect -5492 15412 -120 15428
rect -5492 15348 -204 15412
rect -140 15348 -120 15412
rect -5492 15332 -120 15348
rect -5492 15268 -204 15332
rect -140 15268 -120 15332
rect -5492 15252 -120 15268
rect -5492 15188 -204 15252
rect -140 15188 -120 15252
rect -5492 15172 -120 15188
rect -5492 15108 -204 15172
rect -140 15108 -120 15172
rect -5492 15092 -120 15108
rect -5492 15028 -204 15092
rect -140 15028 -120 15092
rect -5492 15012 -120 15028
rect -5492 14948 -204 15012
rect -140 14948 -120 15012
rect -5492 14932 -120 14948
rect -5492 14868 -204 14932
rect -140 14868 -120 14932
rect -5492 14852 -120 14868
rect -5492 14788 -204 14852
rect -140 14788 -120 14852
rect -5492 14772 -120 14788
rect -5492 14708 -204 14772
rect -140 14708 -120 14772
rect -5492 14692 -120 14708
rect -5492 14628 -204 14692
rect -140 14628 -120 14692
rect -5492 14612 -120 14628
rect -5492 14548 -204 14612
rect -140 14548 -120 14612
rect -5492 14532 -120 14548
rect -5492 14468 -204 14532
rect -140 14468 -120 14532
rect -5492 14452 -120 14468
rect -5492 14388 -204 14452
rect -140 14388 -120 14452
rect -5492 14372 -120 14388
rect -5492 14308 -204 14372
rect -140 14308 -120 14372
rect -5492 14292 -120 14308
rect -5492 14228 -204 14292
rect -140 14228 -120 14292
rect -5492 14212 -120 14228
rect -5492 14148 -204 14212
rect -140 14148 -120 14212
rect -5492 14132 -120 14148
rect -5492 14068 -204 14132
rect -140 14068 -120 14132
rect -5492 14052 -120 14068
rect -5492 13988 -204 14052
rect -140 13988 -120 14052
rect -5492 13972 -120 13988
rect -5492 13908 -204 13972
rect -140 13908 -120 13972
rect -5492 13892 -120 13908
rect -5492 13828 -204 13892
rect -140 13828 -120 13892
rect -5492 13812 -120 13828
rect -5492 13748 -204 13812
rect -140 13748 -120 13812
rect -5492 13732 -120 13748
rect -5492 13668 -204 13732
rect -140 13668 -120 13732
rect -5492 13652 -120 13668
rect -5492 13588 -204 13652
rect -140 13588 -120 13652
rect -5492 13572 -120 13588
rect -5492 13508 -204 13572
rect -140 13508 -120 13572
rect -5492 13492 -120 13508
rect -5492 13428 -204 13492
rect -140 13428 -120 13492
rect -5492 13412 -120 13428
rect -5492 13348 -204 13412
rect -140 13348 -120 13412
rect -5492 13332 -120 13348
rect -5492 13268 -204 13332
rect -140 13268 -120 13332
rect -5492 13252 -120 13268
rect -5492 13188 -204 13252
rect -140 13188 -120 13252
rect -5492 13172 -120 13188
rect -5492 13108 -204 13172
rect -140 13108 -120 13172
rect -5492 13092 -120 13108
rect -5492 13028 -204 13092
rect -140 13028 -120 13092
rect -5492 13012 -120 13028
rect -5492 12948 -204 13012
rect -140 12948 -120 13012
rect -5492 12932 -120 12948
rect -5492 12868 -204 12932
rect -140 12868 -120 12932
rect -5492 12852 -120 12868
rect -5492 12788 -204 12852
rect -140 12788 -120 12852
rect -5492 12772 -120 12788
rect -5492 12708 -204 12772
rect -140 12708 -120 12772
rect -5492 12692 -120 12708
rect -5492 12628 -204 12692
rect -140 12628 -120 12692
rect -5492 12612 -120 12628
rect -5492 12548 -204 12612
rect -140 12548 -120 12612
rect -5492 12532 -120 12548
rect -5492 12468 -204 12532
rect -140 12468 -120 12532
rect -5492 12452 -120 12468
rect -5492 12388 -204 12452
rect -140 12388 -120 12452
rect -5492 12372 -120 12388
rect -5492 12308 -204 12372
rect -140 12308 -120 12372
rect -5492 12292 -120 12308
rect -5492 12228 -204 12292
rect -140 12228 -120 12292
rect -5492 12212 -120 12228
rect -5492 12148 -204 12212
rect -140 12148 -120 12212
rect -5492 12132 -120 12148
rect -5492 12068 -204 12132
rect -140 12068 -120 12132
rect -5492 12052 -120 12068
rect -5492 11988 -204 12052
rect -140 11988 -120 12052
rect -5492 11972 -120 11988
rect -5492 11908 -204 11972
rect -140 11908 -120 11972
rect -5492 11892 -120 11908
rect -5492 11828 -204 11892
rect -140 11828 -120 11892
rect -5492 11812 -120 11828
rect -5492 11748 -204 11812
rect -140 11748 -120 11812
rect -5492 11732 -120 11748
rect -5492 11668 -204 11732
rect -140 11668 -120 11732
rect -5492 11652 -120 11668
rect -5492 11588 -204 11652
rect -140 11588 -120 11652
rect -5492 11572 -120 11588
rect -5492 11508 -204 11572
rect -140 11508 -120 11572
rect -5492 11492 -120 11508
rect -5492 11428 -204 11492
rect -140 11428 -120 11492
rect -5492 11412 -120 11428
rect -5492 11348 -204 11412
rect -140 11348 -120 11412
rect -5492 11332 -120 11348
rect -5492 11268 -204 11332
rect -140 11268 -120 11332
rect -5492 11252 -120 11268
rect -5492 11188 -204 11252
rect -140 11188 -120 11252
rect -5492 11172 -120 11188
rect -5492 11108 -204 11172
rect -140 11108 -120 11172
rect -5492 11092 -120 11108
rect -5492 11028 -204 11092
rect -140 11028 -120 11092
rect -5492 11012 -120 11028
rect -5492 10948 -204 11012
rect -140 10948 -120 11012
rect -5492 10932 -120 10948
rect -5492 10868 -204 10932
rect -140 10868 -120 10932
rect -5492 10852 -120 10868
rect -5492 10788 -204 10852
rect -140 10788 -120 10852
rect -5492 10760 -120 10788
rect 120 15812 5492 15840
rect 120 15748 5408 15812
rect 5472 15748 5492 15812
rect 120 15732 5492 15748
rect 120 15668 5408 15732
rect 5472 15668 5492 15732
rect 120 15652 5492 15668
rect 120 15588 5408 15652
rect 5472 15588 5492 15652
rect 120 15572 5492 15588
rect 120 15508 5408 15572
rect 5472 15508 5492 15572
rect 120 15492 5492 15508
rect 120 15428 5408 15492
rect 5472 15428 5492 15492
rect 120 15412 5492 15428
rect 120 15348 5408 15412
rect 5472 15348 5492 15412
rect 120 15332 5492 15348
rect 120 15268 5408 15332
rect 5472 15268 5492 15332
rect 120 15252 5492 15268
rect 120 15188 5408 15252
rect 5472 15188 5492 15252
rect 120 15172 5492 15188
rect 120 15108 5408 15172
rect 5472 15108 5492 15172
rect 120 15092 5492 15108
rect 120 15028 5408 15092
rect 5472 15028 5492 15092
rect 120 15012 5492 15028
rect 120 14948 5408 15012
rect 5472 14948 5492 15012
rect 120 14932 5492 14948
rect 120 14868 5408 14932
rect 5472 14868 5492 14932
rect 120 14852 5492 14868
rect 120 14788 5408 14852
rect 5472 14788 5492 14852
rect 120 14772 5492 14788
rect 120 14708 5408 14772
rect 5472 14708 5492 14772
rect 120 14692 5492 14708
rect 120 14628 5408 14692
rect 5472 14628 5492 14692
rect 120 14612 5492 14628
rect 120 14548 5408 14612
rect 5472 14548 5492 14612
rect 120 14532 5492 14548
rect 120 14468 5408 14532
rect 5472 14468 5492 14532
rect 120 14452 5492 14468
rect 120 14388 5408 14452
rect 5472 14388 5492 14452
rect 120 14372 5492 14388
rect 120 14308 5408 14372
rect 5472 14308 5492 14372
rect 120 14292 5492 14308
rect 120 14228 5408 14292
rect 5472 14228 5492 14292
rect 120 14212 5492 14228
rect 120 14148 5408 14212
rect 5472 14148 5492 14212
rect 120 14132 5492 14148
rect 120 14068 5408 14132
rect 5472 14068 5492 14132
rect 120 14052 5492 14068
rect 120 13988 5408 14052
rect 5472 13988 5492 14052
rect 120 13972 5492 13988
rect 120 13908 5408 13972
rect 5472 13908 5492 13972
rect 120 13892 5492 13908
rect 120 13828 5408 13892
rect 5472 13828 5492 13892
rect 120 13812 5492 13828
rect 120 13748 5408 13812
rect 5472 13748 5492 13812
rect 120 13732 5492 13748
rect 120 13668 5408 13732
rect 5472 13668 5492 13732
rect 120 13652 5492 13668
rect 120 13588 5408 13652
rect 5472 13588 5492 13652
rect 120 13572 5492 13588
rect 120 13508 5408 13572
rect 5472 13508 5492 13572
rect 120 13492 5492 13508
rect 120 13428 5408 13492
rect 5472 13428 5492 13492
rect 120 13412 5492 13428
rect 120 13348 5408 13412
rect 5472 13348 5492 13412
rect 120 13332 5492 13348
rect 120 13268 5408 13332
rect 5472 13268 5492 13332
rect 120 13252 5492 13268
rect 120 13188 5408 13252
rect 5472 13188 5492 13252
rect 120 13172 5492 13188
rect 120 13108 5408 13172
rect 5472 13108 5492 13172
rect 120 13092 5492 13108
rect 120 13028 5408 13092
rect 5472 13028 5492 13092
rect 120 13012 5492 13028
rect 120 12948 5408 13012
rect 5472 12948 5492 13012
rect 120 12932 5492 12948
rect 120 12868 5408 12932
rect 5472 12868 5492 12932
rect 120 12852 5492 12868
rect 120 12788 5408 12852
rect 5472 12788 5492 12852
rect 120 12772 5492 12788
rect 120 12708 5408 12772
rect 5472 12708 5492 12772
rect 120 12692 5492 12708
rect 120 12628 5408 12692
rect 5472 12628 5492 12692
rect 120 12612 5492 12628
rect 120 12548 5408 12612
rect 5472 12548 5492 12612
rect 120 12532 5492 12548
rect 120 12468 5408 12532
rect 5472 12468 5492 12532
rect 120 12452 5492 12468
rect 120 12388 5408 12452
rect 5472 12388 5492 12452
rect 120 12372 5492 12388
rect 120 12308 5408 12372
rect 5472 12308 5492 12372
rect 120 12292 5492 12308
rect 120 12228 5408 12292
rect 5472 12228 5492 12292
rect 120 12212 5492 12228
rect 120 12148 5408 12212
rect 5472 12148 5492 12212
rect 120 12132 5492 12148
rect 120 12068 5408 12132
rect 5472 12068 5492 12132
rect 120 12052 5492 12068
rect 120 11988 5408 12052
rect 5472 11988 5492 12052
rect 120 11972 5492 11988
rect 120 11908 5408 11972
rect 5472 11908 5492 11972
rect 120 11892 5492 11908
rect 120 11828 5408 11892
rect 5472 11828 5492 11892
rect 120 11812 5492 11828
rect 120 11748 5408 11812
rect 5472 11748 5492 11812
rect 120 11732 5492 11748
rect 120 11668 5408 11732
rect 5472 11668 5492 11732
rect 120 11652 5492 11668
rect 120 11588 5408 11652
rect 5472 11588 5492 11652
rect 120 11572 5492 11588
rect 120 11508 5408 11572
rect 5472 11508 5492 11572
rect 120 11492 5492 11508
rect 120 11428 5408 11492
rect 5472 11428 5492 11492
rect 120 11412 5492 11428
rect 120 11348 5408 11412
rect 5472 11348 5492 11412
rect 120 11332 5492 11348
rect 120 11268 5408 11332
rect 5472 11268 5492 11332
rect 120 11252 5492 11268
rect 120 11188 5408 11252
rect 5472 11188 5492 11252
rect 120 11172 5492 11188
rect 120 11108 5408 11172
rect 5472 11108 5492 11172
rect 120 11092 5492 11108
rect 120 11028 5408 11092
rect 5472 11028 5492 11092
rect 120 11012 5492 11028
rect 120 10948 5408 11012
rect 5472 10948 5492 11012
rect 120 10932 5492 10948
rect 120 10868 5408 10932
rect 5472 10868 5492 10932
rect 120 10852 5492 10868
rect 120 10788 5408 10852
rect 5472 10788 5492 10852
rect 120 10760 5492 10788
rect 5732 15812 11104 15840
rect 5732 15748 11020 15812
rect 11084 15748 11104 15812
rect 5732 15732 11104 15748
rect 5732 15668 11020 15732
rect 11084 15668 11104 15732
rect 5732 15652 11104 15668
rect 5732 15588 11020 15652
rect 11084 15588 11104 15652
rect 5732 15572 11104 15588
rect 5732 15508 11020 15572
rect 11084 15508 11104 15572
rect 5732 15492 11104 15508
rect 5732 15428 11020 15492
rect 11084 15428 11104 15492
rect 5732 15412 11104 15428
rect 5732 15348 11020 15412
rect 11084 15348 11104 15412
rect 5732 15332 11104 15348
rect 5732 15268 11020 15332
rect 11084 15268 11104 15332
rect 5732 15252 11104 15268
rect 5732 15188 11020 15252
rect 11084 15188 11104 15252
rect 5732 15172 11104 15188
rect 5732 15108 11020 15172
rect 11084 15108 11104 15172
rect 5732 15092 11104 15108
rect 5732 15028 11020 15092
rect 11084 15028 11104 15092
rect 5732 15012 11104 15028
rect 5732 14948 11020 15012
rect 11084 14948 11104 15012
rect 5732 14932 11104 14948
rect 5732 14868 11020 14932
rect 11084 14868 11104 14932
rect 5732 14852 11104 14868
rect 5732 14788 11020 14852
rect 11084 14788 11104 14852
rect 5732 14772 11104 14788
rect 5732 14708 11020 14772
rect 11084 14708 11104 14772
rect 5732 14692 11104 14708
rect 5732 14628 11020 14692
rect 11084 14628 11104 14692
rect 5732 14612 11104 14628
rect 5732 14548 11020 14612
rect 11084 14548 11104 14612
rect 5732 14532 11104 14548
rect 5732 14468 11020 14532
rect 11084 14468 11104 14532
rect 5732 14452 11104 14468
rect 5732 14388 11020 14452
rect 11084 14388 11104 14452
rect 5732 14372 11104 14388
rect 5732 14308 11020 14372
rect 11084 14308 11104 14372
rect 5732 14292 11104 14308
rect 5732 14228 11020 14292
rect 11084 14228 11104 14292
rect 5732 14212 11104 14228
rect 5732 14148 11020 14212
rect 11084 14148 11104 14212
rect 5732 14132 11104 14148
rect 5732 14068 11020 14132
rect 11084 14068 11104 14132
rect 5732 14052 11104 14068
rect 5732 13988 11020 14052
rect 11084 13988 11104 14052
rect 5732 13972 11104 13988
rect 5732 13908 11020 13972
rect 11084 13908 11104 13972
rect 5732 13892 11104 13908
rect 5732 13828 11020 13892
rect 11084 13828 11104 13892
rect 5732 13812 11104 13828
rect 5732 13748 11020 13812
rect 11084 13748 11104 13812
rect 5732 13732 11104 13748
rect 5732 13668 11020 13732
rect 11084 13668 11104 13732
rect 5732 13652 11104 13668
rect 5732 13588 11020 13652
rect 11084 13588 11104 13652
rect 5732 13572 11104 13588
rect 5732 13508 11020 13572
rect 11084 13508 11104 13572
rect 5732 13492 11104 13508
rect 5732 13428 11020 13492
rect 11084 13428 11104 13492
rect 5732 13412 11104 13428
rect 5732 13348 11020 13412
rect 11084 13348 11104 13412
rect 5732 13332 11104 13348
rect 5732 13268 11020 13332
rect 11084 13268 11104 13332
rect 5732 13252 11104 13268
rect 5732 13188 11020 13252
rect 11084 13188 11104 13252
rect 5732 13172 11104 13188
rect 5732 13108 11020 13172
rect 11084 13108 11104 13172
rect 5732 13092 11104 13108
rect 5732 13028 11020 13092
rect 11084 13028 11104 13092
rect 5732 13012 11104 13028
rect 5732 12948 11020 13012
rect 11084 12948 11104 13012
rect 5732 12932 11104 12948
rect 5732 12868 11020 12932
rect 11084 12868 11104 12932
rect 5732 12852 11104 12868
rect 5732 12788 11020 12852
rect 11084 12788 11104 12852
rect 5732 12772 11104 12788
rect 5732 12708 11020 12772
rect 11084 12708 11104 12772
rect 5732 12692 11104 12708
rect 5732 12628 11020 12692
rect 11084 12628 11104 12692
rect 5732 12612 11104 12628
rect 5732 12548 11020 12612
rect 11084 12548 11104 12612
rect 5732 12532 11104 12548
rect 5732 12468 11020 12532
rect 11084 12468 11104 12532
rect 5732 12452 11104 12468
rect 5732 12388 11020 12452
rect 11084 12388 11104 12452
rect 5732 12372 11104 12388
rect 5732 12308 11020 12372
rect 11084 12308 11104 12372
rect 5732 12292 11104 12308
rect 5732 12228 11020 12292
rect 11084 12228 11104 12292
rect 5732 12212 11104 12228
rect 5732 12148 11020 12212
rect 11084 12148 11104 12212
rect 5732 12132 11104 12148
rect 5732 12068 11020 12132
rect 11084 12068 11104 12132
rect 5732 12052 11104 12068
rect 5732 11988 11020 12052
rect 11084 11988 11104 12052
rect 5732 11972 11104 11988
rect 5732 11908 11020 11972
rect 11084 11908 11104 11972
rect 5732 11892 11104 11908
rect 5732 11828 11020 11892
rect 11084 11828 11104 11892
rect 5732 11812 11104 11828
rect 5732 11748 11020 11812
rect 11084 11748 11104 11812
rect 5732 11732 11104 11748
rect 5732 11668 11020 11732
rect 11084 11668 11104 11732
rect 5732 11652 11104 11668
rect 5732 11588 11020 11652
rect 11084 11588 11104 11652
rect 5732 11572 11104 11588
rect 5732 11508 11020 11572
rect 11084 11508 11104 11572
rect 5732 11492 11104 11508
rect 5732 11428 11020 11492
rect 11084 11428 11104 11492
rect 5732 11412 11104 11428
rect 5732 11348 11020 11412
rect 11084 11348 11104 11412
rect 5732 11332 11104 11348
rect 5732 11268 11020 11332
rect 11084 11268 11104 11332
rect 5732 11252 11104 11268
rect 5732 11188 11020 11252
rect 11084 11188 11104 11252
rect 5732 11172 11104 11188
rect 5732 11108 11020 11172
rect 11084 11108 11104 11172
rect 5732 11092 11104 11108
rect 5732 11028 11020 11092
rect 11084 11028 11104 11092
rect 5732 11012 11104 11028
rect 5732 10948 11020 11012
rect 11084 10948 11104 11012
rect 5732 10932 11104 10948
rect 5732 10868 11020 10932
rect 11084 10868 11104 10932
rect 5732 10852 11104 10868
rect 5732 10788 11020 10852
rect 11084 10788 11104 10852
rect 5732 10760 11104 10788
rect 11344 15812 16716 15840
rect 11344 15748 16632 15812
rect 16696 15748 16716 15812
rect 11344 15732 16716 15748
rect 11344 15668 16632 15732
rect 16696 15668 16716 15732
rect 11344 15652 16716 15668
rect 11344 15588 16632 15652
rect 16696 15588 16716 15652
rect 11344 15572 16716 15588
rect 11344 15508 16632 15572
rect 16696 15508 16716 15572
rect 11344 15492 16716 15508
rect 11344 15428 16632 15492
rect 16696 15428 16716 15492
rect 11344 15412 16716 15428
rect 11344 15348 16632 15412
rect 16696 15348 16716 15412
rect 11344 15332 16716 15348
rect 11344 15268 16632 15332
rect 16696 15268 16716 15332
rect 11344 15252 16716 15268
rect 11344 15188 16632 15252
rect 16696 15188 16716 15252
rect 11344 15172 16716 15188
rect 11344 15108 16632 15172
rect 16696 15108 16716 15172
rect 11344 15092 16716 15108
rect 11344 15028 16632 15092
rect 16696 15028 16716 15092
rect 11344 15012 16716 15028
rect 11344 14948 16632 15012
rect 16696 14948 16716 15012
rect 11344 14932 16716 14948
rect 11344 14868 16632 14932
rect 16696 14868 16716 14932
rect 11344 14852 16716 14868
rect 11344 14788 16632 14852
rect 16696 14788 16716 14852
rect 11344 14772 16716 14788
rect 11344 14708 16632 14772
rect 16696 14708 16716 14772
rect 11344 14692 16716 14708
rect 11344 14628 16632 14692
rect 16696 14628 16716 14692
rect 11344 14612 16716 14628
rect 11344 14548 16632 14612
rect 16696 14548 16716 14612
rect 11344 14532 16716 14548
rect 11344 14468 16632 14532
rect 16696 14468 16716 14532
rect 11344 14452 16716 14468
rect 11344 14388 16632 14452
rect 16696 14388 16716 14452
rect 11344 14372 16716 14388
rect 11344 14308 16632 14372
rect 16696 14308 16716 14372
rect 11344 14292 16716 14308
rect 11344 14228 16632 14292
rect 16696 14228 16716 14292
rect 11344 14212 16716 14228
rect 11344 14148 16632 14212
rect 16696 14148 16716 14212
rect 11344 14132 16716 14148
rect 11344 14068 16632 14132
rect 16696 14068 16716 14132
rect 11344 14052 16716 14068
rect 11344 13988 16632 14052
rect 16696 13988 16716 14052
rect 11344 13972 16716 13988
rect 11344 13908 16632 13972
rect 16696 13908 16716 13972
rect 11344 13892 16716 13908
rect 11344 13828 16632 13892
rect 16696 13828 16716 13892
rect 11344 13812 16716 13828
rect 11344 13748 16632 13812
rect 16696 13748 16716 13812
rect 11344 13732 16716 13748
rect 11344 13668 16632 13732
rect 16696 13668 16716 13732
rect 11344 13652 16716 13668
rect 11344 13588 16632 13652
rect 16696 13588 16716 13652
rect 11344 13572 16716 13588
rect 11344 13508 16632 13572
rect 16696 13508 16716 13572
rect 11344 13492 16716 13508
rect 11344 13428 16632 13492
rect 16696 13428 16716 13492
rect 11344 13412 16716 13428
rect 11344 13348 16632 13412
rect 16696 13348 16716 13412
rect 11344 13332 16716 13348
rect 11344 13268 16632 13332
rect 16696 13268 16716 13332
rect 11344 13252 16716 13268
rect 11344 13188 16632 13252
rect 16696 13188 16716 13252
rect 11344 13172 16716 13188
rect 11344 13108 16632 13172
rect 16696 13108 16716 13172
rect 11344 13092 16716 13108
rect 11344 13028 16632 13092
rect 16696 13028 16716 13092
rect 11344 13012 16716 13028
rect 11344 12948 16632 13012
rect 16696 12948 16716 13012
rect 11344 12932 16716 12948
rect 11344 12868 16632 12932
rect 16696 12868 16716 12932
rect 11344 12852 16716 12868
rect 11344 12788 16632 12852
rect 16696 12788 16716 12852
rect 11344 12772 16716 12788
rect 11344 12708 16632 12772
rect 16696 12708 16716 12772
rect 11344 12692 16716 12708
rect 11344 12628 16632 12692
rect 16696 12628 16716 12692
rect 11344 12612 16716 12628
rect 11344 12548 16632 12612
rect 16696 12548 16716 12612
rect 11344 12532 16716 12548
rect 11344 12468 16632 12532
rect 16696 12468 16716 12532
rect 11344 12452 16716 12468
rect 11344 12388 16632 12452
rect 16696 12388 16716 12452
rect 11344 12372 16716 12388
rect 11344 12308 16632 12372
rect 16696 12308 16716 12372
rect 11344 12292 16716 12308
rect 11344 12228 16632 12292
rect 16696 12228 16716 12292
rect 11344 12212 16716 12228
rect 11344 12148 16632 12212
rect 16696 12148 16716 12212
rect 11344 12132 16716 12148
rect 11344 12068 16632 12132
rect 16696 12068 16716 12132
rect 11344 12052 16716 12068
rect 11344 11988 16632 12052
rect 16696 11988 16716 12052
rect 11344 11972 16716 11988
rect 11344 11908 16632 11972
rect 16696 11908 16716 11972
rect 11344 11892 16716 11908
rect 11344 11828 16632 11892
rect 16696 11828 16716 11892
rect 11344 11812 16716 11828
rect 11344 11748 16632 11812
rect 16696 11748 16716 11812
rect 11344 11732 16716 11748
rect 11344 11668 16632 11732
rect 16696 11668 16716 11732
rect 11344 11652 16716 11668
rect 11344 11588 16632 11652
rect 16696 11588 16716 11652
rect 11344 11572 16716 11588
rect 11344 11508 16632 11572
rect 16696 11508 16716 11572
rect 11344 11492 16716 11508
rect 11344 11428 16632 11492
rect 16696 11428 16716 11492
rect 11344 11412 16716 11428
rect 11344 11348 16632 11412
rect 16696 11348 16716 11412
rect 11344 11332 16716 11348
rect 11344 11268 16632 11332
rect 16696 11268 16716 11332
rect 11344 11252 16716 11268
rect 11344 11188 16632 11252
rect 16696 11188 16716 11252
rect 11344 11172 16716 11188
rect 11344 11108 16632 11172
rect 16696 11108 16716 11172
rect 11344 11092 16716 11108
rect 11344 11028 16632 11092
rect 16696 11028 16716 11092
rect 11344 11012 16716 11028
rect 11344 10948 16632 11012
rect 16696 10948 16716 11012
rect 11344 10932 16716 10948
rect 11344 10868 16632 10932
rect 16696 10868 16716 10932
rect 11344 10852 16716 10868
rect 11344 10788 16632 10852
rect 16696 10788 16716 10852
rect 11344 10760 16716 10788
rect 16956 15812 22328 15840
rect 16956 15748 22244 15812
rect 22308 15748 22328 15812
rect 16956 15732 22328 15748
rect 16956 15668 22244 15732
rect 22308 15668 22328 15732
rect 16956 15652 22328 15668
rect 16956 15588 22244 15652
rect 22308 15588 22328 15652
rect 16956 15572 22328 15588
rect 16956 15508 22244 15572
rect 22308 15508 22328 15572
rect 16956 15492 22328 15508
rect 16956 15428 22244 15492
rect 22308 15428 22328 15492
rect 16956 15412 22328 15428
rect 16956 15348 22244 15412
rect 22308 15348 22328 15412
rect 16956 15332 22328 15348
rect 16956 15268 22244 15332
rect 22308 15268 22328 15332
rect 16956 15252 22328 15268
rect 16956 15188 22244 15252
rect 22308 15188 22328 15252
rect 16956 15172 22328 15188
rect 16956 15108 22244 15172
rect 22308 15108 22328 15172
rect 16956 15092 22328 15108
rect 16956 15028 22244 15092
rect 22308 15028 22328 15092
rect 16956 15012 22328 15028
rect 16956 14948 22244 15012
rect 22308 14948 22328 15012
rect 16956 14932 22328 14948
rect 16956 14868 22244 14932
rect 22308 14868 22328 14932
rect 16956 14852 22328 14868
rect 16956 14788 22244 14852
rect 22308 14788 22328 14852
rect 16956 14772 22328 14788
rect 16956 14708 22244 14772
rect 22308 14708 22328 14772
rect 16956 14692 22328 14708
rect 16956 14628 22244 14692
rect 22308 14628 22328 14692
rect 16956 14612 22328 14628
rect 16956 14548 22244 14612
rect 22308 14548 22328 14612
rect 16956 14532 22328 14548
rect 16956 14468 22244 14532
rect 22308 14468 22328 14532
rect 16956 14452 22328 14468
rect 16956 14388 22244 14452
rect 22308 14388 22328 14452
rect 16956 14372 22328 14388
rect 16956 14308 22244 14372
rect 22308 14308 22328 14372
rect 16956 14292 22328 14308
rect 16956 14228 22244 14292
rect 22308 14228 22328 14292
rect 16956 14212 22328 14228
rect 16956 14148 22244 14212
rect 22308 14148 22328 14212
rect 16956 14132 22328 14148
rect 16956 14068 22244 14132
rect 22308 14068 22328 14132
rect 16956 14052 22328 14068
rect 16956 13988 22244 14052
rect 22308 13988 22328 14052
rect 16956 13972 22328 13988
rect 16956 13908 22244 13972
rect 22308 13908 22328 13972
rect 16956 13892 22328 13908
rect 16956 13828 22244 13892
rect 22308 13828 22328 13892
rect 16956 13812 22328 13828
rect 16956 13748 22244 13812
rect 22308 13748 22328 13812
rect 16956 13732 22328 13748
rect 16956 13668 22244 13732
rect 22308 13668 22328 13732
rect 16956 13652 22328 13668
rect 16956 13588 22244 13652
rect 22308 13588 22328 13652
rect 16956 13572 22328 13588
rect 16956 13508 22244 13572
rect 22308 13508 22328 13572
rect 16956 13492 22328 13508
rect 16956 13428 22244 13492
rect 22308 13428 22328 13492
rect 16956 13412 22328 13428
rect 16956 13348 22244 13412
rect 22308 13348 22328 13412
rect 16956 13332 22328 13348
rect 16956 13268 22244 13332
rect 22308 13268 22328 13332
rect 16956 13252 22328 13268
rect 16956 13188 22244 13252
rect 22308 13188 22328 13252
rect 16956 13172 22328 13188
rect 16956 13108 22244 13172
rect 22308 13108 22328 13172
rect 16956 13092 22328 13108
rect 16956 13028 22244 13092
rect 22308 13028 22328 13092
rect 16956 13012 22328 13028
rect 16956 12948 22244 13012
rect 22308 12948 22328 13012
rect 16956 12932 22328 12948
rect 16956 12868 22244 12932
rect 22308 12868 22328 12932
rect 16956 12852 22328 12868
rect 16956 12788 22244 12852
rect 22308 12788 22328 12852
rect 16956 12772 22328 12788
rect 16956 12708 22244 12772
rect 22308 12708 22328 12772
rect 16956 12692 22328 12708
rect 16956 12628 22244 12692
rect 22308 12628 22328 12692
rect 16956 12612 22328 12628
rect 16956 12548 22244 12612
rect 22308 12548 22328 12612
rect 16956 12532 22328 12548
rect 16956 12468 22244 12532
rect 22308 12468 22328 12532
rect 16956 12452 22328 12468
rect 16956 12388 22244 12452
rect 22308 12388 22328 12452
rect 16956 12372 22328 12388
rect 16956 12308 22244 12372
rect 22308 12308 22328 12372
rect 16956 12292 22328 12308
rect 16956 12228 22244 12292
rect 22308 12228 22328 12292
rect 16956 12212 22328 12228
rect 16956 12148 22244 12212
rect 22308 12148 22328 12212
rect 16956 12132 22328 12148
rect 16956 12068 22244 12132
rect 22308 12068 22328 12132
rect 16956 12052 22328 12068
rect 16956 11988 22244 12052
rect 22308 11988 22328 12052
rect 16956 11972 22328 11988
rect 16956 11908 22244 11972
rect 22308 11908 22328 11972
rect 16956 11892 22328 11908
rect 16956 11828 22244 11892
rect 22308 11828 22328 11892
rect 16956 11812 22328 11828
rect 16956 11748 22244 11812
rect 22308 11748 22328 11812
rect 16956 11732 22328 11748
rect 16956 11668 22244 11732
rect 22308 11668 22328 11732
rect 16956 11652 22328 11668
rect 16956 11588 22244 11652
rect 22308 11588 22328 11652
rect 16956 11572 22328 11588
rect 16956 11508 22244 11572
rect 22308 11508 22328 11572
rect 16956 11492 22328 11508
rect 16956 11428 22244 11492
rect 22308 11428 22328 11492
rect 16956 11412 22328 11428
rect 16956 11348 22244 11412
rect 22308 11348 22328 11412
rect 16956 11332 22328 11348
rect 16956 11268 22244 11332
rect 22308 11268 22328 11332
rect 16956 11252 22328 11268
rect 16956 11188 22244 11252
rect 22308 11188 22328 11252
rect 16956 11172 22328 11188
rect 16956 11108 22244 11172
rect 22308 11108 22328 11172
rect 16956 11092 22328 11108
rect 16956 11028 22244 11092
rect 22308 11028 22328 11092
rect 16956 11012 22328 11028
rect 16956 10948 22244 11012
rect 22308 10948 22328 11012
rect 16956 10932 22328 10948
rect 16956 10868 22244 10932
rect 22308 10868 22328 10932
rect 16956 10852 22328 10868
rect 16956 10788 22244 10852
rect 22308 10788 22328 10852
rect 16956 10760 22328 10788
rect 22568 15812 27940 15840
rect 22568 15748 27856 15812
rect 27920 15748 27940 15812
rect 22568 15732 27940 15748
rect 22568 15668 27856 15732
rect 27920 15668 27940 15732
rect 22568 15652 27940 15668
rect 22568 15588 27856 15652
rect 27920 15588 27940 15652
rect 22568 15572 27940 15588
rect 22568 15508 27856 15572
rect 27920 15508 27940 15572
rect 22568 15492 27940 15508
rect 22568 15428 27856 15492
rect 27920 15428 27940 15492
rect 22568 15412 27940 15428
rect 22568 15348 27856 15412
rect 27920 15348 27940 15412
rect 22568 15332 27940 15348
rect 22568 15268 27856 15332
rect 27920 15268 27940 15332
rect 22568 15252 27940 15268
rect 22568 15188 27856 15252
rect 27920 15188 27940 15252
rect 22568 15172 27940 15188
rect 22568 15108 27856 15172
rect 27920 15108 27940 15172
rect 22568 15092 27940 15108
rect 22568 15028 27856 15092
rect 27920 15028 27940 15092
rect 22568 15012 27940 15028
rect 22568 14948 27856 15012
rect 27920 14948 27940 15012
rect 22568 14932 27940 14948
rect 22568 14868 27856 14932
rect 27920 14868 27940 14932
rect 22568 14852 27940 14868
rect 22568 14788 27856 14852
rect 27920 14788 27940 14852
rect 22568 14772 27940 14788
rect 22568 14708 27856 14772
rect 27920 14708 27940 14772
rect 22568 14692 27940 14708
rect 22568 14628 27856 14692
rect 27920 14628 27940 14692
rect 22568 14612 27940 14628
rect 22568 14548 27856 14612
rect 27920 14548 27940 14612
rect 22568 14532 27940 14548
rect 22568 14468 27856 14532
rect 27920 14468 27940 14532
rect 22568 14452 27940 14468
rect 22568 14388 27856 14452
rect 27920 14388 27940 14452
rect 22568 14372 27940 14388
rect 22568 14308 27856 14372
rect 27920 14308 27940 14372
rect 22568 14292 27940 14308
rect 22568 14228 27856 14292
rect 27920 14228 27940 14292
rect 22568 14212 27940 14228
rect 22568 14148 27856 14212
rect 27920 14148 27940 14212
rect 22568 14132 27940 14148
rect 22568 14068 27856 14132
rect 27920 14068 27940 14132
rect 22568 14052 27940 14068
rect 22568 13988 27856 14052
rect 27920 13988 27940 14052
rect 22568 13972 27940 13988
rect 22568 13908 27856 13972
rect 27920 13908 27940 13972
rect 22568 13892 27940 13908
rect 22568 13828 27856 13892
rect 27920 13828 27940 13892
rect 22568 13812 27940 13828
rect 22568 13748 27856 13812
rect 27920 13748 27940 13812
rect 22568 13732 27940 13748
rect 22568 13668 27856 13732
rect 27920 13668 27940 13732
rect 22568 13652 27940 13668
rect 22568 13588 27856 13652
rect 27920 13588 27940 13652
rect 22568 13572 27940 13588
rect 22568 13508 27856 13572
rect 27920 13508 27940 13572
rect 22568 13492 27940 13508
rect 22568 13428 27856 13492
rect 27920 13428 27940 13492
rect 22568 13412 27940 13428
rect 22568 13348 27856 13412
rect 27920 13348 27940 13412
rect 22568 13332 27940 13348
rect 22568 13268 27856 13332
rect 27920 13268 27940 13332
rect 22568 13252 27940 13268
rect 22568 13188 27856 13252
rect 27920 13188 27940 13252
rect 22568 13172 27940 13188
rect 22568 13108 27856 13172
rect 27920 13108 27940 13172
rect 22568 13092 27940 13108
rect 22568 13028 27856 13092
rect 27920 13028 27940 13092
rect 22568 13012 27940 13028
rect 22568 12948 27856 13012
rect 27920 12948 27940 13012
rect 22568 12932 27940 12948
rect 22568 12868 27856 12932
rect 27920 12868 27940 12932
rect 22568 12852 27940 12868
rect 22568 12788 27856 12852
rect 27920 12788 27940 12852
rect 22568 12772 27940 12788
rect 22568 12708 27856 12772
rect 27920 12708 27940 12772
rect 22568 12692 27940 12708
rect 22568 12628 27856 12692
rect 27920 12628 27940 12692
rect 22568 12612 27940 12628
rect 22568 12548 27856 12612
rect 27920 12548 27940 12612
rect 22568 12532 27940 12548
rect 22568 12468 27856 12532
rect 27920 12468 27940 12532
rect 22568 12452 27940 12468
rect 22568 12388 27856 12452
rect 27920 12388 27940 12452
rect 22568 12372 27940 12388
rect 22568 12308 27856 12372
rect 27920 12308 27940 12372
rect 22568 12292 27940 12308
rect 22568 12228 27856 12292
rect 27920 12228 27940 12292
rect 22568 12212 27940 12228
rect 22568 12148 27856 12212
rect 27920 12148 27940 12212
rect 22568 12132 27940 12148
rect 22568 12068 27856 12132
rect 27920 12068 27940 12132
rect 22568 12052 27940 12068
rect 22568 11988 27856 12052
rect 27920 11988 27940 12052
rect 22568 11972 27940 11988
rect 22568 11908 27856 11972
rect 27920 11908 27940 11972
rect 22568 11892 27940 11908
rect 22568 11828 27856 11892
rect 27920 11828 27940 11892
rect 22568 11812 27940 11828
rect 22568 11748 27856 11812
rect 27920 11748 27940 11812
rect 22568 11732 27940 11748
rect 22568 11668 27856 11732
rect 27920 11668 27940 11732
rect 22568 11652 27940 11668
rect 22568 11588 27856 11652
rect 27920 11588 27940 11652
rect 22568 11572 27940 11588
rect 22568 11508 27856 11572
rect 27920 11508 27940 11572
rect 22568 11492 27940 11508
rect 22568 11428 27856 11492
rect 27920 11428 27940 11492
rect 22568 11412 27940 11428
rect 22568 11348 27856 11412
rect 27920 11348 27940 11412
rect 22568 11332 27940 11348
rect 22568 11268 27856 11332
rect 27920 11268 27940 11332
rect 22568 11252 27940 11268
rect 22568 11188 27856 11252
rect 27920 11188 27940 11252
rect 22568 11172 27940 11188
rect 22568 11108 27856 11172
rect 27920 11108 27940 11172
rect 22568 11092 27940 11108
rect 22568 11028 27856 11092
rect 27920 11028 27940 11092
rect 22568 11012 27940 11028
rect 22568 10948 27856 11012
rect 27920 10948 27940 11012
rect 22568 10932 27940 10948
rect 22568 10868 27856 10932
rect 27920 10868 27940 10932
rect 22568 10852 27940 10868
rect 22568 10788 27856 10852
rect 27920 10788 27940 10852
rect 22568 10760 27940 10788
rect 28180 15812 33552 15840
rect 28180 15748 33468 15812
rect 33532 15748 33552 15812
rect 28180 15732 33552 15748
rect 28180 15668 33468 15732
rect 33532 15668 33552 15732
rect 28180 15652 33552 15668
rect 28180 15588 33468 15652
rect 33532 15588 33552 15652
rect 28180 15572 33552 15588
rect 28180 15508 33468 15572
rect 33532 15508 33552 15572
rect 28180 15492 33552 15508
rect 28180 15428 33468 15492
rect 33532 15428 33552 15492
rect 28180 15412 33552 15428
rect 28180 15348 33468 15412
rect 33532 15348 33552 15412
rect 28180 15332 33552 15348
rect 28180 15268 33468 15332
rect 33532 15268 33552 15332
rect 28180 15252 33552 15268
rect 28180 15188 33468 15252
rect 33532 15188 33552 15252
rect 28180 15172 33552 15188
rect 28180 15108 33468 15172
rect 33532 15108 33552 15172
rect 28180 15092 33552 15108
rect 28180 15028 33468 15092
rect 33532 15028 33552 15092
rect 28180 15012 33552 15028
rect 28180 14948 33468 15012
rect 33532 14948 33552 15012
rect 28180 14932 33552 14948
rect 28180 14868 33468 14932
rect 33532 14868 33552 14932
rect 28180 14852 33552 14868
rect 28180 14788 33468 14852
rect 33532 14788 33552 14852
rect 28180 14772 33552 14788
rect 28180 14708 33468 14772
rect 33532 14708 33552 14772
rect 28180 14692 33552 14708
rect 28180 14628 33468 14692
rect 33532 14628 33552 14692
rect 28180 14612 33552 14628
rect 28180 14548 33468 14612
rect 33532 14548 33552 14612
rect 28180 14532 33552 14548
rect 28180 14468 33468 14532
rect 33532 14468 33552 14532
rect 28180 14452 33552 14468
rect 28180 14388 33468 14452
rect 33532 14388 33552 14452
rect 28180 14372 33552 14388
rect 28180 14308 33468 14372
rect 33532 14308 33552 14372
rect 28180 14292 33552 14308
rect 28180 14228 33468 14292
rect 33532 14228 33552 14292
rect 28180 14212 33552 14228
rect 28180 14148 33468 14212
rect 33532 14148 33552 14212
rect 28180 14132 33552 14148
rect 28180 14068 33468 14132
rect 33532 14068 33552 14132
rect 28180 14052 33552 14068
rect 28180 13988 33468 14052
rect 33532 13988 33552 14052
rect 28180 13972 33552 13988
rect 28180 13908 33468 13972
rect 33532 13908 33552 13972
rect 28180 13892 33552 13908
rect 28180 13828 33468 13892
rect 33532 13828 33552 13892
rect 28180 13812 33552 13828
rect 28180 13748 33468 13812
rect 33532 13748 33552 13812
rect 28180 13732 33552 13748
rect 28180 13668 33468 13732
rect 33532 13668 33552 13732
rect 28180 13652 33552 13668
rect 28180 13588 33468 13652
rect 33532 13588 33552 13652
rect 28180 13572 33552 13588
rect 28180 13508 33468 13572
rect 33532 13508 33552 13572
rect 28180 13492 33552 13508
rect 28180 13428 33468 13492
rect 33532 13428 33552 13492
rect 28180 13412 33552 13428
rect 28180 13348 33468 13412
rect 33532 13348 33552 13412
rect 28180 13332 33552 13348
rect 28180 13268 33468 13332
rect 33532 13268 33552 13332
rect 28180 13252 33552 13268
rect 28180 13188 33468 13252
rect 33532 13188 33552 13252
rect 28180 13172 33552 13188
rect 28180 13108 33468 13172
rect 33532 13108 33552 13172
rect 28180 13092 33552 13108
rect 28180 13028 33468 13092
rect 33532 13028 33552 13092
rect 28180 13012 33552 13028
rect 28180 12948 33468 13012
rect 33532 12948 33552 13012
rect 28180 12932 33552 12948
rect 28180 12868 33468 12932
rect 33532 12868 33552 12932
rect 28180 12852 33552 12868
rect 28180 12788 33468 12852
rect 33532 12788 33552 12852
rect 28180 12772 33552 12788
rect 28180 12708 33468 12772
rect 33532 12708 33552 12772
rect 28180 12692 33552 12708
rect 28180 12628 33468 12692
rect 33532 12628 33552 12692
rect 28180 12612 33552 12628
rect 28180 12548 33468 12612
rect 33532 12548 33552 12612
rect 28180 12532 33552 12548
rect 28180 12468 33468 12532
rect 33532 12468 33552 12532
rect 28180 12452 33552 12468
rect 28180 12388 33468 12452
rect 33532 12388 33552 12452
rect 28180 12372 33552 12388
rect 28180 12308 33468 12372
rect 33532 12308 33552 12372
rect 28180 12292 33552 12308
rect 28180 12228 33468 12292
rect 33532 12228 33552 12292
rect 28180 12212 33552 12228
rect 28180 12148 33468 12212
rect 33532 12148 33552 12212
rect 28180 12132 33552 12148
rect 28180 12068 33468 12132
rect 33532 12068 33552 12132
rect 28180 12052 33552 12068
rect 28180 11988 33468 12052
rect 33532 11988 33552 12052
rect 28180 11972 33552 11988
rect 28180 11908 33468 11972
rect 33532 11908 33552 11972
rect 28180 11892 33552 11908
rect 28180 11828 33468 11892
rect 33532 11828 33552 11892
rect 28180 11812 33552 11828
rect 28180 11748 33468 11812
rect 33532 11748 33552 11812
rect 28180 11732 33552 11748
rect 28180 11668 33468 11732
rect 33532 11668 33552 11732
rect 28180 11652 33552 11668
rect 28180 11588 33468 11652
rect 33532 11588 33552 11652
rect 28180 11572 33552 11588
rect 28180 11508 33468 11572
rect 33532 11508 33552 11572
rect 28180 11492 33552 11508
rect 28180 11428 33468 11492
rect 33532 11428 33552 11492
rect 28180 11412 33552 11428
rect 28180 11348 33468 11412
rect 33532 11348 33552 11412
rect 28180 11332 33552 11348
rect 28180 11268 33468 11332
rect 33532 11268 33552 11332
rect 28180 11252 33552 11268
rect 28180 11188 33468 11252
rect 33532 11188 33552 11252
rect 28180 11172 33552 11188
rect 28180 11108 33468 11172
rect 33532 11108 33552 11172
rect 28180 11092 33552 11108
rect 28180 11028 33468 11092
rect 33532 11028 33552 11092
rect 28180 11012 33552 11028
rect 28180 10948 33468 11012
rect 33532 10948 33552 11012
rect 28180 10932 33552 10948
rect 28180 10868 33468 10932
rect 33532 10868 33552 10932
rect 28180 10852 33552 10868
rect 28180 10788 33468 10852
rect 33532 10788 33552 10852
rect 28180 10760 33552 10788
rect 33792 15812 39164 15840
rect 33792 15748 39080 15812
rect 39144 15748 39164 15812
rect 33792 15732 39164 15748
rect 33792 15668 39080 15732
rect 39144 15668 39164 15732
rect 33792 15652 39164 15668
rect 33792 15588 39080 15652
rect 39144 15588 39164 15652
rect 33792 15572 39164 15588
rect 33792 15508 39080 15572
rect 39144 15508 39164 15572
rect 33792 15492 39164 15508
rect 33792 15428 39080 15492
rect 39144 15428 39164 15492
rect 33792 15412 39164 15428
rect 33792 15348 39080 15412
rect 39144 15348 39164 15412
rect 33792 15332 39164 15348
rect 33792 15268 39080 15332
rect 39144 15268 39164 15332
rect 33792 15252 39164 15268
rect 33792 15188 39080 15252
rect 39144 15188 39164 15252
rect 33792 15172 39164 15188
rect 33792 15108 39080 15172
rect 39144 15108 39164 15172
rect 33792 15092 39164 15108
rect 33792 15028 39080 15092
rect 39144 15028 39164 15092
rect 33792 15012 39164 15028
rect 33792 14948 39080 15012
rect 39144 14948 39164 15012
rect 33792 14932 39164 14948
rect 33792 14868 39080 14932
rect 39144 14868 39164 14932
rect 33792 14852 39164 14868
rect 33792 14788 39080 14852
rect 39144 14788 39164 14852
rect 33792 14772 39164 14788
rect 33792 14708 39080 14772
rect 39144 14708 39164 14772
rect 33792 14692 39164 14708
rect 33792 14628 39080 14692
rect 39144 14628 39164 14692
rect 33792 14612 39164 14628
rect 33792 14548 39080 14612
rect 39144 14548 39164 14612
rect 33792 14532 39164 14548
rect 33792 14468 39080 14532
rect 39144 14468 39164 14532
rect 33792 14452 39164 14468
rect 33792 14388 39080 14452
rect 39144 14388 39164 14452
rect 33792 14372 39164 14388
rect 33792 14308 39080 14372
rect 39144 14308 39164 14372
rect 33792 14292 39164 14308
rect 33792 14228 39080 14292
rect 39144 14228 39164 14292
rect 33792 14212 39164 14228
rect 33792 14148 39080 14212
rect 39144 14148 39164 14212
rect 33792 14132 39164 14148
rect 33792 14068 39080 14132
rect 39144 14068 39164 14132
rect 33792 14052 39164 14068
rect 33792 13988 39080 14052
rect 39144 13988 39164 14052
rect 33792 13972 39164 13988
rect 33792 13908 39080 13972
rect 39144 13908 39164 13972
rect 33792 13892 39164 13908
rect 33792 13828 39080 13892
rect 39144 13828 39164 13892
rect 33792 13812 39164 13828
rect 33792 13748 39080 13812
rect 39144 13748 39164 13812
rect 33792 13732 39164 13748
rect 33792 13668 39080 13732
rect 39144 13668 39164 13732
rect 33792 13652 39164 13668
rect 33792 13588 39080 13652
rect 39144 13588 39164 13652
rect 33792 13572 39164 13588
rect 33792 13508 39080 13572
rect 39144 13508 39164 13572
rect 33792 13492 39164 13508
rect 33792 13428 39080 13492
rect 39144 13428 39164 13492
rect 33792 13412 39164 13428
rect 33792 13348 39080 13412
rect 39144 13348 39164 13412
rect 33792 13332 39164 13348
rect 33792 13268 39080 13332
rect 39144 13268 39164 13332
rect 33792 13252 39164 13268
rect 33792 13188 39080 13252
rect 39144 13188 39164 13252
rect 33792 13172 39164 13188
rect 33792 13108 39080 13172
rect 39144 13108 39164 13172
rect 33792 13092 39164 13108
rect 33792 13028 39080 13092
rect 39144 13028 39164 13092
rect 33792 13012 39164 13028
rect 33792 12948 39080 13012
rect 39144 12948 39164 13012
rect 33792 12932 39164 12948
rect 33792 12868 39080 12932
rect 39144 12868 39164 12932
rect 33792 12852 39164 12868
rect 33792 12788 39080 12852
rect 39144 12788 39164 12852
rect 33792 12772 39164 12788
rect 33792 12708 39080 12772
rect 39144 12708 39164 12772
rect 33792 12692 39164 12708
rect 33792 12628 39080 12692
rect 39144 12628 39164 12692
rect 33792 12612 39164 12628
rect 33792 12548 39080 12612
rect 39144 12548 39164 12612
rect 33792 12532 39164 12548
rect 33792 12468 39080 12532
rect 39144 12468 39164 12532
rect 33792 12452 39164 12468
rect 33792 12388 39080 12452
rect 39144 12388 39164 12452
rect 33792 12372 39164 12388
rect 33792 12308 39080 12372
rect 39144 12308 39164 12372
rect 33792 12292 39164 12308
rect 33792 12228 39080 12292
rect 39144 12228 39164 12292
rect 33792 12212 39164 12228
rect 33792 12148 39080 12212
rect 39144 12148 39164 12212
rect 33792 12132 39164 12148
rect 33792 12068 39080 12132
rect 39144 12068 39164 12132
rect 33792 12052 39164 12068
rect 33792 11988 39080 12052
rect 39144 11988 39164 12052
rect 33792 11972 39164 11988
rect 33792 11908 39080 11972
rect 39144 11908 39164 11972
rect 33792 11892 39164 11908
rect 33792 11828 39080 11892
rect 39144 11828 39164 11892
rect 33792 11812 39164 11828
rect 33792 11748 39080 11812
rect 39144 11748 39164 11812
rect 33792 11732 39164 11748
rect 33792 11668 39080 11732
rect 39144 11668 39164 11732
rect 33792 11652 39164 11668
rect 33792 11588 39080 11652
rect 39144 11588 39164 11652
rect 33792 11572 39164 11588
rect 33792 11508 39080 11572
rect 39144 11508 39164 11572
rect 33792 11492 39164 11508
rect 33792 11428 39080 11492
rect 39144 11428 39164 11492
rect 33792 11412 39164 11428
rect 33792 11348 39080 11412
rect 39144 11348 39164 11412
rect 33792 11332 39164 11348
rect 33792 11268 39080 11332
rect 39144 11268 39164 11332
rect 33792 11252 39164 11268
rect 33792 11188 39080 11252
rect 39144 11188 39164 11252
rect 33792 11172 39164 11188
rect 33792 11108 39080 11172
rect 39144 11108 39164 11172
rect 33792 11092 39164 11108
rect 33792 11028 39080 11092
rect 39144 11028 39164 11092
rect 33792 11012 39164 11028
rect 33792 10948 39080 11012
rect 39144 10948 39164 11012
rect 33792 10932 39164 10948
rect 33792 10868 39080 10932
rect 39144 10868 39164 10932
rect 33792 10852 39164 10868
rect 33792 10788 39080 10852
rect 39144 10788 39164 10852
rect 33792 10760 39164 10788
rect -39164 10492 -33792 10520
rect -39164 10428 -33876 10492
rect -33812 10428 -33792 10492
rect -39164 10412 -33792 10428
rect -39164 10348 -33876 10412
rect -33812 10348 -33792 10412
rect -39164 10332 -33792 10348
rect -39164 10268 -33876 10332
rect -33812 10268 -33792 10332
rect -39164 10252 -33792 10268
rect -39164 10188 -33876 10252
rect -33812 10188 -33792 10252
rect -39164 10172 -33792 10188
rect -39164 10108 -33876 10172
rect -33812 10108 -33792 10172
rect -39164 10092 -33792 10108
rect -39164 10028 -33876 10092
rect -33812 10028 -33792 10092
rect -39164 10012 -33792 10028
rect -39164 9948 -33876 10012
rect -33812 9948 -33792 10012
rect -39164 9932 -33792 9948
rect -39164 9868 -33876 9932
rect -33812 9868 -33792 9932
rect -39164 9852 -33792 9868
rect -39164 9788 -33876 9852
rect -33812 9788 -33792 9852
rect -39164 9772 -33792 9788
rect -39164 9708 -33876 9772
rect -33812 9708 -33792 9772
rect -39164 9692 -33792 9708
rect -39164 9628 -33876 9692
rect -33812 9628 -33792 9692
rect -39164 9612 -33792 9628
rect -39164 9548 -33876 9612
rect -33812 9548 -33792 9612
rect -39164 9532 -33792 9548
rect -39164 9468 -33876 9532
rect -33812 9468 -33792 9532
rect -39164 9452 -33792 9468
rect -39164 9388 -33876 9452
rect -33812 9388 -33792 9452
rect -39164 9372 -33792 9388
rect -39164 9308 -33876 9372
rect -33812 9308 -33792 9372
rect -39164 9292 -33792 9308
rect -39164 9228 -33876 9292
rect -33812 9228 -33792 9292
rect -39164 9212 -33792 9228
rect -39164 9148 -33876 9212
rect -33812 9148 -33792 9212
rect -39164 9132 -33792 9148
rect -39164 9068 -33876 9132
rect -33812 9068 -33792 9132
rect -39164 9052 -33792 9068
rect -39164 8988 -33876 9052
rect -33812 8988 -33792 9052
rect -39164 8972 -33792 8988
rect -39164 8908 -33876 8972
rect -33812 8908 -33792 8972
rect -39164 8892 -33792 8908
rect -39164 8828 -33876 8892
rect -33812 8828 -33792 8892
rect -39164 8812 -33792 8828
rect -39164 8748 -33876 8812
rect -33812 8748 -33792 8812
rect -39164 8732 -33792 8748
rect -39164 8668 -33876 8732
rect -33812 8668 -33792 8732
rect -39164 8652 -33792 8668
rect -39164 8588 -33876 8652
rect -33812 8588 -33792 8652
rect -39164 8572 -33792 8588
rect -39164 8508 -33876 8572
rect -33812 8508 -33792 8572
rect -39164 8492 -33792 8508
rect -39164 8428 -33876 8492
rect -33812 8428 -33792 8492
rect -39164 8412 -33792 8428
rect -39164 8348 -33876 8412
rect -33812 8348 -33792 8412
rect -39164 8332 -33792 8348
rect -39164 8268 -33876 8332
rect -33812 8268 -33792 8332
rect -39164 8252 -33792 8268
rect -39164 8188 -33876 8252
rect -33812 8188 -33792 8252
rect -39164 8172 -33792 8188
rect -39164 8108 -33876 8172
rect -33812 8108 -33792 8172
rect -39164 8092 -33792 8108
rect -39164 8028 -33876 8092
rect -33812 8028 -33792 8092
rect -39164 8012 -33792 8028
rect -39164 7948 -33876 8012
rect -33812 7948 -33792 8012
rect -39164 7932 -33792 7948
rect -39164 7868 -33876 7932
rect -33812 7868 -33792 7932
rect -39164 7852 -33792 7868
rect -39164 7788 -33876 7852
rect -33812 7788 -33792 7852
rect -39164 7772 -33792 7788
rect -39164 7708 -33876 7772
rect -33812 7708 -33792 7772
rect -39164 7692 -33792 7708
rect -39164 7628 -33876 7692
rect -33812 7628 -33792 7692
rect -39164 7612 -33792 7628
rect -39164 7548 -33876 7612
rect -33812 7548 -33792 7612
rect -39164 7532 -33792 7548
rect -39164 7468 -33876 7532
rect -33812 7468 -33792 7532
rect -39164 7452 -33792 7468
rect -39164 7388 -33876 7452
rect -33812 7388 -33792 7452
rect -39164 7372 -33792 7388
rect -39164 7308 -33876 7372
rect -33812 7308 -33792 7372
rect -39164 7292 -33792 7308
rect -39164 7228 -33876 7292
rect -33812 7228 -33792 7292
rect -39164 7212 -33792 7228
rect -39164 7148 -33876 7212
rect -33812 7148 -33792 7212
rect -39164 7132 -33792 7148
rect -39164 7068 -33876 7132
rect -33812 7068 -33792 7132
rect -39164 7052 -33792 7068
rect -39164 6988 -33876 7052
rect -33812 6988 -33792 7052
rect -39164 6972 -33792 6988
rect -39164 6908 -33876 6972
rect -33812 6908 -33792 6972
rect -39164 6892 -33792 6908
rect -39164 6828 -33876 6892
rect -33812 6828 -33792 6892
rect -39164 6812 -33792 6828
rect -39164 6748 -33876 6812
rect -33812 6748 -33792 6812
rect -39164 6732 -33792 6748
rect -39164 6668 -33876 6732
rect -33812 6668 -33792 6732
rect -39164 6652 -33792 6668
rect -39164 6588 -33876 6652
rect -33812 6588 -33792 6652
rect -39164 6572 -33792 6588
rect -39164 6508 -33876 6572
rect -33812 6508 -33792 6572
rect -39164 6492 -33792 6508
rect -39164 6428 -33876 6492
rect -33812 6428 -33792 6492
rect -39164 6412 -33792 6428
rect -39164 6348 -33876 6412
rect -33812 6348 -33792 6412
rect -39164 6332 -33792 6348
rect -39164 6268 -33876 6332
rect -33812 6268 -33792 6332
rect -39164 6252 -33792 6268
rect -39164 6188 -33876 6252
rect -33812 6188 -33792 6252
rect -39164 6172 -33792 6188
rect -39164 6108 -33876 6172
rect -33812 6108 -33792 6172
rect -39164 6092 -33792 6108
rect -39164 6028 -33876 6092
rect -33812 6028 -33792 6092
rect -39164 6012 -33792 6028
rect -39164 5948 -33876 6012
rect -33812 5948 -33792 6012
rect -39164 5932 -33792 5948
rect -39164 5868 -33876 5932
rect -33812 5868 -33792 5932
rect -39164 5852 -33792 5868
rect -39164 5788 -33876 5852
rect -33812 5788 -33792 5852
rect -39164 5772 -33792 5788
rect -39164 5708 -33876 5772
rect -33812 5708 -33792 5772
rect -39164 5692 -33792 5708
rect -39164 5628 -33876 5692
rect -33812 5628 -33792 5692
rect -39164 5612 -33792 5628
rect -39164 5548 -33876 5612
rect -33812 5548 -33792 5612
rect -39164 5532 -33792 5548
rect -39164 5468 -33876 5532
rect -33812 5468 -33792 5532
rect -39164 5440 -33792 5468
rect -33552 10492 -28180 10520
rect -33552 10428 -28264 10492
rect -28200 10428 -28180 10492
rect -33552 10412 -28180 10428
rect -33552 10348 -28264 10412
rect -28200 10348 -28180 10412
rect -33552 10332 -28180 10348
rect -33552 10268 -28264 10332
rect -28200 10268 -28180 10332
rect -33552 10252 -28180 10268
rect -33552 10188 -28264 10252
rect -28200 10188 -28180 10252
rect -33552 10172 -28180 10188
rect -33552 10108 -28264 10172
rect -28200 10108 -28180 10172
rect -33552 10092 -28180 10108
rect -33552 10028 -28264 10092
rect -28200 10028 -28180 10092
rect -33552 10012 -28180 10028
rect -33552 9948 -28264 10012
rect -28200 9948 -28180 10012
rect -33552 9932 -28180 9948
rect -33552 9868 -28264 9932
rect -28200 9868 -28180 9932
rect -33552 9852 -28180 9868
rect -33552 9788 -28264 9852
rect -28200 9788 -28180 9852
rect -33552 9772 -28180 9788
rect -33552 9708 -28264 9772
rect -28200 9708 -28180 9772
rect -33552 9692 -28180 9708
rect -33552 9628 -28264 9692
rect -28200 9628 -28180 9692
rect -33552 9612 -28180 9628
rect -33552 9548 -28264 9612
rect -28200 9548 -28180 9612
rect -33552 9532 -28180 9548
rect -33552 9468 -28264 9532
rect -28200 9468 -28180 9532
rect -33552 9452 -28180 9468
rect -33552 9388 -28264 9452
rect -28200 9388 -28180 9452
rect -33552 9372 -28180 9388
rect -33552 9308 -28264 9372
rect -28200 9308 -28180 9372
rect -33552 9292 -28180 9308
rect -33552 9228 -28264 9292
rect -28200 9228 -28180 9292
rect -33552 9212 -28180 9228
rect -33552 9148 -28264 9212
rect -28200 9148 -28180 9212
rect -33552 9132 -28180 9148
rect -33552 9068 -28264 9132
rect -28200 9068 -28180 9132
rect -33552 9052 -28180 9068
rect -33552 8988 -28264 9052
rect -28200 8988 -28180 9052
rect -33552 8972 -28180 8988
rect -33552 8908 -28264 8972
rect -28200 8908 -28180 8972
rect -33552 8892 -28180 8908
rect -33552 8828 -28264 8892
rect -28200 8828 -28180 8892
rect -33552 8812 -28180 8828
rect -33552 8748 -28264 8812
rect -28200 8748 -28180 8812
rect -33552 8732 -28180 8748
rect -33552 8668 -28264 8732
rect -28200 8668 -28180 8732
rect -33552 8652 -28180 8668
rect -33552 8588 -28264 8652
rect -28200 8588 -28180 8652
rect -33552 8572 -28180 8588
rect -33552 8508 -28264 8572
rect -28200 8508 -28180 8572
rect -33552 8492 -28180 8508
rect -33552 8428 -28264 8492
rect -28200 8428 -28180 8492
rect -33552 8412 -28180 8428
rect -33552 8348 -28264 8412
rect -28200 8348 -28180 8412
rect -33552 8332 -28180 8348
rect -33552 8268 -28264 8332
rect -28200 8268 -28180 8332
rect -33552 8252 -28180 8268
rect -33552 8188 -28264 8252
rect -28200 8188 -28180 8252
rect -33552 8172 -28180 8188
rect -33552 8108 -28264 8172
rect -28200 8108 -28180 8172
rect -33552 8092 -28180 8108
rect -33552 8028 -28264 8092
rect -28200 8028 -28180 8092
rect -33552 8012 -28180 8028
rect -33552 7948 -28264 8012
rect -28200 7948 -28180 8012
rect -33552 7932 -28180 7948
rect -33552 7868 -28264 7932
rect -28200 7868 -28180 7932
rect -33552 7852 -28180 7868
rect -33552 7788 -28264 7852
rect -28200 7788 -28180 7852
rect -33552 7772 -28180 7788
rect -33552 7708 -28264 7772
rect -28200 7708 -28180 7772
rect -33552 7692 -28180 7708
rect -33552 7628 -28264 7692
rect -28200 7628 -28180 7692
rect -33552 7612 -28180 7628
rect -33552 7548 -28264 7612
rect -28200 7548 -28180 7612
rect -33552 7532 -28180 7548
rect -33552 7468 -28264 7532
rect -28200 7468 -28180 7532
rect -33552 7452 -28180 7468
rect -33552 7388 -28264 7452
rect -28200 7388 -28180 7452
rect -33552 7372 -28180 7388
rect -33552 7308 -28264 7372
rect -28200 7308 -28180 7372
rect -33552 7292 -28180 7308
rect -33552 7228 -28264 7292
rect -28200 7228 -28180 7292
rect -33552 7212 -28180 7228
rect -33552 7148 -28264 7212
rect -28200 7148 -28180 7212
rect -33552 7132 -28180 7148
rect -33552 7068 -28264 7132
rect -28200 7068 -28180 7132
rect -33552 7052 -28180 7068
rect -33552 6988 -28264 7052
rect -28200 6988 -28180 7052
rect -33552 6972 -28180 6988
rect -33552 6908 -28264 6972
rect -28200 6908 -28180 6972
rect -33552 6892 -28180 6908
rect -33552 6828 -28264 6892
rect -28200 6828 -28180 6892
rect -33552 6812 -28180 6828
rect -33552 6748 -28264 6812
rect -28200 6748 -28180 6812
rect -33552 6732 -28180 6748
rect -33552 6668 -28264 6732
rect -28200 6668 -28180 6732
rect -33552 6652 -28180 6668
rect -33552 6588 -28264 6652
rect -28200 6588 -28180 6652
rect -33552 6572 -28180 6588
rect -33552 6508 -28264 6572
rect -28200 6508 -28180 6572
rect -33552 6492 -28180 6508
rect -33552 6428 -28264 6492
rect -28200 6428 -28180 6492
rect -33552 6412 -28180 6428
rect -33552 6348 -28264 6412
rect -28200 6348 -28180 6412
rect -33552 6332 -28180 6348
rect -33552 6268 -28264 6332
rect -28200 6268 -28180 6332
rect -33552 6252 -28180 6268
rect -33552 6188 -28264 6252
rect -28200 6188 -28180 6252
rect -33552 6172 -28180 6188
rect -33552 6108 -28264 6172
rect -28200 6108 -28180 6172
rect -33552 6092 -28180 6108
rect -33552 6028 -28264 6092
rect -28200 6028 -28180 6092
rect -33552 6012 -28180 6028
rect -33552 5948 -28264 6012
rect -28200 5948 -28180 6012
rect -33552 5932 -28180 5948
rect -33552 5868 -28264 5932
rect -28200 5868 -28180 5932
rect -33552 5852 -28180 5868
rect -33552 5788 -28264 5852
rect -28200 5788 -28180 5852
rect -33552 5772 -28180 5788
rect -33552 5708 -28264 5772
rect -28200 5708 -28180 5772
rect -33552 5692 -28180 5708
rect -33552 5628 -28264 5692
rect -28200 5628 -28180 5692
rect -33552 5612 -28180 5628
rect -33552 5548 -28264 5612
rect -28200 5548 -28180 5612
rect -33552 5532 -28180 5548
rect -33552 5468 -28264 5532
rect -28200 5468 -28180 5532
rect -33552 5440 -28180 5468
rect -27940 10492 -22568 10520
rect -27940 10428 -22652 10492
rect -22588 10428 -22568 10492
rect -27940 10412 -22568 10428
rect -27940 10348 -22652 10412
rect -22588 10348 -22568 10412
rect -27940 10332 -22568 10348
rect -27940 10268 -22652 10332
rect -22588 10268 -22568 10332
rect -27940 10252 -22568 10268
rect -27940 10188 -22652 10252
rect -22588 10188 -22568 10252
rect -27940 10172 -22568 10188
rect -27940 10108 -22652 10172
rect -22588 10108 -22568 10172
rect -27940 10092 -22568 10108
rect -27940 10028 -22652 10092
rect -22588 10028 -22568 10092
rect -27940 10012 -22568 10028
rect -27940 9948 -22652 10012
rect -22588 9948 -22568 10012
rect -27940 9932 -22568 9948
rect -27940 9868 -22652 9932
rect -22588 9868 -22568 9932
rect -27940 9852 -22568 9868
rect -27940 9788 -22652 9852
rect -22588 9788 -22568 9852
rect -27940 9772 -22568 9788
rect -27940 9708 -22652 9772
rect -22588 9708 -22568 9772
rect -27940 9692 -22568 9708
rect -27940 9628 -22652 9692
rect -22588 9628 -22568 9692
rect -27940 9612 -22568 9628
rect -27940 9548 -22652 9612
rect -22588 9548 -22568 9612
rect -27940 9532 -22568 9548
rect -27940 9468 -22652 9532
rect -22588 9468 -22568 9532
rect -27940 9452 -22568 9468
rect -27940 9388 -22652 9452
rect -22588 9388 -22568 9452
rect -27940 9372 -22568 9388
rect -27940 9308 -22652 9372
rect -22588 9308 -22568 9372
rect -27940 9292 -22568 9308
rect -27940 9228 -22652 9292
rect -22588 9228 -22568 9292
rect -27940 9212 -22568 9228
rect -27940 9148 -22652 9212
rect -22588 9148 -22568 9212
rect -27940 9132 -22568 9148
rect -27940 9068 -22652 9132
rect -22588 9068 -22568 9132
rect -27940 9052 -22568 9068
rect -27940 8988 -22652 9052
rect -22588 8988 -22568 9052
rect -27940 8972 -22568 8988
rect -27940 8908 -22652 8972
rect -22588 8908 -22568 8972
rect -27940 8892 -22568 8908
rect -27940 8828 -22652 8892
rect -22588 8828 -22568 8892
rect -27940 8812 -22568 8828
rect -27940 8748 -22652 8812
rect -22588 8748 -22568 8812
rect -27940 8732 -22568 8748
rect -27940 8668 -22652 8732
rect -22588 8668 -22568 8732
rect -27940 8652 -22568 8668
rect -27940 8588 -22652 8652
rect -22588 8588 -22568 8652
rect -27940 8572 -22568 8588
rect -27940 8508 -22652 8572
rect -22588 8508 -22568 8572
rect -27940 8492 -22568 8508
rect -27940 8428 -22652 8492
rect -22588 8428 -22568 8492
rect -27940 8412 -22568 8428
rect -27940 8348 -22652 8412
rect -22588 8348 -22568 8412
rect -27940 8332 -22568 8348
rect -27940 8268 -22652 8332
rect -22588 8268 -22568 8332
rect -27940 8252 -22568 8268
rect -27940 8188 -22652 8252
rect -22588 8188 -22568 8252
rect -27940 8172 -22568 8188
rect -27940 8108 -22652 8172
rect -22588 8108 -22568 8172
rect -27940 8092 -22568 8108
rect -27940 8028 -22652 8092
rect -22588 8028 -22568 8092
rect -27940 8012 -22568 8028
rect -27940 7948 -22652 8012
rect -22588 7948 -22568 8012
rect -27940 7932 -22568 7948
rect -27940 7868 -22652 7932
rect -22588 7868 -22568 7932
rect -27940 7852 -22568 7868
rect -27940 7788 -22652 7852
rect -22588 7788 -22568 7852
rect -27940 7772 -22568 7788
rect -27940 7708 -22652 7772
rect -22588 7708 -22568 7772
rect -27940 7692 -22568 7708
rect -27940 7628 -22652 7692
rect -22588 7628 -22568 7692
rect -27940 7612 -22568 7628
rect -27940 7548 -22652 7612
rect -22588 7548 -22568 7612
rect -27940 7532 -22568 7548
rect -27940 7468 -22652 7532
rect -22588 7468 -22568 7532
rect -27940 7452 -22568 7468
rect -27940 7388 -22652 7452
rect -22588 7388 -22568 7452
rect -27940 7372 -22568 7388
rect -27940 7308 -22652 7372
rect -22588 7308 -22568 7372
rect -27940 7292 -22568 7308
rect -27940 7228 -22652 7292
rect -22588 7228 -22568 7292
rect -27940 7212 -22568 7228
rect -27940 7148 -22652 7212
rect -22588 7148 -22568 7212
rect -27940 7132 -22568 7148
rect -27940 7068 -22652 7132
rect -22588 7068 -22568 7132
rect -27940 7052 -22568 7068
rect -27940 6988 -22652 7052
rect -22588 6988 -22568 7052
rect -27940 6972 -22568 6988
rect -27940 6908 -22652 6972
rect -22588 6908 -22568 6972
rect -27940 6892 -22568 6908
rect -27940 6828 -22652 6892
rect -22588 6828 -22568 6892
rect -27940 6812 -22568 6828
rect -27940 6748 -22652 6812
rect -22588 6748 -22568 6812
rect -27940 6732 -22568 6748
rect -27940 6668 -22652 6732
rect -22588 6668 -22568 6732
rect -27940 6652 -22568 6668
rect -27940 6588 -22652 6652
rect -22588 6588 -22568 6652
rect -27940 6572 -22568 6588
rect -27940 6508 -22652 6572
rect -22588 6508 -22568 6572
rect -27940 6492 -22568 6508
rect -27940 6428 -22652 6492
rect -22588 6428 -22568 6492
rect -27940 6412 -22568 6428
rect -27940 6348 -22652 6412
rect -22588 6348 -22568 6412
rect -27940 6332 -22568 6348
rect -27940 6268 -22652 6332
rect -22588 6268 -22568 6332
rect -27940 6252 -22568 6268
rect -27940 6188 -22652 6252
rect -22588 6188 -22568 6252
rect -27940 6172 -22568 6188
rect -27940 6108 -22652 6172
rect -22588 6108 -22568 6172
rect -27940 6092 -22568 6108
rect -27940 6028 -22652 6092
rect -22588 6028 -22568 6092
rect -27940 6012 -22568 6028
rect -27940 5948 -22652 6012
rect -22588 5948 -22568 6012
rect -27940 5932 -22568 5948
rect -27940 5868 -22652 5932
rect -22588 5868 -22568 5932
rect -27940 5852 -22568 5868
rect -27940 5788 -22652 5852
rect -22588 5788 -22568 5852
rect -27940 5772 -22568 5788
rect -27940 5708 -22652 5772
rect -22588 5708 -22568 5772
rect -27940 5692 -22568 5708
rect -27940 5628 -22652 5692
rect -22588 5628 -22568 5692
rect -27940 5612 -22568 5628
rect -27940 5548 -22652 5612
rect -22588 5548 -22568 5612
rect -27940 5532 -22568 5548
rect -27940 5468 -22652 5532
rect -22588 5468 -22568 5532
rect -27940 5440 -22568 5468
rect -22328 10492 -16956 10520
rect -22328 10428 -17040 10492
rect -16976 10428 -16956 10492
rect -22328 10412 -16956 10428
rect -22328 10348 -17040 10412
rect -16976 10348 -16956 10412
rect -22328 10332 -16956 10348
rect -22328 10268 -17040 10332
rect -16976 10268 -16956 10332
rect -22328 10252 -16956 10268
rect -22328 10188 -17040 10252
rect -16976 10188 -16956 10252
rect -22328 10172 -16956 10188
rect -22328 10108 -17040 10172
rect -16976 10108 -16956 10172
rect -22328 10092 -16956 10108
rect -22328 10028 -17040 10092
rect -16976 10028 -16956 10092
rect -22328 10012 -16956 10028
rect -22328 9948 -17040 10012
rect -16976 9948 -16956 10012
rect -22328 9932 -16956 9948
rect -22328 9868 -17040 9932
rect -16976 9868 -16956 9932
rect -22328 9852 -16956 9868
rect -22328 9788 -17040 9852
rect -16976 9788 -16956 9852
rect -22328 9772 -16956 9788
rect -22328 9708 -17040 9772
rect -16976 9708 -16956 9772
rect -22328 9692 -16956 9708
rect -22328 9628 -17040 9692
rect -16976 9628 -16956 9692
rect -22328 9612 -16956 9628
rect -22328 9548 -17040 9612
rect -16976 9548 -16956 9612
rect -22328 9532 -16956 9548
rect -22328 9468 -17040 9532
rect -16976 9468 -16956 9532
rect -22328 9452 -16956 9468
rect -22328 9388 -17040 9452
rect -16976 9388 -16956 9452
rect -22328 9372 -16956 9388
rect -22328 9308 -17040 9372
rect -16976 9308 -16956 9372
rect -22328 9292 -16956 9308
rect -22328 9228 -17040 9292
rect -16976 9228 -16956 9292
rect -22328 9212 -16956 9228
rect -22328 9148 -17040 9212
rect -16976 9148 -16956 9212
rect -22328 9132 -16956 9148
rect -22328 9068 -17040 9132
rect -16976 9068 -16956 9132
rect -22328 9052 -16956 9068
rect -22328 8988 -17040 9052
rect -16976 8988 -16956 9052
rect -22328 8972 -16956 8988
rect -22328 8908 -17040 8972
rect -16976 8908 -16956 8972
rect -22328 8892 -16956 8908
rect -22328 8828 -17040 8892
rect -16976 8828 -16956 8892
rect -22328 8812 -16956 8828
rect -22328 8748 -17040 8812
rect -16976 8748 -16956 8812
rect -22328 8732 -16956 8748
rect -22328 8668 -17040 8732
rect -16976 8668 -16956 8732
rect -22328 8652 -16956 8668
rect -22328 8588 -17040 8652
rect -16976 8588 -16956 8652
rect -22328 8572 -16956 8588
rect -22328 8508 -17040 8572
rect -16976 8508 -16956 8572
rect -22328 8492 -16956 8508
rect -22328 8428 -17040 8492
rect -16976 8428 -16956 8492
rect -22328 8412 -16956 8428
rect -22328 8348 -17040 8412
rect -16976 8348 -16956 8412
rect -22328 8332 -16956 8348
rect -22328 8268 -17040 8332
rect -16976 8268 -16956 8332
rect -22328 8252 -16956 8268
rect -22328 8188 -17040 8252
rect -16976 8188 -16956 8252
rect -22328 8172 -16956 8188
rect -22328 8108 -17040 8172
rect -16976 8108 -16956 8172
rect -22328 8092 -16956 8108
rect -22328 8028 -17040 8092
rect -16976 8028 -16956 8092
rect -22328 8012 -16956 8028
rect -22328 7948 -17040 8012
rect -16976 7948 -16956 8012
rect -22328 7932 -16956 7948
rect -22328 7868 -17040 7932
rect -16976 7868 -16956 7932
rect -22328 7852 -16956 7868
rect -22328 7788 -17040 7852
rect -16976 7788 -16956 7852
rect -22328 7772 -16956 7788
rect -22328 7708 -17040 7772
rect -16976 7708 -16956 7772
rect -22328 7692 -16956 7708
rect -22328 7628 -17040 7692
rect -16976 7628 -16956 7692
rect -22328 7612 -16956 7628
rect -22328 7548 -17040 7612
rect -16976 7548 -16956 7612
rect -22328 7532 -16956 7548
rect -22328 7468 -17040 7532
rect -16976 7468 -16956 7532
rect -22328 7452 -16956 7468
rect -22328 7388 -17040 7452
rect -16976 7388 -16956 7452
rect -22328 7372 -16956 7388
rect -22328 7308 -17040 7372
rect -16976 7308 -16956 7372
rect -22328 7292 -16956 7308
rect -22328 7228 -17040 7292
rect -16976 7228 -16956 7292
rect -22328 7212 -16956 7228
rect -22328 7148 -17040 7212
rect -16976 7148 -16956 7212
rect -22328 7132 -16956 7148
rect -22328 7068 -17040 7132
rect -16976 7068 -16956 7132
rect -22328 7052 -16956 7068
rect -22328 6988 -17040 7052
rect -16976 6988 -16956 7052
rect -22328 6972 -16956 6988
rect -22328 6908 -17040 6972
rect -16976 6908 -16956 6972
rect -22328 6892 -16956 6908
rect -22328 6828 -17040 6892
rect -16976 6828 -16956 6892
rect -22328 6812 -16956 6828
rect -22328 6748 -17040 6812
rect -16976 6748 -16956 6812
rect -22328 6732 -16956 6748
rect -22328 6668 -17040 6732
rect -16976 6668 -16956 6732
rect -22328 6652 -16956 6668
rect -22328 6588 -17040 6652
rect -16976 6588 -16956 6652
rect -22328 6572 -16956 6588
rect -22328 6508 -17040 6572
rect -16976 6508 -16956 6572
rect -22328 6492 -16956 6508
rect -22328 6428 -17040 6492
rect -16976 6428 -16956 6492
rect -22328 6412 -16956 6428
rect -22328 6348 -17040 6412
rect -16976 6348 -16956 6412
rect -22328 6332 -16956 6348
rect -22328 6268 -17040 6332
rect -16976 6268 -16956 6332
rect -22328 6252 -16956 6268
rect -22328 6188 -17040 6252
rect -16976 6188 -16956 6252
rect -22328 6172 -16956 6188
rect -22328 6108 -17040 6172
rect -16976 6108 -16956 6172
rect -22328 6092 -16956 6108
rect -22328 6028 -17040 6092
rect -16976 6028 -16956 6092
rect -22328 6012 -16956 6028
rect -22328 5948 -17040 6012
rect -16976 5948 -16956 6012
rect -22328 5932 -16956 5948
rect -22328 5868 -17040 5932
rect -16976 5868 -16956 5932
rect -22328 5852 -16956 5868
rect -22328 5788 -17040 5852
rect -16976 5788 -16956 5852
rect -22328 5772 -16956 5788
rect -22328 5708 -17040 5772
rect -16976 5708 -16956 5772
rect -22328 5692 -16956 5708
rect -22328 5628 -17040 5692
rect -16976 5628 -16956 5692
rect -22328 5612 -16956 5628
rect -22328 5548 -17040 5612
rect -16976 5548 -16956 5612
rect -22328 5532 -16956 5548
rect -22328 5468 -17040 5532
rect -16976 5468 -16956 5532
rect -22328 5440 -16956 5468
rect -16716 10492 -11344 10520
rect -16716 10428 -11428 10492
rect -11364 10428 -11344 10492
rect -16716 10412 -11344 10428
rect -16716 10348 -11428 10412
rect -11364 10348 -11344 10412
rect -16716 10332 -11344 10348
rect -16716 10268 -11428 10332
rect -11364 10268 -11344 10332
rect -16716 10252 -11344 10268
rect -16716 10188 -11428 10252
rect -11364 10188 -11344 10252
rect -16716 10172 -11344 10188
rect -16716 10108 -11428 10172
rect -11364 10108 -11344 10172
rect -16716 10092 -11344 10108
rect -16716 10028 -11428 10092
rect -11364 10028 -11344 10092
rect -16716 10012 -11344 10028
rect -16716 9948 -11428 10012
rect -11364 9948 -11344 10012
rect -16716 9932 -11344 9948
rect -16716 9868 -11428 9932
rect -11364 9868 -11344 9932
rect -16716 9852 -11344 9868
rect -16716 9788 -11428 9852
rect -11364 9788 -11344 9852
rect -16716 9772 -11344 9788
rect -16716 9708 -11428 9772
rect -11364 9708 -11344 9772
rect -16716 9692 -11344 9708
rect -16716 9628 -11428 9692
rect -11364 9628 -11344 9692
rect -16716 9612 -11344 9628
rect -16716 9548 -11428 9612
rect -11364 9548 -11344 9612
rect -16716 9532 -11344 9548
rect -16716 9468 -11428 9532
rect -11364 9468 -11344 9532
rect -16716 9452 -11344 9468
rect -16716 9388 -11428 9452
rect -11364 9388 -11344 9452
rect -16716 9372 -11344 9388
rect -16716 9308 -11428 9372
rect -11364 9308 -11344 9372
rect -16716 9292 -11344 9308
rect -16716 9228 -11428 9292
rect -11364 9228 -11344 9292
rect -16716 9212 -11344 9228
rect -16716 9148 -11428 9212
rect -11364 9148 -11344 9212
rect -16716 9132 -11344 9148
rect -16716 9068 -11428 9132
rect -11364 9068 -11344 9132
rect -16716 9052 -11344 9068
rect -16716 8988 -11428 9052
rect -11364 8988 -11344 9052
rect -16716 8972 -11344 8988
rect -16716 8908 -11428 8972
rect -11364 8908 -11344 8972
rect -16716 8892 -11344 8908
rect -16716 8828 -11428 8892
rect -11364 8828 -11344 8892
rect -16716 8812 -11344 8828
rect -16716 8748 -11428 8812
rect -11364 8748 -11344 8812
rect -16716 8732 -11344 8748
rect -16716 8668 -11428 8732
rect -11364 8668 -11344 8732
rect -16716 8652 -11344 8668
rect -16716 8588 -11428 8652
rect -11364 8588 -11344 8652
rect -16716 8572 -11344 8588
rect -16716 8508 -11428 8572
rect -11364 8508 -11344 8572
rect -16716 8492 -11344 8508
rect -16716 8428 -11428 8492
rect -11364 8428 -11344 8492
rect -16716 8412 -11344 8428
rect -16716 8348 -11428 8412
rect -11364 8348 -11344 8412
rect -16716 8332 -11344 8348
rect -16716 8268 -11428 8332
rect -11364 8268 -11344 8332
rect -16716 8252 -11344 8268
rect -16716 8188 -11428 8252
rect -11364 8188 -11344 8252
rect -16716 8172 -11344 8188
rect -16716 8108 -11428 8172
rect -11364 8108 -11344 8172
rect -16716 8092 -11344 8108
rect -16716 8028 -11428 8092
rect -11364 8028 -11344 8092
rect -16716 8012 -11344 8028
rect -16716 7948 -11428 8012
rect -11364 7948 -11344 8012
rect -16716 7932 -11344 7948
rect -16716 7868 -11428 7932
rect -11364 7868 -11344 7932
rect -16716 7852 -11344 7868
rect -16716 7788 -11428 7852
rect -11364 7788 -11344 7852
rect -16716 7772 -11344 7788
rect -16716 7708 -11428 7772
rect -11364 7708 -11344 7772
rect -16716 7692 -11344 7708
rect -16716 7628 -11428 7692
rect -11364 7628 -11344 7692
rect -16716 7612 -11344 7628
rect -16716 7548 -11428 7612
rect -11364 7548 -11344 7612
rect -16716 7532 -11344 7548
rect -16716 7468 -11428 7532
rect -11364 7468 -11344 7532
rect -16716 7452 -11344 7468
rect -16716 7388 -11428 7452
rect -11364 7388 -11344 7452
rect -16716 7372 -11344 7388
rect -16716 7308 -11428 7372
rect -11364 7308 -11344 7372
rect -16716 7292 -11344 7308
rect -16716 7228 -11428 7292
rect -11364 7228 -11344 7292
rect -16716 7212 -11344 7228
rect -16716 7148 -11428 7212
rect -11364 7148 -11344 7212
rect -16716 7132 -11344 7148
rect -16716 7068 -11428 7132
rect -11364 7068 -11344 7132
rect -16716 7052 -11344 7068
rect -16716 6988 -11428 7052
rect -11364 6988 -11344 7052
rect -16716 6972 -11344 6988
rect -16716 6908 -11428 6972
rect -11364 6908 -11344 6972
rect -16716 6892 -11344 6908
rect -16716 6828 -11428 6892
rect -11364 6828 -11344 6892
rect -16716 6812 -11344 6828
rect -16716 6748 -11428 6812
rect -11364 6748 -11344 6812
rect -16716 6732 -11344 6748
rect -16716 6668 -11428 6732
rect -11364 6668 -11344 6732
rect -16716 6652 -11344 6668
rect -16716 6588 -11428 6652
rect -11364 6588 -11344 6652
rect -16716 6572 -11344 6588
rect -16716 6508 -11428 6572
rect -11364 6508 -11344 6572
rect -16716 6492 -11344 6508
rect -16716 6428 -11428 6492
rect -11364 6428 -11344 6492
rect -16716 6412 -11344 6428
rect -16716 6348 -11428 6412
rect -11364 6348 -11344 6412
rect -16716 6332 -11344 6348
rect -16716 6268 -11428 6332
rect -11364 6268 -11344 6332
rect -16716 6252 -11344 6268
rect -16716 6188 -11428 6252
rect -11364 6188 -11344 6252
rect -16716 6172 -11344 6188
rect -16716 6108 -11428 6172
rect -11364 6108 -11344 6172
rect -16716 6092 -11344 6108
rect -16716 6028 -11428 6092
rect -11364 6028 -11344 6092
rect -16716 6012 -11344 6028
rect -16716 5948 -11428 6012
rect -11364 5948 -11344 6012
rect -16716 5932 -11344 5948
rect -16716 5868 -11428 5932
rect -11364 5868 -11344 5932
rect -16716 5852 -11344 5868
rect -16716 5788 -11428 5852
rect -11364 5788 -11344 5852
rect -16716 5772 -11344 5788
rect -16716 5708 -11428 5772
rect -11364 5708 -11344 5772
rect -16716 5692 -11344 5708
rect -16716 5628 -11428 5692
rect -11364 5628 -11344 5692
rect -16716 5612 -11344 5628
rect -16716 5548 -11428 5612
rect -11364 5548 -11344 5612
rect -16716 5532 -11344 5548
rect -16716 5468 -11428 5532
rect -11364 5468 -11344 5532
rect -16716 5440 -11344 5468
rect -11104 10492 -5732 10520
rect -11104 10428 -5816 10492
rect -5752 10428 -5732 10492
rect -11104 10412 -5732 10428
rect -11104 10348 -5816 10412
rect -5752 10348 -5732 10412
rect -11104 10332 -5732 10348
rect -11104 10268 -5816 10332
rect -5752 10268 -5732 10332
rect -11104 10252 -5732 10268
rect -11104 10188 -5816 10252
rect -5752 10188 -5732 10252
rect -11104 10172 -5732 10188
rect -11104 10108 -5816 10172
rect -5752 10108 -5732 10172
rect -11104 10092 -5732 10108
rect -11104 10028 -5816 10092
rect -5752 10028 -5732 10092
rect -11104 10012 -5732 10028
rect -11104 9948 -5816 10012
rect -5752 9948 -5732 10012
rect -11104 9932 -5732 9948
rect -11104 9868 -5816 9932
rect -5752 9868 -5732 9932
rect -11104 9852 -5732 9868
rect -11104 9788 -5816 9852
rect -5752 9788 -5732 9852
rect -11104 9772 -5732 9788
rect -11104 9708 -5816 9772
rect -5752 9708 -5732 9772
rect -11104 9692 -5732 9708
rect -11104 9628 -5816 9692
rect -5752 9628 -5732 9692
rect -11104 9612 -5732 9628
rect -11104 9548 -5816 9612
rect -5752 9548 -5732 9612
rect -11104 9532 -5732 9548
rect -11104 9468 -5816 9532
rect -5752 9468 -5732 9532
rect -11104 9452 -5732 9468
rect -11104 9388 -5816 9452
rect -5752 9388 -5732 9452
rect -11104 9372 -5732 9388
rect -11104 9308 -5816 9372
rect -5752 9308 -5732 9372
rect -11104 9292 -5732 9308
rect -11104 9228 -5816 9292
rect -5752 9228 -5732 9292
rect -11104 9212 -5732 9228
rect -11104 9148 -5816 9212
rect -5752 9148 -5732 9212
rect -11104 9132 -5732 9148
rect -11104 9068 -5816 9132
rect -5752 9068 -5732 9132
rect -11104 9052 -5732 9068
rect -11104 8988 -5816 9052
rect -5752 8988 -5732 9052
rect -11104 8972 -5732 8988
rect -11104 8908 -5816 8972
rect -5752 8908 -5732 8972
rect -11104 8892 -5732 8908
rect -11104 8828 -5816 8892
rect -5752 8828 -5732 8892
rect -11104 8812 -5732 8828
rect -11104 8748 -5816 8812
rect -5752 8748 -5732 8812
rect -11104 8732 -5732 8748
rect -11104 8668 -5816 8732
rect -5752 8668 -5732 8732
rect -11104 8652 -5732 8668
rect -11104 8588 -5816 8652
rect -5752 8588 -5732 8652
rect -11104 8572 -5732 8588
rect -11104 8508 -5816 8572
rect -5752 8508 -5732 8572
rect -11104 8492 -5732 8508
rect -11104 8428 -5816 8492
rect -5752 8428 -5732 8492
rect -11104 8412 -5732 8428
rect -11104 8348 -5816 8412
rect -5752 8348 -5732 8412
rect -11104 8332 -5732 8348
rect -11104 8268 -5816 8332
rect -5752 8268 -5732 8332
rect -11104 8252 -5732 8268
rect -11104 8188 -5816 8252
rect -5752 8188 -5732 8252
rect -11104 8172 -5732 8188
rect -11104 8108 -5816 8172
rect -5752 8108 -5732 8172
rect -11104 8092 -5732 8108
rect -11104 8028 -5816 8092
rect -5752 8028 -5732 8092
rect -11104 8012 -5732 8028
rect -11104 7948 -5816 8012
rect -5752 7948 -5732 8012
rect -11104 7932 -5732 7948
rect -11104 7868 -5816 7932
rect -5752 7868 -5732 7932
rect -11104 7852 -5732 7868
rect -11104 7788 -5816 7852
rect -5752 7788 -5732 7852
rect -11104 7772 -5732 7788
rect -11104 7708 -5816 7772
rect -5752 7708 -5732 7772
rect -11104 7692 -5732 7708
rect -11104 7628 -5816 7692
rect -5752 7628 -5732 7692
rect -11104 7612 -5732 7628
rect -11104 7548 -5816 7612
rect -5752 7548 -5732 7612
rect -11104 7532 -5732 7548
rect -11104 7468 -5816 7532
rect -5752 7468 -5732 7532
rect -11104 7452 -5732 7468
rect -11104 7388 -5816 7452
rect -5752 7388 -5732 7452
rect -11104 7372 -5732 7388
rect -11104 7308 -5816 7372
rect -5752 7308 -5732 7372
rect -11104 7292 -5732 7308
rect -11104 7228 -5816 7292
rect -5752 7228 -5732 7292
rect -11104 7212 -5732 7228
rect -11104 7148 -5816 7212
rect -5752 7148 -5732 7212
rect -11104 7132 -5732 7148
rect -11104 7068 -5816 7132
rect -5752 7068 -5732 7132
rect -11104 7052 -5732 7068
rect -11104 6988 -5816 7052
rect -5752 6988 -5732 7052
rect -11104 6972 -5732 6988
rect -11104 6908 -5816 6972
rect -5752 6908 -5732 6972
rect -11104 6892 -5732 6908
rect -11104 6828 -5816 6892
rect -5752 6828 -5732 6892
rect -11104 6812 -5732 6828
rect -11104 6748 -5816 6812
rect -5752 6748 -5732 6812
rect -11104 6732 -5732 6748
rect -11104 6668 -5816 6732
rect -5752 6668 -5732 6732
rect -11104 6652 -5732 6668
rect -11104 6588 -5816 6652
rect -5752 6588 -5732 6652
rect -11104 6572 -5732 6588
rect -11104 6508 -5816 6572
rect -5752 6508 -5732 6572
rect -11104 6492 -5732 6508
rect -11104 6428 -5816 6492
rect -5752 6428 -5732 6492
rect -11104 6412 -5732 6428
rect -11104 6348 -5816 6412
rect -5752 6348 -5732 6412
rect -11104 6332 -5732 6348
rect -11104 6268 -5816 6332
rect -5752 6268 -5732 6332
rect -11104 6252 -5732 6268
rect -11104 6188 -5816 6252
rect -5752 6188 -5732 6252
rect -11104 6172 -5732 6188
rect -11104 6108 -5816 6172
rect -5752 6108 -5732 6172
rect -11104 6092 -5732 6108
rect -11104 6028 -5816 6092
rect -5752 6028 -5732 6092
rect -11104 6012 -5732 6028
rect -11104 5948 -5816 6012
rect -5752 5948 -5732 6012
rect -11104 5932 -5732 5948
rect -11104 5868 -5816 5932
rect -5752 5868 -5732 5932
rect -11104 5852 -5732 5868
rect -11104 5788 -5816 5852
rect -5752 5788 -5732 5852
rect -11104 5772 -5732 5788
rect -11104 5708 -5816 5772
rect -5752 5708 -5732 5772
rect -11104 5692 -5732 5708
rect -11104 5628 -5816 5692
rect -5752 5628 -5732 5692
rect -11104 5612 -5732 5628
rect -11104 5548 -5816 5612
rect -5752 5548 -5732 5612
rect -11104 5532 -5732 5548
rect -11104 5468 -5816 5532
rect -5752 5468 -5732 5532
rect -11104 5440 -5732 5468
rect -5492 10492 -120 10520
rect -5492 10428 -204 10492
rect -140 10428 -120 10492
rect -5492 10412 -120 10428
rect -5492 10348 -204 10412
rect -140 10348 -120 10412
rect -5492 10332 -120 10348
rect -5492 10268 -204 10332
rect -140 10268 -120 10332
rect -5492 10252 -120 10268
rect -5492 10188 -204 10252
rect -140 10188 -120 10252
rect -5492 10172 -120 10188
rect -5492 10108 -204 10172
rect -140 10108 -120 10172
rect -5492 10092 -120 10108
rect -5492 10028 -204 10092
rect -140 10028 -120 10092
rect -5492 10012 -120 10028
rect -5492 9948 -204 10012
rect -140 9948 -120 10012
rect -5492 9932 -120 9948
rect -5492 9868 -204 9932
rect -140 9868 -120 9932
rect -5492 9852 -120 9868
rect -5492 9788 -204 9852
rect -140 9788 -120 9852
rect -5492 9772 -120 9788
rect -5492 9708 -204 9772
rect -140 9708 -120 9772
rect -5492 9692 -120 9708
rect -5492 9628 -204 9692
rect -140 9628 -120 9692
rect -5492 9612 -120 9628
rect -5492 9548 -204 9612
rect -140 9548 -120 9612
rect -5492 9532 -120 9548
rect -5492 9468 -204 9532
rect -140 9468 -120 9532
rect -5492 9452 -120 9468
rect -5492 9388 -204 9452
rect -140 9388 -120 9452
rect -5492 9372 -120 9388
rect -5492 9308 -204 9372
rect -140 9308 -120 9372
rect -5492 9292 -120 9308
rect -5492 9228 -204 9292
rect -140 9228 -120 9292
rect -5492 9212 -120 9228
rect -5492 9148 -204 9212
rect -140 9148 -120 9212
rect -5492 9132 -120 9148
rect -5492 9068 -204 9132
rect -140 9068 -120 9132
rect -5492 9052 -120 9068
rect -5492 8988 -204 9052
rect -140 8988 -120 9052
rect -5492 8972 -120 8988
rect -5492 8908 -204 8972
rect -140 8908 -120 8972
rect -5492 8892 -120 8908
rect -5492 8828 -204 8892
rect -140 8828 -120 8892
rect -5492 8812 -120 8828
rect -5492 8748 -204 8812
rect -140 8748 -120 8812
rect -5492 8732 -120 8748
rect -5492 8668 -204 8732
rect -140 8668 -120 8732
rect -5492 8652 -120 8668
rect -5492 8588 -204 8652
rect -140 8588 -120 8652
rect -5492 8572 -120 8588
rect -5492 8508 -204 8572
rect -140 8508 -120 8572
rect -5492 8492 -120 8508
rect -5492 8428 -204 8492
rect -140 8428 -120 8492
rect -5492 8412 -120 8428
rect -5492 8348 -204 8412
rect -140 8348 -120 8412
rect -5492 8332 -120 8348
rect -5492 8268 -204 8332
rect -140 8268 -120 8332
rect -5492 8252 -120 8268
rect -5492 8188 -204 8252
rect -140 8188 -120 8252
rect -5492 8172 -120 8188
rect -5492 8108 -204 8172
rect -140 8108 -120 8172
rect -5492 8092 -120 8108
rect -5492 8028 -204 8092
rect -140 8028 -120 8092
rect -5492 8012 -120 8028
rect -5492 7948 -204 8012
rect -140 7948 -120 8012
rect -5492 7932 -120 7948
rect -5492 7868 -204 7932
rect -140 7868 -120 7932
rect -5492 7852 -120 7868
rect -5492 7788 -204 7852
rect -140 7788 -120 7852
rect -5492 7772 -120 7788
rect -5492 7708 -204 7772
rect -140 7708 -120 7772
rect -5492 7692 -120 7708
rect -5492 7628 -204 7692
rect -140 7628 -120 7692
rect -5492 7612 -120 7628
rect -5492 7548 -204 7612
rect -140 7548 -120 7612
rect -5492 7532 -120 7548
rect -5492 7468 -204 7532
rect -140 7468 -120 7532
rect -5492 7452 -120 7468
rect -5492 7388 -204 7452
rect -140 7388 -120 7452
rect -5492 7372 -120 7388
rect -5492 7308 -204 7372
rect -140 7308 -120 7372
rect -5492 7292 -120 7308
rect -5492 7228 -204 7292
rect -140 7228 -120 7292
rect -5492 7212 -120 7228
rect -5492 7148 -204 7212
rect -140 7148 -120 7212
rect -5492 7132 -120 7148
rect -5492 7068 -204 7132
rect -140 7068 -120 7132
rect -5492 7052 -120 7068
rect -5492 6988 -204 7052
rect -140 6988 -120 7052
rect -5492 6972 -120 6988
rect -5492 6908 -204 6972
rect -140 6908 -120 6972
rect -5492 6892 -120 6908
rect -5492 6828 -204 6892
rect -140 6828 -120 6892
rect -5492 6812 -120 6828
rect -5492 6748 -204 6812
rect -140 6748 -120 6812
rect -5492 6732 -120 6748
rect -5492 6668 -204 6732
rect -140 6668 -120 6732
rect -5492 6652 -120 6668
rect -5492 6588 -204 6652
rect -140 6588 -120 6652
rect -5492 6572 -120 6588
rect -5492 6508 -204 6572
rect -140 6508 -120 6572
rect -5492 6492 -120 6508
rect -5492 6428 -204 6492
rect -140 6428 -120 6492
rect -5492 6412 -120 6428
rect -5492 6348 -204 6412
rect -140 6348 -120 6412
rect -5492 6332 -120 6348
rect -5492 6268 -204 6332
rect -140 6268 -120 6332
rect -5492 6252 -120 6268
rect -5492 6188 -204 6252
rect -140 6188 -120 6252
rect -5492 6172 -120 6188
rect -5492 6108 -204 6172
rect -140 6108 -120 6172
rect -5492 6092 -120 6108
rect -5492 6028 -204 6092
rect -140 6028 -120 6092
rect -5492 6012 -120 6028
rect -5492 5948 -204 6012
rect -140 5948 -120 6012
rect -5492 5932 -120 5948
rect -5492 5868 -204 5932
rect -140 5868 -120 5932
rect -5492 5852 -120 5868
rect -5492 5788 -204 5852
rect -140 5788 -120 5852
rect -5492 5772 -120 5788
rect -5492 5708 -204 5772
rect -140 5708 -120 5772
rect -5492 5692 -120 5708
rect -5492 5628 -204 5692
rect -140 5628 -120 5692
rect -5492 5612 -120 5628
rect -5492 5548 -204 5612
rect -140 5548 -120 5612
rect -5492 5532 -120 5548
rect -5492 5468 -204 5532
rect -140 5468 -120 5532
rect -5492 5440 -120 5468
rect 120 10492 5492 10520
rect 120 10428 5408 10492
rect 5472 10428 5492 10492
rect 120 10412 5492 10428
rect 120 10348 5408 10412
rect 5472 10348 5492 10412
rect 120 10332 5492 10348
rect 120 10268 5408 10332
rect 5472 10268 5492 10332
rect 120 10252 5492 10268
rect 120 10188 5408 10252
rect 5472 10188 5492 10252
rect 120 10172 5492 10188
rect 120 10108 5408 10172
rect 5472 10108 5492 10172
rect 120 10092 5492 10108
rect 120 10028 5408 10092
rect 5472 10028 5492 10092
rect 120 10012 5492 10028
rect 120 9948 5408 10012
rect 5472 9948 5492 10012
rect 120 9932 5492 9948
rect 120 9868 5408 9932
rect 5472 9868 5492 9932
rect 120 9852 5492 9868
rect 120 9788 5408 9852
rect 5472 9788 5492 9852
rect 120 9772 5492 9788
rect 120 9708 5408 9772
rect 5472 9708 5492 9772
rect 120 9692 5492 9708
rect 120 9628 5408 9692
rect 5472 9628 5492 9692
rect 120 9612 5492 9628
rect 120 9548 5408 9612
rect 5472 9548 5492 9612
rect 120 9532 5492 9548
rect 120 9468 5408 9532
rect 5472 9468 5492 9532
rect 120 9452 5492 9468
rect 120 9388 5408 9452
rect 5472 9388 5492 9452
rect 120 9372 5492 9388
rect 120 9308 5408 9372
rect 5472 9308 5492 9372
rect 120 9292 5492 9308
rect 120 9228 5408 9292
rect 5472 9228 5492 9292
rect 120 9212 5492 9228
rect 120 9148 5408 9212
rect 5472 9148 5492 9212
rect 120 9132 5492 9148
rect 120 9068 5408 9132
rect 5472 9068 5492 9132
rect 120 9052 5492 9068
rect 120 8988 5408 9052
rect 5472 8988 5492 9052
rect 120 8972 5492 8988
rect 120 8908 5408 8972
rect 5472 8908 5492 8972
rect 120 8892 5492 8908
rect 120 8828 5408 8892
rect 5472 8828 5492 8892
rect 120 8812 5492 8828
rect 120 8748 5408 8812
rect 5472 8748 5492 8812
rect 120 8732 5492 8748
rect 120 8668 5408 8732
rect 5472 8668 5492 8732
rect 120 8652 5492 8668
rect 120 8588 5408 8652
rect 5472 8588 5492 8652
rect 120 8572 5492 8588
rect 120 8508 5408 8572
rect 5472 8508 5492 8572
rect 120 8492 5492 8508
rect 120 8428 5408 8492
rect 5472 8428 5492 8492
rect 120 8412 5492 8428
rect 120 8348 5408 8412
rect 5472 8348 5492 8412
rect 120 8332 5492 8348
rect 120 8268 5408 8332
rect 5472 8268 5492 8332
rect 120 8252 5492 8268
rect 120 8188 5408 8252
rect 5472 8188 5492 8252
rect 120 8172 5492 8188
rect 120 8108 5408 8172
rect 5472 8108 5492 8172
rect 120 8092 5492 8108
rect 120 8028 5408 8092
rect 5472 8028 5492 8092
rect 120 8012 5492 8028
rect 120 7948 5408 8012
rect 5472 7948 5492 8012
rect 120 7932 5492 7948
rect 120 7868 5408 7932
rect 5472 7868 5492 7932
rect 120 7852 5492 7868
rect 120 7788 5408 7852
rect 5472 7788 5492 7852
rect 120 7772 5492 7788
rect 120 7708 5408 7772
rect 5472 7708 5492 7772
rect 120 7692 5492 7708
rect 120 7628 5408 7692
rect 5472 7628 5492 7692
rect 120 7612 5492 7628
rect 120 7548 5408 7612
rect 5472 7548 5492 7612
rect 120 7532 5492 7548
rect 120 7468 5408 7532
rect 5472 7468 5492 7532
rect 120 7452 5492 7468
rect 120 7388 5408 7452
rect 5472 7388 5492 7452
rect 120 7372 5492 7388
rect 120 7308 5408 7372
rect 5472 7308 5492 7372
rect 120 7292 5492 7308
rect 120 7228 5408 7292
rect 5472 7228 5492 7292
rect 120 7212 5492 7228
rect 120 7148 5408 7212
rect 5472 7148 5492 7212
rect 120 7132 5492 7148
rect 120 7068 5408 7132
rect 5472 7068 5492 7132
rect 120 7052 5492 7068
rect 120 6988 5408 7052
rect 5472 6988 5492 7052
rect 120 6972 5492 6988
rect 120 6908 5408 6972
rect 5472 6908 5492 6972
rect 120 6892 5492 6908
rect 120 6828 5408 6892
rect 5472 6828 5492 6892
rect 120 6812 5492 6828
rect 120 6748 5408 6812
rect 5472 6748 5492 6812
rect 120 6732 5492 6748
rect 120 6668 5408 6732
rect 5472 6668 5492 6732
rect 120 6652 5492 6668
rect 120 6588 5408 6652
rect 5472 6588 5492 6652
rect 120 6572 5492 6588
rect 120 6508 5408 6572
rect 5472 6508 5492 6572
rect 120 6492 5492 6508
rect 120 6428 5408 6492
rect 5472 6428 5492 6492
rect 120 6412 5492 6428
rect 120 6348 5408 6412
rect 5472 6348 5492 6412
rect 120 6332 5492 6348
rect 120 6268 5408 6332
rect 5472 6268 5492 6332
rect 120 6252 5492 6268
rect 120 6188 5408 6252
rect 5472 6188 5492 6252
rect 120 6172 5492 6188
rect 120 6108 5408 6172
rect 5472 6108 5492 6172
rect 120 6092 5492 6108
rect 120 6028 5408 6092
rect 5472 6028 5492 6092
rect 120 6012 5492 6028
rect 120 5948 5408 6012
rect 5472 5948 5492 6012
rect 120 5932 5492 5948
rect 120 5868 5408 5932
rect 5472 5868 5492 5932
rect 120 5852 5492 5868
rect 120 5788 5408 5852
rect 5472 5788 5492 5852
rect 120 5772 5492 5788
rect 120 5708 5408 5772
rect 5472 5708 5492 5772
rect 120 5692 5492 5708
rect 120 5628 5408 5692
rect 5472 5628 5492 5692
rect 120 5612 5492 5628
rect 120 5548 5408 5612
rect 5472 5548 5492 5612
rect 120 5532 5492 5548
rect 120 5468 5408 5532
rect 5472 5468 5492 5532
rect 120 5440 5492 5468
rect 5732 10492 11104 10520
rect 5732 10428 11020 10492
rect 11084 10428 11104 10492
rect 5732 10412 11104 10428
rect 5732 10348 11020 10412
rect 11084 10348 11104 10412
rect 5732 10332 11104 10348
rect 5732 10268 11020 10332
rect 11084 10268 11104 10332
rect 5732 10252 11104 10268
rect 5732 10188 11020 10252
rect 11084 10188 11104 10252
rect 5732 10172 11104 10188
rect 5732 10108 11020 10172
rect 11084 10108 11104 10172
rect 5732 10092 11104 10108
rect 5732 10028 11020 10092
rect 11084 10028 11104 10092
rect 5732 10012 11104 10028
rect 5732 9948 11020 10012
rect 11084 9948 11104 10012
rect 5732 9932 11104 9948
rect 5732 9868 11020 9932
rect 11084 9868 11104 9932
rect 5732 9852 11104 9868
rect 5732 9788 11020 9852
rect 11084 9788 11104 9852
rect 5732 9772 11104 9788
rect 5732 9708 11020 9772
rect 11084 9708 11104 9772
rect 5732 9692 11104 9708
rect 5732 9628 11020 9692
rect 11084 9628 11104 9692
rect 5732 9612 11104 9628
rect 5732 9548 11020 9612
rect 11084 9548 11104 9612
rect 5732 9532 11104 9548
rect 5732 9468 11020 9532
rect 11084 9468 11104 9532
rect 5732 9452 11104 9468
rect 5732 9388 11020 9452
rect 11084 9388 11104 9452
rect 5732 9372 11104 9388
rect 5732 9308 11020 9372
rect 11084 9308 11104 9372
rect 5732 9292 11104 9308
rect 5732 9228 11020 9292
rect 11084 9228 11104 9292
rect 5732 9212 11104 9228
rect 5732 9148 11020 9212
rect 11084 9148 11104 9212
rect 5732 9132 11104 9148
rect 5732 9068 11020 9132
rect 11084 9068 11104 9132
rect 5732 9052 11104 9068
rect 5732 8988 11020 9052
rect 11084 8988 11104 9052
rect 5732 8972 11104 8988
rect 5732 8908 11020 8972
rect 11084 8908 11104 8972
rect 5732 8892 11104 8908
rect 5732 8828 11020 8892
rect 11084 8828 11104 8892
rect 5732 8812 11104 8828
rect 5732 8748 11020 8812
rect 11084 8748 11104 8812
rect 5732 8732 11104 8748
rect 5732 8668 11020 8732
rect 11084 8668 11104 8732
rect 5732 8652 11104 8668
rect 5732 8588 11020 8652
rect 11084 8588 11104 8652
rect 5732 8572 11104 8588
rect 5732 8508 11020 8572
rect 11084 8508 11104 8572
rect 5732 8492 11104 8508
rect 5732 8428 11020 8492
rect 11084 8428 11104 8492
rect 5732 8412 11104 8428
rect 5732 8348 11020 8412
rect 11084 8348 11104 8412
rect 5732 8332 11104 8348
rect 5732 8268 11020 8332
rect 11084 8268 11104 8332
rect 5732 8252 11104 8268
rect 5732 8188 11020 8252
rect 11084 8188 11104 8252
rect 5732 8172 11104 8188
rect 5732 8108 11020 8172
rect 11084 8108 11104 8172
rect 5732 8092 11104 8108
rect 5732 8028 11020 8092
rect 11084 8028 11104 8092
rect 5732 8012 11104 8028
rect 5732 7948 11020 8012
rect 11084 7948 11104 8012
rect 5732 7932 11104 7948
rect 5732 7868 11020 7932
rect 11084 7868 11104 7932
rect 5732 7852 11104 7868
rect 5732 7788 11020 7852
rect 11084 7788 11104 7852
rect 5732 7772 11104 7788
rect 5732 7708 11020 7772
rect 11084 7708 11104 7772
rect 5732 7692 11104 7708
rect 5732 7628 11020 7692
rect 11084 7628 11104 7692
rect 5732 7612 11104 7628
rect 5732 7548 11020 7612
rect 11084 7548 11104 7612
rect 5732 7532 11104 7548
rect 5732 7468 11020 7532
rect 11084 7468 11104 7532
rect 5732 7452 11104 7468
rect 5732 7388 11020 7452
rect 11084 7388 11104 7452
rect 5732 7372 11104 7388
rect 5732 7308 11020 7372
rect 11084 7308 11104 7372
rect 5732 7292 11104 7308
rect 5732 7228 11020 7292
rect 11084 7228 11104 7292
rect 5732 7212 11104 7228
rect 5732 7148 11020 7212
rect 11084 7148 11104 7212
rect 5732 7132 11104 7148
rect 5732 7068 11020 7132
rect 11084 7068 11104 7132
rect 5732 7052 11104 7068
rect 5732 6988 11020 7052
rect 11084 6988 11104 7052
rect 5732 6972 11104 6988
rect 5732 6908 11020 6972
rect 11084 6908 11104 6972
rect 5732 6892 11104 6908
rect 5732 6828 11020 6892
rect 11084 6828 11104 6892
rect 5732 6812 11104 6828
rect 5732 6748 11020 6812
rect 11084 6748 11104 6812
rect 5732 6732 11104 6748
rect 5732 6668 11020 6732
rect 11084 6668 11104 6732
rect 5732 6652 11104 6668
rect 5732 6588 11020 6652
rect 11084 6588 11104 6652
rect 5732 6572 11104 6588
rect 5732 6508 11020 6572
rect 11084 6508 11104 6572
rect 5732 6492 11104 6508
rect 5732 6428 11020 6492
rect 11084 6428 11104 6492
rect 5732 6412 11104 6428
rect 5732 6348 11020 6412
rect 11084 6348 11104 6412
rect 5732 6332 11104 6348
rect 5732 6268 11020 6332
rect 11084 6268 11104 6332
rect 5732 6252 11104 6268
rect 5732 6188 11020 6252
rect 11084 6188 11104 6252
rect 5732 6172 11104 6188
rect 5732 6108 11020 6172
rect 11084 6108 11104 6172
rect 5732 6092 11104 6108
rect 5732 6028 11020 6092
rect 11084 6028 11104 6092
rect 5732 6012 11104 6028
rect 5732 5948 11020 6012
rect 11084 5948 11104 6012
rect 5732 5932 11104 5948
rect 5732 5868 11020 5932
rect 11084 5868 11104 5932
rect 5732 5852 11104 5868
rect 5732 5788 11020 5852
rect 11084 5788 11104 5852
rect 5732 5772 11104 5788
rect 5732 5708 11020 5772
rect 11084 5708 11104 5772
rect 5732 5692 11104 5708
rect 5732 5628 11020 5692
rect 11084 5628 11104 5692
rect 5732 5612 11104 5628
rect 5732 5548 11020 5612
rect 11084 5548 11104 5612
rect 5732 5532 11104 5548
rect 5732 5468 11020 5532
rect 11084 5468 11104 5532
rect 5732 5440 11104 5468
rect 11344 10492 16716 10520
rect 11344 10428 16632 10492
rect 16696 10428 16716 10492
rect 11344 10412 16716 10428
rect 11344 10348 16632 10412
rect 16696 10348 16716 10412
rect 11344 10332 16716 10348
rect 11344 10268 16632 10332
rect 16696 10268 16716 10332
rect 11344 10252 16716 10268
rect 11344 10188 16632 10252
rect 16696 10188 16716 10252
rect 11344 10172 16716 10188
rect 11344 10108 16632 10172
rect 16696 10108 16716 10172
rect 11344 10092 16716 10108
rect 11344 10028 16632 10092
rect 16696 10028 16716 10092
rect 11344 10012 16716 10028
rect 11344 9948 16632 10012
rect 16696 9948 16716 10012
rect 11344 9932 16716 9948
rect 11344 9868 16632 9932
rect 16696 9868 16716 9932
rect 11344 9852 16716 9868
rect 11344 9788 16632 9852
rect 16696 9788 16716 9852
rect 11344 9772 16716 9788
rect 11344 9708 16632 9772
rect 16696 9708 16716 9772
rect 11344 9692 16716 9708
rect 11344 9628 16632 9692
rect 16696 9628 16716 9692
rect 11344 9612 16716 9628
rect 11344 9548 16632 9612
rect 16696 9548 16716 9612
rect 11344 9532 16716 9548
rect 11344 9468 16632 9532
rect 16696 9468 16716 9532
rect 11344 9452 16716 9468
rect 11344 9388 16632 9452
rect 16696 9388 16716 9452
rect 11344 9372 16716 9388
rect 11344 9308 16632 9372
rect 16696 9308 16716 9372
rect 11344 9292 16716 9308
rect 11344 9228 16632 9292
rect 16696 9228 16716 9292
rect 11344 9212 16716 9228
rect 11344 9148 16632 9212
rect 16696 9148 16716 9212
rect 11344 9132 16716 9148
rect 11344 9068 16632 9132
rect 16696 9068 16716 9132
rect 11344 9052 16716 9068
rect 11344 8988 16632 9052
rect 16696 8988 16716 9052
rect 11344 8972 16716 8988
rect 11344 8908 16632 8972
rect 16696 8908 16716 8972
rect 11344 8892 16716 8908
rect 11344 8828 16632 8892
rect 16696 8828 16716 8892
rect 11344 8812 16716 8828
rect 11344 8748 16632 8812
rect 16696 8748 16716 8812
rect 11344 8732 16716 8748
rect 11344 8668 16632 8732
rect 16696 8668 16716 8732
rect 11344 8652 16716 8668
rect 11344 8588 16632 8652
rect 16696 8588 16716 8652
rect 11344 8572 16716 8588
rect 11344 8508 16632 8572
rect 16696 8508 16716 8572
rect 11344 8492 16716 8508
rect 11344 8428 16632 8492
rect 16696 8428 16716 8492
rect 11344 8412 16716 8428
rect 11344 8348 16632 8412
rect 16696 8348 16716 8412
rect 11344 8332 16716 8348
rect 11344 8268 16632 8332
rect 16696 8268 16716 8332
rect 11344 8252 16716 8268
rect 11344 8188 16632 8252
rect 16696 8188 16716 8252
rect 11344 8172 16716 8188
rect 11344 8108 16632 8172
rect 16696 8108 16716 8172
rect 11344 8092 16716 8108
rect 11344 8028 16632 8092
rect 16696 8028 16716 8092
rect 11344 8012 16716 8028
rect 11344 7948 16632 8012
rect 16696 7948 16716 8012
rect 11344 7932 16716 7948
rect 11344 7868 16632 7932
rect 16696 7868 16716 7932
rect 11344 7852 16716 7868
rect 11344 7788 16632 7852
rect 16696 7788 16716 7852
rect 11344 7772 16716 7788
rect 11344 7708 16632 7772
rect 16696 7708 16716 7772
rect 11344 7692 16716 7708
rect 11344 7628 16632 7692
rect 16696 7628 16716 7692
rect 11344 7612 16716 7628
rect 11344 7548 16632 7612
rect 16696 7548 16716 7612
rect 11344 7532 16716 7548
rect 11344 7468 16632 7532
rect 16696 7468 16716 7532
rect 11344 7452 16716 7468
rect 11344 7388 16632 7452
rect 16696 7388 16716 7452
rect 11344 7372 16716 7388
rect 11344 7308 16632 7372
rect 16696 7308 16716 7372
rect 11344 7292 16716 7308
rect 11344 7228 16632 7292
rect 16696 7228 16716 7292
rect 11344 7212 16716 7228
rect 11344 7148 16632 7212
rect 16696 7148 16716 7212
rect 11344 7132 16716 7148
rect 11344 7068 16632 7132
rect 16696 7068 16716 7132
rect 11344 7052 16716 7068
rect 11344 6988 16632 7052
rect 16696 6988 16716 7052
rect 11344 6972 16716 6988
rect 11344 6908 16632 6972
rect 16696 6908 16716 6972
rect 11344 6892 16716 6908
rect 11344 6828 16632 6892
rect 16696 6828 16716 6892
rect 11344 6812 16716 6828
rect 11344 6748 16632 6812
rect 16696 6748 16716 6812
rect 11344 6732 16716 6748
rect 11344 6668 16632 6732
rect 16696 6668 16716 6732
rect 11344 6652 16716 6668
rect 11344 6588 16632 6652
rect 16696 6588 16716 6652
rect 11344 6572 16716 6588
rect 11344 6508 16632 6572
rect 16696 6508 16716 6572
rect 11344 6492 16716 6508
rect 11344 6428 16632 6492
rect 16696 6428 16716 6492
rect 11344 6412 16716 6428
rect 11344 6348 16632 6412
rect 16696 6348 16716 6412
rect 11344 6332 16716 6348
rect 11344 6268 16632 6332
rect 16696 6268 16716 6332
rect 11344 6252 16716 6268
rect 11344 6188 16632 6252
rect 16696 6188 16716 6252
rect 11344 6172 16716 6188
rect 11344 6108 16632 6172
rect 16696 6108 16716 6172
rect 11344 6092 16716 6108
rect 11344 6028 16632 6092
rect 16696 6028 16716 6092
rect 11344 6012 16716 6028
rect 11344 5948 16632 6012
rect 16696 5948 16716 6012
rect 11344 5932 16716 5948
rect 11344 5868 16632 5932
rect 16696 5868 16716 5932
rect 11344 5852 16716 5868
rect 11344 5788 16632 5852
rect 16696 5788 16716 5852
rect 11344 5772 16716 5788
rect 11344 5708 16632 5772
rect 16696 5708 16716 5772
rect 11344 5692 16716 5708
rect 11344 5628 16632 5692
rect 16696 5628 16716 5692
rect 11344 5612 16716 5628
rect 11344 5548 16632 5612
rect 16696 5548 16716 5612
rect 11344 5532 16716 5548
rect 11344 5468 16632 5532
rect 16696 5468 16716 5532
rect 11344 5440 16716 5468
rect 16956 10492 22328 10520
rect 16956 10428 22244 10492
rect 22308 10428 22328 10492
rect 16956 10412 22328 10428
rect 16956 10348 22244 10412
rect 22308 10348 22328 10412
rect 16956 10332 22328 10348
rect 16956 10268 22244 10332
rect 22308 10268 22328 10332
rect 16956 10252 22328 10268
rect 16956 10188 22244 10252
rect 22308 10188 22328 10252
rect 16956 10172 22328 10188
rect 16956 10108 22244 10172
rect 22308 10108 22328 10172
rect 16956 10092 22328 10108
rect 16956 10028 22244 10092
rect 22308 10028 22328 10092
rect 16956 10012 22328 10028
rect 16956 9948 22244 10012
rect 22308 9948 22328 10012
rect 16956 9932 22328 9948
rect 16956 9868 22244 9932
rect 22308 9868 22328 9932
rect 16956 9852 22328 9868
rect 16956 9788 22244 9852
rect 22308 9788 22328 9852
rect 16956 9772 22328 9788
rect 16956 9708 22244 9772
rect 22308 9708 22328 9772
rect 16956 9692 22328 9708
rect 16956 9628 22244 9692
rect 22308 9628 22328 9692
rect 16956 9612 22328 9628
rect 16956 9548 22244 9612
rect 22308 9548 22328 9612
rect 16956 9532 22328 9548
rect 16956 9468 22244 9532
rect 22308 9468 22328 9532
rect 16956 9452 22328 9468
rect 16956 9388 22244 9452
rect 22308 9388 22328 9452
rect 16956 9372 22328 9388
rect 16956 9308 22244 9372
rect 22308 9308 22328 9372
rect 16956 9292 22328 9308
rect 16956 9228 22244 9292
rect 22308 9228 22328 9292
rect 16956 9212 22328 9228
rect 16956 9148 22244 9212
rect 22308 9148 22328 9212
rect 16956 9132 22328 9148
rect 16956 9068 22244 9132
rect 22308 9068 22328 9132
rect 16956 9052 22328 9068
rect 16956 8988 22244 9052
rect 22308 8988 22328 9052
rect 16956 8972 22328 8988
rect 16956 8908 22244 8972
rect 22308 8908 22328 8972
rect 16956 8892 22328 8908
rect 16956 8828 22244 8892
rect 22308 8828 22328 8892
rect 16956 8812 22328 8828
rect 16956 8748 22244 8812
rect 22308 8748 22328 8812
rect 16956 8732 22328 8748
rect 16956 8668 22244 8732
rect 22308 8668 22328 8732
rect 16956 8652 22328 8668
rect 16956 8588 22244 8652
rect 22308 8588 22328 8652
rect 16956 8572 22328 8588
rect 16956 8508 22244 8572
rect 22308 8508 22328 8572
rect 16956 8492 22328 8508
rect 16956 8428 22244 8492
rect 22308 8428 22328 8492
rect 16956 8412 22328 8428
rect 16956 8348 22244 8412
rect 22308 8348 22328 8412
rect 16956 8332 22328 8348
rect 16956 8268 22244 8332
rect 22308 8268 22328 8332
rect 16956 8252 22328 8268
rect 16956 8188 22244 8252
rect 22308 8188 22328 8252
rect 16956 8172 22328 8188
rect 16956 8108 22244 8172
rect 22308 8108 22328 8172
rect 16956 8092 22328 8108
rect 16956 8028 22244 8092
rect 22308 8028 22328 8092
rect 16956 8012 22328 8028
rect 16956 7948 22244 8012
rect 22308 7948 22328 8012
rect 16956 7932 22328 7948
rect 16956 7868 22244 7932
rect 22308 7868 22328 7932
rect 16956 7852 22328 7868
rect 16956 7788 22244 7852
rect 22308 7788 22328 7852
rect 16956 7772 22328 7788
rect 16956 7708 22244 7772
rect 22308 7708 22328 7772
rect 16956 7692 22328 7708
rect 16956 7628 22244 7692
rect 22308 7628 22328 7692
rect 16956 7612 22328 7628
rect 16956 7548 22244 7612
rect 22308 7548 22328 7612
rect 16956 7532 22328 7548
rect 16956 7468 22244 7532
rect 22308 7468 22328 7532
rect 16956 7452 22328 7468
rect 16956 7388 22244 7452
rect 22308 7388 22328 7452
rect 16956 7372 22328 7388
rect 16956 7308 22244 7372
rect 22308 7308 22328 7372
rect 16956 7292 22328 7308
rect 16956 7228 22244 7292
rect 22308 7228 22328 7292
rect 16956 7212 22328 7228
rect 16956 7148 22244 7212
rect 22308 7148 22328 7212
rect 16956 7132 22328 7148
rect 16956 7068 22244 7132
rect 22308 7068 22328 7132
rect 16956 7052 22328 7068
rect 16956 6988 22244 7052
rect 22308 6988 22328 7052
rect 16956 6972 22328 6988
rect 16956 6908 22244 6972
rect 22308 6908 22328 6972
rect 16956 6892 22328 6908
rect 16956 6828 22244 6892
rect 22308 6828 22328 6892
rect 16956 6812 22328 6828
rect 16956 6748 22244 6812
rect 22308 6748 22328 6812
rect 16956 6732 22328 6748
rect 16956 6668 22244 6732
rect 22308 6668 22328 6732
rect 16956 6652 22328 6668
rect 16956 6588 22244 6652
rect 22308 6588 22328 6652
rect 16956 6572 22328 6588
rect 16956 6508 22244 6572
rect 22308 6508 22328 6572
rect 16956 6492 22328 6508
rect 16956 6428 22244 6492
rect 22308 6428 22328 6492
rect 16956 6412 22328 6428
rect 16956 6348 22244 6412
rect 22308 6348 22328 6412
rect 16956 6332 22328 6348
rect 16956 6268 22244 6332
rect 22308 6268 22328 6332
rect 16956 6252 22328 6268
rect 16956 6188 22244 6252
rect 22308 6188 22328 6252
rect 16956 6172 22328 6188
rect 16956 6108 22244 6172
rect 22308 6108 22328 6172
rect 16956 6092 22328 6108
rect 16956 6028 22244 6092
rect 22308 6028 22328 6092
rect 16956 6012 22328 6028
rect 16956 5948 22244 6012
rect 22308 5948 22328 6012
rect 16956 5932 22328 5948
rect 16956 5868 22244 5932
rect 22308 5868 22328 5932
rect 16956 5852 22328 5868
rect 16956 5788 22244 5852
rect 22308 5788 22328 5852
rect 16956 5772 22328 5788
rect 16956 5708 22244 5772
rect 22308 5708 22328 5772
rect 16956 5692 22328 5708
rect 16956 5628 22244 5692
rect 22308 5628 22328 5692
rect 16956 5612 22328 5628
rect 16956 5548 22244 5612
rect 22308 5548 22328 5612
rect 16956 5532 22328 5548
rect 16956 5468 22244 5532
rect 22308 5468 22328 5532
rect 16956 5440 22328 5468
rect 22568 10492 27940 10520
rect 22568 10428 27856 10492
rect 27920 10428 27940 10492
rect 22568 10412 27940 10428
rect 22568 10348 27856 10412
rect 27920 10348 27940 10412
rect 22568 10332 27940 10348
rect 22568 10268 27856 10332
rect 27920 10268 27940 10332
rect 22568 10252 27940 10268
rect 22568 10188 27856 10252
rect 27920 10188 27940 10252
rect 22568 10172 27940 10188
rect 22568 10108 27856 10172
rect 27920 10108 27940 10172
rect 22568 10092 27940 10108
rect 22568 10028 27856 10092
rect 27920 10028 27940 10092
rect 22568 10012 27940 10028
rect 22568 9948 27856 10012
rect 27920 9948 27940 10012
rect 22568 9932 27940 9948
rect 22568 9868 27856 9932
rect 27920 9868 27940 9932
rect 22568 9852 27940 9868
rect 22568 9788 27856 9852
rect 27920 9788 27940 9852
rect 22568 9772 27940 9788
rect 22568 9708 27856 9772
rect 27920 9708 27940 9772
rect 22568 9692 27940 9708
rect 22568 9628 27856 9692
rect 27920 9628 27940 9692
rect 22568 9612 27940 9628
rect 22568 9548 27856 9612
rect 27920 9548 27940 9612
rect 22568 9532 27940 9548
rect 22568 9468 27856 9532
rect 27920 9468 27940 9532
rect 22568 9452 27940 9468
rect 22568 9388 27856 9452
rect 27920 9388 27940 9452
rect 22568 9372 27940 9388
rect 22568 9308 27856 9372
rect 27920 9308 27940 9372
rect 22568 9292 27940 9308
rect 22568 9228 27856 9292
rect 27920 9228 27940 9292
rect 22568 9212 27940 9228
rect 22568 9148 27856 9212
rect 27920 9148 27940 9212
rect 22568 9132 27940 9148
rect 22568 9068 27856 9132
rect 27920 9068 27940 9132
rect 22568 9052 27940 9068
rect 22568 8988 27856 9052
rect 27920 8988 27940 9052
rect 22568 8972 27940 8988
rect 22568 8908 27856 8972
rect 27920 8908 27940 8972
rect 22568 8892 27940 8908
rect 22568 8828 27856 8892
rect 27920 8828 27940 8892
rect 22568 8812 27940 8828
rect 22568 8748 27856 8812
rect 27920 8748 27940 8812
rect 22568 8732 27940 8748
rect 22568 8668 27856 8732
rect 27920 8668 27940 8732
rect 22568 8652 27940 8668
rect 22568 8588 27856 8652
rect 27920 8588 27940 8652
rect 22568 8572 27940 8588
rect 22568 8508 27856 8572
rect 27920 8508 27940 8572
rect 22568 8492 27940 8508
rect 22568 8428 27856 8492
rect 27920 8428 27940 8492
rect 22568 8412 27940 8428
rect 22568 8348 27856 8412
rect 27920 8348 27940 8412
rect 22568 8332 27940 8348
rect 22568 8268 27856 8332
rect 27920 8268 27940 8332
rect 22568 8252 27940 8268
rect 22568 8188 27856 8252
rect 27920 8188 27940 8252
rect 22568 8172 27940 8188
rect 22568 8108 27856 8172
rect 27920 8108 27940 8172
rect 22568 8092 27940 8108
rect 22568 8028 27856 8092
rect 27920 8028 27940 8092
rect 22568 8012 27940 8028
rect 22568 7948 27856 8012
rect 27920 7948 27940 8012
rect 22568 7932 27940 7948
rect 22568 7868 27856 7932
rect 27920 7868 27940 7932
rect 22568 7852 27940 7868
rect 22568 7788 27856 7852
rect 27920 7788 27940 7852
rect 22568 7772 27940 7788
rect 22568 7708 27856 7772
rect 27920 7708 27940 7772
rect 22568 7692 27940 7708
rect 22568 7628 27856 7692
rect 27920 7628 27940 7692
rect 22568 7612 27940 7628
rect 22568 7548 27856 7612
rect 27920 7548 27940 7612
rect 22568 7532 27940 7548
rect 22568 7468 27856 7532
rect 27920 7468 27940 7532
rect 22568 7452 27940 7468
rect 22568 7388 27856 7452
rect 27920 7388 27940 7452
rect 22568 7372 27940 7388
rect 22568 7308 27856 7372
rect 27920 7308 27940 7372
rect 22568 7292 27940 7308
rect 22568 7228 27856 7292
rect 27920 7228 27940 7292
rect 22568 7212 27940 7228
rect 22568 7148 27856 7212
rect 27920 7148 27940 7212
rect 22568 7132 27940 7148
rect 22568 7068 27856 7132
rect 27920 7068 27940 7132
rect 22568 7052 27940 7068
rect 22568 6988 27856 7052
rect 27920 6988 27940 7052
rect 22568 6972 27940 6988
rect 22568 6908 27856 6972
rect 27920 6908 27940 6972
rect 22568 6892 27940 6908
rect 22568 6828 27856 6892
rect 27920 6828 27940 6892
rect 22568 6812 27940 6828
rect 22568 6748 27856 6812
rect 27920 6748 27940 6812
rect 22568 6732 27940 6748
rect 22568 6668 27856 6732
rect 27920 6668 27940 6732
rect 22568 6652 27940 6668
rect 22568 6588 27856 6652
rect 27920 6588 27940 6652
rect 22568 6572 27940 6588
rect 22568 6508 27856 6572
rect 27920 6508 27940 6572
rect 22568 6492 27940 6508
rect 22568 6428 27856 6492
rect 27920 6428 27940 6492
rect 22568 6412 27940 6428
rect 22568 6348 27856 6412
rect 27920 6348 27940 6412
rect 22568 6332 27940 6348
rect 22568 6268 27856 6332
rect 27920 6268 27940 6332
rect 22568 6252 27940 6268
rect 22568 6188 27856 6252
rect 27920 6188 27940 6252
rect 22568 6172 27940 6188
rect 22568 6108 27856 6172
rect 27920 6108 27940 6172
rect 22568 6092 27940 6108
rect 22568 6028 27856 6092
rect 27920 6028 27940 6092
rect 22568 6012 27940 6028
rect 22568 5948 27856 6012
rect 27920 5948 27940 6012
rect 22568 5932 27940 5948
rect 22568 5868 27856 5932
rect 27920 5868 27940 5932
rect 22568 5852 27940 5868
rect 22568 5788 27856 5852
rect 27920 5788 27940 5852
rect 22568 5772 27940 5788
rect 22568 5708 27856 5772
rect 27920 5708 27940 5772
rect 22568 5692 27940 5708
rect 22568 5628 27856 5692
rect 27920 5628 27940 5692
rect 22568 5612 27940 5628
rect 22568 5548 27856 5612
rect 27920 5548 27940 5612
rect 22568 5532 27940 5548
rect 22568 5468 27856 5532
rect 27920 5468 27940 5532
rect 22568 5440 27940 5468
rect 28180 10492 33552 10520
rect 28180 10428 33468 10492
rect 33532 10428 33552 10492
rect 28180 10412 33552 10428
rect 28180 10348 33468 10412
rect 33532 10348 33552 10412
rect 28180 10332 33552 10348
rect 28180 10268 33468 10332
rect 33532 10268 33552 10332
rect 28180 10252 33552 10268
rect 28180 10188 33468 10252
rect 33532 10188 33552 10252
rect 28180 10172 33552 10188
rect 28180 10108 33468 10172
rect 33532 10108 33552 10172
rect 28180 10092 33552 10108
rect 28180 10028 33468 10092
rect 33532 10028 33552 10092
rect 28180 10012 33552 10028
rect 28180 9948 33468 10012
rect 33532 9948 33552 10012
rect 28180 9932 33552 9948
rect 28180 9868 33468 9932
rect 33532 9868 33552 9932
rect 28180 9852 33552 9868
rect 28180 9788 33468 9852
rect 33532 9788 33552 9852
rect 28180 9772 33552 9788
rect 28180 9708 33468 9772
rect 33532 9708 33552 9772
rect 28180 9692 33552 9708
rect 28180 9628 33468 9692
rect 33532 9628 33552 9692
rect 28180 9612 33552 9628
rect 28180 9548 33468 9612
rect 33532 9548 33552 9612
rect 28180 9532 33552 9548
rect 28180 9468 33468 9532
rect 33532 9468 33552 9532
rect 28180 9452 33552 9468
rect 28180 9388 33468 9452
rect 33532 9388 33552 9452
rect 28180 9372 33552 9388
rect 28180 9308 33468 9372
rect 33532 9308 33552 9372
rect 28180 9292 33552 9308
rect 28180 9228 33468 9292
rect 33532 9228 33552 9292
rect 28180 9212 33552 9228
rect 28180 9148 33468 9212
rect 33532 9148 33552 9212
rect 28180 9132 33552 9148
rect 28180 9068 33468 9132
rect 33532 9068 33552 9132
rect 28180 9052 33552 9068
rect 28180 8988 33468 9052
rect 33532 8988 33552 9052
rect 28180 8972 33552 8988
rect 28180 8908 33468 8972
rect 33532 8908 33552 8972
rect 28180 8892 33552 8908
rect 28180 8828 33468 8892
rect 33532 8828 33552 8892
rect 28180 8812 33552 8828
rect 28180 8748 33468 8812
rect 33532 8748 33552 8812
rect 28180 8732 33552 8748
rect 28180 8668 33468 8732
rect 33532 8668 33552 8732
rect 28180 8652 33552 8668
rect 28180 8588 33468 8652
rect 33532 8588 33552 8652
rect 28180 8572 33552 8588
rect 28180 8508 33468 8572
rect 33532 8508 33552 8572
rect 28180 8492 33552 8508
rect 28180 8428 33468 8492
rect 33532 8428 33552 8492
rect 28180 8412 33552 8428
rect 28180 8348 33468 8412
rect 33532 8348 33552 8412
rect 28180 8332 33552 8348
rect 28180 8268 33468 8332
rect 33532 8268 33552 8332
rect 28180 8252 33552 8268
rect 28180 8188 33468 8252
rect 33532 8188 33552 8252
rect 28180 8172 33552 8188
rect 28180 8108 33468 8172
rect 33532 8108 33552 8172
rect 28180 8092 33552 8108
rect 28180 8028 33468 8092
rect 33532 8028 33552 8092
rect 28180 8012 33552 8028
rect 28180 7948 33468 8012
rect 33532 7948 33552 8012
rect 28180 7932 33552 7948
rect 28180 7868 33468 7932
rect 33532 7868 33552 7932
rect 28180 7852 33552 7868
rect 28180 7788 33468 7852
rect 33532 7788 33552 7852
rect 28180 7772 33552 7788
rect 28180 7708 33468 7772
rect 33532 7708 33552 7772
rect 28180 7692 33552 7708
rect 28180 7628 33468 7692
rect 33532 7628 33552 7692
rect 28180 7612 33552 7628
rect 28180 7548 33468 7612
rect 33532 7548 33552 7612
rect 28180 7532 33552 7548
rect 28180 7468 33468 7532
rect 33532 7468 33552 7532
rect 28180 7452 33552 7468
rect 28180 7388 33468 7452
rect 33532 7388 33552 7452
rect 28180 7372 33552 7388
rect 28180 7308 33468 7372
rect 33532 7308 33552 7372
rect 28180 7292 33552 7308
rect 28180 7228 33468 7292
rect 33532 7228 33552 7292
rect 28180 7212 33552 7228
rect 28180 7148 33468 7212
rect 33532 7148 33552 7212
rect 28180 7132 33552 7148
rect 28180 7068 33468 7132
rect 33532 7068 33552 7132
rect 28180 7052 33552 7068
rect 28180 6988 33468 7052
rect 33532 6988 33552 7052
rect 28180 6972 33552 6988
rect 28180 6908 33468 6972
rect 33532 6908 33552 6972
rect 28180 6892 33552 6908
rect 28180 6828 33468 6892
rect 33532 6828 33552 6892
rect 28180 6812 33552 6828
rect 28180 6748 33468 6812
rect 33532 6748 33552 6812
rect 28180 6732 33552 6748
rect 28180 6668 33468 6732
rect 33532 6668 33552 6732
rect 28180 6652 33552 6668
rect 28180 6588 33468 6652
rect 33532 6588 33552 6652
rect 28180 6572 33552 6588
rect 28180 6508 33468 6572
rect 33532 6508 33552 6572
rect 28180 6492 33552 6508
rect 28180 6428 33468 6492
rect 33532 6428 33552 6492
rect 28180 6412 33552 6428
rect 28180 6348 33468 6412
rect 33532 6348 33552 6412
rect 28180 6332 33552 6348
rect 28180 6268 33468 6332
rect 33532 6268 33552 6332
rect 28180 6252 33552 6268
rect 28180 6188 33468 6252
rect 33532 6188 33552 6252
rect 28180 6172 33552 6188
rect 28180 6108 33468 6172
rect 33532 6108 33552 6172
rect 28180 6092 33552 6108
rect 28180 6028 33468 6092
rect 33532 6028 33552 6092
rect 28180 6012 33552 6028
rect 28180 5948 33468 6012
rect 33532 5948 33552 6012
rect 28180 5932 33552 5948
rect 28180 5868 33468 5932
rect 33532 5868 33552 5932
rect 28180 5852 33552 5868
rect 28180 5788 33468 5852
rect 33532 5788 33552 5852
rect 28180 5772 33552 5788
rect 28180 5708 33468 5772
rect 33532 5708 33552 5772
rect 28180 5692 33552 5708
rect 28180 5628 33468 5692
rect 33532 5628 33552 5692
rect 28180 5612 33552 5628
rect 28180 5548 33468 5612
rect 33532 5548 33552 5612
rect 28180 5532 33552 5548
rect 28180 5468 33468 5532
rect 33532 5468 33552 5532
rect 28180 5440 33552 5468
rect 33792 10492 39164 10520
rect 33792 10428 39080 10492
rect 39144 10428 39164 10492
rect 33792 10412 39164 10428
rect 33792 10348 39080 10412
rect 39144 10348 39164 10412
rect 33792 10332 39164 10348
rect 33792 10268 39080 10332
rect 39144 10268 39164 10332
rect 33792 10252 39164 10268
rect 33792 10188 39080 10252
rect 39144 10188 39164 10252
rect 33792 10172 39164 10188
rect 33792 10108 39080 10172
rect 39144 10108 39164 10172
rect 33792 10092 39164 10108
rect 33792 10028 39080 10092
rect 39144 10028 39164 10092
rect 33792 10012 39164 10028
rect 33792 9948 39080 10012
rect 39144 9948 39164 10012
rect 33792 9932 39164 9948
rect 33792 9868 39080 9932
rect 39144 9868 39164 9932
rect 33792 9852 39164 9868
rect 33792 9788 39080 9852
rect 39144 9788 39164 9852
rect 33792 9772 39164 9788
rect 33792 9708 39080 9772
rect 39144 9708 39164 9772
rect 33792 9692 39164 9708
rect 33792 9628 39080 9692
rect 39144 9628 39164 9692
rect 33792 9612 39164 9628
rect 33792 9548 39080 9612
rect 39144 9548 39164 9612
rect 33792 9532 39164 9548
rect 33792 9468 39080 9532
rect 39144 9468 39164 9532
rect 33792 9452 39164 9468
rect 33792 9388 39080 9452
rect 39144 9388 39164 9452
rect 33792 9372 39164 9388
rect 33792 9308 39080 9372
rect 39144 9308 39164 9372
rect 33792 9292 39164 9308
rect 33792 9228 39080 9292
rect 39144 9228 39164 9292
rect 33792 9212 39164 9228
rect 33792 9148 39080 9212
rect 39144 9148 39164 9212
rect 33792 9132 39164 9148
rect 33792 9068 39080 9132
rect 39144 9068 39164 9132
rect 33792 9052 39164 9068
rect 33792 8988 39080 9052
rect 39144 8988 39164 9052
rect 33792 8972 39164 8988
rect 33792 8908 39080 8972
rect 39144 8908 39164 8972
rect 33792 8892 39164 8908
rect 33792 8828 39080 8892
rect 39144 8828 39164 8892
rect 33792 8812 39164 8828
rect 33792 8748 39080 8812
rect 39144 8748 39164 8812
rect 33792 8732 39164 8748
rect 33792 8668 39080 8732
rect 39144 8668 39164 8732
rect 33792 8652 39164 8668
rect 33792 8588 39080 8652
rect 39144 8588 39164 8652
rect 33792 8572 39164 8588
rect 33792 8508 39080 8572
rect 39144 8508 39164 8572
rect 33792 8492 39164 8508
rect 33792 8428 39080 8492
rect 39144 8428 39164 8492
rect 33792 8412 39164 8428
rect 33792 8348 39080 8412
rect 39144 8348 39164 8412
rect 33792 8332 39164 8348
rect 33792 8268 39080 8332
rect 39144 8268 39164 8332
rect 33792 8252 39164 8268
rect 33792 8188 39080 8252
rect 39144 8188 39164 8252
rect 33792 8172 39164 8188
rect 33792 8108 39080 8172
rect 39144 8108 39164 8172
rect 33792 8092 39164 8108
rect 33792 8028 39080 8092
rect 39144 8028 39164 8092
rect 33792 8012 39164 8028
rect 33792 7948 39080 8012
rect 39144 7948 39164 8012
rect 33792 7932 39164 7948
rect 33792 7868 39080 7932
rect 39144 7868 39164 7932
rect 33792 7852 39164 7868
rect 33792 7788 39080 7852
rect 39144 7788 39164 7852
rect 33792 7772 39164 7788
rect 33792 7708 39080 7772
rect 39144 7708 39164 7772
rect 33792 7692 39164 7708
rect 33792 7628 39080 7692
rect 39144 7628 39164 7692
rect 33792 7612 39164 7628
rect 33792 7548 39080 7612
rect 39144 7548 39164 7612
rect 33792 7532 39164 7548
rect 33792 7468 39080 7532
rect 39144 7468 39164 7532
rect 33792 7452 39164 7468
rect 33792 7388 39080 7452
rect 39144 7388 39164 7452
rect 33792 7372 39164 7388
rect 33792 7308 39080 7372
rect 39144 7308 39164 7372
rect 33792 7292 39164 7308
rect 33792 7228 39080 7292
rect 39144 7228 39164 7292
rect 33792 7212 39164 7228
rect 33792 7148 39080 7212
rect 39144 7148 39164 7212
rect 33792 7132 39164 7148
rect 33792 7068 39080 7132
rect 39144 7068 39164 7132
rect 33792 7052 39164 7068
rect 33792 6988 39080 7052
rect 39144 6988 39164 7052
rect 33792 6972 39164 6988
rect 33792 6908 39080 6972
rect 39144 6908 39164 6972
rect 33792 6892 39164 6908
rect 33792 6828 39080 6892
rect 39144 6828 39164 6892
rect 33792 6812 39164 6828
rect 33792 6748 39080 6812
rect 39144 6748 39164 6812
rect 33792 6732 39164 6748
rect 33792 6668 39080 6732
rect 39144 6668 39164 6732
rect 33792 6652 39164 6668
rect 33792 6588 39080 6652
rect 39144 6588 39164 6652
rect 33792 6572 39164 6588
rect 33792 6508 39080 6572
rect 39144 6508 39164 6572
rect 33792 6492 39164 6508
rect 33792 6428 39080 6492
rect 39144 6428 39164 6492
rect 33792 6412 39164 6428
rect 33792 6348 39080 6412
rect 39144 6348 39164 6412
rect 33792 6332 39164 6348
rect 33792 6268 39080 6332
rect 39144 6268 39164 6332
rect 33792 6252 39164 6268
rect 33792 6188 39080 6252
rect 39144 6188 39164 6252
rect 33792 6172 39164 6188
rect 33792 6108 39080 6172
rect 39144 6108 39164 6172
rect 33792 6092 39164 6108
rect 33792 6028 39080 6092
rect 39144 6028 39164 6092
rect 33792 6012 39164 6028
rect 33792 5948 39080 6012
rect 39144 5948 39164 6012
rect 33792 5932 39164 5948
rect 33792 5868 39080 5932
rect 39144 5868 39164 5932
rect 33792 5852 39164 5868
rect 33792 5788 39080 5852
rect 39144 5788 39164 5852
rect 33792 5772 39164 5788
rect 33792 5708 39080 5772
rect 39144 5708 39164 5772
rect 33792 5692 39164 5708
rect 33792 5628 39080 5692
rect 39144 5628 39164 5692
rect 33792 5612 39164 5628
rect 33792 5548 39080 5612
rect 39144 5548 39164 5612
rect 33792 5532 39164 5548
rect 33792 5468 39080 5532
rect 39144 5468 39164 5532
rect 33792 5440 39164 5468
rect -39164 5172 -33792 5200
rect -39164 5108 -33876 5172
rect -33812 5108 -33792 5172
rect -39164 5092 -33792 5108
rect -39164 5028 -33876 5092
rect -33812 5028 -33792 5092
rect -39164 5012 -33792 5028
rect -39164 4948 -33876 5012
rect -33812 4948 -33792 5012
rect -39164 4932 -33792 4948
rect -39164 4868 -33876 4932
rect -33812 4868 -33792 4932
rect -39164 4852 -33792 4868
rect -39164 4788 -33876 4852
rect -33812 4788 -33792 4852
rect -39164 4772 -33792 4788
rect -39164 4708 -33876 4772
rect -33812 4708 -33792 4772
rect -39164 4692 -33792 4708
rect -39164 4628 -33876 4692
rect -33812 4628 -33792 4692
rect -39164 4612 -33792 4628
rect -39164 4548 -33876 4612
rect -33812 4548 -33792 4612
rect -39164 4532 -33792 4548
rect -39164 4468 -33876 4532
rect -33812 4468 -33792 4532
rect -39164 4452 -33792 4468
rect -39164 4388 -33876 4452
rect -33812 4388 -33792 4452
rect -39164 4372 -33792 4388
rect -39164 4308 -33876 4372
rect -33812 4308 -33792 4372
rect -39164 4292 -33792 4308
rect -39164 4228 -33876 4292
rect -33812 4228 -33792 4292
rect -39164 4212 -33792 4228
rect -39164 4148 -33876 4212
rect -33812 4148 -33792 4212
rect -39164 4132 -33792 4148
rect -39164 4068 -33876 4132
rect -33812 4068 -33792 4132
rect -39164 4052 -33792 4068
rect -39164 3988 -33876 4052
rect -33812 3988 -33792 4052
rect -39164 3972 -33792 3988
rect -39164 3908 -33876 3972
rect -33812 3908 -33792 3972
rect -39164 3892 -33792 3908
rect -39164 3828 -33876 3892
rect -33812 3828 -33792 3892
rect -39164 3812 -33792 3828
rect -39164 3748 -33876 3812
rect -33812 3748 -33792 3812
rect -39164 3732 -33792 3748
rect -39164 3668 -33876 3732
rect -33812 3668 -33792 3732
rect -39164 3652 -33792 3668
rect -39164 3588 -33876 3652
rect -33812 3588 -33792 3652
rect -39164 3572 -33792 3588
rect -39164 3508 -33876 3572
rect -33812 3508 -33792 3572
rect -39164 3492 -33792 3508
rect -39164 3428 -33876 3492
rect -33812 3428 -33792 3492
rect -39164 3412 -33792 3428
rect -39164 3348 -33876 3412
rect -33812 3348 -33792 3412
rect -39164 3332 -33792 3348
rect -39164 3268 -33876 3332
rect -33812 3268 -33792 3332
rect -39164 3252 -33792 3268
rect -39164 3188 -33876 3252
rect -33812 3188 -33792 3252
rect -39164 3172 -33792 3188
rect -39164 3108 -33876 3172
rect -33812 3108 -33792 3172
rect -39164 3092 -33792 3108
rect -39164 3028 -33876 3092
rect -33812 3028 -33792 3092
rect -39164 3012 -33792 3028
rect -39164 2948 -33876 3012
rect -33812 2948 -33792 3012
rect -39164 2932 -33792 2948
rect -39164 2868 -33876 2932
rect -33812 2868 -33792 2932
rect -39164 2852 -33792 2868
rect -39164 2788 -33876 2852
rect -33812 2788 -33792 2852
rect -39164 2772 -33792 2788
rect -39164 2708 -33876 2772
rect -33812 2708 -33792 2772
rect -39164 2692 -33792 2708
rect -39164 2628 -33876 2692
rect -33812 2628 -33792 2692
rect -39164 2612 -33792 2628
rect -39164 2548 -33876 2612
rect -33812 2548 -33792 2612
rect -39164 2532 -33792 2548
rect -39164 2468 -33876 2532
rect -33812 2468 -33792 2532
rect -39164 2452 -33792 2468
rect -39164 2388 -33876 2452
rect -33812 2388 -33792 2452
rect -39164 2372 -33792 2388
rect -39164 2308 -33876 2372
rect -33812 2308 -33792 2372
rect -39164 2292 -33792 2308
rect -39164 2228 -33876 2292
rect -33812 2228 -33792 2292
rect -39164 2212 -33792 2228
rect -39164 2148 -33876 2212
rect -33812 2148 -33792 2212
rect -39164 2132 -33792 2148
rect -39164 2068 -33876 2132
rect -33812 2068 -33792 2132
rect -39164 2052 -33792 2068
rect -39164 1988 -33876 2052
rect -33812 1988 -33792 2052
rect -39164 1972 -33792 1988
rect -39164 1908 -33876 1972
rect -33812 1908 -33792 1972
rect -39164 1892 -33792 1908
rect -39164 1828 -33876 1892
rect -33812 1828 -33792 1892
rect -39164 1812 -33792 1828
rect -39164 1748 -33876 1812
rect -33812 1748 -33792 1812
rect -39164 1732 -33792 1748
rect -39164 1668 -33876 1732
rect -33812 1668 -33792 1732
rect -39164 1652 -33792 1668
rect -39164 1588 -33876 1652
rect -33812 1588 -33792 1652
rect -39164 1572 -33792 1588
rect -39164 1508 -33876 1572
rect -33812 1508 -33792 1572
rect -39164 1492 -33792 1508
rect -39164 1428 -33876 1492
rect -33812 1428 -33792 1492
rect -39164 1412 -33792 1428
rect -39164 1348 -33876 1412
rect -33812 1348 -33792 1412
rect -39164 1332 -33792 1348
rect -39164 1268 -33876 1332
rect -33812 1268 -33792 1332
rect -39164 1252 -33792 1268
rect -39164 1188 -33876 1252
rect -33812 1188 -33792 1252
rect -39164 1172 -33792 1188
rect -39164 1108 -33876 1172
rect -33812 1108 -33792 1172
rect -39164 1092 -33792 1108
rect -39164 1028 -33876 1092
rect -33812 1028 -33792 1092
rect -39164 1012 -33792 1028
rect -39164 948 -33876 1012
rect -33812 948 -33792 1012
rect -39164 932 -33792 948
rect -39164 868 -33876 932
rect -33812 868 -33792 932
rect -39164 852 -33792 868
rect -39164 788 -33876 852
rect -33812 788 -33792 852
rect -39164 772 -33792 788
rect -39164 708 -33876 772
rect -33812 708 -33792 772
rect -39164 692 -33792 708
rect -39164 628 -33876 692
rect -33812 628 -33792 692
rect -39164 612 -33792 628
rect -39164 548 -33876 612
rect -33812 548 -33792 612
rect -39164 532 -33792 548
rect -39164 468 -33876 532
rect -33812 468 -33792 532
rect -39164 452 -33792 468
rect -39164 388 -33876 452
rect -33812 388 -33792 452
rect -39164 372 -33792 388
rect -39164 308 -33876 372
rect -33812 308 -33792 372
rect -39164 292 -33792 308
rect -39164 228 -33876 292
rect -33812 228 -33792 292
rect -39164 212 -33792 228
rect -39164 148 -33876 212
rect -33812 148 -33792 212
rect -39164 120 -33792 148
rect -33552 5172 -28180 5200
rect -33552 5108 -28264 5172
rect -28200 5108 -28180 5172
rect -33552 5092 -28180 5108
rect -33552 5028 -28264 5092
rect -28200 5028 -28180 5092
rect -33552 5012 -28180 5028
rect -33552 4948 -28264 5012
rect -28200 4948 -28180 5012
rect -33552 4932 -28180 4948
rect -33552 4868 -28264 4932
rect -28200 4868 -28180 4932
rect -33552 4852 -28180 4868
rect -33552 4788 -28264 4852
rect -28200 4788 -28180 4852
rect -33552 4772 -28180 4788
rect -33552 4708 -28264 4772
rect -28200 4708 -28180 4772
rect -33552 4692 -28180 4708
rect -33552 4628 -28264 4692
rect -28200 4628 -28180 4692
rect -33552 4612 -28180 4628
rect -33552 4548 -28264 4612
rect -28200 4548 -28180 4612
rect -33552 4532 -28180 4548
rect -33552 4468 -28264 4532
rect -28200 4468 -28180 4532
rect -33552 4452 -28180 4468
rect -33552 4388 -28264 4452
rect -28200 4388 -28180 4452
rect -33552 4372 -28180 4388
rect -33552 4308 -28264 4372
rect -28200 4308 -28180 4372
rect -33552 4292 -28180 4308
rect -33552 4228 -28264 4292
rect -28200 4228 -28180 4292
rect -33552 4212 -28180 4228
rect -33552 4148 -28264 4212
rect -28200 4148 -28180 4212
rect -33552 4132 -28180 4148
rect -33552 4068 -28264 4132
rect -28200 4068 -28180 4132
rect -33552 4052 -28180 4068
rect -33552 3988 -28264 4052
rect -28200 3988 -28180 4052
rect -33552 3972 -28180 3988
rect -33552 3908 -28264 3972
rect -28200 3908 -28180 3972
rect -33552 3892 -28180 3908
rect -33552 3828 -28264 3892
rect -28200 3828 -28180 3892
rect -33552 3812 -28180 3828
rect -33552 3748 -28264 3812
rect -28200 3748 -28180 3812
rect -33552 3732 -28180 3748
rect -33552 3668 -28264 3732
rect -28200 3668 -28180 3732
rect -33552 3652 -28180 3668
rect -33552 3588 -28264 3652
rect -28200 3588 -28180 3652
rect -33552 3572 -28180 3588
rect -33552 3508 -28264 3572
rect -28200 3508 -28180 3572
rect -33552 3492 -28180 3508
rect -33552 3428 -28264 3492
rect -28200 3428 -28180 3492
rect -33552 3412 -28180 3428
rect -33552 3348 -28264 3412
rect -28200 3348 -28180 3412
rect -33552 3332 -28180 3348
rect -33552 3268 -28264 3332
rect -28200 3268 -28180 3332
rect -33552 3252 -28180 3268
rect -33552 3188 -28264 3252
rect -28200 3188 -28180 3252
rect -33552 3172 -28180 3188
rect -33552 3108 -28264 3172
rect -28200 3108 -28180 3172
rect -33552 3092 -28180 3108
rect -33552 3028 -28264 3092
rect -28200 3028 -28180 3092
rect -33552 3012 -28180 3028
rect -33552 2948 -28264 3012
rect -28200 2948 -28180 3012
rect -33552 2932 -28180 2948
rect -33552 2868 -28264 2932
rect -28200 2868 -28180 2932
rect -33552 2852 -28180 2868
rect -33552 2788 -28264 2852
rect -28200 2788 -28180 2852
rect -33552 2772 -28180 2788
rect -33552 2708 -28264 2772
rect -28200 2708 -28180 2772
rect -33552 2692 -28180 2708
rect -33552 2628 -28264 2692
rect -28200 2628 -28180 2692
rect -33552 2612 -28180 2628
rect -33552 2548 -28264 2612
rect -28200 2548 -28180 2612
rect -33552 2532 -28180 2548
rect -33552 2468 -28264 2532
rect -28200 2468 -28180 2532
rect -33552 2452 -28180 2468
rect -33552 2388 -28264 2452
rect -28200 2388 -28180 2452
rect -33552 2372 -28180 2388
rect -33552 2308 -28264 2372
rect -28200 2308 -28180 2372
rect -33552 2292 -28180 2308
rect -33552 2228 -28264 2292
rect -28200 2228 -28180 2292
rect -33552 2212 -28180 2228
rect -33552 2148 -28264 2212
rect -28200 2148 -28180 2212
rect -33552 2132 -28180 2148
rect -33552 2068 -28264 2132
rect -28200 2068 -28180 2132
rect -33552 2052 -28180 2068
rect -33552 1988 -28264 2052
rect -28200 1988 -28180 2052
rect -33552 1972 -28180 1988
rect -33552 1908 -28264 1972
rect -28200 1908 -28180 1972
rect -33552 1892 -28180 1908
rect -33552 1828 -28264 1892
rect -28200 1828 -28180 1892
rect -33552 1812 -28180 1828
rect -33552 1748 -28264 1812
rect -28200 1748 -28180 1812
rect -33552 1732 -28180 1748
rect -33552 1668 -28264 1732
rect -28200 1668 -28180 1732
rect -33552 1652 -28180 1668
rect -33552 1588 -28264 1652
rect -28200 1588 -28180 1652
rect -33552 1572 -28180 1588
rect -33552 1508 -28264 1572
rect -28200 1508 -28180 1572
rect -33552 1492 -28180 1508
rect -33552 1428 -28264 1492
rect -28200 1428 -28180 1492
rect -33552 1412 -28180 1428
rect -33552 1348 -28264 1412
rect -28200 1348 -28180 1412
rect -33552 1332 -28180 1348
rect -33552 1268 -28264 1332
rect -28200 1268 -28180 1332
rect -33552 1252 -28180 1268
rect -33552 1188 -28264 1252
rect -28200 1188 -28180 1252
rect -33552 1172 -28180 1188
rect -33552 1108 -28264 1172
rect -28200 1108 -28180 1172
rect -33552 1092 -28180 1108
rect -33552 1028 -28264 1092
rect -28200 1028 -28180 1092
rect -33552 1012 -28180 1028
rect -33552 948 -28264 1012
rect -28200 948 -28180 1012
rect -33552 932 -28180 948
rect -33552 868 -28264 932
rect -28200 868 -28180 932
rect -33552 852 -28180 868
rect -33552 788 -28264 852
rect -28200 788 -28180 852
rect -33552 772 -28180 788
rect -33552 708 -28264 772
rect -28200 708 -28180 772
rect -33552 692 -28180 708
rect -33552 628 -28264 692
rect -28200 628 -28180 692
rect -33552 612 -28180 628
rect -33552 548 -28264 612
rect -28200 548 -28180 612
rect -33552 532 -28180 548
rect -33552 468 -28264 532
rect -28200 468 -28180 532
rect -33552 452 -28180 468
rect -33552 388 -28264 452
rect -28200 388 -28180 452
rect -33552 372 -28180 388
rect -33552 308 -28264 372
rect -28200 308 -28180 372
rect -33552 292 -28180 308
rect -33552 228 -28264 292
rect -28200 228 -28180 292
rect -33552 212 -28180 228
rect -33552 148 -28264 212
rect -28200 148 -28180 212
rect -33552 120 -28180 148
rect -27940 5172 -22568 5200
rect -27940 5108 -22652 5172
rect -22588 5108 -22568 5172
rect -27940 5092 -22568 5108
rect -27940 5028 -22652 5092
rect -22588 5028 -22568 5092
rect -27940 5012 -22568 5028
rect -27940 4948 -22652 5012
rect -22588 4948 -22568 5012
rect -27940 4932 -22568 4948
rect -27940 4868 -22652 4932
rect -22588 4868 -22568 4932
rect -27940 4852 -22568 4868
rect -27940 4788 -22652 4852
rect -22588 4788 -22568 4852
rect -27940 4772 -22568 4788
rect -27940 4708 -22652 4772
rect -22588 4708 -22568 4772
rect -27940 4692 -22568 4708
rect -27940 4628 -22652 4692
rect -22588 4628 -22568 4692
rect -27940 4612 -22568 4628
rect -27940 4548 -22652 4612
rect -22588 4548 -22568 4612
rect -27940 4532 -22568 4548
rect -27940 4468 -22652 4532
rect -22588 4468 -22568 4532
rect -27940 4452 -22568 4468
rect -27940 4388 -22652 4452
rect -22588 4388 -22568 4452
rect -27940 4372 -22568 4388
rect -27940 4308 -22652 4372
rect -22588 4308 -22568 4372
rect -27940 4292 -22568 4308
rect -27940 4228 -22652 4292
rect -22588 4228 -22568 4292
rect -27940 4212 -22568 4228
rect -27940 4148 -22652 4212
rect -22588 4148 -22568 4212
rect -27940 4132 -22568 4148
rect -27940 4068 -22652 4132
rect -22588 4068 -22568 4132
rect -27940 4052 -22568 4068
rect -27940 3988 -22652 4052
rect -22588 3988 -22568 4052
rect -27940 3972 -22568 3988
rect -27940 3908 -22652 3972
rect -22588 3908 -22568 3972
rect -27940 3892 -22568 3908
rect -27940 3828 -22652 3892
rect -22588 3828 -22568 3892
rect -27940 3812 -22568 3828
rect -27940 3748 -22652 3812
rect -22588 3748 -22568 3812
rect -27940 3732 -22568 3748
rect -27940 3668 -22652 3732
rect -22588 3668 -22568 3732
rect -27940 3652 -22568 3668
rect -27940 3588 -22652 3652
rect -22588 3588 -22568 3652
rect -27940 3572 -22568 3588
rect -27940 3508 -22652 3572
rect -22588 3508 -22568 3572
rect -27940 3492 -22568 3508
rect -27940 3428 -22652 3492
rect -22588 3428 -22568 3492
rect -27940 3412 -22568 3428
rect -27940 3348 -22652 3412
rect -22588 3348 -22568 3412
rect -27940 3332 -22568 3348
rect -27940 3268 -22652 3332
rect -22588 3268 -22568 3332
rect -27940 3252 -22568 3268
rect -27940 3188 -22652 3252
rect -22588 3188 -22568 3252
rect -27940 3172 -22568 3188
rect -27940 3108 -22652 3172
rect -22588 3108 -22568 3172
rect -27940 3092 -22568 3108
rect -27940 3028 -22652 3092
rect -22588 3028 -22568 3092
rect -27940 3012 -22568 3028
rect -27940 2948 -22652 3012
rect -22588 2948 -22568 3012
rect -27940 2932 -22568 2948
rect -27940 2868 -22652 2932
rect -22588 2868 -22568 2932
rect -27940 2852 -22568 2868
rect -27940 2788 -22652 2852
rect -22588 2788 -22568 2852
rect -27940 2772 -22568 2788
rect -27940 2708 -22652 2772
rect -22588 2708 -22568 2772
rect -27940 2692 -22568 2708
rect -27940 2628 -22652 2692
rect -22588 2628 -22568 2692
rect -27940 2612 -22568 2628
rect -27940 2548 -22652 2612
rect -22588 2548 -22568 2612
rect -27940 2532 -22568 2548
rect -27940 2468 -22652 2532
rect -22588 2468 -22568 2532
rect -27940 2452 -22568 2468
rect -27940 2388 -22652 2452
rect -22588 2388 -22568 2452
rect -27940 2372 -22568 2388
rect -27940 2308 -22652 2372
rect -22588 2308 -22568 2372
rect -27940 2292 -22568 2308
rect -27940 2228 -22652 2292
rect -22588 2228 -22568 2292
rect -27940 2212 -22568 2228
rect -27940 2148 -22652 2212
rect -22588 2148 -22568 2212
rect -27940 2132 -22568 2148
rect -27940 2068 -22652 2132
rect -22588 2068 -22568 2132
rect -27940 2052 -22568 2068
rect -27940 1988 -22652 2052
rect -22588 1988 -22568 2052
rect -27940 1972 -22568 1988
rect -27940 1908 -22652 1972
rect -22588 1908 -22568 1972
rect -27940 1892 -22568 1908
rect -27940 1828 -22652 1892
rect -22588 1828 -22568 1892
rect -27940 1812 -22568 1828
rect -27940 1748 -22652 1812
rect -22588 1748 -22568 1812
rect -27940 1732 -22568 1748
rect -27940 1668 -22652 1732
rect -22588 1668 -22568 1732
rect -27940 1652 -22568 1668
rect -27940 1588 -22652 1652
rect -22588 1588 -22568 1652
rect -27940 1572 -22568 1588
rect -27940 1508 -22652 1572
rect -22588 1508 -22568 1572
rect -27940 1492 -22568 1508
rect -27940 1428 -22652 1492
rect -22588 1428 -22568 1492
rect -27940 1412 -22568 1428
rect -27940 1348 -22652 1412
rect -22588 1348 -22568 1412
rect -27940 1332 -22568 1348
rect -27940 1268 -22652 1332
rect -22588 1268 -22568 1332
rect -27940 1252 -22568 1268
rect -27940 1188 -22652 1252
rect -22588 1188 -22568 1252
rect -27940 1172 -22568 1188
rect -27940 1108 -22652 1172
rect -22588 1108 -22568 1172
rect -27940 1092 -22568 1108
rect -27940 1028 -22652 1092
rect -22588 1028 -22568 1092
rect -27940 1012 -22568 1028
rect -27940 948 -22652 1012
rect -22588 948 -22568 1012
rect -27940 932 -22568 948
rect -27940 868 -22652 932
rect -22588 868 -22568 932
rect -27940 852 -22568 868
rect -27940 788 -22652 852
rect -22588 788 -22568 852
rect -27940 772 -22568 788
rect -27940 708 -22652 772
rect -22588 708 -22568 772
rect -27940 692 -22568 708
rect -27940 628 -22652 692
rect -22588 628 -22568 692
rect -27940 612 -22568 628
rect -27940 548 -22652 612
rect -22588 548 -22568 612
rect -27940 532 -22568 548
rect -27940 468 -22652 532
rect -22588 468 -22568 532
rect -27940 452 -22568 468
rect -27940 388 -22652 452
rect -22588 388 -22568 452
rect -27940 372 -22568 388
rect -27940 308 -22652 372
rect -22588 308 -22568 372
rect -27940 292 -22568 308
rect -27940 228 -22652 292
rect -22588 228 -22568 292
rect -27940 212 -22568 228
rect -27940 148 -22652 212
rect -22588 148 -22568 212
rect -27940 120 -22568 148
rect -22328 5172 -16956 5200
rect -22328 5108 -17040 5172
rect -16976 5108 -16956 5172
rect -22328 5092 -16956 5108
rect -22328 5028 -17040 5092
rect -16976 5028 -16956 5092
rect -22328 5012 -16956 5028
rect -22328 4948 -17040 5012
rect -16976 4948 -16956 5012
rect -22328 4932 -16956 4948
rect -22328 4868 -17040 4932
rect -16976 4868 -16956 4932
rect -22328 4852 -16956 4868
rect -22328 4788 -17040 4852
rect -16976 4788 -16956 4852
rect -22328 4772 -16956 4788
rect -22328 4708 -17040 4772
rect -16976 4708 -16956 4772
rect -22328 4692 -16956 4708
rect -22328 4628 -17040 4692
rect -16976 4628 -16956 4692
rect -22328 4612 -16956 4628
rect -22328 4548 -17040 4612
rect -16976 4548 -16956 4612
rect -22328 4532 -16956 4548
rect -22328 4468 -17040 4532
rect -16976 4468 -16956 4532
rect -22328 4452 -16956 4468
rect -22328 4388 -17040 4452
rect -16976 4388 -16956 4452
rect -22328 4372 -16956 4388
rect -22328 4308 -17040 4372
rect -16976 4308 -16956 4372
rect -22328 4292 -16956 4308
rect -22328 4228 -17040 4292
rect -16976 4228 -16956 4292
rect -22328 4212 -16956 4228
rect -22328 4148 -17040 4212
rect -16976 4148 -16956 4212
rect -22328 4132 -16956 4148
rect -22328 4068 -17040 4132
rect -16976 4068 -16956 4132
rect -22328 4052 -16956 4068
rect -22328 3988 -17040 4052
rect -16976 3988 -16956 4052
rect -22328 3972 -16956 3988
rect -22328 3908 -17040 3972
rect -16976 3908 -16956 3972
rect -22328 3892 -16956 3908
rect -22328 3828 -17040 3892
rect -16976 3828 -16956 3892
rect -22328 3812 -16956 3828
rect -22328 3748 -17040 3812
rect -16976 3748 -16956 3812
rect -22328 3732 -16956 3748
rect -22328 3668 -17040 3732
rect -16976 3668 -16956 3732
rect -22328 3652 -16956 3668
rect -22328 3588 -17040 3652
rect -16976 3588 -16956 3652
rect -22328 3572 -16956 3588
rect -22328 3508 -17040 3572
rect -16976 3508 -16956 3572
rect -22328 3492 -16956 3508
rect -22328 3428 -17040 3492
rect -16976 3428 -16956 3492
rect -22328 3412 -16956 3428
rect -22328 3348 -17040 3412
rect -16976 3348 -16956 3412
rect -22328 3332 -16956 3348
rect -22328 3268 -17040 3332
rect -16976 3268 -16956 3332
rect -22328 3252 -16956 3268
rect -22328 3188 -17040 3252
rect -16976 3188 -16956 3252
rect -22328 3172 -16956 3188
rect -22328 3108 -17040 3172
rect -16976 3108 -16956 3172
rect -22328 3092 -16956 3108
rect -22328 3028 -17040 3092
rect -16976 3028 -16956 3092
rect -22328 3012 -16956 3028
rect -22328 2948 -17040 3012
rect -16976 2948 -16956 3012
rect -22328 2932 -16956 2948
rect -22328 2868 -17040 2932
rect -16976 2868 -16956 2932
rect -22328 2852 -16956 2868
rect -22328 2788 -17040 2852
rect -16976 2788 -16956 2852
rect -22328 2772 -16956 2788
rect -22328 2708 -17040 2772
rect -16976 2708 -16956 2772
rect -22328 2692 -16956 2708
rect -22328 2628 -17040 2692
rect -16976 2628 -16956 2692
rect -22328 2612 -16956 2628
rect -22328 2548 -17040 2612
rect -16976 2548 -16956 2612
rect -22328 2532 -16956 2548
rect -22328 2468 -17040 2532
rect -16976 2468 -16956 2532
rect -22328 2452 -16956 2468
rect -22328 2388 -17040 2452
rect -16976 2388 -16956 2452
rect -22328 2372 -16956 2388
rect -22328 2308 -17040 2372
rect -16976 2308 -16956 2372
rect -22328 2292 -16956 2308
rect -22328 2228 -17040 2292
rect -16976 2228 -16956 2292
rect -22328 2212 -16956 2228
rect -22328 2148 -17040 2212
rect -16976 2148 -16956 2212
rect -22328 2132 -16956 2148
rect -22328 2068 -17040 2132
rect -16976 2068 -16956 2132
rect -22328 2052 -16956 2068
rect -22328 1988 -17040 2052
rect -16976 1988 -16956 2052
rect -22328 1972 -16956 1988
rect -22328 1908 -17040 1972
rect -16976 1908 -16956 1972
rect -22328 1892 -16956 1908
rect -22328 1828 -17040 1892
rect -16976 1828 -16956 1892
rect -22328 1812 -16956 1828
rect -22328 1748 -17040 1812
rect -16976 1748 -16956 1812
rect -22328 1732 -16956 1748
rect -22328 1668 -17040 1732
rect -16976 1668 -16956 1732
rect -22328 1652 -16956 1668
rect -22328 1588 -17040 1652
rect -16976 1588 -16956 1652
rect -22328 1572 -16956 1588
rect -22328 1508 -17040 1572
rect -16976 1508 -16956 1572
rect -22328 1492 -16956 1508
rect -22328 1428 -17040 1492
rect -16976 1428 -16956 1492
rect -22328 1412 -16956 1428
rect -22328 1348 -17040 1412
rect -16976 1348 -16956 1412
rect -22328 1332 -16956 1348
rect -22328 1268 -17040 1332
rect -16976 1268 -16956 1332
rect -22328 1252 -16956 1268
rect -22328 1188 -17040 1252
rect -16976 1188 -16956 1252
rect -22328 1172 -16956 1188
rect -22328 1108 -17040 1172
rect -16976 1108 -16956 1172
rect -22328 1092 -16956 1108
rect -22328 1028 -17040 1092
rect -16976 1028 -16956 1092
rect -22328 1012 -16956 1028
rect -22328 948 -17040 1012
rect -16976 948 -16956 1012
rect -22328 932 -16956 948
rect -22328 868 -17040 932
rect -16976 868 -16956 932
rect -22328 852 -16956 868
rect -22328 788 -17040 852
rect -16976 788 -16956 852
rect -22328 772 -16956 788
rect -22328 708 -17040 772
rect -16976 708 -16956 772
rect -22328 692 -16956 708
rect -22328 628 -17040 692
rect -16976 628 -16956 692
rect -22328 612 -16956 628
rect -22328 548 -17040 612
rect -16976 548 -16956 612
rect -22328 532 -16956 548
rect -22328 468 -17040 532
rect -16976 468 -16956 532
rect -22328 452 -16956 468
rect -22328 388 -17040 452
rect -16976 388 -16956 452
rect -22328 372 -16956 388
rect -22328 308 -17040 372
rect -16976 308 -16956 372
rect -22328 292 -16956 308
rect -22328 228 -17040 292
rect -16976 228 -16956 292
rect -22328 212 -16956 228
rect -22328 148 -17040 212
rect -16976 148 -16956 212
rect -22328 120 -16956 148
rect -16716 5172 -11344 5200
rect -16716 5108 -11428 5172
rect -11364 5108 -11344 5172
rect -16716 5092 -11344 5108
rect -16716 5028 -11428 5092
rect -11364 5028 -11344 5092
rect -16716 5012 -11344 5028
rect -16716 4948 -11428 5012
rect -11364 4948 -11344 5012
rect -16716 4932 -11344 4948
rect -16716 4868 -11428 4932
rect -11364 4868 -11344 4932
rect -16716 4852 -11344 4868
rect -16716 4788 -11428 4852
rect -11364 4788 -11344 4852
rect -16716 4772 -11344 4788
rect -16716 4708 -11428 4772
rect -11364 4708 -11344 4772
rect -16716 4692 -11344 4708
rect -16716 4628 -11428 4692
rect -11364 4628 -11344 4692
rect -16716 4612 -11344 4628
rect -16716 4548 -11428 4612
rect -11364 4548 -11344 4612
rect -16716 4532 -11344 4548
rect -16716 4468 -11428 4532
rect -11364 4468 -11344 4532
rect -16716 4452 -11344 4468
rect -16716 4388 -11428 4452
rect -11364 4388 -11344 4452
rect -16716 4372 -11344 4388
rect -16716 4308 -11428 4372
rect -11364 4308 -11344 4372
rect -16716 4292 -11344 4308
rect -16716 4228 -11428 4292
rect -11364 4228 -11344 4292
rect -16716 4212 -11344 4228
rect -16716 4148 -11428 4212
rect -11364 4148 -11344 4212
rect -16716 4132 -11344 4148
rect -16716 4068 -11428 4132
rect -11364 4068 -11344 4132
rect -16716 4052 -11344 4068
rect -16716 3988 -11428 4052
rect -11364 3988 -11344 4052
rect -16716 3972 -11344 3988
rect -16716 3908 -11428 3972
rect -11364 3908 -11344 3972
rect -16716 3892 -11344 3908
rect -16716 3828 -11428 3892
rect -11364 3828 -11344 3892
rect -16716 3812 -11344 3828
rect -16716 3748 -11428 3812
rect -11364 3748 -11344 3812
rect -16716 3732 -11344 3748
rect -16716 3668 -11428 3732
rect -11364 3668 -11344 3732
rect -16716 3652 -11344 3668
rect -16716 3588 -11428 3652
rect -11364 3588 -11344 3652
rect -16716 3572 -11344 3588
rect -16716 3508 -11428 3572
rect -11364 3508 -11344 3572
rect -16716 3492 -11344 3508
rect -16716 3428 -11428 3492
rect -11364 3428 -11344 3492
rect -16716 3412 -11344 3428
rect -16716 3348 -11428 3412
rect -11364 3348 -11344 3412
rect -16716 3332 -11344 3348
rect -16716 3268 -11428 3332
rect -11364 3268 -11344 3332
rect -16716 3252 -11344 3268
rect -16716 3188 -11428 3252
rect -11364 3188 -11344 3252
rect -16716 3172 -11344 3188
rect -16716 3108 -11428 3172
rect -11364 3108 -11344 3172
rect -16716 3092 -11344 3108
rect -16716 3028 -11428 3092
rect -11364 3028 -11344 3092
rect -16716 3012 -11344 3028
rect -16716 2948 -11428 3012
rect -11364 2948 -11344 3012
rect -16716 2932 -11344 2948
rect -16716 2868 -11428 2932
rect -11364 2868 -11344 2932
rect -16716 2852 -11344 2868
rect -16716 2788 -11428 2852
rect -11364 2788 -11344 2852
rect -16716 2772 -11344 2788
rect -16716 2708 -11428 2772
rect -11364 2708 -11344 2772
rect -16716 2692 -11344 2708
rect -16716 2628 -11428 2692
rect -11364 2628 -11344 2692
rect -16716 2612 -11344 2628
rect -16716 2548 -11428 2612
rect -11364 2548 -11344 2612
rect -16716 2532 -11344 2548
rect -16716 2468 -11428 2532
rect -11364 2468 -11344 2532
rect -16716 2452 -11344 2468
rect -16716 2388 -11428 2452
rect -11364 2388 -11344 2452
rect -16716 2372 -11344 2388
rect -16716 2308 -11428 2372
rect -11364 2308 -11344 2372
rect -16716 2292 -11344 2308
rect -16716 2228 -11428 2292
rect -11364 2228 -11344 2292
rect -16716 2212 -11344 2228
rect -16716 2148 -11428 2212
rect -11364 2148 -11344 2212
rect -16716 2132 -11344 2148
rect -16716 2068 -11428 2132
rect -11364 2068 -11344 2132
rect -16716 2052 -11344 2068
rect -16716 1988 -11428 2052
rect -11364 1988 -11344 2052
rect -16716 1972 -11344 1988
rect -16716 1908 -11428 1972
rect -11364 1908 -11344 1972
rect -16716 1892 -11344 1908
rect -16716 1828 -11428 1892
rect -11364 1828 -11344 1892
rect -16716 1812 -11344 1828
rect -16716 1748 -11428 1812
rect -11364 1748 -11344 1812
rect -16716 1732 -11344 1748
rect -16716 1668 -11428 1732
rect -11364 1668 -11344 1732
rect -16716 1652 -11344 1668
rect -16716 1588 -11428 1652
rect -11364 1588 -11344 1652
rect -16716 1572 -11344 1588
rect -16716 1508 -11428 1572
rect -11364 1508 -11344 1572
rect -16716 1492 -11344 1508
rect -16716 1428 -11428 1492
rect -11364 1428 -11344 1492
rect -16716 1412 -11344 1428
rect -16716 1348 -11428 1412
rect -11364 1348 -11344 1412
rect -16716 1332 -11344 1348
rect -16716 1268 -11428 1332
rect -11364 1268 -11344 1332
rect -16716 1252 -11344 1268
rect -16716 1188 -11428 1252
rect -11364 1188 -11344 1252
rect -16716 1172 -11344 1188
rect -16716 1108 -11428 1172
rect -11364 1108 -11344 1172
rect -16716 1092 -11344 1108
rect -16716 1028 -11428 1092
rect -11364 1028 -11344 1092
rect -16716 1012 -11344 1028
rect -16716 948 -11428 1012
rect -11364 948 -11344 1012
rect -16716 932 -11344 948
rect -16716 868 -11428 932
rect -11364 868 -11344 932
rect -16716 852 -11344 868
rect -16716 788 -11428 852
rect -11364 788 -11344 852
rect -16716 772 -11344 788
rect -16716 708 -11428 772
rect -11364 708 -11344 772
rect -16716 692 -11344 708
rect -16716 628 -11428 692
rect -11364 628 -11344 692
rect -16716 612 -11344 628
rect -16716 548 -11428 612
rect -11364 548 -11344 612
rect -16716 532 -11344 548
rect -16716 468 -11428 532
rect -11364 468 -11344 532
rect -16716 452 -11344 468
rect -16716 388 -11428 452
rect -11364 388 -11344 452
rect -16716 372 -11344 388
rect -16716 308 -11428 372
rect -11364 308 -11344 372
rect -16716 292 -11344 308
rect -16716 228 -11428 292
rect -11364 228 -11344 292
rect -16716 212 -11344 228
rect -16716 148 -11428 212
rect -11364 148 -11344 212
rect -16716 120 -11344 148
rect -11104 5172 -5732 5200
rect -11104 5108 -5816 5172
rect -5752 5108 -5732 5172
rect -11104 5092 -5732 5108
rect -11104 5028 -5816 5092
rect -5752 5028 -5732 5092
rect -11104 5012 -5732 5028
rect -11104 4948 -5816 5012
rect -5752 4948 -5732 5012
rect -11104 4932 -5732 4948
rect -11104 4868 -5816 4932
rect -5752 4868 -5732 4932
rect -11104 4852 -5732 4868
rect -11104 4788 -5816 4852
rect -5752 4788 -5732 4852
rect -11104 4772 -5732 4788
rect -11104 4708 -5816 4772
rect -5752 4708 -5732 4772
rect -11104 4692 -5732 4708
rect -11104 4628 -5816 4692
rect -5752 4628 -5732 4692
rect -11104 4612 -5732 4628
rect -11104 4548 -5816 4612
rect -5752 4548 -5732 4612
rect -11104 4532 -5732 4548
rect -11104 4468 -5816 4532
rect -5752 4468 -5732 4532
rect -11104 4452 -5732 4468
rect -11104 4388 -5816 4452
rect -5752 4388 -5732 4452
rect -11104 4372 -5732 4388
rect -11104 4308 -5816 4372
rect -5752 4308 -5732 4372
rect -11104 4292 -5732 4308
rect -11104 4228 -5816 4292
rect -5752 4228 -5732 4292
rect -11104 4212 -5732 4228
rect -11104 4148 -5816 4212
rect -5752 4148 -5732 4212
rect -11104 4132 -5732 4148
rect -11104 4068 -5816 4132
rect -5752 4068 -5732 4132
rect -11104 4052 -5732 4068
rect -11104 3988 -5816 4052
rect -5752 3988 -5732 4052
rect -11104 3972 -5732 3988
rect -11104 3908 -5816 3972
rect -5752 3908 -5732 3972
rect -11104 3892 -5732 3908
rect -11104 3828 -5816 3892
rect -5752 3828 -5732 3892
rect -11104 3812 -5732 3828
rect -11104 3748 -5816 3812
rect -5752 3748 -5732 3812
rect -11104 3732 -5732 3748
rect -11104 3668 -5816 3732
rect -5752 3668 -5732 3732
rect -11104 3652 -5732 3668
rect -11104 3588 -5816 3652
rect -5752 3588 -5732 3652
rect -11104 3572 -5732 3588
rect -11104 3508 -5816 3572
rect -5752 3508 -5732 3572
rect -11104 3492 -5732 3508
rect -11104 3428 -5816 3492
rect -5752 3428 -5732 3492
rect -11104 3412 -5732 3428
rect -11104 3348 -5816 3412
rect -5752 3348 -5732 3412
rect -11104 3332 -5732 3348
rect -11104 3268 -5816 3332
rect -5752 3268 -5732 3332
rect -11104 3252 -5732 3268
rect -11104 3188 -5816 3252
rect -5752 3188 -5732 3252
rect -11104 3172 -5732 3188
rect -11104 3108 -5816 3172
rect -5752 3108 -5732 3172
rect -11104 3092 -5732 3108
rect -11104 3028 -5816 3092
rect -5752 3028 -5732 3092
rect -11104 3012 -5732 3028
rect -11104 2948 -5816 3012
rect -5752 2948 -5732 3012
rect -11104 2932 -5732 2948
rect -11104 2868 -5816 2932
rect -5752 2868 -5732 2932
rect -11104 2852 -5732 2868
rect -11104 2788 -5816 2852
rect -5752 2788 -5732 2852
rect -11104 2772 -5732 2788
rect -11104 2708 -5816 2772
rect -5752 2708 -5732 2772
rect -11104 2692 -5732 2708
rect -11104 2628 -5816 2692
rect -5752 2628 -5732 2692
rect -11104 2612 -5732 2628
rect -11104 2548 -5816 2612
rect -5752 2548 -5732 2612
rect -11104 2532 -5732 2548
rect -11104 2468 -5816 2532
rect -5752 2468 -5732 2532
rect -11104 2452 -5732 2468
rect -11104 2388 -5816 2452
rect -5752 2388 -5732 2452
rect -11104 2372 -5732 2388
rect -11104 2308 -5816 2372
rect -5752 2308 -5732 2372
rect -11104 2292 -5732 2308
rect -11104 2228 -5816 2292
rect -5752 2228 -5732 2292
rect -11104 2212 -5732 2228
rect -11104 2148 -5816 2212
rect -5752 2148 -5732 2212
rect -11104 2132 -5732 2148
rect -11104 2068 -5816 2132
rect -5752 2068 -5732 2132
rect -11104 2052 -5732 2068
rect -11104 1988 -5816 2052
rect -5752 1988 -5732 2052
rect -11104 1972 -5732 1988
rect -11104 1908 -5816 1972
rect -5752 1908 -5732 1972
rect -11104 1892 -5732 1908
rect -11104 1828 -5816 1892
rect -5752 1828 -5732 1892
rect -11104 1812 -5732 1828
rect -11104 1748 -5816 1812
rect -5752 1748 -5732 1812
rect -11104 1732 -5732 1748
rect -11104 1668 -5816 1732
rect -5752 1668 -5732 1732
rect -11104 1652 -5732 1668
rect -11104 1588 -5816 1652
rect -5752 1588 -5732 1652
rect -11104 1572 -5732 1588
rect -11104 1508 -5816 1572
rect -5752 1508 -5732 1572
rect -11104 1492 -5732 1508
rect -11104 1428 -5816 1492
rect -5752 1428 -5732 1492
rect -11104 1412 -5732 1428
rect -11104 1348 -5816 1412
rect -5752 1348 -5732 1412
rect -11104 1332 -5732 1348
rect -11104 1268 -5816 1332
rect -5752 1268 -5732 1332
rect -11104 1252 -5732 1268
rect -11104 1188 -5816 1252
rect -5752 1188 -5732 1252
rect -11104 1172 -5732 1188
rect -11104 1108 -5816 1172
rect -5752 1108 -5732 1172
rect -11104 1092 -5732 1108
rect -11104 1028 -5816 1092
rect -5752 1028 -5732 1092
rect -11104 1012 -5732 1028
rect -11104 948 -5816 1012
rect -5752 948 -5732 1012
rect -11104 932 -5732 948
rect -11104 868 -5816 932
rect -5752 868 -5732 932
rect -11104 852 -5732 868
rect -11104 788 -5816 852
rect -5752 788 -5732 852
rect -11104 772 -5732 788
rect -11104 708 -5816 772
rect -5752 708 -5732 772
rect -11104 692 -5732 708
rect -11104 628 -5816 692
rect -5752 628 -5732 692
rect -11104 612 -5732 628
rect -11104 548 -5816 612
rect -5752 548 -5732 612
rect -11104 532 -5732 548
rect -11104 468 -5816 532
rect -5752 468 -5732 532
rect -11104 452 -5732 468
rect -11104 388 -5816 452
rect -5752 388 -5732 452
rect -11104 372 -5732 388
rect -11104 308 -5816 372
rect -5752 308 -5732 372
rect -11104 292 -5732 308
rect -11104 228 -5816 292
rect -5752 228 -5732 292
rect -11104 212 -5732 228
rect -11104 148 -5816 212
rect -5752 148 -5732 212
rect -11104 120 -5732 148
rect -5492 5172 -120 5200
rect -5492 5108 -204 5172
rect -140 5108 -120 5172
rect -5492 5092 -120 5108
rect -5492 5028 -204 5092
rect -140 5028 -120 5092
rect -5492 5012 -120 5028
rect -5492 4948 -204 5012
rect -140 4948 -120 5012
rect -5492 4932 -120 4948
rect -5492 4868 -204 4932
rect -140 4868 -120 4932
rect -5492 4852 -120 4868
rect -5492 4788 -204 4852
rect -140 4788 -120 4852
rect -5492 4772 -120 4788
rect -5492 4708 -204 4772
rect -140 4708 -120 4772
rect -5492 4692 -120 4708
rect -5492 4628 -204 4692
rect -140 4628 -120 4692
rect -5492 4612 -120 4628
rect -5492 4548 -204 4612
rect -140 4548 -120 4612
rect -5492 4532 -120 4548
rect -5492 4468 -204 4532
rect -140 4468 -120 4532
rect -5492 4452 -120 4468
rect -5492 4388 -204 4452
rect -140 4388 -120 4452
rect -5492 4372 -120 4388
rect -5492 4308 -204 4372
rect -140 4308 -120 4372
rect -5492 4292 -120 4308
rect -5492 4228 -204 4292
rect -140 4228 -120 4292
rect -5492 4212 -120 4228
rect -5492 4148 -204 4212
rect -140 4148 -120 4212
rect -5492 4132 -120 4148
rect -5492 4068 -204 4132
rect -140 4068 -120 4132
rect -5492 4052 -120 4068
rect -5492 3988 -204 4052
rect -140 3988 -120 4052
rect -5492 3972 -120 3988
rect -5492 3908 -204 3972
rect -140 3908 -120 3972
rect -5492 3892 -120 3908
rect -5492 3828 -204 3892
rect -140 3828 -120 3892
rect -5492 3812 -120 3828
rect -5492 3748 -204 3812
rect -140 3748 -120 3812
rect -5492 3732 -120 3748
rect -5492 3668 -204 3732
rect -140 3668 -120 3732
rect -5492 3652 -120 3668
rect -5492 3588 -204 3652
rect -140 3588 -120 3652
rect -5492 3572 -120 3588
rect -5492 3508 -204 3572
rect -140 3508 -120 3572
rect -5492 3492 -120 3508
rect -5492 3428 -204 3492
rect -140 3428 -120 3492
rect -5492 3412 -120 3428
rect -5492 3348 -204 3412
rect -140 3348 -120 3412
rect -5492 3332 -120 3348
rect -5492 3268 -204 3332
rect -140 3268 -120 3332
rect -5492 3252 -120 3268
rect -5492 3188 -204 3252
rect -140 3188 -120 3252
rect -5492 3172 -120 3188
rect -5492 3108 -204 3172
rect -140 3108 -120 3172
rect -5492 3092 -120 3108
rect -5492 3028 -204 3092
rect -140 3028 -120 3092
rect -5492 3012 -120 3028
rect -5492 2948 -204 3012
rect -140 2948 -120 3012
rect -5492 2932 -120 2948
rect -5492 2868 -204 2932
rect -140 2868 -120 2932
rect -5492 2852 -120 2868
rect -5492 2788 -204 2852
rect -140 2788 -120 2852
rect -5492 2772 -120 2788
rect -5492 2708 -204 2772
rect -140 2708 -120 2772
rect -5492 2692 -120 2708
rect -5492 2628 -204 2692
rect -140 2628 -120 2692
rect -5492 2612 -120 2628
rect -5492 2548 -204 2612
rect -140 2548 -120 2612
rect -5492 2532 -120 2548
rect -5492 2468 -204 2532
rect -140 2468 -120 2532
rect -5492 2452 -120 2468
rect -5492 2388 -204 2452
rect -140 2388 -120 2452
rect -5492 2372 -120 2388
rect -5492 2308 -204 2372
rect -140 2308 -120 2372
rect -5492 2292 -120 2308
rect -5492 2228 -204 2292
rect -140 2228 -120 2292
rect -5492 2212 -120 2228
rect -5492 2148 -204 2212
rect -140 2148 -120 2212
rect -5492 2132 -120 2148
rect -5492 2068 -204 2132
rect -140 2068 -120 2132
rect -5492 2052 -120 2068
rect -5492 1988 -204 2052
rect -140 1988 -120 2052
rect -5492 1972 -120 1988
rect -5492 1908 -204 1972
rect -140 1908 -120 1972
rect -5492 1892 -120 1908
rect -5492 1828 -204 1892
rect -140 1828 -120 1892
rect -5492 1812 -120 1828
rect -5492 1748 -204 1812
rect -140 1748 -120 1812
rect -5492 1732 -120 1748
rect -5492 1668 -204 1732
rect -140 1668 -120 1732
rect -5492 1652 -120 1668
rect -5492 1588 -204 1652
rect -140 1588 -120 1652
rect -5492 1572 -120 1588
rect -5492 1508 -204 1572
rect -140 1508 -120 1572
rect -5492 1492 -120 1508
rect -5492 1428 -204 1492
rect -140 1428 -120 1492
rect -5492 1412 -120 1428
rect -5492 1348 -204 1412
rect -140 1348 -120 1412
rect -5492 1332 -120 1348
rect -5492 1268 -204 1332
rect -140 1268 -120 1332
rect -5492 1252 -120 1268
rect -5492 1188 -204 1252
rect -140 1188 -120 1252
rect -5492 1172 -120 1188
rect -5492 1108 -204 1172
rect -140 1108 -120 1172
rect -5492 1092 -120 1108
rect -5492 1028 -204 1092
rect -140 1028 -120 1092
rect -5492 1012 -120 1028
rect -5492 948 -204 1012
rect -140 948 -120 1012
rect -5492 932 -120 948
rect -5492 868 -204 932
rect -140 868 -120 932
rect -5492 852 -120 868
rect -5492 788 -204 852
rect -140 788 -120 852
rect -5492 772 -120 788
rect -5492 708 -204 772
rect -140 708 -120 772
rect -5492 692 -120 708
rect -5492 628 -204 692
rect -140 628 -120 692
rect -5492 612 -120 628
rect -5492 548 -204 612
rect -140 548 -120 612
rect -5492 532 -120 548
rect -5492 468 -204 532
rect -140 468 -120 532
rect -5492 452 -120 468
rect -5492 388 -204 452
rect -140 388 -120 452
rect -5492 372 -120 388
rect -5492 308 -204 372
rect -140 308 -120 372
rect -5492 292 -120 308
rect -5492 228 -204 292
rect -140 228 -120 292
rect -5492 212 -120 228
rect -5492 148 -204 212
rect -140 148 -120 212
rect -5492 120 -120 148
rect 120 5172 5492 5200
rect 120 5108 5408 5172
rect 5472 5108 5492 5172
rect 120 5092 5492 5108
rect 120 5028 5408 5092
rect 5472 5028 5492 5092
rect 120 5012 5492 5028
rect 120 4948 5408 5012
rect 5472 4948 5492 5012
rect 120 4932 5492 4948
rect 120 4868 5408 4932
rect 5472 4868 5492 4932
rect 120 4852 5492 4868
rect 120 4788 5408 4852
rect 5472 4788 5492 4852
rect 120 4772 5492 4788
rect 120 4708 5408 4772
rect 5472 4708 5492 4772
rect 120 4692 5492 4708
rect 120 4628 5408 4692
rect 5472 4628 5492 4692
rect 120 4612 5492 4628
rect 120 4548 5408 4612
rect 5472 4548 5492 4612
rect 120 4532 5492 4548
rect 120 4468 5408 4532
rect 5472 4468 5492 4532
rect 120 4452 5492 4468
rect 120 4388 5408 4452
rect 5472 4388 5492 4452
rect 120 4372 5492 4388
rect 120 4308 5408 4372
rect 5472 4308 5492 4372
rect 120 4292 5492 4308
rect 120 4228 5408 4292
rect 5472 4228 5492 4292
rect 120 4212 5492 4228
rect 120 4148 5408 4212
rect 5472 4148 5492 4212
rect 120 4132 5492 4148
rect 120 4068 5408 4132
rect 5472 4068 5492 4132
rect 120 4052 5492 4068
rect 120 3988 5408 4052
rect 5472 3988 5492 4052
rect 120 3972 5492 3988
rect 120 3908 5408 3972
rect 5472 3908 5492 3972
rect 120 3892 5492 3908
rect 120 3828 5408 3892
rect 5472 3828 5492 3892
rect 120 3812 5492 3828
rect 120 3748 5408 3812
rect 5472 3748 5492 3812
rect 120 3732 5492 3748
rect 120 3668 5408 3732
rect 5472 3668 5492 3732
rect 120 3652 5492 3668
rect 120 3588 5408 3652
rect 5472 3588 5492 3652
rect 120 3572 5492 3588
rect 120 3508 5408 3572
rect 5472 3508 5492 3572
rect 120 3492 5492 3508
rect 120 3428 5408 3492
rect 5472 3428 5492 3492
rect 120 3412 5492 3428
rect 120 3348 5408 3412
rect 5472 3348 5492 3412
rect 120 3332 5492 3348
rect 120 3268 5408 3332
rect 5472 3268 5492 3332
rect 120 3252 5492 3268
rect 120 3188 5408 3252
rect 5472 3188 5492 3252
rect 120 3172 5492 3188
rect 120 3108 5408 3172
rect 5472 3108 5492 3172
rect 120 3092 5492 3108
rect 120 3028 5408 3092
rect 5472 3028 5492 3092
rect 120 3012 5492 3028
rect 120 2948 5408 3012
rect 5472 2948 5492 3012
rect 120 2932 5492 2948
rect 120 2868 5408 2932
rect 5472 2868 5492 2932
rect 120 2852 5492 2868
rect 120 2788 5408 2852
rect 5472 2788 5492 2852
rect 120 2772 5492 2788
rect 120 2708 5408 2772
rect 5472 2708 5492 2772
rect 120 2692 5492 2708
rect 120 2628 5408 2692
rect 5472 2628 5492 2692
rect 120 2612 5492 2628
rect 120 2548 5408 2612
rect 5472 2548 5492 2612
rect 120 2532 5492 2548
rect 120 2468 5408 2532
rect 5472 2468 5492 2532
rect 120 2452 5492 2468
rect 120 2388 5408 2452
rect 5472 2388 5492 2452
rect 120 2372 5492 2388
rect 120 2308 5408 2372
rect 5472 2308 5492 2372
rect 120 2292 5492 2308
rect 120 2228 5408 2292
rect 5472 2228 5492 2292
rect 120 2212 5492 2228
rect 120 2148 5408 2212
rect 5472 2148 5492 2212
rect 120 2132 5492 2148
rect 120 2068 5408 2132
rect 5472 2068 5492 2132
rect 120 2052 5492 2068
rect 120 1988 5408 2052
rect 5472 1988 5492 2052
rect 120 1972 5492 1988
rect 120 1908 5408 1972
rect 5472 1908 5492 1972
rect 120 1892 5492 1908
rect 120 1828 5408 1892
rect 5472 1828 5492 1892
rect 120 1812 5492 1828
rect 120 1748 5408 1812
rect 5472 1748 5492 1812
rect 120 1732 5492 1748
rect 120 1668 5408 1732
rect 5472 1668 5492 1732
rect 120 1652 5492 1668
rect 120 1588 5408 1652
rect 5472 1588 5492 1652
rect 120 1572 5492 1588
rect 120 1508 5408 1572
rect 5472 1508 5492 1572
rect 120 1492 5492 1508
rect 120 1428 5408 1492
rect 5472 1428 5492 1492
rect 120 1412 5492 1428
rect 120 1348 5408 1412
rect 5472 1348 5492 1412
rect 120 1332 5492 1348
rect 120 1268 5408 1332
rect 5472 1268 5492 1332
rect 120 1252 5492 1268
rect 120 1188 5408 1252
rect 5472 1188 5492 1252
rect 120 1172 5492 1188
rect 120 1108 5408 1172
rect 5472 1108 5492 1172
rect 120 1092 5492 1108
rect 120 1028 5408 1092
rect 5472 1028 5492 1092
rect 120 1012 5492 1028
rect 120 948 5408 1012
rect 5472 948 5492 1012
rect 120 932 5492 948
rect 120 868 5408 932
rect 5472 868 5492 932
rect 120 852 5492 868
rect 120 788 5408 852
rect 5472 788 5492 852
rect 120 772 5492 788
rect 120 708 5408 772
rect 5472 708 5492 772
rect 120 692 5492 708
rect 120 628 5408 692
rect 5472 628 5492 692
rect 120 612 5492 628
rect 120 548 5408 612
rect 5472 548 5492 612
rect 120 532 5492 548
rect 120 468 5408 532
rect 5472 468 5492 532
rect 120 452 5492 468
rect 120 388 5408 452
rect 5472 388 5492 452
rect 120 372 5492 388
rect 120 308 5408 372
rect 5472 308 5492 372
rect 120 292 5492 308
rect 120 228 5408 292
rect 5472 228 5492 292
rect 120 212 5492 228
rect 120 148 5408 212
rect 5472 148 5492 212
rect 120 120 5492 148
rect 5732 5172 11104 5200
rect 5732 5108 11020 5172
rect 11084 5108 11104 5172
rect 5732 5092 11104 5108
rect 5732 5028 11020 5092
rect 11084 5028 11104 5092
rect 5732 5012 11104 5028
rect 5732 4948 11020 5012
rect 11084 4948 11104 5012
rect 5732 4932 11104 4948
rect 5732 4868 11020 4932
rect 11084 4868 11104 4932
rect 5732 4852 11104 4868
rect 5732 4788 11020 4852
rect 11084 4788 11104 4852
rect 5732 4772 11104 4788
rect 5732 4708 11020 4772
rect 11084 4708 11104 4772
rect 5732 4692 11104 4708
rect 5732 4628 11020 4692
rect 11084 4628 11104 4692
rect 5732 4612 11104 4628
rect 5732 4548 11020 4612
rect 11084 4548 11104 4612
rect 5732 4532 11104 4548
rect 5732 4468 11020 4532
rect 11084 4468 11104 4532
rect 5732 4452 11104 4468
rect 5732 4388 11020 4452
rect 11084 4388 11104 4452
rect 5732 4372 11104 4388
rect 5732 4308 11020 4372
rect 11084 4308 11104 4372
rect 5732 4292 11104 4308
rect 5732 4228 11020 4292
rect 11084 4228 11104 4292
rect 5732 4212 11104 4228
rect 5732 4148 11020 4212
rect 11084 4148 11104 4212
rect 5732 4132 11104 4148
rect 5732 4068 11020 4132
rect 11084 4068 11104 4132
rect 5732 4052 11104 4068
rect 5732 3988 11020 4052
rect 11084 3988 11104 4052
rect 5732 3972 11104 3988
rect 5732 3908 11020 3972
rect 11084 3908 11104 3972
rect 5732 3892 11104 3908
rect 5732 3828 11020 3892
rect 11084 3828 11104 3892
rect 5732 3812 11104 3828
rect 5732 3748 11020 3812
rect 11084 3748 11104 3812
rect 5732 3732 11104 3748
rect 5732 3668 11020 3732
rect 11084 3668 11104 3732
rect 5732 3652 11104 3668
rect 5732 3588 11020 3652
rect 11084 3588 11104 3652
rect 5732 3572 11104 3588
rect 5732 3508 11020 3572
rect 11084 3508 11104 3572
rect 5732 3492 11104 3508
rect 5732 3428 11020 3492
rect 11084 3428 11104 3492
rect 5732 3412 11104 3428
rect 5732 3348 11020 3412
rect 11084 3348 11104 3412
rect 5732 3332 11104 3348
rect 5732 3268 11020 3332
rect 11084 3268 11104 3332
rect 5732 3252 11104 3268
rect 5732 3188 11020 3252
rect 11084 3188 11104 3252
rect 5732 3172 11104 3188
rect 5732 3108 11020 3172
rect 11084 3108 11104 3172
rect 5732 3092 11104 3108
rect 5732 3028 11020 3092
rect 11084 3028 11104 3092
rect 5732 3012 11104 3028
rect 5732 2948 11020 3012
rect 11084 2948 11104 3012
rect 5732 2932 11104 2948
rect 5732 2868 11020 2932
rect 11084 2868 11104 2932
rect 5732 2852 11104 2868
rect 5732 2788 11020 2852
rect 11084 2788 11104 2852
rect 5732 2772 11104 2788
rect 5732 2708 11020 2772
rect 11084 2708 11104 2772
rect 5732 2692 11104 2708
rect 5732 2628 11020 2692
rect 11084 2628 11104 2692
rect 5732 2612 11104 2628
rect 5732 2548 11020 2612
rect 11084 2548 11104 2612
rect 5732 2532 11104 2548
rect 5732 2468 11020 2532
rect 11084 2468 11104 2532
rect 5732 2452 11104 2468
rect 5732 2388 11020 2452
rect 11084 2388 11104 2452
rect 5732 2372 11104 2388
rect 5732 2308 11020 2372
rect 11084 2308 11104 2372
rect 5732 2292 11104 2308
rect 5732 2228 11020 2292
rect 11084 2228 11104 2292
rect 5732 2212 11104 2228
rect 5732 2148 11020 2212
rect 11084 2148 11104 2212
rect 5732 2132 11104 2148
rect 5732 2068 11020 2132
rect 11084 2068 11104 2132
rect 5732 2052 11104 2068
rect 5732 1988 11020 2052
rect 11084 1988 11104 2052
rect 5732 1972 11104 1988
rect 5732 1908 11020 1972
rect 11084 1908 11104 1972
rect 5732 1892 11104 1908
rect 5732 1828 11020 1892
rect 11084 1828 11104 1892
rect 5732 1812 11104 1828
rect 5732 1748 11020 1812
rect 11084 1748 11104 1812
rect 5732 1732 11104 1748
rect 5732 1668 11020 1732
rect 11084 1668 11104 1732
rect 5732 1652 11104 1668
rect 5732 1588 11020 1652
rect 11084 1588 11104 1652
rect 5732 1572 11104 1588
rect 5732 1508 11020 1572
rect 11084 1508 11104 1572
rect 5732 1492 11104 1508
rect 5732 1428 11020 1492
rect 11084 1428 11104 1492
rect 5732 1412 11104 1428
rect 5732 1348 11020 1412
rect 11084 1348 11104 1412
rect 5732 1332 11104 1348
rect 5732 1268 11020 1332
rect 11084 1268 11104 1332
rect 5732 1252 11104 1268
rect 5732 1188 11020 1252
rect 11084 1188 11104 1252
rect 5732 1172 11104 1188
rect 5732 1108 11020 1172
rect 11084 1108 11104 1172
rect 5732 1092 11104 1108
rect 5732 1028 11020 1092
rect 11084 1028 11104 1092
rect 5732 1012 11104 1028
rect 5732 948 11020 1012
rect 11084 948 11104 1012
rect 5732 932 11104 948
rect 5732 868 11020 932
rect 11084 868 11104 932
rect 5732 852 11104 868
rect 5732 788 11020 852
rect 11084 788 11104 852
rect 5732 772 11104 788
rect 5732 708 11020 772
rect 11084 708 11104 772
rect 5732 692 11104 708
rect 5732 628 11020 692
rect 11084 628 11104 692
rect 5732 612 11104 628
rect 5732 548 11020 612
rect 11084 548 11104 612
rect 5732 532 11104 548
rect 5732 468 11020 532
rect 11084 468 11104 532
rect 5732 452 11104 468
rect 5732 388 11020 452
rect 11084 388 11104 452
rect 5732 372 11104 388
rect 5732 308 11020 372
rect 11084 308 11104 372
rect 5732 292 11104 308
rect 5732 228 11020 292
rect 11084 228 11104 292
rect 5732 212 11104 228
rect 5732 148 11020 212
rect 11084 148 11104 212
rect 5732 120 11104 148
rect 11344 5172 16716 5200
rect 11344 5108 16632 5172
rect 16696 5108 16716 5172
rect 11344 5092 16716 5108
rect 11344 5028 16632 5092
rect 16696 5028 16716 5092
rect 11344 5012 16716 5028
rect 11344 4948 16632 5012
rect 16696 4948 16716 5012
rect 11344 4932 16716 4948
rect 11344 4868 16632 4932
rect 16696 4868 16716 4932
rect 11344 4852 16716 4868
rect 11344 4788 16632 4852
rect 16696 4788 16716 4852
rect 11344 4772 16716 4788
rect 11344 4708 16632 4772
rect 16696 4708 16716 4772
rect 11344 4692 16716 4708
rect 11344 4628 16632 4692
rect 16696 4628 16716 4692
rect 11344 4612 16716 4628
rect 11344 4548 16632 4612
rect 16696 4548 16716 4612
rect 11344 4532 16716 4548
rect 11344 4468 16632 4532
rect 16696 4468 16716 4532
rect 11344 4452 16716 4468
rect 11344 4388 16632 4452
rect 16696 4388 16716 4452
rect 11344 4372 16716 4388
rect 11344 4308 16632 4372
rect 16696 4308 16716 4372
rect 11344 4292 16716 4308
rect 11344 4228 16632 4292
rect 16696 4228 16716 4292
rect 11344 4212 16716 4228
rect 11344 4148 16632 4212
rect 16696 4148 16716 4212
rect 11344 4132 16716 4148
rect 11344 4068 16632 4132
rect 16696 4068 16716 4132
rect 11344 4052 16716 4068
rect 11344 3988 16632 4052
rect 16696 3988 16716 4052
rect 11344 3972 16716 3988
rect 11344 3908 16632 3972
rect 16696 3908 16716 3972
rect 11344 3892 16716 3908
rect 11344 3828 16632 3892
rect 16696 3828 16716 3892
rect 11344 3812 16716 3828
rect 11344 3748 16632 3812
rect 16696 3748 16716 3812
rect 11344 3732 16716 3748
rect 11344 3668 16632 3732
rect 16696 3668 16716 3732
rect 11344 3652 16716 3668
rect 11344 3588 16632 3652
rect 16696 3588 16716 3652
rect 11344 3572 16716 3588
rect 11344 3508 16632 3572
rect 16696 3508 16716 3572
rect 11344 3492 16716 3508
rect 11344 3428 16632 3492
rect 16696 3428 16716 3492
rect 11344 3412 16716 3428
rect 11344 3348 16632 3412
rect 16696 3348 16716 3412
rect 11344 3332 16716 3348
rect 11344 3268 16632 3332
rect 16696 3268 16716 3332
rect 11344 3252 16716 3268
rect 11344 3188 16632 3252
rect 16696 3188 16716 3252
rect 11344 3172 16716 3188
rect 11344 3108 16632 3172
rect 16696 3108 16716 3172
rect 11344 3092 16716 3108
rect 11344 3028 16632 3092
rect 16696 3028 16716 3092
rect 11344 3012 16716 3028
rect 11344 2948 16632 3012
rect 16696 2948 16716 3012
rect 11344 2932 16716 2948
rect 11344 2868 16632 2932
rect 16696 2868 16716 2932
rect 11344 2852 16716 2868
rect 11344 2788 16632 2852
rect 16696 2788 16716 2852
rect 11344 2772 16716 2788
rect 11344 2708 16632 2772
rect 16696 2708 16716 2772
rect 11344 2692 16716 2708
rect 11344 2628 16632 2692
rect 16696 2628 16716 2692
rect 11344 2612 16716 2628
rect 11344 2548 16632 2612
rect 16696 2548 16716 2612
rect 11344 2532 16716 2548
rect 11344 2468 16632 2532
rect 16696 2468 16716 2532
rect 11344 2452 16716 2468
rect 11344 2388 16632 2452
rect 16696 2388 16716 2452
rect 11344 2372 16716 2388
rect 11344 2308 16632 2372
rect 16696 2308 16716 2372
rect 11344 2292 16716 2308
rect 11344 2228 16632 2292
rect 16696 2228 16716 2292
rect 11344 2212 16716 2228
rect 11344 2148 16632 2212
rect 16696 2148 16716 2212
rect 11344 2132 16716 2148
rect 11344 2068 16632 2132
rect 16696 2068 16716 2132
rect 11344 2052 16716 2068
rect 11344 1988 16632 2052
rect 16696 1988 16716 2052
rect 11344 1972 16716 1988
rect 11344 1908 16632 1972
rect 16696 1908 16716 1972
rect 11344 1892 16716 1908
rect 11344 1828 16632 1892
rect 16696 1828 16716 1892
rect 11344 1812 16716 1828
rect 11344 1748 16632 1812
rect 16696 1748 16716 1812
rect 11344 1732 16716 1748
rect 11344 1668 16632 1732
rect 16696 1668 16716 1732
rect 11344 1652 16716 1668
rect 11344 1588 16632 1652
rect 16696 1588 16716 1652
rect 11344 1572 16716 1588
rect 11344 1508 16632 1572
rect 16696 1508 16716 1572
rect 11344 1492 16716 1508
rect 11344 1428 16632 1492
rect 16696 1428 16716 1492
rect 11344 1412 16716 1428
rect 11344 1348 16632 1412
rect 16696 1348 16716 1412
rect 11344 1332 16716 1348
rect 11344 1268 16632 1332
rect 16696 1268 16716 1332
rect 11344 1252 16716 1268
rect 11344 1188 16632 1252
rect 16696 1188 16716 1252
rect 11344 1172 16716 1188
rect 11344 1108 16632 1172
rect 16696 1108 16716 1172
rect 11344 1092 16716 1108
rect 11344 1028 16632 1092
rect 16696 1028 16716 1092
rect 11344 1012 16716 1028
rect 11344 948 16632 1012
rect 16696 948 16716 1012
rect 11344 932 16716 948
rect 11344 868 16632 932
rect 16696 868 16716 932
rect 11344 852 16716 868
rect 11344 788 16632 852
rect 16696 788 16716 852
rect 11344 772 16716 788
rect 11344 708 16632 772
rect 16696 708 16716 772
rect 11344 692 16716 708
rect 11344 628 16632 692
rect 16696 628 16716 692
rect 11344 612 16716 628
rect 11344 548 16632 612
rect 16696 548 16716 612
rect 11344 532 16716 548
rect 11344 468 16632 532
rect 16696 468 16716 532
rect 11344 452 16716 468
rect 11344 388 16632 452
rect 16696 388 16716 452
rect 11344 372 16716 388
rect 11344 308 16632 372
rect 16696 308 16716 372
rect 11344 292 16716 308
rect 11344 228 16632 292
rect 16696 228 16716 292
rect 11344 212 16716 228
rect 11344 148 16632 212
rect 16696 148 16716 212
rect 11344 120 16716 148
rect 16956 5172 22328 5200
rect 16956 5108 22244 5172
rect 22308 5108 22328 5172
rect 16956 5092 22328 5108
rect 16956 5028 22244 5092
rect 22308 5028 22328 5092
rect 16956 5012 22328 5028
rect 16956 4948 22244 5012
rect 22308 4948 22328 5012
rect 16956 4932 22328 4948
rect 16956 4868 22244 4932
rect 22308 4868 22328 4932
rect 16956 4852 22328 4868
rect 16956 4788 22244 4852
rect 22308 4788 22328 4852
rect 16956 4772 22328 4788
rect 16956 4708 22244 4772
rect 22308 4708 22328 4772
rect 16956 4692 22328 4708
rect 16956 4628 22244 4692
rect 22308 4628 22328 4692
rect 16956 4612 22328 4628
rect 16956 4548 22244 4612
rect 22308 4548 22328 4612
rect 16956 4532 22328 4548
rect 16956 4468 22244 4532
rect 22308 4468 22328 4532
rect 16956 4452 22328 4468
rect 16956 4388 22244 4452
rect 22308 4388 22328 4452
rect 16956 4372 22328 4388
rect 16956 4308 22244 4372
rect 22308 4308 22328 4372
rect 16956 4292 22328 4308
rect 16956 4228 22244 4292
rect 22308 4228 22328 4292
rect 16956 4212 22328 4228
rect 16956 4148 22244 4212
rect 22308 4148 22328 4212
rect 16956 4132 22328 4148
rect 16956 4068 22244 4132
rect 22308 4068 22328 4132
rect 16956 4052 22328 4068
rect 16956 3988 22244 4052
rect 22308 3988 22328 4052
rect 16956 3972 22328 3988
rect 16956 3908 22244 3972
rect 22308 3908 22328 3972
rect 16956 3892 22328 3908
rect 16956 3828 22244 3892
rect 22308 3828 22328 3892
rect 16956 3812 22328 3828
rect 16956 3748 22244 3812
rect 22308 3748 22328 3812
rect 16956 3732 22328 3748
rect 16956 3668 22244 3732
rect 22308 3668 22328 3732
rect 16956 3652 22328 3668
rect 16956 3588 22244 3652
rect 22308 3588 22328 3652
rect 16956 3572 22328 3588
rect 16956 3508 22244 3572
rect 22308 3508 22328 3572
rect 16956 3492 22328 3508
rect 16956 3428 22244 3492
rect 22308 3428 22328 3492
rect 16956 3412 22328 3428
rect 16956 3348 22244 3412
rect 22308 3348 22328 3412
rect 16956 3332 22328 3348
rect 16956 3268 22244 3332
rect 22308 3268 22328 3332
rect 16956 3252 22328 3268
rect 16956 3188 22244 3252
rect 22308 3188 22328 3252
rect 16956 3172 22328 3188
rect 16956 3108 22244 3172
rect 22308 3108 22328 3172
rect 16956 3092 22328 3108
rect 16956 3028 22244 3092
rect 22308 3028 22328 3092
rect 16956 3012 22328 3028
rect 16956 2948 22244 3012
rect 22308 2948 22328 3012
rect 16956 2932 22328 2948
rect 16956 2868 22244 2932
rect 22308 2868 22328 2932
rect 16956 2852 22328 2868
rect 16956 2788 22244 2852
rect 22308 2788 22328 2852
rect 16956 2772 22328 2788
rect 16956 2708 22244 2772
rect 22308 2708 22328 2772
rect 16956 2692 22328 2708
rect 16956 2628 22244 2692
rect 22308 2628 22328 2692
rect 16956 2612 22328 2628
rect 16956 2548 22244 2612
rect 22308 2548 22328 2612
rect 16956 2532 22328 2548
rect 16956 2468 22244 2532
rect 22308 2468 22328 2532
rect 16956 2452 22328 2468
rect 16956 2388 22244 2452
rect 22308 2388 22328 2452
rect 16956 2372 22328 2388
rect 16956 2308 22244 2372
rect 22308 2308 22328 2372
rect 16956 2292 22328 2308
rect 16956 2228 22244 2292
rect 22308 2228 22328 2292
rect 16956 2212 22328 2228
rect 16956 2148 22244 2212
rect 22308 2148 22328 2212
rect 16956 2132 22328 2148
rect 16956 2068 22244 2132
rect 22308 2068 22328 2132
rect 16956 2052 22328 2068
rect 16956 1988 22244 2052
rect 22308 1988 22328 2052
rect 16956 1972 22328 1988
rect 16956 1908 22244 1972
rect 22308 1908 22328 1972
rect 16956 1892 22328 1908
rect 16956 1828 22244 1892
rect 22308 1828 22328 1892
rect 16956 1812 22328 1828
rect 16956 1748 22244 1812
rect 22308 1748 22328 1812
rect 16956 1732 22328 1748
rect 16956 1668 22244 1732
rect 22308 1668 22328 1732
rect 16956 1652 22328 1668
rect 16956 1588 22244 1652
rect 22308 1588 22328 1652
rect 16956 1572 22328 1588
rect 16956 1508 22244 1572
rect 22308 1508 22328 1572
rect 16956 1492 22328 1508
rect 16956 1428 22244 1492
rect 22308 1428 22328 1492
rect 16956 1412 22328 1428
rect 16956 1348 22244 1412
rect 22308 1348 22328 1412
rect 16956 1332 22328 1348
rect 16956 1268 22244 1332
rect 22308 1268 22328 1332
rect 16956 1252 22328 1268
rect 16956 1188 22244 1252
rect 22308 1188 22328 1252
rect 16956 1172 22328 1188
rect 16956 1108 22244 1172
rect 22308 1108 22328 1172
rect 16956 1092 22328 1108
rect 16956 1028 22244 1092
rect 22308 1028 22328 1092
rect 16956 1012 22328 1028
rect 16956 948 22244 1012
rect 22308 948 22328 1012
rect 16956 932 22328 948
rect 16956 868 22244 932
rect 22308 868 22328 932
rect 16956 852 22328 868
rect 16956 788 22244 852
rect 22308 788 22328 852
rect 16956 772 22328 788
rect 16956 708 22244 772
rect 22308 708 22328 772
rect 16956 692 22328 708
rect 16956 628 22244 692
rect 22308 628 22328 692
rect 16956 612 22328 628
rect 16956 548 22244 612
rect 22308 548 22328 612
rect 16956 532 22328 548
rect 16956 468 22244 532
rect 22308 468 22328 532
rect 16956 452 22328 468
rect 16956 388 22244 452
rect 22308 388 22328 452
rect 16956 372 22328 388
rect 16956 308 22244 372
rect 22308 308 22328 372
rect 16956 292 22328 308
rect 16956 228 22244 292
rect 22308 228 22328 292
rect 16956 212 22328 228
rect 16956 148 22244 212
rect 22308 148 22328 212
rect 16956 120 22328 148
rect 22568 5172 27940 5200
rect 22568 5108 27856 5172
rect 27920 5108 27940 5172
rect 22568 5092 27940 5108
rect 22568 5028 27856 5092
rect 27920 5028 27940 5092
rect 22568 5012 27940 5028
rect 22568 4948 27856 5012
rect 27920 4948 27940 5012
rect 22568 4932 27940 4948
rect 22568 4868 27856 4932
rect 27920 4868 27940 4932
rect 22568 4852 27940 4868
rect 22568 4788 27856 4852
rect 27920 4788 27940 4852
rect 22568 4772 27940 4788
rect 22568 4708 27856 4772
rect 27920 4708 27940 4772
rect 22568 4692 27940 4708
rect 22568 4628 27856 4692
rect 27920 4628 27940 4692
rect 22568 4612 27940 4628
rect 22568 4548 27856 4612
rect 27920 4548 27940 4612
rect 22568 4532 27940 4548
rect 22568 4468 27856 4532
rect 27920 4468 27940 4532
rect 22568 4452 27940 4468
rect 22568 4388 27856 4452
rect 27920 4388 27940 4452
rect 22568 4372 27940 4388
rect 22568 4308 27856 4372
rect 27920 4308 27940 4372
rect 22568 4292 27940 4308
rect 22568 4228 27856 4292
rect 27920 4228 27940 4292
rect 22568 4212 27940 4228
rect 22568 4148 27856 4212
rect 27920 4148 27940 4212
rect 22568 4132 27940 4148
rect 22568 4068 27856 4132
rect 27920 4068 27940 4132
rect 22568 4052 27940 4068
rect 22568 3988 27856 4052
rect 27920 3988 27940 4052
rect 22568 3972 27940 3988
rect 22568 3908 27856 3972
rect 27920 3908 27940 3972
rect 22568 3892 27940 3908
rect 22568 3828 27856 3892
rect 27920 3828 27940 3892
rect 22568 3812 27940 3828
rect 22568 3748 27856 3812
rect 27920 3748 27940 3812
rect 22568 3732 27940 3748
rect 22568 3668 27856 3732
rect 27920 3668 27940 3732
rect 22568 3652 27940 3668
rect 22568 3588 27856 3652
rect 27920 3588 27940 3652
rect 22568 3572 27940 3588
rect 22568 3508 27856 3572
rect 27920 3508 27940 3572
rect 22568 3492 27940 3508
rect 22568 3428 27856 3492
rect 27920 3428 27940 3492
rect 22568 3412 27940 3428
rect 22568 3348 27856 3412
rect 27920 3348 27940 3412
rect 22568 3332 27940 3348
rect 22568 3268 27856 3332
rect 27920 3268 27940 3332
rect 22568 3252 27940 3268
rect 22568 3188 27856 3252
rect 27920 3188 27940 3252
rect 22568 3172 27940 3188
rect 22568 3108 27856 3172
rect 27920 3108 27940 3172
rect 22568 3092 27940 3108
rect 22568 3028 27856 3092
rect 27920 3028 27940 3092
rect 22568 3012 27940 3028
rect 22568 2948 27856 3012
rect 27920 2948 27940 3012
rect 22568 2932 27940 2948
rect 22568 2868 27856 2932
rect 27920 2868 27940 2932
rect 22568 2852 27940 2868
rect 22568 2788 27856 2852
rect 27920 2788 27940 2852
rect 22568 2772 27940 2788
rect 22568 2708 27856 2772
rect 27920 2708 27940 2772
rect 22568 2692 27940 2708
rect 22568 2628 27856 2692
rect 27920 2628 27940 2692
rect 22568 2612 27940 2628
rect 22568 2548 27856 2612
rect 27920 2548 27940 2612
rect 22568 2532 27940 2548
rect 22568 2468 27856 2532
rect 27920 2468 27940 2532
rect 22568 2452 27940 2468
rect 22568 2388 27856 2452
rect 27920 2388 27940 2452
rect 22568 2372 27940 2388
rect 22568 2308 27856 2372
rect 27920 2308 27940 2372
rect 22568 2292 27940 2308
rect 22568 2228 27856 2292
rect 27920 2228 27940 2292
rect 22568 2212 27940 2228
rect 22568 2148 27856 2212
rect 27920 2148 27940 2212
rect 22568 2132 27940 2148
rect 22568 2068 27856 2132
rect 27920 2068 27940 2132
rect 22568 2052 27940 2068
rect 22568 1988 27856 2052
rect 27920 1988 27940 2052
rect 22568 1972 27940 1988
rect 22568 1908 27856 1972
rect 27920 1908 27940 1972
rect 22568 1892 27940 1908
rect 22568 1828 27856 1892
rect 27920 1828 27940 1892
rect 22568 1812 27940 1828
rect 22568 1748 27856 1812
rect 27920 1748 27940 1812
rect 22568 1732 27940 1748
rect 22568 1668 27856 1732
rect 27920 1668 27940 1732
rect 22568 1652 27940 1668
rect 22568 1588 27856 1652
rect 27920 1588 27940 1652
rect 22568 1572 27940 1588
rect 22568 1508 27856 1572
rect 27920 1508 27940 1572
rect 22568 1492 27940 1508
rect 22568 1428 27856 1492
rect 27920 1428 27940 1492
rect 22568 1412 27940 1428
rect 22568 1348 27856 1412
rect 27920 1348 27940 1412
rect 22568 1332 27940 1348
rect 22568 1268 27856 1332
rect 27920 1268 27940 1332
rect 22568 1252 27940 1268
rect 22568 1188 27856 1252
rect 27920 1188 27940 1252
rect 22568 1172 27940 1188
rect 22568 1108 27856 1172
rect 27920 1108 27940 1172
rect 22568 1092 27940 1108
rect 22568 1028 27856 1092
rect 27920 1028 27940 1092
rect 22568 1012 27940 1028
rect 22568 948 27856 1012
rect 27920 948 27940 1012
rect 22568 932 27940 948
rect 22568 868 27856 932
rect 27920 868 27940 932
rect 22568 852 27940 868
rect 22568 788 27856 852
rect 27920 788 27940 852
rect 22568 772 27940 788
rect 22568 708 27856 772
rect 27920 708 27940 772
rect 22568 692 27940 708
rect 22568 628 27856 692
rect 27920 628 27940 692
rect 22568 612 27940 628
rect 22568 548 27856 612
rect 27920 548 27940 612
rect 22568 532 27940 548
rect 22568 468 27856 532
rect 27920 468 27940 532
rect 22568 452 27940 468
rect 22568 388 27856 452
rect 27920 388 27940 452
rect 22568 372 27940 388
rect 22568 308 27856 372
rect 27920 308 27940 372
rect 22568 292 27940 308
rect 22568 228 27856 292
rect 27920 228 27940 292
rect 22568 212 27940 228
rect 22568 148 27856 212
rect 27920 148 27940 212
rect 22568 120 27940 148
rect 28180 5172 33552 5200
rect 28180 5108 33468 5172
rect 33532 5108 33552 5172
rect 28180 5092 33552 5108
rect 28180 5028 33468 5092
rect 33532 5028 33552 5092
rect 28180 5012 33552 5028
rect 28180 4948 33468 5012
rect 33532 4948 33552 5012
rect 28180 4932 33552 4948
rect 28180 4868 33468 4932
rect 33532 4868 33552 4932
rect 28180 4852 33552 4868
rect 28180 4788 33468 4852
rect 33532 4788 33552 4852
rect 28180 4772 33552 4788
rect 28180 4708 33468 4772
rect 33532 4708 33552 4772
rect 28180 4692 33552 4708
rect 28180 4628 33468 4692
rect 33532 4628 33552 4692
rect 28180 4612 33552 4628
rect 28180 4548 33468 4612
rect 33532 4548 33552 4612
rect 28180 4532 33552 4548
rect 28180 4468 33468 4532
rect 33532 4468 33552 4532
rect 28180 4452 33552 4468
rect 28180 4388 33468 4452
rect 33532 4388 33552 4452
rect 28180 4372 33552 4388
rect 28180 4308 33468 4372
rect 33532 4308 33552 4372
rect 28180 4292 33552 4308
rect 28180 4228 33468 4292
rect 33532 4228 33552 4292
rect 28180 4212 33552 4228
rect 28180 4148 33468 4212
rect 33532 4148 33552 4212
rect 28180 4132 33552 4148
rect 28180 4068 33468 4132
rect 33532 4068 33552 4132
rect 28180 4052 33552 4068
rect 28180 3988 33468 4052
rect 33532 3988 33552 4052
rect 28180 3972 33552 3988
rect 28180 3908 33468 3972
rect 33532 3908 33552 3972
rect 28180 3892 33552 3908
rect 28180 3828 33468 3892
rect 33532 3828 33552 3892
rect 28180 3812 33552 3828
rect 28180 3748 33468 3812
rect 33532 3748 33552 3812
rect 28180 3732 33552 3748
rect 28180 3668 33468 3732
rect 33532 3668 33552 3732
rect 28180 3652 33552 3668
rect 28180 3588 33468 3652
rect 33532 3588 33552 3652
rect 28180 3572 33552 3588
rect 28180 3508 33468 3572
rect 33532 3508 33552 3572
rect 28180 3492 33552 3508
rect 28180 3428 33468 3492
rect 33532 3428 33552 3492
rect 28180 3412 33552 3428
rect 28180 3348 33468 3412
rect 33532 3348 33552 3412
rect 28180 3332 33552 3348
rect 28180 3268 33468 3332
rect 33532 3268 33552 3332
rect 28180 3252 33552 3268
rect 28180 3188 33468 3252
rect 33532 3188 33552 3252
rect 28180 3172 33552 3188
rect 28180 3108 33468 3172
rect 33532 3108 33552 3172
rect 28180 3092 33552 3108
rect 28180 3028 33468 3092
rect 33532 3028 33552 3092
rect 28180 3012 33552 3028
rect 28180 2948 33468 3012
rect 33532 2948 33552 3012
rect 28180 2932 33552 2948
rect 28180 2868 33468 2932
rect 33532 2868 33552 2932
rect 28180 2852 33552 2868
rect 28180 2788 33468 2852
rect 33532 2788 33552 2852
rect 28180 2772 33552 2788
rect 28180 2708 33468 2772
rect 33532 2708 33552 2772
rect 28180 2692 33552 2708
rect 28180 2628 33468 2692
rect 33532 2628 33552 2692
rect 28180 2612 33552 2628
rect 28180 2548 33468 2612
rect 33532 2548 33552 2612
rect 28180 2532 33552 2548
rect 28180 2468 33468 2532
rect 33532 2468 33552 2532
rect 28180 2452 33552 2468
rect 28180 2388 33468 2452
rect 33532 2388 33552 2452
rect 28180 2372 33552 2388
rect 28180 2308 33468 2372
rect 33532 2308 33552 2372
rect 28180 2292 33552 2308
rect 28180 2228 33468 2292
rect 33532 2228 33552 2292
rect 28180 2212 33552 2228
rect 28180 2148 33468 2212
rect 33532 2148 33552 2212
rect 28180 2132 33552 2148
rect 28180 2068 33468 2132
rect 33532 2068 33552 2132
rect 28180 2052 33552 2068
rect 28180 1988 33468 2052
rect 33532 1988 33552 2052
rect 28180 1972 33552 1988
rect 28180 1908 33468 1972
rect 33532 1908 33552 1972
rect 28180 1892 33552 1908
rect 28180 1828 33468 1892
rect 33532 1828 33552 1892
rect 28180 1812 33552 1828
rect 28180 1748 33468 1812
rect 33532 1748 33552 1812
rect 28180 1732 33552 1748
rect 28180 1668 33468 1732
rect 33532 1668 33552 1732
rect 28180 1652 33552 1668
rect 28180 1588 33468 1652
rect 33532 1588 33552 1652
rect 28180 1572 33552 1588
rect 28180 1508 33468 1572
rect 33532 1508 33552 1572
rect 28180 1492 33552 1508
rect 28180 1428 33468 1492
rect 33532 1428 33552 1492
rect 28180 1412 33552 1428
rect 28180 1348 33468 1412
rect 33532 1348 33552 1412
rect 28180 1332 33552 1348
rect 28180 1268 33468 1332
rect 33532 1268 33552 1332
rect 28180 1252 33552 1268
rect 28180 1188 33468 1252
rect 33532 1188 33552 1252
rect 28180 1172 33552 1188
rect 28180 1108 33468 1172
rect 33532 1108 33552 1172
rect 28180 1092 33552 1108
rect 28180 1028 33468 1092
rect 33532 1028 33552 1092
rect 28180 1012 33552 1028
rect 28180 948 33468 1012
rect 33532 948 33552 1012
rect 28180 932 33552 948
rect 28180 868 33468 932
rect 33532 868 33552 932
rect 28180 852 33552 868
rect 28180 788 33468 852
rect 33532 788 33552 852
rect 28180 772 33552 788
rect 28180 708 33468 772
rect 33532 708 33552 772
rect 28180 692 33552 708
rect 28180 628 33468 692
rect 33532 628 33552 692
rect 28180 612 33552 628
rect 28180 548 33468 612
rect 33532 548 33552 612
rect 28180 532 33552 548
rect 28180 468 33468 532
rect 33532 468 33552 532
rect 28180 452 33552 468
rect 28180 388 33468 452
rect 33532 388 33552 452
rect 28180 372 33552 388
rect 28180 308 33468 372
rect 33532 308 33552 372
rect 28180 292 33552 308
rect 28180 228 33468 292
rect 33532 228 33552 292
rect 28180 212 33552 228
rect 28180 148 33468 212
rect 33532 148 33552 212
rect 28180 120 33552 148
rect 33792 5172 39164 5200
rect 33792 5108 39080 5172
rect 39144 5108 39164 5172
rect 33792 5092 39164 5108
rect 33792 5028 39080 5092
rect 39144 5028 39164 5092
rect 33792 5012 39164 5028
rect 33792 4948 39080 5012
rect 39144 4948 39164 5012
rect 33792 4932 39164 4948
rect 33792 4868 39080 4932
rect 39144 4868 39164 4932
rect 33792 4852 39164 4868
rect 33792 4788 39080 4852
rect 39144 4788 39164 4852
rect 33792 4772 39164 4788
rect 33792 4708 39080 4772
rect 39144 4708 39164 4772
rect 33792 4692 39164 4708
rect 33792 4628 39080 4692
rect 39144 4628 39164 4692
rect 33792 4612 39164 4628
rect 33792 4548 39080 4612
rect 39144 4548 39164 4612
rect 33792 4532 39164 4548
rect 33792 4468 39080 4532
rect 39144 4468 39164 4532
rect 33792 4452 39164 4468
rect 33792 4388 39080 4452
rect 39144 4388 39164 4452
rect 33792 4372 39164 4388
rect 33792 4308 39080 4372
rect 39144 4308 39164 4372
rect 33792 4292 39164 4308
rect 33792 4228 39080 4292
rect 39144 4228 39164 4292
rect 33792 4212 39164 4228
rect 33792 4148 39080 4212
rect 39144 4148 39164 4212
rect 33792 4132 39164 4148
rect 33792 4068 39080 4132
rect 39144 4068 39164 4132
rect 33792 4052 39164 4068
rect 33792 3988 39080 4052
rect 39144 3988 39164 4052
rect 33792 3972 39164 3988
rect 33792 3908 39080 3972
rect 39144 3908 39164 3972
rect 33792 3892 39164 3908
rect 33792 3828 39080 3892
rect 39144 3828 39164 3892
rect 33792 3812 39164 3828
rect 33792 3748 39080 3812
rect 39144 3748 39164 3812
rect 33792 3732 39164 3748
rect 33792 3668 39080 3732
rect 39144 3668 39164 3732
rect 33792 3652 39164 3668
rect 33792 3588 39080 3652
rect 39144 3588 39164 3652
rect 33792 3572 39164 3588
rect 33792 3508 39080 3572
rect 39144 3508 39164 3572
rect 33792 3492 39164 3508
rect 33792 3428 39080 3492
rect 39144 3428 39164 3492
rect 33792 3412 39164 3428
rect 33792 3348 39080 3412
rect 39144 3348 39164 3412
rect 33792 3332 39164 3348
rect 33792 3268 39080 3332
rect 39144 3268 39164 3332
rect 33792 3252 39164 3268
rect 33792 3188 39080 3252
rect 39144 3188 39164 3252
rect 33792 3172 39164 3188
rect 33792 3108 39080 3172
rect 39144 3108 39164 3172
rect 33792 3092 39164 3108
rect 33792 3028 39080 3092
rect 39144 3028 39164 3092
rect 33792 3012 39164 3028
rect 33792 2948 39080 3012
rect 39144 2948 39164 3012
rect 33792 2932 39164 2948
rect 33792 2868 39080 2932
rect 39144 2868 39164 2932
rect 33792 2852 39164 2868
rect 33792 2788 39080 2852
rect 39144 2788 39164 2852
rect 33792 2772 39164 2788
rect 33792 2708 39080 2772
rect 39144 2708 39164 2772
rect 33792 2692 39164 2708
rect 33792 2628 39080 2692
rect 39144 2628 39164 2692
rect 33792 2612 39164 2628
rect 33792 2548 39080 2612
rect 39144 2548 39164 2612
rect 33792 2532 39164 2548
rect 33792 2468 39080 2532
rect 39144 2468 39164 2532
rect 33792 2452 39164 2468
rect 33792 2388 39080 2452
rect 39144 2388 39164 2452
rect 33792 2372 39164 2388
rect 33792 2308 39080 2372
rect 39144 2308 39164 2372
rect 33792 2292 39164 2308
rect 33792 2228 39080 2292
rect 39144 2228 39164 2292
rect 33792 2212 39164 2228
rect 33792 2148 39080 2212
rect 39144 2148 39164 2212
rect 33792 2132 39164 2148
rect 33792 2068 39080 2132
rect 39144 2068 39164 2132
rect 33792 2052 39164 2068
rect 33792 1988 39080 2052
rect 39144 1988 39164 2052
rect 33792 1972 39164 1988
rect 33792 1908 39080 1972
rect 39144 1908 39164 1972
rect 33792 1892 39164 1908
rect 33792 1828 39080 1892
rect 39144 1828 39164 1892
rect 33792 1812 39164 1828
rect 33792 1748 39080 1812
rect 39144 1748 39164 1812
rect 33792 1732 39164 1748
rect 33792 1668 39080 1732
rect 39144 1668 39164 1732
rect 33792 1652 39164 1668
rect 33792 1588 39080 1652
rect 39144 1588 39164 1652
rect 33792 1572 39164 1588
rect 33792 1508 39080 1572
rect 39144 1508 39164 1572
rect 33792 1492 39164 1508
rect 33792 1428 39080 1492
rect 39144 1428 39164 1492
rect 33792 1412 39164 1428
rect 33792 1348 39080 1412
rect 39144 1348 39164 1412
rect 33792 1332 39164 1348
rect 33792 1268 39080 1332
rect 39144 1268 39164 1332
rect 33792 1252 39164 1268
rect 33792 1188 39080 1252
rect 39144 1188 39164 1252
rect 33792 1172 39164 1188
rect 33792 1108 39080 1172
rect 39144 1108 39164 1172
rect 33792 1092 39164 1108
rect 33792 1028 39080 1092
rect 39144 1028 39164 1092
rect 33792 1012 39164 1028
rect 33792 948 39080 1012
rect 39144 948 39164 1012
rect 33792 932 39164 948
rect 33792 868 39080 932
rect 39144 868 39164 932
rect 33792 852 39164 868
rect 33792 788 39080 852
rect 39144 788 39164 852
rect 33792 772 39164 788
rect 33792 708 39080 772
rect 39144 708 39164 772
rect 33792 692 39164 708
rect 33792 628 39080 692
rect 39144 628 39164 692
rect 33792 612 39164 628
rect 33792 548 39080 612
rect 39144 548 39164 612
rect 33792 532 39164 548
rect 33792 468 39080 532
rect 39144 468 39164 532
rect 33792 452 39164 468
rect 33792 388 39080 452
rect 39144 388 39164 452
rect 33792 372 39164 388
rect 33792 308 39080 372
rect 39144 308 39164 372
rect 33792 292 39164 308
rect 33792 228 39080 292
rect 39144 228 39164 292
rect 33792 212 39164 228
rect 33792 148 39080 212
rect 39144 148 39164 212
rect 33792 120 39164 148
rect -39164 -148 -33792 -120
rect -39164 -212 -33876 -148
rect -33812 -212 -33792 -148
rect -39164 -228 -33792 -212
rect -39164 -292 -33876 -228
rect -33812 -292 -33792 -228
rect -39164 -308 -33792 -292
rect -39164 -372 -33876 -308
rect -33812 -372 -33792 -308
rect -39164 -388 -33792 -372
rect -39164 -452 -33876 -388
rect -33812 -452 -33792 -388
rect -39164 -468 -33792 -452
rect -39164 -532 -33876 -468
rect -33812 -532 -33792 -468
rect -39164 -548 -33792 -532
rect -39164 -612 -33876 -548
rect -33812 -612 -33792 -548
rect -39164 -628 -33792 -612
rect -39164 -692 -33876 -628
rect -33812 -692 -33792 -628
rect -39164 -708 -33792 -692
rect -39164 -772 -33876 -708
rect -33812 -772 -33792 -708
rect -39164 -788 -33792 -772
rect -39164 -852 -33876 -788
rect -33812 -852 -33792 -788
rect -39164 -868 -33792 -852
rect -39164 -932 -33876 -868
rect -33812 -932 -33792 -868
rect -39164 -948 -33792 -932
rect -39164 -1012 -33876 -948
rect -33812 -1012 -33792 -948
rect -39164 -1028 -33792 -1012
rect -39164 -1092 -33876 -1028
rect -33812 -1092 -33792 -1028
rect -39164 -1108 -33792 -1092
rect -39164 -1172 -33876 -1108
rect -33812 -1172 -33792 -1108
rect -39164 -1188 -33792 -1172
rect -39164 -1252 -33876 -1188
rect -33812 -1252 -33792 -1188
rect -39164 -1268 -33792 -1252
rect -39164 -1332 -33876 -1268
rect -33812 -1332 -33792 -1268
rect -39164 -1348 -33792 -1332
rect -39164 -1412 -33876 -1348
rect -33812 -1412 -33792 -1348
rect -39164 -1428 -33792 -1412
rect -39164 -1492 -33876 -1428
rect -33812 -1492 -33792 -1428
rect -39164 -1508 -33792 -1492
rect -39164 -1572 -33876 -1508
rect -33812 -1572 -33792 -1508
rect -39164 -1588 -33792 -1572
rect -39164 -1652 -33876 -1588
rect -33812 -1652 -33792 -1588
rect -39164 -1668 -33792 -1652
rect -39164 -1732 -33876 -1668
rect -33812 -1732 -33792 -1668
rect -39164 -1748 -33792 -1732
rect -39164 -1812 -33876 -1748
rect -33812 -1812 -33792 -1748
rect -39164 -1828 -33792 -1812
rect -39164 -1892 -33876 -1828
rect -33812 -1892 -33792 -1828
rect -39164 -1908 -33792 -1892
rect -39164 -1972 -33876 -1908
rect -33812 -1972 -33792 -1908
rect -39164 -1988 -33792 -1972
rect -39164 -2052 -33876 -1988
rect -33812 -2052 -33792 -1988
rect -39164 -2068 -33792 -2052
rect -39164 -2132 -33876 -2068
rect -33812 -2132 -33792 -2068
rect -39164 -2148 -33792 -2132
rect -39164 -2212 -33876 -2148
rect -33812 -2212 -33792 -2148
rect -39164 -2228 -33792 -2212
rect -39164 -2292 -33876 -2228
rect -33812 -2292 -33792 -2228
rect -39164 -2308 -33792 -2292
rect -39164 -2372 -33876 -2308
rect -33812 -2372 -33792 -2308
rect -39164 -2388 -33792 -2372
rect -39164 -2452 -33876 -2388
rect -33812 -2452 -33792 -2388
rect -39164 -2468 -33792 -2452
rect -39164 -2532 -33876 -2468
rect -33812 -2532 -33792 -2468
rect -39164 -2548 -33792 -2532
rect -39164 -2612 -33876 -2548
rect -33812 -2612 -33792 -2548
rect -39164 -2628 -33792 -2612
rect -39164 -2692 -33876 -2628
rect -33812 -2692 -33792 -2628
rect -39164 -2708 -33792 -2692
rect -39164 -2772 -33876 -2708
rect -33812 -2772 -33792 -2708
rect -39164 -2788 -33792 -2772
rect -39164 -2852 -33876 -2788
rect -33812 -2852 -33792 -2788
rect -39164 -2868 -33792 -2852
rect -39164 -2932 -33876 -2868
rect -33812 -2932 -33792 -2868
rect -39164 -2948 -33792 -2932
rect -39164 -3012 -33876 -2948
rect -33812 -3012 -33792 -2948
rect -39164 -3028 -33792 -3012
rect -39164 -3092 -33876 -3028
rect -33812 -3092 -33792 -3028
rect -39164 -3108 -33792 -3092
rect -39164 -3172 -33876 -3108
rect -33812 -3172 -33792 -3108
rect -39164 -3188 -33792 -3172
rect -39164 -3252 -33876 -3188
rect -33812 -3252 -33792 -3188
rect -39164 -3268 -33792 -3252
rect -39164 -3332 -33876 -3268
rect -33812 -3332 -33792 -3268
rect -39164 -3348 -33792 -3332
rect -39164 -3412 -33876 -3348
rect -33812 -3412 -33792 -3348
rect -39164 -3428 -33792 -3412
rect -39164 -3492 -33876 -3428
rect -33812 -3492 -33792 -3428
rect -39164 -3508 -33792 -3492
rect -39164 -3572 -33876 -3508
rect -33812 -3572 -33792 -3508
rect -39164 -3588 -33792 -3572
rect -39164 -3652 -33876 -3588
rect -33812 -3652 -33792 -3588
rect -39164 -3668 -33792 -3652
rect -39164 -3732 -33876 -3668
rect -33812 -3732 -33792 -3668
rect -39164 -3748 -33792 -3732
rect -39164 -3812 -33876 -3748
rect -33812 -3812 -33792 -3748
rect -39164 -3828 -33792 -3812
rect -39164 -3892 -33876 -3828
rect -33812 -3892 -33792 -3828
rect -39164 -3908 -33792 -3892
rect -39164 -3972 -33876 -3908
rect -33812 -3972 -33792 -3908
rect -39164 -3988 -33792 -3972
rect -39164 -4052 -33876 -3988
rect -33812 -4052 -33792 -3988
rect -39164 -4068 -33792 -4052
rect -39164 -4132 -33876 -4068
rect -33812 -4132 -33792 -4068
rect -39164 -4148 -33792 -4132
rect -39164 -4212 -33876 -4148
rect -33812 -4212 -33792 -4148
rect -39164 -4228 -33792 -4212
rect -39164 -4292 -33876 -4228
rect -33812 -4292 -33792 -4228
rect -39164 -4308 -33792 -4292
rect -39164 -4372 -33876 -4308
rect -33812 -4372 -33792 -4308
rect -39164 -4388 -33792 -4372
rect -39164 -4452 -33876 -4388
rect -33812 -4452 -33792 -4388
rect -39164 -4468 -33792 -4452
rect -39164 -4532 -33876 -4468
rect -33812 -4532 -33792 -4468
rect -39164 -4548 -33792 -4532
rect -39164 -4612 -33876 -4548
rect -33812 -4612 -33792 -4548
rect -39164 -4628 -33792 -4612
rect -39164 -4692 -33876 -4628
rect -33812 -4692 -33792 -4628
rect -39164 -4708 -33792 -4692
rect -39164 -4772 -33876 -4708
rect -33812 -4772 -33792 -4708
rect -39164 -4788 -33792 -4772
rect -39164 -4852 -33876 -4788
rect -33812 -4852 -33792 -4788
rect -39164 -4868 -33792 -4852
rect -39164 -4932 -33876 -4868
rect -33812 -4932 -33792 -4868
rect -39164 -4948 -33792 -4932
rect -39164 -5012 -33876 -4948
rect -33812 -5012 -33792 -4948
rect -39164 -5028 -33792 -5012
rect -39164 -5092 -33876 -5028
rect -33812 -5092 -33792 -5028
rect -39164 -5108 -33792 -5092
rect -39164 -5172 -33876 -5108
rect -33812 -5172 -33792 -5108
rect -39164 -5200 -33792 -5172
rect -33552 -148 -28180 -120
rect -33552 -212 -28264 -148
rect -28200 -212 -28180 -148
rect -33552 -228 -28180 -212
rect -33552 -292 -28264 -228
rect -28200 -292 -28180 -228
rect -33552 -308 -28180 -292
rect -33552 -372 -28264 -308
rect -28200 -372 -28180 -308
rect -33552 -388 -28180 -372
rect -33552 -452 -28264 -388
rect -28200 -452 -28180 -388
rect -33552 -468 -28180 -452
rect -33552 -532 -28264 -468
rect -28200 -532 -28180 -468
rect -33552 -548 -28180 -532
rect -33552 -612 -28264 -548
rect -28200 -612 -28180 -548
rect -33552 -628 -28180 -612
rect -33552 -692 -28264 -628
rect -28200 -692 -28180 -628
rect -33552 -708 -28180 -692
rect -33552 -772 -28264 -708
rect -28200 -772 -28180 -708
rect -33552 -788 -28180 -772
rect -33552 -852 -28264 -788
rect -28200 -852 -28180 -788
rect -33552 -868 -28180 -852
rect -33552 -932 -28264 -868
rect -28200 -932 -28180 -868
rect -33552 -948 -28180 -932
rect -33552 -1012 -28264 -948
rect -28200 -1012 -28180 -948
rect -33552 -1028 -28180 -1012
rect -33552 -1092 -28264 -1028
rect -28200 -1092 -28180 -1028
rect -33552 -1108 -28180 -1092
rect -33552 -1172 -28264 -1108
rect -28200 -1172 -28180 -1108
rect -33552 -1188 -28180 -1172
rect -33552 -1252 -28264 -1188
rect -28200 -1252 -28180 -1188
rect -33552 -1268 -28180 -1252
rect -33552 -1332 -28264 -1268
rect -28200 -1332 -28180 -1268
rect -33552 -1348 -28180 -1332
rect -33552 -1412 -28264 -1348
rect -28200 -1412 -28180 -1348
rect -33552 -1428 -28180 -1412
rect -33552 -1492 -28264 -1428
rect -28200 -1492 -28180 -1428
rect -33552 -1508 -28180 -1492
rect -33552 -1572 -28264 -1508
rect -28200 -1572 -28180 -1508
rect -33552 -1588 -28180 -1572
rect -33552 -1652 -28264 -1588
rect -28200 -1652 -28180 -1588
rect -33552 -1668 -28180 -1652
rect -33552 -1732 -28264 -1668
rect -28200 -1732 -28180 -1668
rect -33552 -1748 -28180 -1732
rect -33552 -1812 -28264 -1748
rect -28200 -1812 -28180 -1748
rect -33552 -1828 -28180 -1812
rect -33552 -1892 -28264 -1828
rect -28200 -1892 -28180 -1828
rect -33552 -1908 -28180 -1892
rect -33552 -1972 -28264 -1908
rect -28200 -1972 -28180 -1908
rect -33552 -1988 -28180 -1972
rect -33552 -2052 -28264 -1988
rect -28200 -2052 -28180 -1988
rect -33552 -2068 -28180 -2052
rect -33552 -2132 -28264 -2068
rect -28200 -2132 -28180 -2068
rect -33552 -2148 -28180 -2132
rect -33552 -2212 -28264 -2148
rect -28200 -2212 -28180 -2148
rect -33552 -2228 -28180 -2212
rect -33552 -2292 -28264 -2228
rect -28200 -2292 -28180 -2228
rect -33552 -2308 -28180 -2292
rect -33552 -2372 -28264 -2308
rect -28200 -2372 -28180 -2308
rect -33552 -2388 -28180 -2372
rect -33552 -2452 -28264 -2388
rect -28200 -2452 -28180 -2388
rect -33552 -2468 -28180 -2452
rect -33552 -2532 -28264 -2468
rect -28200 -2532 -28180 -2468
rect -33552 -2548 -28180 -2532
rect -33552 -2612 -28264 -2548
rect -28200 -2612 -28180 -2548
rect -33552 -2628 -28180 -2612
rect -33552 -2692 -28264 -2628
rect -28200 -2692 -28180 -2628
rect -33552 -2708 -28180 -2692
rect -33552 -2772 -28264 -2708
rect -28200 -2772 -28180 -2708
rect -33552 -2788 -28180 -2772
rect -33552 -2852 -28264 -2788
rect -28200 -2852 -28180 -2788
rect -33552 -2868 -28180 -2852
rect -33552 -2932 -28264 -2868
rect -28200 -2932 -28180 -2868
rect -33552 -2948 -28180 -2932
rect -33552 -3012 -28264 -2948
rect -28200 -3012 -28180 -2948
rect -33552 -3028 -28180 -3012
rect -33552 -3092 -28264 -3028
rect -28200 -3092 -28180 -3028
rect -33552 -3108 -28180 -3092
rect -33552 -3172 -28264 -3108
rect -28200 -3172 -28180 -3108
rect -33552 -3188 -28180 -3172
rect -33552 -3252 -28264 -3188
rect -28200 -3252 -28180 -3188
rect -33552 -3268 -28180 -3252
rect -33552 -3332 -28264 -3268
rect -28200 -3332 -28180 -3268
rect -33552 -3348 -28180 -3332
rect -33552 -3412 -28264 -3348
rect -28200 -3412 -28180 -3348
rect -33552 -3428 -28180 -3412
rect -33552 -3492 -28264 -3428
rect -28200 -3492 -28180 -3428
rect -33552 -3508 -28180 -3492
rect -33552 -3572 -28264 -3508
rect -28200 -3572 -28180 -3508
rect -33552 -3588 -28180 -3572
rect -33552 -3652 -28264 -3588
rect -28200 -3652 -28180 -3588
rect -33552 -3668 -28180 -3652
rect -33552 -3732 -28264 -3668
rect -28200 -3732 -28180 -3668
rect -33552 -3748 -28180 -3732
rect -33552 -3812 -28264 -3748
rect -28200 -3812 -28180 -3748
rect -33552 -3828 -28180 -3812
rect -33552 -3892 -28264 -3828
rect -28200 -3892 -28180 -3828
rect -33552 -3908 -28180 -3892
rect -33552 -3972 -28264 -3908
rect -28200 -3972 -28180 -3908
rect -33552 -3988 -28180 -3972
rect -33552 -4052 -28264 -3988
rect -28200 -4052 -28180 -3988
rect -33552 -4068 -28180 -4052
rect -33552 -4132 -28264 -4068
rect -28200 -4132 -28180 -4068
rect -33552 -4148 -28180 -4132
rect -33552 -4212 -28264 -4148
rect -28200 -4212 -28180 -4148
rect -33552 -4228 -28180 -4212
rect -33552 -4292 -28264 -4228
rect -28200 -4292 -28180 -4228
rect -33552 -4308 -28180 -4292
rect -33552 -4372 -28264 -4308
rect -28200 -4372 -28180 -4308
rect -33552 -4388 -28180 -4372
rect -33552 -4452 -28264 -4388
rect -28200 -4452 -28180 -4388
rect -33552 -4468 -28180 -4452
rect -33552 -4532 -28264 -4468
rect -28200 -4532 -28180 -4468
rect -33552 -4548 -28180 -4532
rect -33552 -4612 -28264 -4548
rect -28200 -4612 -28180 -4548
rect -33552 -4628 -28180 -4612
rect -33552 -4692 -28264 -4628
rect -28200 -4692 -28180 -4628
rect -33552 -4708 -28180 -4692
rect -33552 -4772 -28264 -4708
rect -28200 -4772 -28180 -4708
rect -33552 -4788 -28180 -4772
rect -33552 -4852 -28264 -4788
rect -28200 -4852 -28180 -4788
rect -33552 -4868 -28180 -4852
rect -33552 -4932 -28264 -4868
rect -28200 -4932 -28180 -4868
rect -33552 -4948 -28180 -4932
rect -33552 -5012 -28264 -4948
rect -28200 -5012 -28180 -4948
rect -33552 -5028 -28180 -5012
rect -33552 -5092 -28264 -5028
rect -28200 -5092 -28180 -5028
rect -33552 -5108 -28180 -5092
rect -33552 -5172 -28264 -5108
rect -28200 -5172 -28180 -5108
rect -33552 -5200 -28180 -5172
rect -27940 -148 -22568 -120
rect -27940 -212 -22652 -148
rect -22588 -212 -22568 -148
rect -27940 -228 -22568 -212
rect -27940 -292 -22652 -228
rect -22588 -292 -22568 -228
rect -27940 -308 -22568 -292
rect -27940 -372 -22652 -308
rect -22588 -372 -22568 -308
rect -27940 -388 -22568 -372
rect -27940 -452 -22652 -388
rect -22588 -452 -22568 -388
rect -27940 -468 -22568 -452
rect -27940 -532 -22652 -468
rect -22588 -532 -22568 -468
rect -27940 -548 -22568 -532
rect -27940 -612 -22652 -548
rect -22588 -612 -22568 -548
rect -27940 -628 -22568 -612
rect -27940 -692 -22652 -628
rect -22588 -692 -22568 -628
rect -27940 -708 -22568 -692
rect -27940 -772 -22652 -708
rect -22588 -772 -22568 -708
rect -27940 -788 -22568 -772
rect -27940 -852 -22652 -788
rect -22588 -852 -22568 -788
rect -27940 -868 -22568 -852
rect -27940 -932 -22652 -868
rect -22588 -932 -22568 -868
rect -27940 -948 -22568 -932
rect -27940 -1012 -22652 -948
rect -22588 -1012 -22568 -948
rect -27940 -1028 -22568 -1012
rect -27940 -1092 -22652 -1028
rect -22588 -1092 -22568 -1028
rect -27940 -1108 -22568 -1092
rect -27940 -1172 -22652 -1108
rect -22588 -1172 -22568 -1108
rect -27940 -1188 -22568 -1172
rect -27940 -1252 -22652 -1188
rect -22588 -1252 -22568 -1188
rect -27940 -1268 -22568 -1252
rect -27940 -1332 -22652 -1268
rect -22588 -1332 -22568 -1268
rect -27940 -1348 -22568 -1332
rect -27940 -1412 -22652 -1348
rect -22588 -1412 -22568 -1348
rect -27940 -1428 -22568 -1412
rect -27940 -1492 -22652 -1428
rect -22588 -1492 -22568 -1428
rect -27940 -1508 -22568 -1492
rect -27940 -1572 -22652 -1508
rect -22588 -1572 -22568 -1508
rect -27940 -1588 -22568 -1572
rect -27940 -1652 -22652 -1588
rect -22588 -1652 -22568 -1588
rect -27940 -1668 -22568 -1652
rect -27940 -1732 -22652 -1668
rect -22588 -1732 -22568 -1668
rect -27940 -1748 -22568 -1732
rect -27940 -1812 -22652 -1748
rect -22588 -1812 -22568 -1748
rect -27940 -1828 -22568 -1812
rect -27940 -1892 -22652 -1828
rect -22588 -1892 -22568 -1828
rect -27940 -1908 -22568 -1892
rect -27940 -1972 -22652 -1908
rect -22588 -1972 -22568 -1908
rect -27940 -1988 -22568 -1972
rect -27940 -2052 -22652 -1988
rect -22588 -2052 -22568 -1988
rect -27940 -2068 -22568 -2052
rect -27940 -2132 -22652 -2068
rect -22588 -2132 -22568 -2068
rect -27940 -2148 -22568 -2132
rect -27940 -2212 -22652 -2148
rect -22588 -2212 -22568 -2148
rect -27940 -2228 -22568 -2212
rect -27940 -2292 -22652 -2228
rect -22588 -2292 -22568 -2228
rect -27940 -2308 -22568 -2292
rect -27940 -2372 -22652 -2308
rect -22588 -2372 -22568 -2308
rect -27940 -2388 -22568 -2372
rect -27940 -2452 -22652 -2388
rect -22588 -2452 -22568 -2388
rect -27940 -2468 -22568 -2452
rect -27940 -2532 -22652 -2468
rect -22588 -2532 -22568 -2468
rect -27940 -2548 -22568 -2532
rect -27940 -2612 -22652 -2548
rect -22588 -2612 -22568 -2548
rect -27940 -2628 -22568 -2612
rect -27940 -2692 -22652 -2628
rect -22588 -2692 -22568 -2628
rect -27940 -2708 -22568 -2692
rect -27940 -2772 -22652 -2708
rect -22588 -2772 -22568 -2708
rect -27940 -2788 -22568 -2772
rect -27940 -2852 -22652 -2788
rect -22588 -2852 -22568 -2788
rect -27940 -2868 -22568 -2852
rect -27940 -2932 -22652 -2868
rect -22588 -2932 -22568 -2868
rect -27940 -2948 -22568 -2932
rect -27940 -3012 -22652 -2948
rect -22588 -3012 -22568 -2948
rect -27940 -3028 -22568 -3012
rect -27940 -3092 -22652 -3028
rect -22588 -3092 -22568 -3028
rect -27940 -3108 -22568 -3092
rect -27940 -3172 -22652 -3108
rect -22588 -3172 -22568 -3108
rect -27940 -3188 -22568 -3172
rect -27940 -3252 -22652 -3188
rect -22588 -3252 -22568 -3188
rect -27940 -3268 -22568 -3252
rect -27940 -3332 -22652 -3268
rect -22588 -3332 -22568 -3268
rect -27940 -3348 -22568 -3332
rect -27940 -3412 -22652 -3348
rect -22588 -3412 -22568 -3348
rect -27940 -3428 -22568 -3412
rect -27940 -3492 -22652 -3428
rect -22588 -3492 -22568 -3428
rect -27940 -3508 -22568 -3492
rect -27940 -3572 -22652 -3508
rect -22588 -3572 -22568 -3508
rect -27940 -3588 -22568 -3572
rect -27940 -3652 -22652 -3588
rect -22588 -3652 -22568 -3588
rect -27940 -3668 -22568 -3652
rect -27940 -3732 -22652 -3668
rect -22588 -3732 -22568 -3668
rect -27940 -3748 -22568 -3732
rect -27940 -3812 -22652 -3748
rect -22588 -3812 -22568 -3748
rect -27940 -3828 -22568 -3812
rect -27940 -3892 -22652 -3828
rect -22588 -3892 -22568 -3828
rect -27940 -3908 -22568 -3892
rect -27940 -3972 -22652 -3908
rect -22588 -3972 -22568 -3908
rect -27940 -3988 -22568 -3972
rect -27940 -4052 -22652 -3988
rect -22588 -4052 -22568 -3988
rect -27940 -4068 -22568 -4052
rect -27940 -4132 -22652 -4068
rect -22588 -4132 -22568 -4068
rect -27940 -4148 -22568 -4132
rect -27940 -4212 -22652 -4148
rect -22588 -4212 -22568 -4148
rect -27940 -4228 -22568 -4212
rect -27940 -4292 -22652 -4228
rect -22588 -4292 -22568 -4228
rect -27940 -4308 -22568 -4292
rect -27940 -4372 -22652 -4308
rect -22588 -4372 -22568 -4308
rect -27940 -4388 -22568 -4372
rect -27940 -4452 -22652 -4388
rect -22588 -4452 -22568 -4388
rect -27940 -4468 -22568 -4452
rect -27940 -4532 -22652 -4468
rect -22588 -4532 -22568 -4468
rect -27940 -4548 -22568 -4532
rect -27940 -4612 -22652 -4548
rect -22588 -4612 -22568 -4548
rect -27940 -4628 -22568 -4612
rect -27940 -4692 -22652 -4628
rect -22588 -4692 -22568 -4628
rect -27940 -4708 -22568 -4692
rect -27940 -4772 -22652 -4708
rect -22588 -4772 -22568 -4708
rect -27940 -4788 -22568 -4772
rect -27940 -4852 -22652 -4788
rect -22588 -4852 -22568 -4788
rect -27940 -4868 -22568 -4852
rect -27940 -4932 -22652 -4868
rect -22588 -4932 -22568 -4868
rect -27940 -4948 -22568 -4932
rect -27940 -5012 -22652 -4948
rect -22588 -5012 -22568 -4948
rect -27940 -5028 -22568 -5012
rect -27940 -5092 -22652 -5028
rect -22588 -5092 -22568 -5028
rect -27940 -5108 -22568 -5092
rect -27940 -5172 -22652 -5108
rect -22588 -5172 -22568 -5108
rect -27940 -5200 -22568 -5172
rect -22328 -148 -16956 -120
rect -22328 -212 -17040 -148
rect -16976 -212 -16956 -148
rect -22328 -228 -16956 -212
rect -22328 -292 -17040 -228
rect -16976 -292 -16956 -228
rect -22328 -308 -16956 -292
rect -22328 -372 -17040 -308
rect -16976 -372 -16956 -308
rect -22328 -388 -16956 -372
rect -22328 -452 -17040 -388
rect -16976 -452 -16956 -388
rect -22328 -468 -16956 -452
rect -22328 -532 -17040 -468
rect -16976 -532 -16956 -468
rect -22328 -548 -16956 -532
rect -22328 -612 -17040 -548
rect -16976 -612 -16956 -548
rect -22328 -628 -16956 -612
rect -22328 -692 -17040 -628
rect -16976 -692 -16956 -628
rect -22328 -708 -16956 -692
rect -22328 -772 -17040 -708
rect -16976 -772 -16956 -708
rect -22328 -788 -16956 -772
rect -22328 -852 -17040 -788
rect -16976 -852 -16956 -788
rect -22328 -868 -16956 -852
rect -22328 -932 -17040 -868
rect -16976 -932 -16956 -868
rect -22328 -948 -16956 -932
rect -22328 -1012 -17040 -948
rect -16976 -1012 -16956 -948
rect -22328 -1028 -16956 -1012
rect -22328 -1092 -17040 -1028
rect -16976 -1092 -16956 -1028
rect -22328 -1108 -16956 -1092
rect -22328 -1172 -17040 -1108
rect -16976 -1172 -16956 -1108
rect -22328 -1188 -16956 -1172
rect -22328 -1252 -17040 -1188
rect -16976 -1252 -16956 -1188
rect -22328 -1268 -16956 -1252
rect -22328 -1332 -17040 -1268
rect -16976 -1332 -16956 -1268
rect -22328 -1348 -16956 -1332
rect -22328 -1412 -17040 -1348
rect -16976 -1412 -16956 -1348
rect -22328 -1428 -16956 -1412
rect -22328 -1492 -17040 -1428
rect -16976 -1492 -16956 -1428
rect -22328 -1508 -16956 -1492
rect -22328 -1572 -17040 -1508
rect -16976 -1572 -16956 -1508
rect -22328 -1588 -16956 -1572
rect -22328 -1652 -17040 -1588
rect -16976 -1652 -16956 -1588
rect -22328 -1668 -16956 -1652
rect -22328 -1732 -17040 -1668
rect -16976 -1732 -16956 -1668
rect -22328 -1748 -16956 -1732
rect -22328 -1812 -17040 -1748
rect -16976 -1812 -16956 -1748
rect -22328 -1828 -16956 -1812
rect -22328 -1892 -17040 -1828
rect -16976 -1892 -16956 -1828
rect -22328 -1908 -16956 -1892
rect -22328 -1972 -17040 -1908
rect -16976 -1972 -16956 -1908
rect -22328 -1988 -16956 -1972
rect -22328 -2052 -17040 -1988
rect -16976 -2052 -16956 -1988
rect -22328 -2068 -16956 -2052
rect -22328 -2132 -17040 -2068
rect -16976 -2132 -16956 -2068
rect -22328 -2148 -16956 -2132
rect -22328 -2212 -17040 -2148
rect -16976 -2212 -16956 -2148
rect -22328 -2228 -16956 -2212
rect -22328 -2292 -17040 -2228
rect -16976 -2292 -16956 -2228
rect -22328 -2308 -16956 -2292
rect -22328 -2372 -17040 -2308
rect -16976 -2372 -16956 -2308
rect -22328 -2388 -16956 -2372
rect -22328 -2452 -17040 -2388
rect -16976 -2452 -16956 -2388
rect -22328 -2468 -16956 -2452
rect -22328 -2532 -17040 -2468
rect -16976 -2532 -16956 -2468
rect -22328 -2548 -16956 -2532
rect -22328 -2612 -17040 -2548
rect -16976 -2612 -16956 -2548
rect -22328 -2628 -16956 -2612
rect -22328 -2692 -17040 -2628
rect -16976 -2692 -16956 -2628
rect -22328 -2708 -16956 -2692
rect -22328 -2772 -17040 -2708
rect -16976 -2772 -16956 -2708
rect -22328 -2788 -16956 -2772
rect -22328 -2852 -17040 -2788
rect -16976 -2852 -16956 -2788
rect -22328 -2868 -16956 -2852
rect -22328 -2932 -17040 -2868
rect -16976 -2932 -16956 -2868
rect -22328 -2948 -16956 -2932
rect -22328 -3012 -17040 -2948
rect -16976 -3012 -16956 -2948
rect -22328 -3028 -16956 -3012
rect -22328 -3092 -17040 -3028
rect -16976 -3092 -16956 -3028
rect -22328 -3108 -16956 -3092
rect -22328 -3172 -17040 -3108
rect -16976 -3172 -16956 -3108
rect -22328 -3188 -16956 -3172
rect -22328 -3252 -17040 -3188
rect -16976 -3252 -16956 -3188
rect -22328 -3268 -16956 -3252
rect -22328 -3332 -17040 -3268
rect -16976 -3332 -16956 -3268
rect -22328 -3348 -16956 -3332
rect -22328 -3412 -17040 -3348
rect -16976 -3412 -16956 -3348
rect -22328 -3428 -16956 -3412
rect -22328 -3492 -17040 -3428
rect -16976 -3492 -16956 -3428
rect -22328 -3508 -16956 -3492
rect -22328 -3572 -17040 -3508
rect -16976 -3572 -16956 -3508
rect -22328 -3588 -16956 -3572
rect -22328 -3652 -17040 -3588
rect -16976 -3652 -16956 -3588
rect -22328 -3668 -16956 -3652
rect -22328 -3732 -17040 -3668
rect -16976 -3732 -16956 -3668
rect -22328 -3748 -16956 -3732
rect -22328 -3812 -17040 -3748
rect -16976 -3812 -16956 -3748
rect -22328 -3828 -16956 -3812
rect -22328 -3892 -17040 -3828
rect -16976 -3892 -16956 -3828
rect -22328 -3908 -16956 -3892
rect -22328 -3972 -17040 -3908
rect -16976 -3972 -16956 -3908
rect -22328 -3988 -16956 -3972
rect -22328 -4052 -17040 -3988
rect -16976 -4052 -16956 -3988
rect -22328 -4068 -16956 -4052
rect -22328 -4132 -17040 -4068
rect -16976 -4132 -16956 -4068
rect -22328 -4148 -16956 -4132
rect -22328 -4212 -17040 -4148
rect -16976 -4212 -16956 -4148
rect -22328 -4228 -16956 -4212
rect -22328 -4292 -17040 -4228
rect -16976 -4292 -16956 -4228
rect -22328 -4308 -16956 -4292
rect -22328 -4372 -17040 -4308
rect -16976 -4372 -16956 -4308
rect -22328 -4388 -16956 -4372
rect -22328 -4452 -17040 -4388
rect -16976 -4452 -16956 -4388
rect -22328 -4468 -16956 -4452
rect -22328 -4532 -17040 -4468
rect -16976 -4532 -16956 -4468
rect -22328 -4548 -16956 -4532
rect -22328 -4612 -17040 -4548
rect -16976 -4612 -16956 -4548
rect -22328 -4628 -16956 -4612
rect -22328 -4692 -17040 -4628
rect -16976 -4692 -16956 -4628
rect -22328 -4708 -16956 -4692
rect -22328 -4772 -17040 -4708
rect -16976 -4772 -16956 -4708
rect -22328 -4788 -16956 -4772
rect -22328 -4852 -17040 -4788
rect -16976 -4852 -16956 -4788
rect -22328 -4868 -16956 -4852
rect -22328 -4932 -17040 -4868
rect -16976 -4932 -16956 -4868
rect -22328 -4948 -16956 -4932
rect -22328 -5012 -17040 -4948
rect -16976 -5012 -16956 -4948
rect -22328 -5028 -16956 -5012
rect -22328 -5092 -17040 -5028
rect -16976 -5092 -16956 -5028
rect -22328 -5108 -16956 -5092
rect -22328 -5172 -17040 -5108
rect -16976 -5172 -16956 -5108
rect -22328 -5200 -16956 -5172
rect -16716 -148 -11344 -120
rect -16716 -212 -11428 -148
rect -11364 -212 -11344 -148
rect -16716 -228 -11344 -212
rect -16716 -292 -11428 -228
rect -11364 -292 -11344 -228
rect -16716 -308 -11344 -292
rect -16716 -372 -11428 -308
rect -11364 -372 -11344 -308
rect -16716 -388 -11344 -372
rect -16716 -452 -11428 -388
rect -11364 -452 -11344 -388
rect -16716 -468 -11344 -452
rect -16716 -532 -11428 -468
rect -11364 -532 -11344 -468
rect -16716 -548 -11344 -532
rect -16716 -612 -11428 -548
rect -11364 -612 -11344 -548
rect -16716 -628 -11344 -612
rect -16716 -692 -11428 -628
rect -11364 -692 -11344 -628
rect -16716 -708 -11344 -692
rect -16716 -772 -11428 -708
rect -11364 -772 -11344 -708
rect -16716 -788 -11344 -772
rect -16716 -852 -11428 -788
rect -11364 -852 -11344 -788
rect -16716 -868 -11344 -852
rect -16716 -932 -11428 -868
rect -11364 -932 -11344 -868
rect -16716 -948 -11344 -932
rect -16716 -1012 -11428 -948
rect -11364 -1012 -11344 -948
rect -16716 -1028 -11344 -1012
rect -16716 -1092 -11428 -1028
rect -11364 -1092 -11344 -1028
rect -16716 -1108 -11344 -1092
rect -16716 -1172 -11428 -1108
rect -11364 -1172 -11344 -1108
rect -16716 -1188 -11344 -1172
rect -16716 -1252 -11428 -1188
rect -11364 -1252 -11344 -1188
rect -16716 -1268 -11344 -1252
rect -16716 -1332 -11428 -1268
rect -11364 -1332 -11344 -1268
rect -16716 -1348 -11344 -1332
rect -16716 -1412 -11428 -1348
rect -11364 -1412 -11344 -1348
rect -16716 -1428 -11344 -1412
rect -16716 -1492 -11428 -1428
rect -11364 -1492 -11344 -1428
rect -16716 -1508 -11344 -1492
rect -16716 -1572 -11428 -1508
rect -11364 -1572 -11344 -1508
rect -16716 -1588 -11344 -1572
rect -16716 -1652 -11428 -1588
rect -11364 -1652 -11344 -1588
rect -16716 -1668 -11344 -1652
rect -16716 -1732 -11428 -1668
rect -11364 -1732 -11344 -1668
rect -16716 -1748 -11344 -1732
rect -16716 -1812 -11428 -1748
rect -11364 -1812 -11344 -1748
rect -16716 -1828 -11344 -1812
rect -16716 -1892 -11428 -1828
rect -11364 -1892 -11344 -1828
rect -16716 -1908 -11344 -1892
rect -16716 -1972 -11428 -1908
rect -11364 -1972 -11344 -1908
rect -16716 -1988 -11344 -1972
rect -16716 -2052 -11428 -1988
rect -11364 -2052 -11344 -1988
rect -16716 -2068 -11344 -2052
rect -16716 -2132 -11428 -2068
rect -11364 -2132 -11344 -2068
rect -16716 -2148 -11344 -2132
rect -16716 -2212 -11428 -2148
rect -11364 -2212 -11344 -2148
rect -16716 -2228 -11344 -2212
rect -16716 -2292 -11428 -2228
rect -11364 -2292 -11344 -2228
rect -16716 -2308 -11344 -2292
rect -16716 -2372 -11428 -2308
rect -11364 -2372 -11344 -2308
rect -16716 -2388 -11344 -2372
rect -16716 -2452 -11428 -2388
rect -11364 -2452 -11344 -2388
rect -16716 -2468 -11344 -2452
rect -16716 -2532 -11428 -2468
rect -11364 -2532 -11344 -2468
rect -16716 -2548 -11344 -2532
rect -16716 -2612 -11428 -2548
rect -11364 -2612 -11344 -2548
rect -16716 -2628 -11344 -2612
rect -16716 -2692 -11428 -2628
rect -11364 -2692 -11344 -2628
rect -16716 -2708 -11344 -2692
rect -16716 -2772 -11428 -2708
rect -11364 -2772 -11344 -2708
rect -16716 -2788 -11344 -2772
rect -16716 -2852 -11428 -2788
rect -11364 -2852 -11344 -2788
rect -16716 -2868 -11344 -2852
rect -16716 -2932 -11428 -2868
rect -11364 -2932 -11344 -2868
rect -16716 -2948 -11344 -2932
rect -16716 -3012 -11428 -2948
rect -11364 -3012 -11344 -2948
rect -16716 -3028 -11344 -3012
rect -16716 -3092 -11428 -3028
rect -11364 -3092 -11344 -3028
rect -16716 -3108 -11344 -3092
rect -16716 -3172 -11428 -3108
rect -11364 -3172 -11344 -3108
rect -16716 -3188 -11344 -3172
rect -16716 -3252 -11428 -3188
rect -11364 -3252 -11344 -3188
rect -16716 -3268 -11344 -3252
rect -16716 -3332 -11428 -3268
rect -11364 -3332 -11344 -3268
rect -16716 -3348 -11344 -3332
rect -16716 -3412 -11428 -3348
rect -11364 -3412 -11344 -3348
rect -16716 -3428 -11344 -3412
rect -16716 -3492 -11428 -3428
rect -11364 -3492 -11344 -3428
rect -16716 -3508 -11344 -3492
rect -16716 -3572 -11428 -3508
rect -11364 -3572 -11344 -3508
rect -16716 -3588 -11344 -3572
rect -16716 -3652 -11428 -3588
rect -11364 -3652 -11344 -3588
rect -16716 -3668 -11344 -3652
rect -16716 -3732 -11428 -3668
rect -11364 -3732 -11344 -3668
rect -16716 -3748 -11344 -3732
rect -16716 -3812 -11428 -3748
rect -11364 -3812 -11344 -3748
rect -16716 -3828 -11344 -3812
rect -16716 -3892 -11428 -3828
rect -11364 -3892 -11344 -3828
rect -16716 -3908 -11344 -3892
rect -16716 -3972 -11428 -3908
rect -11364 -3972 -11344 -3908
rect -16716 -3988 -11344 -3972
rect -16716 -4052 -11428 -3988
rect -11364 -4052 -11344 -3988
rect -16716 -4068 -11344 -4052
rect -16716 -4132 -11428 -4068
rect -11364 -4132 -11344 -4068
rect -16716 -4148 -11344 -4132
rect -16716 -4212 -11428 -4148
rect -11364 -4212 -11344 -4148
rect -16716 -4228 -11344 -4212
rect -16716 -4292 -11428 -4228
rect -11364 -4292 -11344 -4228
rect -16716 -4308 -11344 -4292
rect -16716 -4372 -11428 -4308
rect -11364 -4372 -11344 -4308
rect -16716 -4388 -11344 -4372
rect -16716 -4452 -11428 -4388
rect -11364 -4452 -11344 -4388
rect -16716 -4468 -11344 -4452
rect -16716 -4532 -11428 -4468
rect -11364 -4532 -11344 -4468
rect -16716 -4548 -11344 -4532
rect -16716 -4612 -11428 -4548
rect -11364 -4612 -11344 -4548
rect -16716 -4628 -11344 -4612
rect -16716 -4692 -11428 -4628
rect -11364 -4692 -11344 -4628
rect -16716 -4708 -11344 -4692
rect -16716 -4772 -11428 -4708
rect -11364 -4772 -11344 -4708
rect -16716 -4788 -11344 -4772
rect -16716 -4852 -11428 -4788
rect -11364 -4852 -11344 -4788
rect -16716 -4868 -11344 -4852
rect -16716 -4932 -11428 -4868
rect -11364 -4932 -11344 -4868
rect -16716 -4948 -11344 -4932
rect -16716 -5012 -11428 -4948
rect -11364 -5012 -11344 -4948
rect -16716 -5028 -11344 -5012
rect -16716 -5092 -11428 -5028
rect -11364 -5092 -11344 -5028
rect -16716 -5108 -11344 -5092
rect -16716 -5172 -11428 -5108
rect -11364 -5172 -11344 -5108
rect -16716 -5200 -11344 -5172
rect -11104 -148 -5732 -120
rect -11104 -212 -5816 -148
rect -5752 -212 -5732 -148
rect -11104 -228 -5732 -212
rect -11104 -292 -5816 -228
rect -5752 -292 -5732 -228
rect -11104 -308 -5732 -292
rect -11104 -372 -5816 -308
rect -5752 -372 -5732 -308
rect -11104 -388 -5732 -372
rect -11104 -452 -5816 -388
rect -5752 -452 -5732 -388
rect -11104 -468 -5732 -452
rect -11104 -532 -5816 -468
rect -5752 -532 -5732 -468
rect -11104 -548 -5732 -532
rect -11104 -612 -5816 -548
rect -5752 -612 -5732 -548
rect -11104 -628 -5732 -612
rect -11104 -692 -5816 -628
rect -5752 -692 -5732 -628
rect -11104 -708 -5732 -692
rect -11104 -772 -5816 -708
rect -5752 -772 -5732 -708
rect -11104 -788 -5732 -772
rect -11104 -852 -5816 -788
rect -5752 -852 -5732 -788
rect -11104 -868 -5732 -852
rect -11104 -932 -5816 -868
rect -5752 -932 -5732 -868
rect -11104 -948 -5732 -932
rect -11104 -1012 -5816 -948
rect -5752 -1012 -5732 -948
rect -11104 -1028 -5732 -1012
rect -11104 -1092 -5816 -1028
rect -5752 -1092 -5732 -1028
rect -11104 -1108 -5732 -1092
rect -11104 -1172 -5816 -1108
rect -5752 -1172 -5732 -1108
rect -11104 -1188 -5732 -1172
rect -11104 -1252 -5816 -1188
rect -5752 -1252 -5732 -1188
rect -11104 -1268 -5732 -1252
rect -11104 -1332 -5816 -1268
rect -5752 -1332 -5732 -1268
rect -11104 -1348 -5732 -1332
rect -11104 -1412 -5816 -1348
rect -5752 -1412 -5732 -1348
rect -11104 -1428 -5732 -1412
rect -11104 -1492 -5816 -1428
rect -5752 -1492 -5732 -1428
rect -11104 -1508 -5732 -1492
rect -11104 -1572 -5816 -1508
rect -5752 -1572 -5732 -1508
rect -11104 -1588 -5732 -1572
rect -11104 -1652 -5816 -1588
rect -5752 -1652 -5732 -1588
rect -11104 -1668 -5732 -1652
rect -11104 -1732 -5816 -1668
rect -5752 -1732 -5732 -1668
rect -11104 -1748 -5732 -1732
rect -11104 -1812 -5816 -1748
rect -5752 -1812 -5732 -1748
rect -11104 -1828 -5732 -1812
rect -11104 -1892 -5816 -1828
rect -5752 -1892 -5732 -1828
rect -11104 -1908 -5732 -1892
rect -11104 -1972 -5816 -1908
rect -5752 -1972 -5732 -1908
rect -11104 -1988 -5732 -1972
rect -11104 -2052 -5816 -1988
rect -5752 -2052 -5732 -1988
rect -11104 -2068 -5732 -2052
rect -11104 -2132 -5816 -2068
rect -5752 -2132 -5732 -2068
rect -11104 -2148 -5732 -2132
rect -11104 -2212 -5816 -2148
rect -5752 -2212 -5732 -2148
rect -11104 -2228 -5732 -2212
rect -11104 -2292 -5816 -2228
rect -5752 -2292 -5732 -2228
rect -11104 -2308 -5732 -2292
rect -11104 -2372 -5816 -2308
rect -5752 -2372 -5732 -2308
rect -11104 -2388 -5732 -2372
rect -11104 -2452 -5816 -2388
rect -5752 -2452 -5732 -2388
rect -11104 -2468 -5732 -2452
rect -11104 -2532 -5816 -2468
rect -5752 -2532 -5732 -2468
rect -11104 -2548 -5732 -2532
rect -11104 -2612 -5816 -2548
rect -5752 -2612 -5732 -2548
rect -11104 -2628 -5732 -2612
rect -11104 -2692 -5816 -2628
rect -5752 -2692 -5732 -2628
rect -11104 -2708 -5732 -2692
rect -11104 -2772 -5816 -2708
rect -5752 -2772 -5732 -2708
rect -11104 -2788 -5732 -2772
rect -11104 -2852 -5816 -2788
rect -5752 -2852 -5732 -2788
rect -11104 -2868 -5732 -2852
rect -11104 -2932 -5816 -2868
rect -5752 -2932 -5732 -2868
rect -11104 -2948 -5732 -2932
rect -11104 -3012 -5816 -2948
rect -5752 -3012 -5732 -2948
rect -11104 -3028 -5732 -3012
rect -11104 -3092 -5816 -3028
rect -5752 -3092 -5732 -3028
rect -11104 -3108 -5732 -3092
rect -11104 -3172 -5816 -3108
rect -5752 -3172 -5732 -3108
rect -11104 -3188 -5732 -3172
rect -11104 -3252 -5816 -3188
rect -5752 -3252 -5732 -3188
rect -11104 -3268 -5732 -3252
rect -11104 -3332 -5816 -3268
rect -5752 -3332 -5732 -3268
rect -11104 -3348 -5732 -3332
rect -11104 -3412 -5816 -3348
rect -5752 -3412 -5732 -3348
rect -11104 -3428 -5732 -3412
rect -11104 -3492 -5816 -3428
rect -5752 -3492 -5732 -3428
rect -11104 -3508 -5732 -3492
rect -11104 -3572 -5816 -3508
rect -5752 -3572 -5732 -3508
rect -11104 -3588 -5732 -3572
rect -11104 -3652 -5816 -3588
rect -5752 -3652 -5732 -3588
rect -11104 -3668 -5732 -3652
rect -11104 -3732 -5816 -3668
rect -5752 -3732 -5732 -3668
rect -11104 -3748 -5732 -3732
rect -11104 -3812 -5816 -3748
rect -5752 -3812 -5732 -3748
rect -11104 -3828 -5732 -3812
rect -11104 -3892 -5816 -3828
rect -5752 -3892 -5732 -3828
rect -11104 -3908 -5732 -3892
rect -11104 -3972 -5816 -3908
rect -5752 -3972 -5732 -3908
rect -11104 -3988 -5732 -3972
rect -11104 -4052 -5816 -3988
rect -5752 -4052 -5732 -3988
rect -11104 -4068 -5732 -4052
rect -11104 -4132 -5816 -4068
rect -5752 -4132 -5732 -4068
rect -11104 -4148 -5732 -4132
rect -11104 -4212 -5816 -4148
rect -5752 -4212 -5732 -4148
rect -11104 -4228 -5732 -4212
rect -11104 -4292 -5816 -4228
rect -5752 -4292 -5732 -4228
rect -11104 -4308 -5732 -4292
rect -11104 -4372 -5816 -4308
rect -5752 -4372 -5732 -4308
rect -11104 -4388 -5732 -4372
rect -11104 -4452 -5816 -4388
rect -5752 -4452 -5732 -4388
rect -11104 -4468 -5732 -4452
rect -11104 -4532 -5816 -4468
rect -5752 -4532 -5732 -4468
rect -11104 -4548 -5732 -4532
rect -11104 -4612 -5816 -4548
rect -5752 -4612 -5732 -4548
rect -11104 -4628 -5732 -4612
rect -11104 -4692 -5816 -4628
rect -5752 -4692 -5732 -4628
rect -11104 -4708 -5732 -4692
rect -11104 -4772 -5816 -4708
rect -5752 -4772 -5732 -4708
rect -11104 -4788 -5732 -4772
rect -11104 -4852 -5816 -4788
rect -5752 -4852 -5732 -4788
rect -11104 -4868 -5732 -4852
rect -11104 -4932 -5816 -4868
rect -5752 -4932 -5732 -4868
rect -11104 -4948 -5732 -4932
rect -11104 -5012 -5816 -4948
rect -5752 -5012 -5732 -4948
rect -11104 -5028 -5732 -5012
rect -11104 -5092 -5816 -5028
rect -5752 -5092 -5732 -5028
rect -11104 -5108 -5732 -5092
rect -11104 -5172 -5816 -5108
rect -5752 -5172 -5732 -5108
rect -11104 -5200 -5732 -5172
rect -5492 -148 -120 -120
rect -5492 -212 -204 -148
rect -140 -212 -120 -148
rect -5492 -228 -120 -212
rect -5492 -292 -204 -228
rect -140 -292 -120 -228
rect -5492 -308 -120 -292
rect -5492 -372 -204 -308
rect -140 -372 -120 -308
rect -5492 -388 -120 -372
rect -5492 -452 -204 -388
rect -140 -452 -120 -388
rect -5492 -468 -120 -452
rect -5492 -532 -204 -468
rect -140 -532 -120 -468
rect -5492 -548 -120 -532
rect -5492 -612 -204 -548
rect -140 -612 -120 -548
rect -5492 -628 -120 -612
rect -5492 -692 -204 -628
rect -140 -692 -120 -628
rect -5492 -708 -120 -692
rect -5492 -772 -204 -708
rect -140 -772 -120 -708
rect -5492 -788 -120 -772
rect -5492 -852 -204 -788
rect -140 -852 -120 -788
rect -5492 -868 -120 -852
rect -5492 -932 -204 -868
rect -140 -932 -120 -868
rect -5492 -948 -120 -932
rect -5492 -1012 -204 -948
rect -140 -1012 -120 -948
rect -5492 -1028 -120 -1012
rect -5492 -1092 -204 -1028
rect -140 -1092 -120 -1028
rect -5492 -1108 -120 -1092
rect -5492 -1172 -204 -1108
rect -140 -1172 -120 -1108
rect -5492 -1188 -120 -1172
rect -5492 -1252 -204 -1188
rect -140 -1252 -120 -1188
rect -5492 -1268 -120 -1252
rect -5492 -1332 -204 -1268
rect -140 -1332 -120 -1268
rect -5492 -1348 -120 -1332
rect -5492 -1412 -204 -1348
rect -140 -1412 -120 -1348
rect -5492 -1428 -120 -1412
rect -5492 -1492 -204 -1428
rect -140 -1492 -120 -1428
rect -5492 -1508 -120 -1492
rect -5492 -1572 -204 -1508
rect -140 -1572 -120 -1508
rect -5492 -1588 -120 -1572
rect -5492 -1652 -204 -1588
rect -140 -1652 -120 -1588
rect -5492 -1668 -120 -1652
rect -5492 -1732 -204 -1668
rect -140 -1732 -120 -1668
rect -5492 -1748 -120 -1732
rect -5492 -1812 -204 -1748
rect -140 -1812 -120 -1748
rect -5492 -1828 -120 -1812
rect -5492 -1892 -204 -1828
rect -140 -1892 -120 -1828
rect -5492 -1908 -120 -1892
rect -5492 -1972 -204 -1908
rect -140 -1972 -120 -1908
rect -5492 -1988 -120 -1972
rect -5492 -2052 -204 -1988
rect -140 -2052 -120 -1988
rect -5492 -2068 -120 -2052
rect -5492 -2132 -204 -2068
rect -140 -2132 -120 -2068
rect -5492 -2148 -120 -2132
rect -5492 -2212 -204 -2148
rect -140 -2212 -120 -2148
rect -5492 -2228 -120 -2212
rect -5492 -2292 -204 -2228
rect -140 -2292 -120 -2228
rect -5492 -2308 -120 -2292
rect -5492 -2372 -204 -2308
rect -140 -2372 -120 -2308
rect -5492 -2388 -120 -2372
rect -5492 -2452 -204 -2388
rect -140 -2452 -120 -2388
rect -5492 -2468 -120 -2452
rect -5492 -2532 -204 -2468
rect -140 -2532 -120 -2468
rect -5492 -2548 -120 -2532
rect -5492 -2612 -204 -2548
rect -140 -2612 -120 -2548
rect -5492 -2628 -120 -2612
rect -5492 -2692 -204 -2628
rect -140 -2692 -120 -2628
rect -5492 -2708 -120 -2692
rect -5492 -2772 -204 -2708
rect -140 -2772 -120 -2708
rect -5492 -2788 -120 -2772
rect -5492 -2852 -204 -2788
rect -140 -2852 -120 -2788
rect -5492 -2868 -120 -2852
rect -5492 -2932 -204 -2868
rect -140 -2932 -120 -2868
rect -5492 -2948 -120 -2932
rect -5492 -3012 -204 -2948
rect -140 -3012 -120 -2948
rect -5492 -3028 -120 -3012
rect -5492 -3092 -204 -3028
rect -140 -3092 -120 -3028
rect -5492 -3108 -120 -3092
rect -5492 -3172 -204 -3108
rect -140 -3172 -120 -3108
rect -5492 -3188 -120 -3172
rect -5492 -3252 -204 -3188
rect -140 -3252 -120 -3188
rect -5492 -3268 -120 -3252
rect -5492 -3332 -204 -3268
rect -140 -3332 -120 -3268
rect -5492 -3348 -120 -3332
rect -5492 -3412 -204 -3348
rect -140 -3412 -120 -3348
rect -5492 -3428 -120 -3412
rect -5492 -3492 -204 -3428
rect -140 -3492 -120 -3428
rect -5492 -3508 -120 -3492
rect -5492 -3572 -204 -3508
rect -140 -3572 -120 -3508
rect -5492 -3588 -120 -3572
rect -5492 -3652 -204 -3588
rect -140 -3652 -120 -3588
rect -5492 -3668 -120 -3652
rect -5492 -3732 -204 -3668
rect -140 -3732 -120 -3668
rect -5492 -3748 -120 -3732
rect -5492 -3812 -204 -3748
rect -140 -3812 -120 -3748
rect -5492 -3828 -120 -3812
rect -5492 -3892 -204 -3828
rect -140 -3892 -120 -3828
rect -5492 -3908 -120 -3892
rect -5492 -3972 -204 -3908
rect -140 -3972 -120 -3908
rect -5492 -3988 -120 -3972
rect -5492 -4052 -204 -3988
rect -140 -4052 -120 -3988
rect -5492 -4068 -120 -4052
rect -5492 -4132 -204 -4068
rect -140 -4132 -120 -4068
rect -5492 -4148 -120 -4132
rect -5492 -4212 -204 -4148
rect -140 -4212 -120 -4148
rect -5492 -4228 -120 -4212
rect -5492 -4292 -204 -4228
rect -140 -4292 -120 -4228
rect -5492 -4308 -120 -4292
rect -5492 -4372 -204 -4308
rect -140 -4372 -120 -4308
rect -5492 -4388 -120 -4372
rect -5492 -4452 -204 -4388
rect -140 -4452 -120 -4388
rect -5492 -4468 -120 -4452
rect -5492 -4532 -204 -4468
rect -140 -4532 -120 -4468
rect -5492 -4548 -120 -4532
rect -5492 -4612 -204 -4548
rect -140 -4612 -120 -4548
rect -5492 -4628 -120 -4612
rect -5492 -4692 -204 -4628
rect -140 -4692 -120 -4628
rect -5492 -4708 -120 -4692
rect -5492 -4772 -204 -4708
rect -140 -4772 -120 -4708
rect -5492 -4788 -120 -4772
rect -5492 -4852 -204 -4788
rect -140 -4852 -120 -4788
rect -5492 -4868 -120 -4852
rect -5492 -4932 -204 -4868
rect -140 -4932 -120 -4868
rect -5492 -4948 -120 -4932
rect -5492 -5012 -204 -4948
rect -140 -5012 -120 -4948
rect -5492 -5028 -120 -5012
rect -5492 -5092 -204 -5028
rect -140 -5092 -120 -5028
rect -5492 -5108 -120 -5092
rect -5492 -5172 -204 -5108
rect -140 -5172 -120 -5108
rect -5492 -5200 -120 -5172
rect 120 -148 5492 -120
rect 120 -212 5408 -148
rect 5472 -212 5492 -148
rect 120 -228 5492 -212
rect 120 -292 5408 -228
rect 5472 -292 5492 -228
rect 120 -308 5492 -292
rect 120 -372 5408 -308
rect 5472 -372 5492 -308
rect 120 -388 5492 -372
rect 120 -452 5408 -388
rect 5472 -452 5492 -388
rect 120 -468 5492 -452
rect 120 -532 5408 -468
rect 5472 -532 5492 -468
rect 120 -548 5492 -532
rect 120 -612 5408 -548
rect 5472 -612 5492 -548
rect 120 -628 5492 -612
rect 120 -692 5408 -628
rect 5472 -692 5492 -628
rect 120 -708 5492 -692
rect 120 -772 5408 -708
rect 5472 -772 5492 -708
rect 120 -788 5492 -772
rect 120 -852 5408 -788
rect 5472 -852 5492 -788
rect 120 -868 5492 -852
rect 120 -932 5408 -868
rect 5472 -932 5492 -868
rect 120 -948 5492 -932
rect 120 -1012 5408 -948
rect 5472 -1012 5492 -948
rect 120 -1028 5492 -1012
rect 120 -1092 5408 -1028
rect 5472 -1092 5492 -1028
rect 120 -1108 5492 -1092
rect 120 -1172 5408 -1108
rect 5472 -1172 5492 -1108
rect 120 -1188 5492 -1172
rect 120 -1252 5408 -1188
rect 5472 -1252 5492 -1188
rect 120 -1268 5492 -1252
rect 120 -1332 5408 -1268
rect 5472 -1332 5492 -1268
rect 120 -1348 5492 -1332
rect 120 -1412 5408 -1348
rect 5472 -1412 5492 -1348
rect 120 -1428 5492 -1412
rect 120 -1492 5408 -1428
rect 5472 -1492 5492 -1428
rect 120 -1508 5492 -1492
rect 120 -1572 5408 -1508
rect 5472 -1572 5492 -1508
rect 120 -1588 5492 -1572
rect 120 -1652 5408 -1588
rect 5472 -1652 5492 -1588
rect 120 -1668 5492 -1652
rect 120 -1732 5408 -1668
rect 5472 -1732 5492 -1668
rect 120 -1748 5492 -1732
rect 120 -1812 5408 -1748
rect 5472 -1812 5492 -1748
rect 120 -1828 5492 -1812
rect 120 -1892 5408 -1828
rect 5472 -1892 5492 -1828
rect 120 -1908 5492 -1892
rect 120 -1972 5408 -1908
rect 5472 -1972 5492 -1908
rect 120 -1988 5492 -1972
rect 120 -2052 5408 -1988
rect 5472 -2052 5492 -1988
rect 120 -2068 5492 -2052
rect 120 -2132 5408 -2068
rect 5472 -2132 5492 -2068
rect 120 -2148 5492 -2132
rect 120 -2212 5408 -2148
rect 5472 -2212 5492 -2148
rect 120 -2228 5492 -2212
rect 120 -2292 5408 -2228
rect 5472 -2292 5492 -2228
rect 120 -2308 5492 -2292
rect 120 -2372 5408 -2308
rect 5472 -2372 5492 -2308
rect 120 -2388 5492 -2372
rect 120 -2452 5408 -2388
rect 5472 -2452 5492 -2388
rect 120 -2468 5492 -2452
rect 120 -2532 5408 -2468
rect 5472 -2532 5492 -2468
rect 120 -2548 5492 -2532
rect 120 -2612 5408 -2548
rect 5472 -2612 5492 -2548
rect 120 -2628 5492 -2612
rect 120 -2692 5408 -2628
rect 5472 -2692 5492 -2628
rect 120 -2708 5492 -2692
rect 120 -2772 5408 -2708
rect 5472 -2772 5492 -2708
rect 120 -2788 5492 -2772
rect 120 -2852 5408 -2788
rect 5472 -2852 5492 -2788
rect 120 -2868 5492 -2852
rect 120 -2932 5408 -2868
rect 5472 -2932 5492 -2868
rect 120 -2948 5492 -2932
rect 120 -3012 5408 -2948
rect 5472 -3012 5492 -2948
rect 120 -3028 5492 -3012
rect 120 -3092 5408 -3028
rect 5472 -3092 5492 -3028
rect 120 -3108 5492 -3092
rect 120 -3172 5408 -3108
rect 5472 -3172 5492 -3108
rect 120 -3188 5492 -3172
rect 120 -3252 5408 -3188
rect 5472 -3252 5492 -3188
rect 120 -3268 5492 -3252
rect 120 -3332 5408 -3268
rect 5472 -3332 5492 -3268
rect 120 -3348 5492 -3332
rect 120 -3412 5408 -3348
rect 5472 -3412 5492 -3348
rect 120 -3428 5492 -3412
rect 120 -3492 5408 -3428
rect 5472 -3492 5492 -3428
rect 120 -3508 5492 -3492
rect 120 -3572 5408 -3508
rect 5472 -3572 5492 -3508
rect 120 -3588 5492 -3572
rect 120 -3652 5408 -3588
rect 5472 -3652 5492 -3588
rect 120 -3668 5492 -3652
rect 120 -3732 5408 -3668
rect 5472 -3732 5492 -3668
rect 120 -3748 5492 -3732
rect 120 -3812 5408 -3748
rect 5472 -3812 5492 -3748
rect 120 -3828 5492 -3812
rect 120 -3892 5408 -3828
rect 5472 -3892 5492 -3828
rect 120 -3908 5492 -3892
rect 120 -3972 5408 -3908
rect 5472 -3972 5492 -3908
rect 120 -3988 5492 -3972
rect 120 -4052 5408 -3988
rect 5472 -4052 5492 -3988
rect 120 -4068 5492 -4052
rect 120 -4132 5408 -4068
rect 5472 -4132 5492 -4068
rect 120 -4148 5492 -4132
rect 120 -4212 5408 -4148
rect 5472 -4212 5492 -4148
rect 120 -4228 5492 -4212
rect 120 -4292 5408 -4228
rect 5472 -4292 5492 -4228
rect 120 -4308 5492 -4292
rect 120 -4372 5408 -4308
rect 5472 -4372 5492 -4308
rect 120 -4388 5492 -4372
rect 120 -4452 5408 -4388
rect 5472 -4452 5492 -4388
rect 120 -4468 5492 -4452
rect 120 -4532 5408 -4468
rect 5472 -4532 5492 -4468
rect 120 -4548 5492 -4532
rect 120 -4612 5408 -4548
rect 5472 -4612 5492 -4548
rect 120 -4628 5492 -4612
rect 120 -4692 5408 -4628
rect 5472 -4692 5492 -4628
rect 120 -4708 5492 -4692
rect 120 -4772 5408 -4708
rect 5472 -4772 5492 -4708
rect 120 -4788 5492 -4772
rect 120 -4852 5408 -4788
rect 5472 -4852 5492 -4788
rect 120 -4868 5492 -4852
rect 120 -4932 5408 -4868
rect 5472 -4932 5492 -4868
rect 120 -4948 5492 -4932
rect 120 -5012 5408 -4948
rect 5472 -5012 5492 -4948
rect 120 -5028 5492 -5012
rect 120 -5092 5408 -5028
rect 5472 -5092 5492 -5028
rect 120 -5108 5492 -5092
rect 120 -5172 5408 -5108
rect 5472 -5172 5492 -5108
rect 120 -5200 5492 -5172
rect 5732 -148 11104 -120
rect 5732 -212 11020 -148
rect 11084 -212 11104 -148
rect 5732 -228 11104 -212
rect 5732 -292 11020 -228
rect 11084 -292 11104 -228
rect 5732 -308 11104 -292
rect 5732 -372 11020 -308
rect 11084 -372 11104 -308
rect 5732 -388 11104 -372
rect 5732 -452 11020 -388
rect 11084 -452 11104 -388
rect 5732 -468 11104 -452
rect 5732 -532 11020 -468
rect 11084 -532 11104 -468
rect 5732 -548 11104 -532
rect 5732 -612 11020 -548
rect 11084 -612 11104 -548
rect 5732 -628 11104 -612
rect 5732 -692 11020 -628
rect 11084 -692 11104 -628
rect 5732 -708 11104 -692
rect 5732 -772 11020 -708
rect 11084 -772 11104 -708
rect 5732 -788 11104 -772
rect 5732 -852 11020 -788
rect 11084 -852 11104 -788
rect 5732 -868 11104 -852
rect 5732 -932 11020 -868
rect 11084 -932 11104 -868
rect 5732 -948 11104 -932
rect 5732 -1012 11020 -948
rect 11084 -1012 11104 -948
rect 5732 -1028 11104 -1012
rect 5732 -1092 11020 -1028
rect 11084 -1092 11104 -1028
rect 5732 -1108 11104 -1092
rect 5732 -1172 11020 -1108
rect 11084 -1172 11104 -1108
rect 5732 -1188 11104 -1172
rect 5732 -1252 11020 -1188
rect 11084 -1252 11104 -1188
rect 5732 -1268 11104 -1252
rect 5732 -1332 11020 -1268
rect 11084 -1332 11104 -1268
rect 5732 -1348 11104 -1332
rect 5732 -1412 11020 -1348
rect 11084 -1412 11104 -1348
rect 5732 -1428 11104 -1412
rect 5732 -1492 11020 -1428
rect 11084 -1492 11104 -1428
rect 5732 -1508 11104 -1492
rect 5732 -1572 11020 -1508
rect 11084 -1572 11104 -1508
rect 5732 -1588 11104 -1572
rect 5732 -1652 11020 -1588
rect 11084 -1652 11104 -1588
rect 5732 -1668 11104 -1652
rect 5732 -1732 11020 -1668
rect 11084 -1732 11104 -1668
rect 5732 -1748 11104 -1732
rect 5732 -1812 11020 -1748
rect 11084 -1812 11104 -1748
rect 5732 -1828 11104 -1812
rect 5732 -1892 11020 -1828
rect 11084 -1892 11104 -1828
rect 5732 -1908 11104 -1892
rect 5732 -1972 11020 -1908
rect 11084 -1972 11104 -1908
rect 5732 -1988 11104 -1972
rect 5732 -2052 11020 -1988
rect 11084 -2052 11104 -1988
rect 5732 -2068 11104 -2052
rect 5732 -2132 11020 -2068
rect 11084 -2132 11104 -2068
rect 5732 -2148 11104 -2132
rect 5732 -2212 11020 -2148
rect 11084 -2212 11104 -2148
rect 5732 -2228 11104 -2212
rect 5732 -2292 11020 -2228
rect 11084 -2292 11104 -2228
rect 5732 -2308 11104 -2292
rect 5732 -2372 11020 -2308
rect 11084 -2372 11104 -2308
rect 5732 -2388 11104 -2372
rect 5732 -2452 11020 -2388
rect 11084 -2452 11104 -2388
rect 5732 -2468 11104 -2452
rect 5732 -2532 11020 -2468
rect 11084 -2532 11104 -2468
rect 5732 -2548 11104 -2532
rect 5732 -2612 11020 -2548
rect 11084 -2612 11104 -2548
rect 5732 -2628 11104 -2612
rect 5732 -2692 11020 -2628
rect 11084 -2692 11104 -2628
rect 5732 -2708 11104 -2692
rect 5732 -2772 11020 -2708
rect 11084 -2772 11104 -2708
rect 5732 -2788 11104 -2772
rect 5732 -2852 11020 -2788
rect 11084 -2852 11104 -2788
rect 5732 -2868 11104 -2852
rect 5732 -2932 11020 -2868
rect 11084 -2932 11104 -2868
rect 5732 -2948 11104 -2932
rect 5732 -3012 11020 -2948
rect 11084 -3012 11104 -2948
rect 5732 -3028 11104 -3012
rect 5732 -3092 11020 -3028
rect 11084 -3092 11104 -3028
rect 5732 -3108 11104 -3092
rect 5732 -3172 11020 -3108
rect 11084 -3172 11104 -3108
rect 5732 -3188 11104 -3172
rect 5732 -3252 11020 -3188
rect 11084 -3252 11104 -3188
rect 5732 -3268 11104 -3252
rect 5732 -3332 11020 -3268
rect 11084 -3332 11104 -3268
rect 5732 -3348 11104 -3332
rect 5732 -3412 11020 -3348
rect 11084 -3412 11104 -3348
rect 5732 -3428 11104 -3412
rect 5732 -3492 11020 -3428
rect 11084 -3492 11104 -3428
rect 5732 -3508 11104 -3492
rect 5732 -3572 11020 -3508
rect 11084 -3572 11104 -3508
rect 5732 -3588 11104 -3572
rect 5732 -3652 11020 -3588
rect 11084 -3652 11104 -3588
rect 5732 -3668 11104 -3652
rect 5732 -3732 11020 -3668
rect 11084 -3732 11104 -3668
rect 5732 -3748 11104 -3732
rect 5732 -3812 11020 -3748
rect 11084 -3812 11104 -3748
rect 5732 -3828 11104 -3812
rect 5732 -3892 11020 -3828
rect 11084 -3892 11104 -3828
rect 5732 -3908 11104 -3892
rect 5732 -3972 11020 -3908
rect 11084 -3972 11104 -3908
rect 5732 -3988 11104 -3972
rect 5732 -4052 11020 -3988
rect 11084 -4052 11104 -3988
rect 5732 -4068 11104 -4052
rect 5732 -4132 11020 -4068
rect 11084 -4132 11104 -4068
rect 5732 -4148 11104 -4132
rect 5732 -4212 11020 -4148
rect 11084 -4212 11104 -4148
rect 5732 -4228 11104 -4212
rect 5732 -4292 11020 -4228
rect 11084 -4292 11104 -4228
rect 5732 -4308 11104 -4292
rect 5732 -4372 11020 -4308
rect 11084 -4372 11104 -4308
rect 5732 -4388 11104 -4372
rect 5732 -4452 11020 -4388
rect 11084 -4452 11104 -4388
rect 5732 -4468 11104 -4452
rect 5732 -4532 11020 -4468
rect 11084 -4532 11104 -4468
rect 5732 -4548 11104 -4532
rect 5732 -4612 11020 -4548
rect 11084 -4612 11104 -4548
rect 5732 -4628 11104 -4612
rect 5732 -4692 11020 -4628
rect 11084 -4692 11104 -4628
rect 5732 -4708 11104 -4692
rect 5732 -4772 11020 -4708
rect 11084 -4772 11104 -4708
rect 5732 -4788 11104 -4772
rect 5732 -4852 11020 -4788
rect 11084 -4852 11104 -4788
rect 5732 -4868 11104 -4852
rect 5732 -4932 11020 -4868
rect 11084 -4932 11104 -4868
rect 5732 -4948 11104 -4932
rect 5732 -5012 11020 -4948
rect 11084 -5012 11104 -4948
rect 5732 -5028 11104 -5012
rect 5732 -5092 11020 -5028
rect 11084 -5092 11104 -5028
rect 5732 -5108 11104 -5092
rect 5732 -5172 11020 -5108
rect 11084 -5172 11104 -5108
rect 5732 -5200 11104 -5172
rect 11344 -148 16716 -120
rect 11344 -212 16632 -148
rect 16696 -212 16716 -148
rect 11344 -228 16716 -212
rect 11344 -292 16632 -228
rect 16696 -292 16716 -228
rect 11344 -308 16716 -292
rect 11344 -372 16632 -308
rect 16696 -372 16716 -308
rect 11344 -388 16716 -372
rect 11344 -452 16632 -388
rect 16696 -452 16716 -388
rect 11344 -468 16716 -452
rect 11344 -532 16632 -468
rect 16696 -532 16716 -468
rect 11344 -548 16716 -532
rect 11344 -612 16632 -548
rect 16696 -612 16716 -548
rect 11344 -628 16716 -612
rect 11344 -692 16632 -628
rect 16696 -692 16716 -628
rect 11344 -708 16716 -692
rect 11344 -772 16632 -708
rect 16696 -772 16716 -708
rect 11344 -788 16716 -772
rect 11344 -852 16632 -788
rect 16696 -852 16716 -788
rect 11344 -868 16716 -852
rect 11344 -932 16632 -868
rect 16696 -932 16716 -868
rect 11344 -948 16716 -932
rect 11344 -1012 16632 -948
rect 16696 -1012 16716 -948
rect 11344 -1028 16716 -1012
rect 11344 -1092 16632 -1028
rect 16696 -1092 16716 -1028
rect 11344 -1108 16716 -1092
rect 11344 -1172 16632 -1108
rect 16696 -1172 16716 -1108
rect 11344 -1188 16716 -1172
rect 11344 -1252 16632 -1188
rect 16696 -1252 16716 -1188
rect 11344 -1268 16716 -1252
rect 11344 -1332 16632 -1268
rect 16696 -1332 16716 -1268
rect 11344 -1348 16716 -1332
rect 11344 -1412 16632 -1348
rect 16696 -1412 16716 -1348
rect 11344 -1428 16716 -1412
rect 11344 -1492 16632 -1428
rect 16696 -1492 16716 -1428
rect 11344 -1508 16716 -1492
rect 11344 -1572 16632 -1508
rect 16696 -1572 16716 -1508
rect 11344 -1588 16716 -1572
rect 11344 -1652 16632 -1588
rect 16696 -1652 16716 -1588
rect 11344 -1668 16716 -1652
rect 11344 -1732 16632 -1668
rect 16696 -1732 16716 -1668
rect 11344 -1748 16716 -1732
rect 11344 -1812 16632 -1748
rect 16696 -1812 16716 -1748
rect 11344 -1828 16716 -1812
rect 11344 -1892 16632 -1828
rect 16696 -1892 16716 -1828
rect 11344 -1908 16716 -1892
rect 11344 -1972 16632 -1908
rect 16696 -1972 16716 -1908
rect 11344 -1988 16716 -1972
rect 11344 -2052 16632 -1988
rect 16696 -2052 16716 -1988
rect 11344 -2068 16716 -2052
rect 11344 -2132 16632 -2068
rect 16696 -2132 16716 -2068
rect 11344 -2148 16716 -2132
rect 11344 -2212 16632 -2148
rect 16696 -2212 16716 -2148
rect 11344 -2228 16716 -2212
rect 11344 -2292 16632 -2228
rect 16696 -2292 16716 -2228
rect 11344 -2308 16716 -2292
rect 11344 -2372 16632 -2308
rect 16696 -2372 16716 -2308
rect 11344 -2388 16716 -2372
rect 11344 -2452 16632 -2388
rect 16696 -2452 16716 -2388
rect 11344 -2468 16716 -2452
rect 11344 -2532 16632 -2468
rect 16696 -2532 16716 -2468
rect 11344 -2548 16716 -2532
rect 11344 -2612 16632 -2548
rect 16696 -2612 16716 -2548
rect 11344 -2628 16716 -2612
rect 11344 -2692 16632 -2628
rect 16696 -2692 16716 -2628
rect 11344 -2708 16716 -2692
rect 11344 -2772 16632 -2708
rect 16696 -2772 16716 -2708
rect 11344 -2788 16716 -2772
rect 11344 -2852 16632 -2788
rect 16696 -2852 16716 -2788
rect 11344 -2868 16716 -2852
rect 11344 -2932 16632 -2868
rect 16696 -2932 16716 -2868
rect 11344 -2948 16716 -2932
rect 11344 -3012 16632 -2948
rect 16696 -3012 16716 -2948
rect 11344 -3028 16716 -3012
rect 11344 -3092 16632 -3028
rect 16696 -3092 16716 -3028
rect 11344 -3108 16716 -3092
rect 11344 -3172 16632 -3108
rect 16696 -3172 16716 -3108
rect 11344 -3188 16716 -3172
rect 11344 -3252 16632 -3188
rect 16696 -3252 16716 -3188
rect 11344 -3268 16716 -3252
rect 11344 -3332 16632 -3268
rect 16696 -3332 16716 -3268
rect 11344 -3348 16716 -3332
rect 11344 -3412 16632 -3348
rect 16696 -3412 16716 -3348
rect 11344 -3428 16716 -3412
rect 11344 -3492 16632 -3428
rect 16696 -3492 16716 -3428
rect 11344 -3508 16716 -3492
rect 11344 -3572 16632 -3508
rect 16696 -3572 16716 -3508
rect 11344 -3588 16716 -3572
rect 11344 -3652 16632 -3588
rect 16696 -3652 16716 -3588
rect 11344 -3668 16716 -3652
rect 11344 -3732 16632 -3668
rect 16696 -3732 16716 -3668
rect 11344 -3748 16716 -3732
rect 11344 -3812 16632 -3748
rect 16696 -3812 16716 -3748
rect 11344 -3828 16716 -3812
rect 11344 -3892 16632 -3828
rect 16696 -3892 16716 -3828
rect 11344 -3908 16716 -3892
rect 11344 -3972 16632 -3908
rect 16696 -3972 16716 -3908
rect 11344 -3988 16716 -3972
rect 11344 -4052 16632 -3988
rect 16696 -4052 16716 -3988
rect 11344 -4068 16716 -4052
rect 11344 -4132 16632 -4068
rect 16696 -4132 16716 -4068
rect 11344 -4148 16716 -4132
rect 11344 -4212 16632 -4148
rect 16696 -4212 16716 -4148
rect 11344 -4228 16716 -4212
rect 11344 -4292 16632 -4228
rect 16696 -4292 16716 -4228
rect 11344 -4308 16716 -4292
rect 11344 -4372 16632 -4308
rect 16696 -4372 16716 -4308
rect 11344 -4388 16716 -4372
rect 11344 -4452 16632 -4388
rect 16696 -4452 16716 -4388
rect 11344 -4468 16716 -4452
rect 11344 -4532 16632 -4468
rect 16696 -4532 16716 -4468
rect 11344 -4548 16716 -4532
rect 11344 -4612 16632 -4548
rect 16696 -4612 16716 -4548
rect 11344 -4628 16716 -4612
rect 11344 -4692 16632 -4628
rect 16696 -4692 16716 -4628
rect 11344 -4708 16716 -4692
rect 11344 -4772 16632 -4708
rect 16696 -4772 16716 -4708
rect 11344 -4788 16716 -4772
rect 11344 -4852 16632 -4788
rect 16696 -4852 16716 -4788
rect 11344 -4868 16716 -4852
rect 11344 -4932 16632 -4868
rect 16696 -4932 16716 -4868
rect 11344 -4948 16716 -4932
rect 11344 -5012 16632 -4948
rect 16696 -5012 16716 -4948
rect 11344 -5028 16716 -5012
rect 11344 -5092 16632 -5028
rect 16696 -5092 16716 -5028
rect 11344 -5108 16716 -5092
rect 11344 -5172 16632 -5108
rect 16696 -5172 16716 -5108
rect 11344 -5200 16716 -5172
rect 16956 -148 22328 -120
rect 16956 -212 22244 -148
rect 22308 -212 22328 -148
rect 16956 -228 22328 -212
rect 16956 -292 22244 -228
rect 22308 -292 22328 -228
rect 16956 -308 22328 -292
rect 16956 -372 22244 -308
rect 22308 -372 22328 -308
rect 16956 -388 22328 -372
rect 16956 -452 22244 -388
rect 22308 -452 22328 -388
rect 16956 -468 22328 -452
rect 16956 -532 22244 -468
rect 22308 -532 22328 -468
rect 16956 -548 22328 -532
rect 16956 -612 22244 -548
rect 22308 -612 22328 -548
rect 16956 -628 22328 -612
rect 16956 -692 22244 -628
rect 22308 -692 22328 -628
rect 16956 -708 22328 -692
rect 16956 -772 22244 -708
rect 22308 -772 22328 -708
rect 16956 -788 22328 -772
rect 16956 -852 22244 -788
rect 22308 -852 22328 -788
rect 16956 -868 22328 -852
rect 16956 -932 22244 -868
rect 22308 -932 22328 -868
rect 16956 -948 22328 -932
rect 16956 -1012 22244 -948
rect 22308 -1012 22328 -948
rect 16956 -1028 22328 -1012
rect 16956 -1092 22244 -1028
rect 22308 -1092 22328 -1028
rect 16956 -1108 22328 -1092
rect 16956 -1172 22244 -1108
rect 22308 -1172 22328 -1108
rect 16956 -1188 22328 -1172
rect 16956 -1252 22244 -1188
rect 22308 -1252 22328 -1188
rect 16956 -1268 22328 -1252
rect 16956 -1332 22244 -1268
rect 22308 -1332 22328 -1268
rect 16956 -1348 22328 -1332
rect 16956 -1412 22244 -1348
rect 22308 -1412 22328 -1348
rect 16956 -1428 22328 -1412
rect 16956 -1492 22244 -1428
rect 22308 -1492 22328 -1428
rect 16956 -1508 22328 -1492
rect 16956 -1572 22244 -1508
rect 22308 -1572 22328 -1508
rect 16956 -1588 22328 -1572
rect 16956 -1652 22244 -1588
rect 22308 -1652 22328 -1588
rect 16956 -1668 22328 -1652
rect 16956 -1732 22244 -1668
rect 22308 -1732 22328 -1668
rect 16956 -1748 22328 -1732
rect 16956 -1812 22244 -1748
rect 22308 -1812 22328 -1748
rect 16956 -1828 22328 -1812
rect 16956 -1892 22244 -1828
rect 22308 -1892 22328 -1828
rect 16956 -1908 22328 -1892
rect 16956 -1972 22244 -1908
rect 22308 -1972 22328 -1908
rect 16956 -1988 22328 -1972
rect 16956 -2052 22244 -1988
rect 22308 -2052 22328 -1988
rect 16956 -2068 22328 -2052
rect 16956 -2132 22244 -2068
rect 22308 -2132 22328 -2068
rect 16956 -2148 22328 -2132
rect 16956 -2212 22244 -2148
rect 22308 -2212 22328 -2148
rect 16956 -2228 22328 -2212
rect 16956 -2292 22244 -2228
rect 22308 -2292 22328 -2228
rect 16956 -2308 22328 -2292
rect 16956 -2372 22244 -2308
rect 22308 -2372 22328 -2308
rect 16956 -2388 22328 -2372
rect 16956 -2452 22244 -2388
rect 22308 -2452 22328 -2388
rect 16956 -2468 22328 -2452
rect 16956 -2532 22244 -2468
rect 22308 -2532 22328 -2468
rect 16956 -2548 22328 -2532
rect 16956 -2612 22244 -2548
rect 22308 -2612 22328 -2548
rect 16956 -2628 22328 -2612
rect 16956 -2692 22244 -2628
rect 22308 -2692 22328 -2628
rect 16956 -2708 22328 -2692
rect 16956 -2772 22244 -2708
rect 22308 -2772 22328 -2708
rect 16956 -2788 22328 -2772
rect 16956 -2852 22244 -2788
rect 22308 -2852 22328 -2788
rect 16956 -2868 22328 -2852
rect 16956 -2932 22244 -2868
rect 22308 -2932 22328 -2868
rect 16956 -2948 22328 -2932
rect 16956 -3012 22244 -2948
rect 22308 -3012 22328 -2948
rect 16956 -3028 22328 -3012
rect 16956 -3092 22244 -3028
rect 22308 -3092 22328 -3028
rect 16956 -3108 22328 -3092
rect 16956 -3172 22244 -3108
rect 22308 -3172 22328 -3108
rect 16956 -3188 22328 -3172
rect 16956 -3252 22244 -3188
rect 22308 -3252 22328 -3188
rect 16956 -3268 22328 -3252
rect 16956 -3332 22244 -3268
rect 22308 -3332 22328 -3268
rect 16956 -3348 22328 -3332
rect 16956 -3412 22244 -3348
rect 22308 -3412 22328 -3348
rect 16956 -3428 22328 -3412
rect 16956 -3492 22244 -3428
rect 22308 -3492 22328 -3428
rect 16956 -3508 22328 -3492
rect 16956 -3572 22244 -3508
rect 22308 -3572 22328 -3508
rect 16956 -3588 22328 -3572
rect 16956 -3652 22244 -3588
rect 22308 -3652 22328 -3588
rect 16956 -3668 22328 -3652
rect 16956 -3732 22244 -3668
rect 22308 -3732 22328 -3668
rect 16956 -3748 22328 -3732
rect 16956 -3812 22244 -3748
rect 22308 -3812 22328 -3748
rect 16956 -3828 22328 -3812
rect 16956 -3892 22244 -3828
rect 22308 -3892 22328 -3828
rect 16956 -3908 22328 -3892
rect 16956 -3972 22244 -3908
rect 22308 -3972 22328 -3908
rect 16956 -3988 22328 -3972
rect 16956 -4052 22244 -3988
rect 22308 -4052 22328 -3988
rect 16956 -4068 22328 -4052
rect 16956 -4132 22244 -4068
rect 22308 -4132 22328 -4068
rect 16956 -4148 22328 -4132
rect 16956 -4212 22244 -4148
rect 22308 -4212 22328 -4148
rect 16956 -4228 22328 -4212
rect 16956 -4292 22244 -4228
rect 22308 -4292 22328 -4228
rect 16956 -4308 22328 -4292
rect 16956 -4372 22244 -4308
rect 22308 -4372 22328 -4308
rect 16956 -4388 22328 -4372
rect 16956 -4452 22244 -4388
rect 22308 -4452 22328 -4388
rect 16956 -4468 22328 -4452
rect 16956 -4532 22244 -4468
rect 22308 -4532 22328 -4468
rect 16956 -4548 22328 -4532
rect 16956 -4612 22244 -4548
rect 22308 -4612 22328 -4548
rect 16956 -4628 22328 -4612
rect 16956 -4692 22244 -4628
rect 22308 -4692 22328 -4628
rect 16956 -4708 22328 -4692
rect 16956 -4772 22244 -4708
rect 22308 -4772 22328 -4708
rect 16956 -4788 22328 -4772
rect 16956 -4852 22244 -4788
rect 22308 -4852 22328 -4788
rect 16956 -4868 22328 -4852
rect 16956 -4932 22244 -4868
rect 22308 -4932 22328 -4868
rect 16956 -4948 22328 -4932
rect 16956 -5012 22244 -4948
rect 22308 -5012 22328 -4948
rect 16956 -5028 22328 -5012
rect 16956 -5092 22244 -5028
rect 22308 -5092 22328 -5028
rect 16956 -5108 22328 -5092
rect 16956 -5172 22244 -5108
rect 22308 -5172 22328 -5108
rect 16956 -5200 22328 -5172
rect 22568 -148 27940 -120
rect 22568 -212 27856 -148
rect 27920 -212 27940 -148
rect 22568 -228 27940 -212
rect 22568 -292 27856 -228
rect 27920 -292 27940 -228
rect 22568 -308 27940 -292
rect 22568 -372 27856 -308
rect 27920 -372 27940 -308
rect 22568 -388 27940 -372
rect 22568 -452 27856 -388
rect 27920 -452 27940 -388
rect 22568 -468 27940 -452
rect 22568 -532 27856 -468
rect 27920 -532 27940 -468
rect 22568 -548 27940 -532
rect 22568 -612 27856 -548
rect 27920 -612 27940 -548
rect 22568 -628 27940 -612
rect 22568 -692 27856 -628
rect 27920 -692 27940 -628
rect 22568 -708 27940 -692
rect 22568 -772 27856 -708
rect 27920 -772 27940 -708
rect 22568 -788 27940 -772
rect 22568 -852 27856 -788
rect 27920 -852 27940 -788
rect 22568 -868 27940 -852
rect 22568 -932 27856 -868
rect 27920 -932 27940 -868
rect 22568 -948 27940 -932
rect 22568 -1012 27856 -948
rect 27920 -1012 27940 -948
rect 22568 -1028 27940 -1012
rect 22568 -1092 27856 -1028
rect 27920 -1092 27940 -1028
rect 22568 -1108 27940 -1092
rect 22568 -1172 27856 -1108
rect 27920 -1172 27940 -1108
rect 22568 -1188 27940 -1172
rect 22568 -1252 27856 -1188
rect 27920 -1252 27940 -1188
rect 22568 -1268 27940 -1252
rect 22568 -1332 27856 -1268
rect 27920 -1332 27940 -1268
rect 22568 -1348 27940 -1332
rect 22568 -1412 27856 -1348
rect 27920 -1412 27940 -1348
rect 22568 -1428 27940 -1412
rect 22568 -1492 27856 -1428
rect 27920 -1492 27940 -1428
rect 22568 -1508 27940 -1492
rect 22568 -1572 27856 -1508
rect 27920 -1572 27940 -1508
rect 22568 -1588 27940 -1572
rect 22568 -1652 27856 -1588
rect 27920 -1652 27940 -1588
rect 22568 -1668 27940 -1652
rect 22568 -1732 27856 -1668
rect 27920 -1732 27940 -1668
rect 22568 -1748 27940 -1732
rect 22568 -1812 27856 -1748
rect 27920 -1812 27940 -1748
rect 22568 -1828 27940 -1812
rect 22568 -1892 27856 -1828
rect 27920 -1892 27940 -1828
rect 22568 -1908 27940 -1892
rect 22568 -1972 27856 -1908
rect 27920 -1972 27940 -1908
rect 22568 -1988 27940 -1972
rect 22568 -2052 27856 -1988
rect 27920 -2052 27940 -1988
rect 22568 -2068 27940 -2052
rect 22568 -2132 27856 -2068
rect 27920 -2132 27940 -2068
rect 22568 -2148 27940 -2132
rect 22568 -2212 27856 -2148
rect 27920 -2212 27940 -2148
rect 22568 -2228 27940 -2212
rect 22568 -2292 27856 -2228
rect 27920 -2292 27940 -2228
rect 22568 -2308 27940 -2292
rect 22568 -2372 27856 -2308
rect 27920 -2372 27940 -2308
rect 22568 -2388 27940 -2372
rect 22568 -2452 27856 -2388
rect 27920 -2452 27940 -2388
rect 22568 -2468 27940 -2452
rect 22568 -2532 27856 -2468
rect 27920 -2532 27940 -2468
rect 22568 -2548 27940 -2532
rect 22568 -2612 27856 -2548
rect 27920 -2612 27940 -2548
rect 22568 -2628 27940 -2612
rect 22568 -2692 27856 -2628
rect 27920 -2692 27940 -2628
rect 22568 -2708 27940 -2692
rect 22568 -2772 27856 -2708
rect 27920 -2772 27940 -2708
rect 22568 -2788 27940 -2772
rect 22568 -2852 27856 -2788
rect 27920 -2852 27940 -2788
rect 22568 -2868 27940 -2852
rect 22568 -2932 27856 -2868
rect 27920 -2932 27940 -2868
rect 22568 -2948 27940 -2932
rect 22568 -3012 27856 -2948
rect 27920 -3012 27940 -2948
rect 22568 -3028 27940 -3012
rect 22568 -3092 27856 -3028
rect 27920 -3092 27940 -3028
rect 22568 -3108 27940 -3092
rect 22568 -3172 27856 -3108
rect 27920 -3172 27940 -3108
rect 22568 -3188 27940 -3172
rect 22568 -3252 27856 -3188
rect 27920 -3252 27940 -3188
rect 22568 -3268 27940 -3252
rect 22568 -3332 27856 -3268
rect 27920 -3332 27940 -3268
rect 22568 -3348 27940 -3332
rect 22568 -3412 27856 -3348
rect 27920 -3412 27940 -3348
rect 22568 -3428 27940 -3412
rect 22568 -3492 27856 -3428
rect 27920 -3492 27940 -3428
rect 22568 -3508 27940 -3492
rect 22568 -3572 27856 -3508
rect 27920 -3572 27940 -3508
rect 22568 -3588 27940 -3572
rect 22568 -3652 27856 -3588
rect 27920 -3652 27940 -3588
rect 22568 -3668 27940 -3652
rect 22568 -3732 27856 -3668
rect 27920 -3732 27940 -3668
rect 22568 -3748 27940 -3732
rect 22568 -3812 27856 -3748
rect 27920 -3812 27940 -3748
rect 22568 -3828 27940 -3812
rect 22568 -3892 27856 -3828
rect 27920 -3892 27940 -3828
rect 22568 -3908 27940 -3892
rect 22568 -3972 27856 -3908
rect 27920 -3972 27940 -3908
rect 22568 -3988 27940 -3972
rect 22568 -4052 27856 -3988
rect 27920 -4052 27940 -3988
rect 22568 -4068 27940 -4052
rect 22568 -4132 27856 -4068
rect 27920 -4132 27940 -4068
rect 22568 -4148 27940 -4132
rect 22568 -4212 27856 -4148
rect 27920 -4212 27940 -4148
rect 22568 -4228 27940 -4212
rect 22568 -4292 27856 -4228
rect 27920 -4292 27940 -4228
rect 22568 -4308 27940 -4292
rect 22568 -4372 27856 -4308
rect 27920 -4372 27940 -4308
rect 22568 -4388 27940 -4372
rect 22568 -4452 27856 -4388
rect 27920 -4452 27940 -4388
rect 22568 -4468 27940 -4452
rect 22568 -4532 27856 -4468
rect 27920 -4532 27940 -4468
rect 22568 -4548 27940 -4532
rect 22568 -4612 27856 -4548
rect 27920 -4612 27940 -4548
rect 22568 -4628 27940 -4612
rect 22568 -4692 27856 -4628
rect 27920 -4692 27940 -4628
rect 22568 -4708 27940 -4692
rect 22568 -4772 27856 -4708
rect 27920 -4772 27940 -4708
rect 22568 -4788 27940 -4772
rect 22568 -4852 27856 -4788
rect 27920 -4852 27940 -4788
rect 22568 -4868 27940 -4852
rect 22568 -4932 27856 -4868
rect 27920 -4932 27940 -4868
rect 22568 -4948 27940 -4932
rect 22568 -5012 27856 -4948
rect 27920 -5012 27940 -4948
rect 22568 -5028 27940 -5012
rect 22568 -5092 27856 -5028
rect 27920 -5092 27940 -5028
rect 22568 -5108 27940 -5092
rect 22568 -5172 27856 -5108
rect 27920 -5172 27940 -5108
rect 22568 -5200 27940 -5172
rect 28180 -148 33552 -120
rect 28180 -212 33468 -148
rect 33532 -212 33552 -148
rect 28180 -228 33552 -212
rect 28180 -292 33468 -228
rect 33532 -292 33552 -228
rect 28180 -308 33552 -292
rect 28180 -372 33468 -308
rect 33532 -372 33552 -308
rect 28180 -388 33552 -372
rect 28180 -452 33468 -388
rect 33532 -452 33552 -388
rect 28180 -468 33552 -452
rect 28180 -532 33468 -468
rect 33532 -532 33552 -468
rect 28180 -548 33552 -532
rect 28180 -612 33468 -548
rect 33532 -612 33552 -548
rect 28180 -628 33552 -612
rect 28180 -692 33468 -628
rect 33532 -692 33552 -628
rect 28180 -708 33552 -692
rect 28180 -772 33468 -708
rect 33532 -772 33552 -708
rect 28180 -788 33552 -772
rect 28180 -852 33468 -788
rect 33532 -852 33552 -788
rect 28180 -868 33552 -852
rect 28180 -932 33468 -868
rect 33532 -932 33552 -868
rect 28180 -948 33552 -932
rect 28180 -1012 33468 -948
rect 33532 -1012 33552 -948
rect 28180 -1028 33552 -1012
rect 28180 -1092 33468 -1028
rect 33532 -1092 33552 -1028
rect 28180 -1108 33552 -1092
rect 28180 -1172 33468 -1108
rect 33532 -1172 33552 -1108
rect 28180 -1188 33552 -1172
rect 28180 -1252 33468 -1188
rect 33532 -1252 33552 -1188
rect 28180 -1268 33552 -1252
rect 28180 -1332 33468 -1268
rect 33532 -1332 33552 -1268
rect 28180 -1348 33552 -1332
rect 28180 -1412 33468 -1348
rect 33532 -1412 33552 -1348
rect 28180 -1428 33552 -1412
rect 28180 -1492 33468 -1428
rect 33532 -1492 33552 -1428
rect 28180 -1508 33552 -1492
rect 28180 -1572 33468 -1508
rect 33532 -1572 33552 -1508
rect 28180 -1588 33552 -1572
rect 28180 -1652 33468 -1588
rect 33532 -1652 33552 -1588
rect 28180 -1668 33552 -1652
rect 28180 -1732 33468 -1668
rect 33532 -1732 33552 -1668
rect 28180 -1748 33552 -1732
rect 28180 -1812 33468 -1748
rect 33532 -1812 33552 -1748
rect 28180 -1828 33552 -1812
rect 28180 -1892 33468 -1828
rect 33532 -1892 33552 -1828
rect 28180 -1908 33552 -1892
rect 28180 -1972 33468 -1908
rect 33532 -1972 33552 -1908
rect 28180 -1988 33552 -1972
rect 28180 -2052 33468 -1988
rect 33532 -2052 33552 -1988
rect 28180 -2068 33552 -2052
rect 28180 -2132 33468 -2068
rect 33532 -2132 33552 -2068
rect 28180 -2148 33552 -2132
rect 28180 -2212 33468 -2148
rect 33532 -2212 33552 -2148
rect 28180 -2228 33552 -2212
rect 28180 -2292 33468 -2228
rect 33532 -2292 33552 -2228
rect 28180 -2308 33552 -2292
rect 28180 -2372 33468 -2308
rect 33532 -2372 33552 -2308
rect 28180 -2388 33552 -2372
rect 28180 -2452 33468 -2388
rect 33532 -2452 33552 -2388
rect 28180 -2468 33552 -2452
rect 28180 -2532 33468 -2468
rect 33532 -2532 33552 -2468
rect 28180 -2548 33552 -2532
rect 28180 -2612 33468 -2548
rect 33532 -2612 33552 -2548
rect 28180 -2628 33552 -2612
rect 28180 -2692 33468 -2628
rect 33532 -2692 33552 -2628
rect 28180 -2708 33552 -2692
rect 28180 -2772 33468 -2708
rect 33532 -2772 33552 -2708
rect 28180 -2788 33552 -2772
rect 28180 -2852 33468 -2788
rect 33532 -2852 33552 -2788
rect 28180 -2868 33552 -2852
rect 28180 -2932 33468 -2868
rect 33532 -2932 33552 -2868
rect 28180 -2948 33552 -2932
rect 28180 -3012 33468 -2948
rect 33532 -3012 33552 -2948
rect 28180 -3028 33552 -3012
rect 28180 -3092 33468 -3028
rect 33532 -3092 33552 -3028
rect 28180 -3108 33552 -3092
rect 28180 -3172 33468 -3108
rect 33532 -3172 33552 -3108
rect 28180 -3188 33552 -3172
rect 28180 -3252 33468 -3188
rect 33532 -3252 33552 -3188
rect 28180 -3268 33552 -3252
rect 28180 -3332 33468 -3268
rect 33532 -3332 33552 -3268
rect 28180 -3348 33552 -3332
rect 28180 -3412 33468 -3348
rect 33532 -3412 33552 -3348
rect 28180 -3428 33552 -3412
rect 28180 -3492 33468 -3428
rect 33532 -3492 33552 -3428
rect 28180 -3508 33552 -3492
rect 28180 -3572 33468 -3508
rect 33532 -3572 33552 -3508
rect 28180 -3588 33552 -3572
rect 28180 -3652 33468 -3588
rect 33532 -3652 33552 -3588
rect 28180 -3668 33552 -3652
rect 28180 -3732 33468 -3668
rect 33532 -3732 33552 -3668
rect 28180 -3748 33552 -3732
rect 28180 -3812 33468 -3748
rect 33532 -3812 33552 -3748
rect 28180 -3828 33552 -3812
rect 28180 -3892 33468 -3828
rect 33532 -3892 33552 -3828
rect 28180 -3908 33552 -3892
rect 28180 -3972 33468 -3908
rect 33532 -3972 33552 -3908
rect 28180 -3988 33552 -3972
rect 28180 -4052 33468 -3988
rect 33532 -4052 33552 -3988
rect 28180 -4068 33552 -4052
rect 28180 -4132 33468 -4068
rect 33532 -4132 33552 -4068
rect 28180 -4148 33552 -4132
rect 28180 -4212 33468 -4148
rect 33532 -4212 33552 -4148
rect 28180 -4228 33552 -4212
rect 28180 -4292 33468 -4228
rect 33532 -4292 33552 -4228
rect 28180 -4308 33552 -4292
rect 28180 -4372 33468 -4308
rect 33532 -4372 33552 -4308
rect 28180 -4388 33552 -4372
rect 28180 -4452 33468 -4388
rect 33532 -4452 33552 -4388
rect 28180 -4468 33552 -4452
rect 28180 -4532 33468 -4468
rect 33532 -4532 33552 -4468
rect 28180 -4548 33552 -4532
rect 28180 -4612 33468 -4548
rect 33532 -4612 33552 -4548
rect 28180 -4628 33552 -4612
rect 28180 -4692 33468 -4628
rect 33532 -4692 33552 -4628
rect 28180 -4708 33552 -4692
rect 28180 -4772 33468 -4708
rect 33532 -4772 33552 -4708
rect 28180 -4788 33552 -4772
rect 28180 -4852 33468 -4788
rect 33532 -4852 33552 -4788
rect 28180 -4868 33552 -4852
rect 28180 -4932 33468 -4868
rect 33532 -4932 33552 -4868
rect 28180 -4948 33552 -4932
rect 28180 -5012 33468 -4948
rect 33532 -5012 33552 -4948
rect 28180 -5028 33552 -5012
rect 28180 -5092 33468 -5028
rect 33532 -5092 33552 -5028
rect 28180 -5108 33552 -5092
rect 28180 -5172 33468 -5108
rect 33532 -5172 33552 -5108
rect 28180 -5200 33552 -5172
rect 33792 -148 39164 -120
rect 33792 -212 39080 -148
rect 39144 -212 39164 -148
rect 33792 -228 39164 -212
rect 33792 -292 39080 -228
rect 39144 -292 39164 -228
rect 33792 -308 39164 -292
rect 33792 -372 39080 -308
rect 39144 -372 39164 -308
rect 33792 -388 39164 -372
rect 33792 -452 39080 -388
rect 39144 -452 39164 -388
rect 33792 -468 39164 -452
rect 33792 -532 39080 -468
rect 39144 -532 39164 -468
rect 33792 -548 39164 -532
rect 33792 -612 39080 -548
rect 39144 -612 39164 -548
rect 33792 -628 39164 -612
rect 33792 -692 39080 -628
rect 39144 -692 39164 -628
rect 33792 -708 39164 -692
rect 33792 -772 39080 -708
rect 39144 -772 39164 -708
rect 33792 -788 39164 -772
rect 33792 -852 39080 -788
rect 39144 -852 39164 -788
rect 33792 -868 39164 -852
rect 33792 -932 39080 -868
rect 39144 -932 39164 -868
rect 33792 -948 39164 -932
rect 33792 -1012 39080 -948
rect 39144 -1012 39164 -948
rect 33792 -1028 39164 -1012
rect 33792 -1092 39080 -1028
rect 39144 -1092 39164 -1028
rect 33792 -1108 39164 -1092
rect 33792 -1172 39080 -1108
rect 39144 -1172 39164 -1108
rect 33792 -1188 39164 -1172
rect 33792 -1252 39080 -1188
rect 39144 -1252 39164 -1188
rect 33792 -1268 39164 -1252
rect 33792 -1332 39080 -1268
rect 39144 -1332 39164 -1268
rect 33792 -1348 39164 -1332
rect 33792 -1412 39080 -1348
rect 39144 -1412 39164 -1348
rect 33792 -1428 39164 -1412
rect 33792 -1492 39080 -1428
rect 39144 -1492 39164 -1428
rect 33792 -1508 39164 -1492
rect 33792 -1572 39080 -1508
rect 39144 -1572 39164 -1508
rect 33792 -1588 39164 -1572
rect 33792 -1652 39080 -1588
rect 39144 -1652 39164 -1588
rect 33792 -1668 39164 -1652
rect 33792 -1732 39080 -1668
rect 39144 -1732 39164 -1668
rect 33792 -1748 39164 -1732
rect 33792 -1812 39080 -1748
rect 39144 -1812 39164 -1748
rect 33792 -1828 39164 -1812
rect 33792 -1892 39080 -1828
rect 39144 -1892 39164 -1828
rect 33792 -1908 39164 -1892
rect 33792 -1972 39080 -1908
rect 39144 -1972 39164 -1908
rect 33792 -1988 39164 -1972
rect 33792 -2052 39080 -1988
rect 39144 -2052 39164 -1988
rect 33792 -2068 39164 -2052
rect 33792 -2132 39080 -2068
rect 39144 -2132 39164 -2068
rect 33792 -2148 39164 -2132
rect 33792 -2212 39080 -2148
rect 39144 -2212 39164 -2148
rect 33792 -2228 39164 -2212
rect 33792 -2292 39080 -2228
rect 39144 -2292 39164 -2228
rect 33792 -2308 39164 -2292
rect 33792 -2372 39080 -2308
rect 39144 -2372 39164 -2308
rect 33792 -2388 39164 -2372
rect 33792 -2452 39080 -2388
rect 39144 -2452 39164 -2388
rect 33792 -2468 39164 -2452
rect 33792 -2532 39080 -2468
rect 39144 -2532 39164 -2468
rect 33792 -2548 39164 -2532
rect 33792 -2612 39080 -2548
rect 39144 -2612 39164 -2548
rect 33792 -2628 39164 -2612
rect 33792 -2692 39080 -2628
rect 39144 -2692 39164 -2628
rect 33792 -2708 39164 -2692
rect 33792 -2772 39080 -2708
rect 39144 -2772 39164 -2708
rect 33792 -2788 39164 -2772
rect 33792 -2852 39080 -2788
rect 39144 -2852 39164 -2788
rect 33792 -2868 39164 -2852
rect 33792 -2932 39080 -2868
rect 39144 -2932 39164 -2868
rect 33792 -2948 39164 -2932
rect 33792 -3012 39080 -2948
rect 39144 -3012 39164 -2948
rect 33792 -3028 39164 -3012
rect 33792 -3092 39080 -3028
rect 39144 -3092 39164 -3028
rect 33792 -3108 39164 -3092
rect 33792 -3172 39080 -3108
rect 39144 -3172 39164 -3108
rect 33792 -3188 39164 -3172
rect 33792 -3252 39080 -3188
rect 39144 -3252 39164 -3188
rect 33792 -3268 39164 -3252
rect 33792 -3332 39080 -3268
rect 39144 -3332 39164 -3268
rect 33792 -3348 39164 -3332
rect 33792 -3412 39080 -3348
rect 39144 -3412 39164 -3348
rect 33792 -3428 39164 -3412
rect 33792 -3492 39080 -3428
rect 39144 -3492 39164 -3428
rect 33792 -3508 39164 -3492
rect 33792 -3572 39080 -3508
rect 39144 -3572 39164 -3508
rect 33792 -3588 39164 -3572
rect 33792 -3652 39080 -3588
rect 39144 -3652 39164 -3588
rect 33792 -3668 39164 -3652
rect 33792 -3732 39080 -3668
rect 39144 -3732 39164 -3668
rect 33792 -3748 39164 -3732
rect 33792 -3812 39080 -3748
rect 39144 -3812 39164 -3748
rect 33792 -3828 39164 -3812
rect 33792 -3892 39080 -3828
rect 39144 -3892 39164 -3828
rect 33792 -3908 39164 -3892
rect 33792 -3972 39080 -3908
rect 39144 -3972 39164 -3908
rect 33792 -3988 39164 -3972
rect 33792 -4052 39080 -3988
rect 39144 -4052 39164 -3988
rect 33792 -4068 39164 -4052
rect 33792 -4132 39080 -4068
rect 39144 -4132 39164 -4068
rect 33792 -4148 39164 -4132
rect 33792 -4212 39080 -4148
rect 39144 -4212 39164 -4148
rect 33792 -4228 39164 -4212
rect 33792 -4292 39080 -4228
rect 39144 -4292 39164 -4228
rect 33792 -4308 39164 -4292
rect 33792 -4372 39080 -4308
rect 39144 -4372 39164 -4308
rect 33792 -4388 39164 -4372
rect 33792 -4452 39080 -4388
rect 39144 -4452 39164 -4388
rect 33792 -4468 39164 -4452
rect 33792 -4532 39080 -4468
rect 39144 -4532 39164 -4468
rect 33792 -4548 39164 -4532
rect 33792 -4612 39080 -4548
rect 39144 -4612 39164 -4548
rect 33792 -4628 39164 -4612
rect 33792 -4692 39080 -4628
rect 39144 -4692 39164 -4628
rect 33792 -4708 39164 -4692
rect 33792 -4772 39080 -4708
rect 39144 -4772 39164 -4708
rect 33792 -4788 39164 -4772
rect 33792 -4852 39080 -4788
rect 39144 -4852 39164 -4788
rect 33792 -4868 39164 -4852
rect 33792 -4932 39080 -4868
rect 39144 -4932 39164 -4868
rect 33792 -4948 39164 -4932
rect 33792 -5012 39080 -4948
rect 39144 -5012 39164 -4948
rect 33792 -5028 39164 -5012
rect 33792 -5092 39080 -5028
rect 39144 -5092 39164 -5028
rect 33792 -5108 39164 -5092
rect 33792 -5172 39080 -5108
rect 39144 -5172 39164 -5108
rect 33792 -5200 39164 -5172
rect -39164 -5468 -33792 -5440
rect -39164 -5532 -33876 -5468
rect -33812 -5532 -33792 -5468
rect -39164 -5548 -33792 -5532
rect -39164 -5612 -33876 -5548
rect -33812 -5612 -33792 -5548
rect -39164 -5628 -33792 -5612
rect -39164 -5692 -33876 -5628
rect -33812 -5692 -33792 -5628
rect -39164 -5708 -33792 -5692
rect -39164 -5772 -33876 -5708
rect -33812 -5772 -33792 -5708
rect -39164 -5788 -33792 -5772
rect -39164 -5852 -33876 -5788
rect -33812 -5852 -33792 -5788
rect -39164 -5868 -33792 -5852
rect -39164 -5932 -33876 -5868
rect -33812 -5932 -33792 -5868
rect -39164 -5948 -33792 -5932
rect -39164 -6012 -33876 -5948
rect -33812 -6012 -33792 -5948
rect -39164 -6028 -33792 -6012
rect -39164 -6092 -33876 -6028
rect -33812 -6092 -33792 -6028
rect -39164 -6108 -33792 -6092
rect -39164 -6172 -33876 -6108
rect -33812 -6172 -33792 -6108
rect -39164 -6188 -33792 -6172
rect -39164 -6252 -33876 -6188
rect -33812 -6252 -33792 -6188
rect -39164 -6268 -33792 -6252
rect -39164 -6332 -33876 -6268
rect -33812 -6332 -33792 -6268
rect -39164 -6348 -33792 -6332
rect -39164 -6412 -33876 -6348
rect -33812 -6412 -33792 -6348
rect -39164 -6428 -33792 -6412
rect -39164 -6492 -33876 -6428
rect -33812 -6492 -33792 -6428
rect -39164 -6508 -33792 -6492
rect -39164 -6572 -33876 -6508
rect -33812 -6572 -33792 -6508
rect -39164 -6588 -33792 -6572
rect -39164 -6652 -33876 -6588
rect -33812 -6652 -33792 -6588
rect -39164 -6668 -33792 -6652
rect -39164 -6732 -33876 -6668
rect -33812 -6732 -33792 -6668
rect -39164 -6748 -33792 -6732
rect -39164 -6812 -33876 -6748
rect -33812 -6812 -33792 -6748
rect -39164 -6828 -33792 -6812
rect -39164 -6892 -33876 -6828
rect -33812 -6892 -33792 -6828
rect -39164 -6908 -33792 -6892
rect -39164 -6972 -33876 -6908
rect -33812 -6972 -33792 -6908
rect -39164 -6988 -33792 -6972
rect -39164 -7052 -33876 -6988
rect -33812 -7052 -33792 -6988
rect -39164 -7068 -33792 -7052
rect -39164 -7132 -33876 -7068
rect -33812 -7132 -33792 -7068
rect -39164 -7148 -33792 -7132
rect -39164 -7212 -33876 -7148
rect -33812 -7212 -33792 -7148
rect -39164 -7228 -33792 -7212
rect -39164 -7292 -33876 -7228
rect -33812 -7292 -33792 -7228
rect -39164 -7308 -33792 -7292
rect -39164 -7372 -33876 -7308
rect -33812 -7372 -33792 -7308
rect -39164 -7388 -33792 -7372
rect -39164 -7452 -33876 -7388
rect -33812 -7452 -33792 -7388
rect -39164 -7468 -33792 -7452
rect -39164 -7532 -33876 -7468
rect -33812 -7532 -33792 -7468
rect -39164 -7548 -33792 -7532
rect -39164 -7612 -33876 -7548
rect -33812 -7612 -33792 -7548
rect -39164 -7628 -33792 -7612
rect -39164 -7692 -33876 -7628
rect -33812 -7692 -33792 -7628
rect -39164 -7708 -33792 -7692
rect -39164 -7772 -33876 -7708
rect -33812 -7772 -33792 -7708
rect -39164 -7788 -33792 -7772
rect -39164 -7852 -33876 -7788
rect -33812 -7852 -33792 -7788
rect -39164 -7868 -33792 -7852
rect -39164 -7932 -33876 -7868
rect -33812 -7932 -33792 -7868
rect -39164 -7948 -33792 -7932
rect -39164 -8012 -33876 -7948
rect -33812 -8012 -33792 -7948
rect -39164 -8028 -33792 -8012
rect -39164 -8092 -33876 -8028
rect -33812 -8092 -33792 -8028
rect -39164 -8108 -33792 -8092
rect -39164 -8172 -33876 -8108
rect -33812 -8172 -33792 -8108
rect -39164 -8188 -33792 -8172
rect -39164 -8252 -33876 -8188
rect -33812 -8252 -33792 -8188
rect -39164 -8268 -33792 -8252
rect -39164 -8332 -33876 -8268
rect -33812 -8332 -33792 -8268
rect -39164 -8348 -33792 -8332
rect -39164 -8412 -33876 -8348
rect -33812 -8412 -33792 -8348
rect -39164 -8428 -33792 -8412
rect -39164 -8492 -33876 -8428
rect -33812 -8492 -33792 -8428
rect -39164 -8508 -33792 -8492
rect -39164 -8572 -33876 -8508
rect -33812 -8572 -33792 -8508
rect -39164 -8588 -33792 -8572
rect -39164 -8652 -33876 -8588
rect -33812 -8652 -33792 -8588
rect -39164 -8668 -33792 -8652
rect -39164 -8732 -33876 -8668
rect -33812 -8732 -33792 -8668
rect -39164 -8748 -33792 -8732
rect -39164 -8812 -33876 -8748
rect -33812 -8812 -33792 -8748
rect -39164 -8828 -33792 -8812
rect -39164 -8892 -33876 -8828
rect -33812 -8892 -33792 -8828
rect -39164 -8908 -33792 -8892
rect -39164 -8972 -33876 -8908
rect -33812 -8972 -33792 -8908
rect -39164 -8988 -33792 -8972
rect -39164 -9052 -33876 -8988
rect -33812 -9052 -33792 -8988
rect -39164 -9068 -33792 -9052
rect -39164 -9132 -33876 -9068
rect -33812 -9132 -33792 -9068
rect -39164 -9148 -33792 -9132
rect -39164 -9212 -33876 -9148
rect -33812 -9212 -33792 -9148
rect -39164 -9228 -33792 -9212
rect -39164 -9292 -33876 -9228
rect -33812 -9292 -33792 -9228
rect -39164 -9308 -33792 -9292
rect -39164 -9372 -33876 -9308
rect -33812 -9372 -33792 -9308
rect -39164 -9388 -33792 -9372
rect -39164 -9452 -33876 -9388
rect -33812 -9452 -33792 -9388
rect -39164 -9468 -33792 -9452
rect -39164 -9532 -33876 -9468
rect -33812 -9532 -33792 -9468
rect -39164 -9548 -33792 -9532
rect -39164 -9612 -33876 -9548
rect -33812 -9612 -33792 -9548
rect -39164 -9628 -33792 -9612
rect -39164 -9692 -33876 -9628
rect -33812 -9692 -33792 -9628
rect -39164 -9708 -33792 -9692
rect -39164 -9772 -33876 -9708
rect -33812 -9772 -33792 -9708
rect -39164 -9788 -33792 -9772
rect -39164 -9852 -33876 -9788
rect -33812 -9852 -33792 -9788
rect -39164 -9868 -33792 -9852
rect -39164 -9932 -33876 -9868
rect -33812 -9932 -33792 -9868
rect -39164 -9948 -33792 -9932
rect -39164 -10012 -33876 -9948
rect -33812 -10012 -33792 -9948
rect -39164 -10028 -33792 -10012
rect -39164 -10092 -33876 -10028
rect -33812 -10092 -33792 -10028
rect -39164 -10108 -33792 -10092
rect -39164 -10172 -33876 -10108
rect -33812 -10172 -33792 -10108
rect -39164 -10188 -33792 -10172
rect -39164 -10252 -33876 -10188
rect -33812 -10252 -33792 -10188
rect -39164 -10268 -33792 -10252
rect -39164 -10332 -33876 -10268
rect -33812 -10332 -33792 -10268
rect -39164 -10348 -33792 -10332
rect -39164 -10412 -33876 -10348
rect -33812 -10412 -33792 -10348
rect -39164 -10428 -33792 -10412
rect -39164 -10492 -33876 -10428
rect -33812 -10492 -33792 -10428
rect -39164 -10520 -33792 -10492
rect -33552 -5468 -28180 -5440
rect -33552 -5532 -28264 -5468
rect -28200 -5532 -28180 -5468
rect -33552 -5548 -28180 -5532
rect -33552 -5612 -28264 -5548
rect -28200 -5612 -28180 -5548
rect -33552 -5628 -28180 -5612
rect -33552 -5692 -28264 -5628
rect -28200 -5692 -28180 -5628
rect -33552 -5708 -28180 -5692
rect -33552 -5772 -28264 -5708
rect -28200 -5772 -28180 -5708
rect -33552 -5788 -28180 -5772
rect -33552 -5852 -28264 -5788
rect -28200 -5852 -28180 -5788
rect -33552 -5868 -28180 -5852
rect -33552 -5932 -28264 -5868
rect -28200 -5932 -28180 -5868
rect -33552 -5948 -28180 -5932
rect -33552 -6012 -28264 -5948
rect -28200 -6012 -28180 -5948
rect -33552 -6028 -28180 -6012
rect -33552 -6092 -28264 -6028
rect -28200 -6092 -28180 -6028
rect -33552 -6108 -28180 -6092
rect -33552 -6172 -28264 -6108
rect -28200 -6172 -28180 -6108
rect -33552 -6188 -28180 -6172
rect -33552 -6252 -28264 -6188
rect -28200 -6252 -28180 -6188
rect -33552 -6268 -28180 -6252
rect -33552 -6332 -28264 -6268
rect -28200 -6332 -28180 -6268
rect -33552 -6348 -28180 -6332
rect -33552 -6412 -28264 -6348
rect -28200 -6412 -28180 -6348
rect -33552 -6428 -28180 -6412
rect -33552 -6492 -28264 -6428
rect -28200 -6492 -28180 -6428
rect -33552 -6508 -28180 -6492
rect -33552 -6572 -28264 -6508
rect -28200 -6572 -28180 -6508
rect -33552 -6588 -28180 -6572
rect -33552 -6652 -28264 -6588
rect -28200 -6652 -28180 -6588
rect -33552 -6668 -28180 -6652
rect -33552 -6732 -28264 -6668
rect -28200 -6732 -28180 -6668
rect -33552 -6748 -28180 -6732
rect -33552 -6812 -28264 -6748
rect -28200 -6812 -28180 -6748
rect -33552 -6828 -28180 -6812
rect -33552 -6892 -28264 -6828
rect -28200 -6892 -28180 -6828
rect -33552 -6908 -28180 -6892
rect -33552 -6972 -28264 -6908
rect -28200 -6972 -28180 -6908
rect -33552 -6988 -28180 -6972
rect -33552 -7052 -28264 -6988
rect -28200 -7052 -28180 -6988
rect -33552 -7068 -28180 -7052
rect -33552 -7132 -28264 -7068
rect -28200 -7132 -28180 -7068
rect -33552 -7148 -28180 -7132
rect -33552 -7212 -28264 -7148
rect -28200 -7212 -28180 -7148
rect -33552 -7228 -28180 -7212
rect -33552 -7292 -28264 -7228
rect -28200 -7292 -28180 -7228
rect -33552 -7308 -28180 -7292
rect -33552 -7372 -28264 -7308
rect -28200 -7372 -28180 -7308
rect -33552 -7388 -28180 -7372
rect -33552 -7452 -28264 -7388
rect -28200 -7452 -28180 -7388
rect -33552 -7468 -28180 -7452
rect -33552 -7532 -28264 -7468
rect -28200 -7532 -28180 -7468
rect -33552 -7548 -28180 -7532
rect -33552 -7612 -28264 -7548
rect -28200 -7612 -28180 -7548
rect -33552 -7628 -28180 -7612
rect -33552 -7692 -28264 -7628
rect -28200 -7692 -28180 -7628
rect -33552 -7708 -28180 -7692
rect -33552 -7772 -28264 -7708
rect -28200 -7772 -28180 -7708
rect -33552 -7788 -28180 -7772
rect -33552 -7852 -28264 -7788
rect -28200 -7852 -28180 -7788
rect -33552 -7868 -28180 -7852
rect -33552 -7932 -28264 -7868
rect -28200 -7932 -28180 -7868
rect -33552 -7948 -28180 -7932
rect -33552 -8012 -28264 -7948
rect -28200 -8012 -28180 -7948
rect -33552 -8028 -28180 -8012
rect -33552 -8092 -28264 -8028
rect -28200 -8092 -28180 -8028
rect -33552 -8108 -28180 -8092
rect -33552 -8172 -28264 -8108
rect -28200 -8172 -28180 -8108
rect -33552 -8188 -28180 -8172
rect -33552 -8252 -28264 -8188
rect -28200 -8252 -28180 -8188
rect -33552 -8268 -28180 -8252
rect -33552 -8332 -28264 -8268
rect -28200 -8332 -28180 -8268
rect -33552 -8348 -28180 -8332
rect -33552 -8412 -28264 -8348
rect -28200 -8412 -28180 -8348
rect -33552 -8428 -28180 -8412
rect -33552 -8492 -28264 -8428
rect -28200 -8492 -28180 -8428
rect -33552 -8508 -28180 -8492
rect -33552 -8572 -28264 -8508
rect -28200 -8572 -28180 -8508
rect -33552 -8588 -28180 -8572
rect -33552 -8652 -28264 -8588
rect -28200 -8652 -28180 -8588
rect -33552 -8668 -28180 -8652
rect -33552 -8732 -28264 -8668
rect -28200 -8732 -28180 -8668
rect -33552 -8748 -28180 -8732
rect -33552 -8812 -28264 -8748
rect -28200 -8812 -28180 -8748
rect -33552 -8828 -28180 -8812
rect -33552 -8892 -28264 -8828
rect -28200 -8892 -28180 -8828
rect -33552 -8908 -28180 -8892
rect -33552 -8972 -28264 -8908
rect -28200 -8972 -28180 -8908
rect -33552 -8988 -28180 -8972
rect -33552 -9052 -28264 -8988
rect -28200 -9052 -28180 -8988
rect -33552 -9068 -28180 -9052
rect -33552 -9132 -28264 -9068
rect -28200 -9132 -28180 -9068
rect -33552 -9148 -28180 -9132
rect -33552 -9212 -28264 -9148
rect -28200 -9212 -28180 -9148
rect -33552 -9228 -28180 -9212
rect -33552 -9292 -28264 -9228
rect -28200 -9292 -28180 -9228
rect -33552 -9308 -28180 -9292
rect -33552 -9372 -28264 -9308
rect -28200 -9372 -28180 -9308
rect -33552 -9388 -28180 -9372
rect -33552 -9452 -28264 -9388
rect -28200 -9452 -28180 -9388
rect -33552 -9468 -28180 -9452
rect -33552 -9532 -28264 -9468
rect -28200 -9532 -28180 -9468
rect -33552 -9548 -28180 -9532
rect -33552 -9612 -28264 -9548
rect -28200 -9612 -28180 -9548
rect -33552 -9628 -28180 -9612
rect -33552 -9692 -28264 -9628
rect -28200 -9692 -28180 -9628
rect -33552 -9708 -28180 -9692
rect -33552 -9772 -28264 -9708
rect -28200 -9772 -28180 -9708
rect -33552 -9788 -28180 -9772
rect -33552 -9852 -28264 -9788
rect -28200 -9852 -28180 -9788
rect -33552 -9868 -28180 -9852
rect -33552 -9932 -28264 -9868
rect -28200 -9932 -28180 -9868
rect -33552 -9948 -28180 -9932
rect -33552 -10012 -28264 -9948
rect -28200 -10012 -28180 -9948
rect -33552 -10028 -28180 -10012
rect -33552 -10092 -28264 -10028
rect -28200 -10092 -28180 -10028
rect -33552 -10108 -28180 -10092
rect -33552 -10172 -28264 -10108
rect -28200 -10172 -28180 -10108
rect -33552 -10188 -28180 -10172
rect -33552 -10252 -28264 -10188
rect -28200 -10252 -28180 -10188
rect -33552 -10268 -28180 -10252
rect -33552 -10332 -28264 -10268
rect -28200 -10332 -28180 -10268
rect -33552 -10348 -28180 -10332
rect -33552 -10412 -28264 -10348
rect -28200 -10412 -28180 -10348
rect -33552 -10428 -28180 -10412
rect -33552 -10492 -28264 -10428
rect -28200 -10492 -28180 -10428
rect -33552 -10520 -28180 -10492
rect -27940 -5468 -22568 -5440
rect -27940 -5532 -22652 -5468
rect -22588 -5532 -22568 -5468
rect -27940 -5548 -22568 -5532
rect -27940 -5612 -22652 -5548
rect -22588 -5612 -22568 -5548
rect -27940 -5628 -22568 -5612
rect -27940 -5692 -22652 -5628
rect -22588 -5692 -22568 -5628
rect -27940 -5708 -22568 -5692
rect -27940 -5772 -22652 -5708
rect -22588 -5772 -22568 -5708
rect -27940 -5788 -22568 -5772
rect -27940 -5852 -22652 -5788
rect -22588 -5852 -22568 -5788
rect -27940 -5868 -22568 -5852
rect -27940 -5932 -22652 -5868
rect -22588 -5932 -22568 -5868
rect -27940 -5948 -22568 -5932
rect -27940 -6012 -22652 -5948
rect -22588 -6012 -22568 -5948
rect -27940 -6028 -22568 -6012
rect -27940 -6092 -22652 -6028
rect -22588 -6092 -22568 -6028
rect -27940 -6108 -22568 -6092
rect -27940 -6172 -22652 -6108
rect -22588 -6172 -22568 -6108
rect -27940 -6188 -22568 -6172
rect -27940 -6252 -22652 -6188
rect -22588 -6252 -22568 -6188
rect -27940 -6268 -22568 -6252
rect -27940 -6332 -22652 -6268
rect -22588 -6332 -22568 -6268
rect -27940 -6348 -22568 -6332
rect -27940 -6412 -22652 -6348
rect -22588 -6412 -22568 -6348
rect -27940 -6428 -22568 -6412
rect -27940 -6492 -22652 -6428
rect -22588 -6492 -22568 -6428
rect -27940 -6508 -22568 -6492
rect -27940 -6572 -22652 -6508
rect -22588 -6572 -22568 -6508
rect -27940 -6588 -22568 -6572
rect -27940 -6652 -22652 -6588
rect -22588 -6652 -22568 -6588
rect -27940 -6668 -22568 -6652
rect -27940 -6732 -22652 -6668
rect -22588 -6732 -22568 -6668
rect -27940 -6748 -22568 -6732
rect -27940 -6812 -22652 -6748
rect -22588 -6812 -22568 -6748
rect -27940 -6828 -22568 -6812
rect -27940 -6892 -22652 -6828
rect -22588 -6892 -22568 -6828
rect -27940 -6908 -22568 -6892
rect -27940 -6972 -22652 -6908
rect -22588 -6972 -22568 -6908
rect -27940 -6988 -22568 -6972
rect -27940 -7052 -22652 -6988
rect -22588 -7052 -22568 -6988
rect -27940 -7068 -22568 -7052
rect -27940 -7132 -22652 -7068
rect -22588 -7132 -22568 -7068
rect -27940 -7148 -22568 -7132
rect -27940 -7212 -22652 -7148
rect -22588 -7212 -22568 -7148
rect -27940 -7228 -22568 -7212
rect -27940 -7292 -22652 -7228
rect -22588 -7292 -22568 -7228
rect -27940 -7308 -22568 -7292
rect -27940 -7372 -22652 -7308
rect -22588 -7372 -22568 -7308
rect -27940 -7388 -22568 -7372
rect -27940 -7452 -22652 -7388
rect -22588 -7452 -22568 -7388
rect -27940 -7468 -22568 -7452
rect -27940 -7532 -22652 -7468
rect -22588 -7532 -22568 -7468
rect -27940 -7548 -22568 -7532
rect -27940 -7612 -22652 -7548
rect -22588 -7612 -22568 -7548
rect -27940 -7628 -22568 -7612
rect -27940 -7692 -22652 -7628
rect -22588 -7692 -22568 -7628
rect -27940 -7708 -22568 -7692
rect -27940 -7772 -22652 -7708
rect -22588 -7772 -22568 -7708
rect -27940 -7788 -22568 -7772
rect -27940 -7852 -22652 -7788
rect -22588 -7852 -22568 -7788
rect -27940 -7868 -22568 -7852
rect -27940 -7932 -22652 -7868
rect -22588 -7932 -22568 -7868
rect -27940 -7948 -22568 -7932
rect -27940 -8012 -22652 -7948
rect -22588 -8012 -22568 -7948
rect -27940 -8028 -22568 -8012
rect -27940 -8092 -22652 -8028
rect -22588 -8092 -22568 -8028
rect -27940 -8108 -22568 -8092
rect -27940 -8172 -22652 -8108
rect -22588 -8172 -22568 -8108
rect -27940 -8188 -22568 -8172
rect -27940 -8252 -22652 -8188
rect -22588 -8252 -22568 -8188
rect -27940 -8268 -22568 -8252
rect -27940 -8332 -22652 -8268
rect -22588 -8332 -22568 -8268
rect -27940 -8348 -22568 -8332
rect -27940 -8412 -22652 -8348
rect -22588 -8412 -22568 -8348
rect -27940 -8428 -22568 -8412
rect -27940 -8492 -22652 -8428
rect -22588 -8492 -22568 -8428
rect -27940 -8508 -22568 -8492
rect -27940 -8572 -22652 -8508
rect -22588 -8572 -22568 -8508
rect -27940 -8588 -22568 -8572
rect -27940 -8652 -22652 -8588
rect -22588 -8652 -22568 -8588
rect -27940 -8668 -22568 -8652
rect -27940 -8732 -22652 -8668
rect -22588 -8732 -22568 -8668
rect -27940 -8748 -22568 -8732
rect -27940 -8812 -22652 -8748
rect -22588 -8812 -22568 -8748
rect -27940 -8828 -22568 -8812
rect -27940 -8892 -22652 -8828
rect -22588 -8892 -22568 -8828
rect -27940 -8908 -22568 -8892
rect -27940 -8972 -22652 -8908
rect -22588 -8972 -22568 -8908
rect -27940 -8988 -22568 -8972
rect -27940 -9052 -22652 -8988
rect -22588 -9052 -22568 -8988
rect -27940 -9068 -22568 -9052
rect -27940 -9132 -22652 -9068
rect -22588 -9132 -22568 -9068
rect -27940 -9148 -22568 -9132
rect -27940 -9212 -22652 -9148
rect -22588 -9212 -22568 -9148
rect -27940 -9228 -22568 -9212
rect -27940 -9292 -22652 -9228
rect -22588 -9292 -22568 -9228
rect -27940 -9308 -22568 -9292
rect -27940 -9372 -22652 -9308
rect -22588 -9372 -22568 -9308
rect -27940 -9388 -22568 -9372
rect -27940 -9452 -22652 -9388
rect -22588 -9452 -22568 -9388
rect -27940 -9468 -22568 -9452
rect -27940 -9532 -22652 -9468
rect -22588 -9532 -22568 -9468
rect -27940 -9548 -22568 -9532
rect -27940 -9612 -22652 -9548
rect -22588 -9612 -22568 -9548
rect -27940 -9628 -22568 -9612
rect -27940 -9692 -22652 -9628
rect -22588 -9692 -22568 -9628
rect -27940 -9708 -22568 -9692
rect -27940 -9772 -22652 -9708
rect -22588 -9772 -22568 -9708
rect -27940 -9788 -22568 -9772
rect -27940 -9852 -22652 -9788
rect -22588 -9852 -22568 -9788
rect -27940 -9868 -22568 -9852
rect -27940 -9932 -22652 -9868
rect -22588 -9932 -22568 -9868
rect -27940 -9948 -22568 -9932
rect -27940 -10012 -22652 -9948
rect -22588 -10012 -22568 -9948
rect -27940 -10028 -22568 -10012
rect -27940 -10092 -22652 -10028
rect -22588 -10092 -22568 -10028
rect -27940 -10108 -22568 -10092
rect -27940 -10172 -22652 -10108
rect -22588 -10172 -22568 -10108
rect -27940 -10188 -22568 -10172
rect -27940 -10252 -22652 -10188
rect -22588 -10252 -22568 -10188
rect -27940 -10268 -22568 -10252
rect -27940 -10332 -22652 -10268
rect -22588 -10332 -22568 -10268
rect -27940 -10348 -22568 -10332
rect -27940 -10412 -22652 -10348
rect -22588 -10412 -22568 -10348
rect -27940 -10428 -22568 -10412
rect -27940 -10492 -22652 -10428
rect -22588 -10492 -22568 -10428
rect -27940 -10520 -22568 -10492
rect -22328 -5468 -16956 -5440
rect -22328 -5532 -17040 -5468
rect -16976 -5532 -16956 -5468
rect -22328 -5548 -16956 -5532
rect -22328 -5612 -17040 -5548
rect -16976 -5612 -16956 -5548
rect -22328 -5628 -16956 -5612
rect -22328 -5692 -17040 -5628
rect -16976 -5692 -16956 -5628
rect -22328 -5708 -16956 -5692
rect -22328 -5772 -17040 -5708
rect -16976 -5772 -16956 -5708
rect -22328 -5788 -16956 -5772
rect -22328 -5852 -17040 -5788
rect -16976 -5852 -16956 -5788
rect -22328 -5868 -16956 -5852
rect -22328 -5932 -17040 -5868
rect -16976 -5932 -16956 -5868
rect -22328 -5948 -16956 -5932
rect -22328 -6012 -17040 -5948
rect -16976 -6012 -16956 -5948
rect -22328 -6028 -16956 -6012
rect -22328 -6092 -17040 -6028
rect -16976 -6092 -16956 -6028
rect -22328 -6108 -16956 -6092
rect -22328 -6172 -17040 -6108
rect -16976 -6172 -16956 -6108
rect -22328 -6188 -16956 -6172
rect -22328 -6252 -17040 -6188
rect -16976 -6252 -16956 -6188
rect -22328 -6268 -16956 -6252
rect -22328 -6332 -17040 -6268
rect -16976 -6332 -16956 -6268
rect -22328 -6348 -16956 -6332
rect -22328 -6412 -17040 -6348
rect -16976 -6412 -16956 -6348
rect -22328 -6428 -16956 -6412
rect -22328 -6492 -17040 -6428
rect -16976 -6492 -16956 -6428
rect -22328 -6508 -16956 -6492
rect -22328 -6572 -17040 -6508
rect -16976 -6572 -16956 -6508
rect -22328 -6588 -16956 -6572
rect -22328 -6652 -17040 -6588
rect -16976 -6652 -16956 -6588
rect -22328 -6668 -16956 -6652
rect -22328 -6732 -17040 -6668
rect -16976 -6732 -16956 -6668
rect -22328 -6748 -16956 -6732
rect -22328 -6812 -17040 -6748
rect -16976 -6812 -16956 -6748
rect -22328 -6828 -16956 -6812
rect -22328 -6892 -17040 -6828
rect -16976 -6892 -16956 -6828
rect -22328 -6908 -16956 -6892
rect -22328 -6972 -17040 -6908
rect -16976 -6972 -16956 -6908
rect -22328 -6988 -16956 -6972
rect -22328 -7052 -17040 -6988
rect -16976 -7052 -16956 -6988
rect -22328 -7068 -16956 -7052
rect -22328 -7132 -17040 -7068
rect -16976 -7132 -16956 -7068
rect -22328 -7148 -16956 -7132
rect -22328 -7212 -17040 -7148
rect -16976 -7212 -16956 -7148
rect -22328 -7228 -16956 -7212
rect -22328 -7292 -17040 -7228
rect -16976 -7292 -16956 -7228
rect -22328 -7308 -16956 -7292
rect -22328 -7372 -17040 -7308
rect -16976 -7372 -16956 -7308
rect -22328 -7388 -16956 -7372
rect -22328 -7452 -17040 -7388
rect -16976 -7452 -16956 -7388
rect -22328 -7468 -16956 -7452
rect -22328 -7532 -17040 -7468
rect -16976 -7532 -16956 -7468
rect -22328 -7548 -16956 -7532
rect -22328 -7612 -17040 -7548
rect -16976 -7612 -16956 -7548
rect -22328 -7628 -16956 -7612
rect -22328 -7692 -17040 -7628
rect -16976 -7692 -16956 -7628
rect -22328 -7708 -16956 -7692
rect -22328 -7772 -17040 -7708
rect -16976 -7772 -16956 -7708
rect -22328 -7788 -16956 -7772
rect -22328 -7852 -17040 -7788
rect -16976 -7852 -16956 -7788
rect -22328 -7868 -16956 -7852
rect -22328 -7932 -17040 -7868
rect -16976 -7932 -16956 -7868
rect -22328 -7948 -16956 -7932
rect -22328 -8012 -17040 -7948
rect -16976 -8012 -16956 -7948
rect -22328 -8028 -16956 -8012
rect -22328 -8092 -17040 -8028
rect -16976 -8092 -16956 -8028
rect -22328 -8108 -16956 -8092
rect -22328 -8172 -17040 -8108
rect -16976 -8172 -16956 -8108
rect -22328 -8188 -16956 -8172
rect -22328 -8252 -17040 -8188
rect -16976 -8252 -16956 -8188
rect -22328 -8268 -16956 -8252
rect -22328 -8332 -17040 -8268
rect -16976 -8332 -16956 -8268
rect -22328 -8348 -16956 -8332
rect -22328 -8412 -17040 -8348
rect -16976 -8412 -16956 -8348
rect -22328 -8428 -16956 -8412
rect -22328 -8492 -17040 -8428
rect -16976 -8492 -16956 -8428
rect -22328 -8508 -16956 -8492
rect -22328 -8572 -17040 -8508
rect -16976 -8572 -16956 -8508
rect -22328 -8588 -16956 -8572
rect -22328 -8652 -17040 -8588
rect -16976 -8652 -16956 -8588
rect -22328 -8668 -16956 -8652
rect -22328 -8732 -17040 -8668
rect -16976 -8732 -16956 -8668
rect -22328 -8748 -16956 -8732
rect -22328 -8812 -17040 -8748
rect -16976 -8812 -16956 -8748
rect -22328 -8828 -16956 -8812
rect -22328 -8892 -17040 -8828
rect -16976 -8892 -16956 -8828
rect -22328 -8908 -16956 -8892
rect -22328 -8972 -17040 -8908
rect -16976 -8972 -16956 -8908
rect -22328 -8988 -16956 -8972
rect -22328 -9052 -17040 -8988
rect -16976 -9052 -16956 -8988
rect -22328 -9068 -16956 -9052
rect -22328 -9132 -17040 -9068
rect -16976 -9132 -16956 -9068
rect -22328 -9148 -16956 -9132
rect -22328 -9212 -17040 -9148
rect -16976 -9212 -16956 -9148
rect -22328 -9228 -16956 -9212
rect -22328 -9292 -17040 -9228
rect -16976 -9292 -16956 -9228
rect -22328 -9308 -16956 -9292
rect -22328 -9372 -17040 -9308
rect -16976 -9372 -16956 -9308
rect -22328 -9388 -16956 -9372
rect -22328 -9452 -17040 -9388
rect -16976 -9452 -16956 -9388
rect -22328 -9468 -16956 -9452
rect -22328 -9532 -17040 -9468
rect -16976 -9532 -16956 -9468
rect -22328 -9548 -16956 -9532
rect -22328 -9612 -17040 -9548
rect -16976 -9612 -16956 -9548
rect -22328 -9628 -16956 -9612
rect -22328 -9692 -17040 -9628
rect -16976 -9692 -16956 -9628
rect -22328 -9708 -16956 -9692
rect -22328 -9772 -17040 -9708
rect -16976 -9772 -16956 -9708
rect -22328 -9788 -16956 -9772
rect -22328 -9852 -17040 -9788
rect -16976 -9852 -16956 -9788
rect -22328 -9868 -16956 -9852
rect -22328 -9932 -17040 -9868
rect -16976 -9932 -16956 -9868
rect -22328 -9948 -16956 -9932
rect -22328 -10012 -17040 -9948
rect -16976 -10012 -16956 -9948
rect -22328 -10028 -16956 -10012
rect -22328 -10092 -17040 -10028
rect -16976 -10092 -16956 -10028
rect -22328 -10108 -16956 -10092
rect -22328 -10172 -17040 -10108
rect -16976 -10172 -16956 -10108
rect -22328 -10188 -16956 -10172
rect -22328 -10252 -17040 -10188
rect -16976 -10252 -16956 -10188
rect -22328 -10268 -16956 -10252
rect -22328 -10332 -17040 -10268
rect -16976 -10332 -16956 -10268
rect -22328 -10348 -16956 -10332
rect -22328 -10412 -17040 -10348
rect -16976 -10412 -16956 -10348
rect -22328 -10428 -16956 -10412
rect -22328 -10492 -17040 -10428
rect -16976 -10492 -16956 -10428
rect -22328 -10520 -16956 -10492
rect -16716 -5468 -11344 -5440
rect -16716 -5532 -11428 -5468
rect -11364 -5532 -11344 -5468
rect -16716 -5548 -11344 -5532
rect -16716 -5612 -11428 -5548
rect -11364 -5612 -11344 -5548
rect -16716 -5628 -11344 -5612
rect -16716 -5692 -11428 -5628
rect -11364 -5692 -11344 -5628
rect -16716 -5708 -11344 -5692
rect -16716 -5772 -11428 -5708
rect -11364 -5772 -11344 -5708
rect -16716 -5788 -11344 -5772
rect -16716 -5852 -11428 -5788
rect -11364 -5852 -11344 -5788
rect -16716 -5868 -11344 -5852
rect -16716 -5932 -11428 -5868
rect -11364 -5932 -11344 -5868
rect -16716 -5948 -11344 -5932
rect -16716 -6012 -11428 -5948
rect -11364 -6012 -11344 -5948
rect -16716 -6028 -11344 -6012
rect -16716 -6092 -11428 -6028
rect -11364 -6092 -11344 -6028
rect -16716 -6108 -11344 -6092
rect -16716 -6172 -11428 -6108
rect -11364 -6172 -11344 -6108
rect -16716 -6188 -11344 -6172
rect -16716 -6252 -11428 -6188
rect -11364 -6252 -11344 -6188
rect -16716 -6268 -11344 -6252
rect -16716 -6332 -11428 -6268
rect -11364 -6332 -11344 -6268
rect -16716 -6348 -11344 -6332
rect -16716 -6412 -11428 -6348
rect -11364 -6412 -11344 -6348
rect -16716 -6428 -11344 -6412
rect -16716 -6492 -11428 -6428
rect -11364 -6492 -11344 -6428
rect -16716 -6508 -11344 -6492
rect -16716 -6572 -11428 -6508
rect -11364 -6572 -11344 -6508
rect -16716 -6588 -11344 -6572
rect -16716 -6652 -11428 -6588
rect -11364 -6652 -11344 -6588
rect -16716 -6668 -11344 -6652
rect -16716 -6732 -11428 -6668
rect -11364 -6732 -11344 -6668
rect -16716 -6748 -11344 -6732
rect -16716 -6812 -11428 -6748
rect -11364 -6812 -11344 -6748
rect -16716 -6828 -11344 -6812
rect -16716 -6892 -11428 -6828
rect -11364 -6892 -11344 -6828
rect -16716 -6908 -11344 -6892
rect -16716 -6972 -11428 -6908
rect -11364 -6972 -11344 -6908
rect -16716 -6988 -11344 -6972
rect -16716 -7052 -11428 -6988
rect -11364 -7052 -11344 -6988
rect -16716 -7068 -11344 -7052
rect -16716 -7132 -11428 -7068
rect -11364 -7132 -11344 -7068
rect -16716 -7148 -11344 -7132
rect -16716 -7212 -11428 -7148
rect -11364 -7212 -11344 -7148
rect -16716 -7228 -11344 -7212
rect -16716 -7292 -11428 -7228
rect -11364 -7292 -11344 -7228
rect -16716 -7308 -11344 -7292
rect -16716 -7372 -11428 -7308
rect -11364 -7372 -11344 -7308
rect -16716 -7388 -11344 -7372
rect -16716 -7452 -11428 -7388
rect -11364 -7452 -11344 -7388
rect -16716 -7468 -11344 -7452
rect -16716 -7532 -11428 -7468
rect -11364 -7532 -11344 -7468
rect -16716 -7548 -11344 -7532
rect -16716 -7612 -11428 -7548
rect -11364 -7612 -11344 -7548
rect -16716 -7628 -11344 -7612
rect -16716 -7692 -11428 -7628
rect -11364 -7692 -11344 -7628
rect -16716 -7708 -11344 -7692
rect -16716 -7772 -11428 -7708
rect -11364 -7772 -11344 -7708
rect -16716 -7788 -11344 -7772
rect -16716 -7852 -11428 -7788
rect -11364 -7852 -11344 -7788
rect -16716 -7868 -11344 -7852
rect -16716 -7932 -11428 -7868
rect -11364 -7932 -11344 -7868
rect -16716 -7948 -11344 -7932
rect -16716 -8012 -11428 -7948
rect -11364 -8012 -11344 -7948
rect -16716 -8028 -11344 -8012
rect -16716 -8092 -11428 -8028
rect -11364 -8092 -11344 -8028
rect -16716 -8108 -11344 -8092
rect -16716 -8172 -11428 -8108
rect -11364 -8172 -11344 -8108
rect -16716 -8188 -11344 -8172
rect -16716 -8252 -11428 -8188
rect -11364 -8252 -11344 -8188
rect -16716 -8268 -11344 -8252
rect -16716 -8332 -11428 -8268
rect -11364 -8332 -11344 -8268
rect -16716 -8348 -11344 -8332
rect -16716 -8412 -11428 -8348
rect -11364 -8412 -11344 -8348
rect -16716 -8428 -11344 -8412
rect -16716 -8492 -11428 -8428
rect -11364 -8492 -11344 -8428
rect -16716 -8508 -11344 -8492
rect -16716 -8572 -11428 -8508
rect -11364 -8572 -11344 -8508
rect -16716 -8588 -11344 -8572
rect -16716 -8652 -11428 -8588
rect -11364 -8652 -11344 -8588
rect -16716 -8668 -11344 -8652
rect -16716 -8732 -11428 -8668
rect -11364 -8732 -11344 -8668
rect -16716 -8748 -11344 -8732
rect -16716 -8812 -11428 -8748
rect -11364 -8812 -11344 -8748
rect -16716 -8828 -11344 -8812
rect -16716 -8892 -11428 -8828
rect -11364 -8892 -11344 -8828
rect -16716 -8908 -11344 -8892
rect -16716 -8972 -11428 -8908
rect -11364 -8972 -11344 -8908
rect -16716 -8988 -11344 -8972
rect -16716 -9052 -11428 -8988
rect -11364 -9052 -11344 -8988
rect -16716 -9068 -11344 -9052
rect -16716 -9132 -11428 -9068
rect -11364 -9132 -11344 -9068
rect -16716 -9148 -11344 -9132
rect -16716 -9212 -11428 -9148
rect -11364 -9212 -11344 -9148
rect -16716 -9228 -11344 -9212
rect -16716 -9292 -11428 -9228
rect -11364 -9292 -11344 -9228
rect -16716 -9308 -11344 -9292
rect -16716 -9372 -11428 -9308
rect -11364 -9372 -11344 -9308
rect -16716 -9388 -11344 -9372
rect -16716 -9452 -11428 -9388
rect -11364 -9452 -11344 -9388
rect -16716 -9468 -11344 -9452
rect -16716 -9532 -11428 -9468
rect -11364 -9532 -11344 -9468
rect -16716 -9548 -11344 -9532
rect -16716 -9612 -11428 -9548
rect -11364 -9612 -11344 -9548
rect -16716 -9628 -11344 -9612
rect -16716 -9692 -11428 -9628
rect -11364 -9692 -11344 -9628
rect -16716 -9708 -11344 -9692
rect -16716 -9772 -11428 -9708
rect -11364 -9772 -11344 -9708
rect -16716 -9788 -11344 -9772
rect -16716 -9852 -11428 -9788
rect -11364 -9852 -11344 -9788
rect -16716 -9868 -11344 -9852
rect -16716 -9932 -11428 -9868
rect -11364 -9932 -11344 -9868
rect -16716 -9948 -11344 -9932
rect -16716 -10012 -11428 -9948
rect -11364 -10012 -11344 -9948
rect -16716 -10028 -11344 -10012
rect -16716 -10092 -11428 -10028
rect -11364 -10092 -11344 -10028
rect -16716 -10108 -11344 -10092
rect -16716 -10172 -11428 -10108
rect -11364 -10172 -11344 -10108
rect -16716 -10188 -11344 -10172
rect -16716 -10252 -11428 -10188
rect -11364 -10252 -11344 -10188
rect -16716 -10268 -11344 -10252
rect -16716 -10332 -11428 -10268
rect -11364 -10332 -11344 -10268
rect -16716 -10348 -11344 -10332
rect -16716 -10412 -11428 -10348
rect -11364 -10412 -11344 -10348
rect -16716 -10428 -11344 -10412
rect -16716 -10492 -11428 -10428
rect -11364 -10492 -11344 -10428
rect -16716 -10520 -11344 -10492
rect -11104 -5468 -5732 -5440
rect -11104 -5532 -5816 -5468
rect -5752 -5532 -5732 -5468
rect -11104 -5548 -5732 -5532
rect -11104 -5612 -5816 -5548
rect -5752 -5612 -5732 -5548
rect -11104 -5628 -5732 -5612
rect -11104 -5692 -5816 -5628
rect -5752 -5692 -5732 -5628
rect -11104 -5708 -5732 -5692
rect -11104 -5772 -5816 -5708
rect -5752 -5772 -5732 -5708
rect -11104 -5788 -5732 -5772
rect -11104 -5852 -5816 -5788
rect -5752 -5852 -5732 -5788
rect -11104 -5868 -5732 -5852
rect -11104 -5932 -5816 -5868
rect -5752 -5932 -5732 -5868
rect -11104 -5948 -5732 -5932
rect -11104 -6012 -5816 -5948
rect -5752 -6012 -5732 -5948
rect -11104 -6028 -5732 -6012
rect -11104 -6092 -5816 -6028
rect -5752 -6092 -5732 -6028
rect -11104 -6108 -5732 -6092
rect -11104 -6172 -5816 -6108
rect -5752 -6172 -5732 -6108
rect -11104 -6188 -5732 -6172
rect -11104 -6252 -5816 -6188
rect -5752 -6252 -5732 -6188
rect -11104 -6268 -5732 -6252
rect -11104 -6332 -5816 -6268
rect -5752 -6332 -5732 -6268
rect -11104 -6348 -5732 -6332
rect -11104 -6412 -5816 -6348
rect -5752 -6412 -5732 -6348
rect -11104 -6428 -5732 -6412
rect -11104 -6492 -5816 -6428
rect -5752 -6492 -5732 -6428
rect -11104 -6508 -5732 -6492
rect -11104 -6572 -5816 -6508
rect -5752 -6572 -5732 -6508
rect -11104 -6588 -5732 -6572
rect -11104 -6652 -5816 -6588
rect -5752 -6652 -5732 -6588
rect -11104 -6668 -5732 -6652
rect -11104 -6732 -5816 -6668
rect -5752 -6732 -5732 -6668
rect -11104 -6748 -5732 -6732
rect -11104 -6812 -5816 -6748
rect -5752 -6812 -5732 -6748
rect -11104 -6828 -5732 -6812
rect -11104 -6892 -5816 -6828
rect -5752 -6892 -5732 -6828
rect -11104 -6908 -5732 -6892
rect -11104 -6972 -5816 -6908
rect -5752 -6972 -5732 -6908
rect -11104 -6988 -5732 -6972
rect -11104 -7052 -5816 -6988
rect -5752 -7052 -5732 -6988
rect -11104 -7068 -5732 -7052
rect -11104 -7132 -5816 -7068
rect -5752 -7132 -5732 -7068
rect -11104 -7148 -5732 -7132
rect -11104 -7212 -5816 -7148
rect -5752 -7212 -5732 -7148
rect -11104 -7228 -5732 -7212
rect -11104 -7292 -5816 -7228
rect -5752 -7292 -5732 -7228
rect -11104 -7308 -5732 -7292
rect -11104 -7372 -5816 -7308
rect -5752 -7372 -5732 -7308
rect -11104 -7388 -5732 -7372
rect -11104 -7452 -5816 -7388
rect -5752 -7452 -5732 -7388
rect -11104 -7468 -5732 -7452
rect -11104 -7532 -5816 -7468
rect -5752 -7532 -5732 -7468
rect -11104 -7548 -5732 -7532
rect -11104 -7612 -5816 -7548
rect -5752 -7612 -5732 -7548
rect -11104 -7628 -5732 -7612
rect -11104 -7692 -5816 -7628
rect -5752 -7692 -5732 -7628
rect -11104 -7708 -5732 -7692
rect -11104 -7772 -5816 -7708
rect -5752 -7772 -5732 -7708
rect -11104 -7788 -5732 -7772
rect -11104 -7852 -5816 -7788
rect -5752 -7852 -5732 -7788
rect -11104 -7868 -5732 -7852
rect -11104 -7932 -5816 -7868
rect -5752 -7932 -5732 -7868
rect -11104 -7948 -5732 -7932
rect -11104 -8012 -5816 -7948
rect -5752 -8012 -5732 -7948
rect -11104 -8028 -5732 -8012
rect -11104 -8092 -5816 -8028
rect -5752 -8092 -5732 -8028
rect -11104 -8108 -5732 -8092
rect -11104 -8172 -5816 -8108
rect -5752 -8172 -5732 -8108
rect -11104 -8188 -5732 -8172
rect -11104 -8252 -5816 -8188
rect -5752 -8252 -5732 -8188
rect -11104 -8268 -5732 -8252
rect -11104 -8332 -5816 -8268
rect -5752 -8332 -5732 -8268
rect -11104 -8348 -5732 -8332
rect -11104 -8412 -5816 -8348
rect -5752 -8412 -5732 -8348
rect -11104 -8428 -5732 -8412
rect -11104 -8492 -5816 -8428
rect -5752 -8492 -5732 -8428
rect -11104 -8508 -5732 -8492
rect -11104 -8572 -5816 -8508
rect -5752 -8572 -5732 -8508
rect -11104 -8588 -5732 -8572
rect -11104 -8652 -5816 -8588
rect -5752 -8652 -5732 -8588
rect -11104 -8668 -5732 -8652
rect -11104 -8732 -5816 -8668
rect -5752 -8732 -5732 -8668
rect -11104 -8748 -5732 -8732
rect -11104 -8812 -5816 -8748
rect -5752 -8812 -5732 -8748
rect -11104 -8828 -5732 -8812
rect -11104 -8892 -5816 -8828
rect -5752 -8892 -5732 -8828
rect -11104 -8908 -5732 -8892
rect -11104 -8972 -5816 -8908
rect -5752 -8972 -5732 -8908
rect -11104 -8988 -5732 -8972
rect -11104 -9052 -5816 -8988
rect -5752 -9052 -5732 -8988
rect -11104 -9068 -5732 -9052
rect -11104 -9132 -5816 -9068
rect -5752 -9132 -5732 -9068
rect -11104 -9148 -5732 -9132
rect -11104 -9212 -5816 -9148
rect -5752 -9212 -5732 -9148
rect -11104 -9228 -5732 -9212
rect -11104 -9292 -5816 -9228
rect -5752 -9292 -5732 -9228
rect -11104 -9308 -5732 -9292
rect -11104 -9372 -5816 -9308
rect -5752 -9372 -5732 -9308
rect -11104 -9388 -5732 -9372
rect -11104 -9452 -5816 -9388
rect -5752 -9452 -5732 -9388
rect -11104 -9468 -5732 -9452
rect -11104 -9532 -5816 -9468
rect -5752 -9532 -5732 -9468
rect -11104 -9548 -5732 -9532
rect -11104 -9612 -5816 -9548
rect -5752 -9612 -5732 -9548
rect -11104 -9628 -5732 -9612
rect -11104 -9692 -5816 -9628
rect -5752 -9692 -5732 -9628
rect -11104 -9708 -5732 -9692
rect -11104 -9772 -5816 -9708
rect -5752 -9772 -5732 -9708
rect -11104 -9788 -5732 -9772
rect -11104 -9852 -5816 -9788
rect -5752 -9852 -5732 -9788
rect -11104 -9868 -5732 -9852
rect -11104 -9932 -5816 -9868
rect -5752 -9932 -5732 -9868
rect -11104 -9948 -5732 -9932
rect -11104 -10012 -5816 -9948
rect -5752 -10012 -5732 -9948
rect -11104 -10028 -5732 -10012
rect -11104 -10092 -5816 -10028
rect -5752 -10092 -5732 -10028
rect -11104 -10108 -5732 -10092
rect -11104 -10172 -5816 -10108
rect -5752 -10172 -5732 -10108
rect -11104 -10188 -5732 -10172
rect -11104 -10252 -5816 -10188
rect -5752 -10252 -5732 -10188
rect -11104 -10268 -5732 -10252
rect -11104 -10332 -5816 -10268
rect -5752 -10332 -5732 -10268
rect -11104 -10348 -5732 -10332
rect -11104 -10412 -5816 -10348
rect -5752 -10412 -5732 -10348
rect -11104 -10428 -5732 -10412
rect -11104 -10492 -5816 -10428
rect -5752 -10492 -5732 -10428
rect -11104 -10520 -5732 -10492
rect -5492 -5468 -120 -5440
rect -5492 -5532 -204 -5468
rect -140 -5532 -120 -5468
rect -5492 -5548 -120 -5532
rect -5492 -5612 -204 -5548
rect -140 -5612 -120 -5548
rect -5492 -5628 -120 -5612
rect -5492 -5692 -204 -5628
rect -140 -5692 -120 -5628
rect -5492 -5708 -120 -5692
rect -5492 -5772 -204 -5708
rect -140 -5772 -120 -5708
rect -5492 -5788 -120 -5772
rect -5492 -5852 -204 -5788
rect -140 -5852 -120 -5788
rect -5492 -5868 -120 -5852
rect -5492 -5932 -204 -5868
rect -140 -5932 -120 -5868
rect -5492 -5948 -120 -5932
rect -5492 -6012 -204 -5948
rect -140 -6012 -120 -5948
rect -5492 -6028 -120 -6012
rect -5492 -6092 -204 -6028
rect -140 -6092 -120 -6028
rect -5492 -6108 -120 -6092
rect -5492 -6172 -204 -6108
rect -140 -6172 -120 -6108
rect -5492 -6188 -120 -6172
rect -5492 -6252 -204 -6188
rect -140 -6252 -120 -6188
rect -5492 -6268 -120 -6252
rect -5492 -6332 -204 -6268
rect -140 -6332 -120 -6268
rect -5492 -6348 -120 -6332
rect -5492 -6412 -204 -6348
rect -140 -6412 -120 -6348
rect -5492 -6428 -120 -6412
rect -5492 -6492 -204 -6428
rect -140 -6492 -120 -6428
rect -5492 -6508 -120 -6492
rect -5492 -6572 -204 -6508
rect -140 -6572 -120 -6508
rect -5492 -6588 -120 -6572
rect -5492 -6652 -204 -6588
rect -140 -6652 -120 -6588
rect -5492 -6668 -120 -6652
rect -5492 -6732 -204 -6668
rect -140 -6732 -120 -6668
rect -5492 -6748 -120 -6732
rect -5492 -6812 -204 -6748
rect -140 -6812 -120 -6748
rect -5492 -6828 -120 -6812
rect -5492 -6892 -204 -6828
rect -140 -6892 -120 -6828
rect -5492 -6908 -120 -6892
rect -5492 -6972 -204 -6908
rect -140 -6972 -120 -6908
rect -5492 -6988 -120 -6972
rect -5492 -7052 -204 -6988
rect -140 -7052 -120 -6988
rect -5492 -7068 -120 -7052
rect -5492 -7132 -204 -7068
rect -140 -7132 -120 -7068
rect -5492 -7148 -120 -7132
rect -5492 -7212 -204 -7148
rect -140 -7212 -120 -7148
rect -5492 -7228 -120 -7212
rect -5492 -7292 -204 -7228
rect -140 -7292 -120 -7228
rect -5492 -7308 -120 -7292
rect -5492 -7372 -204 -7308
rect -140 -7372 -120 -7308
rect -5492 -7388 -120 -7372
rect -5492 -7452 -204 -7388
rect -140 -7452 -120 -7388
rect -5492 -7468 -120 -7452
rect -5492 -7532 -204 -7468
rect -140 -7532 -120 -7468
rect -5492 -7548 -120 -7532
rect -5492 -7612 -204 -7548
rect -140 -7612 -120 -7548
rect -5492 -7628 -120 -7612
rect -5492 -7692 -204 -7628
rect -140 -7692 -120 -7628
rect -5492 -7708 -120 -7692
rect -5492 -7772 -204 -7708
rect -140 -7772 -120 -7708
rect -5492 -7788 -120 -7772
rect -5492 -7852 -204 -7788
rect -140 -7852 -120 -7788
rect -5492 -7868 -120 -7852
rect -5492 -7932 -204 -7868
rect -140 -7932 -120 -7868
rect -5492 -7948 -120 -7932
rect -5492 -8012 -204 -7948
rect -140 -8012 -120 -7948
rect -5492 -8028 -120 -8012
rect -5492 -8092 -204 -8028
rect -140 -8092 -120 -8028
rect -5492 -8108 -120 -8092
rect -5492 -8172 -204 -8108
rect -140 -8172 -120 -8108
rect -5492 -8188 -120 -8172
rect -5492 -8252 -204 -8188
rect -140 -8252 -120 -8188
rect -5492 -8268 -120 -8252
rect -5492 -8332 -204 -8268
rect -140 -8332 -120 -8268
rect -5492 -8348 -120 -8332
rect -5492 -8412 -204 -8348
rect -140 -8412 -120 -8348
rect -5492 -8428 -120 -8412
rect -5492 -8492 -204 -8428
rect -140 -8492 -120 -8428
rect -5492 -8508 -120 -8492
rect -5492 -8572 -204 -8508
rect -140 -8572 -120 -8508
rect -5492 -8588 -120 -8572
rect -5492 -8652 -204 -8588
rect -140 -8652 -120 -8588
rect -5492 -8668 -120 -8652
rect -5492 -8732 -204 -8668
rect -140 -8732 -120 -8668
rect -5492 -8748 -120 -8732
rect -5492 -8812 -204 -8748
rect -140 -8812 -120 -8748
rect -5492 -8828 -120 -8812
rect -5492 -8892 -204 -8828
rect -140 -8892 -120 -8828
rect -5492 -8908 -120 -8892
rect -5492 -8972 -204 -8908
rect -140 -8972 -120 -8908
rect -5492 -8988 -120 -8972
rect -5492 -9052 -204 -8988
rect -140 -9052 -120 -8988
rect -5492 -9068 -120 -9052
rect -5492 -9132 -204 -9068
rect -140 -9132 -120 -9068
rect -5492 -9148 -120 -9132
rect -5492 -9212 -204 -9148
rect -140 -9212 -120 -9148
rect -5492 -9228 -120 -9212
rect -5492 -9292 -204 -9228
rect -140 -9292 -120 -9228
rect -5492 -9308 -120 -9292
rect -5492 -9372 -204 -9308
rect -140 -9372 -120 -9308
rect -5492 -9388 -120 -9372
rect -5492 -9452 -204 -9388
rect -140 -9452 -120 -9388
rect -5492 -9468 -120 -9452
rect -5492 -9532 -204 -9468
rect -140 -9532 -120 -9468
rect -5492 -9548 -120 -9532
rect -5492 -9612 -204 -9548
rect -140 -9612 -120 -9548
rect -5492 -9628 -120 -9612
rect -5492 -9692 -204 -9628
rect -140 -9692 -120 -9628
rect -5492 -9708 -120 -9692
rect -5492 -9772 -204 -9708
rect -140 -9772 -120 -9708
rect -5492 -9788 -120 -9772
rect -5492 -9852 -204 -9788
rect -140 -9852 -120 -9788
rect -5492 -9868 -120 -9852
rect -5492 -9932 -204 -9868
rect -140 -9932 -120 -9868
rect -5492 -9948 -120 -9932
rect -5492 -10012 -204 -9948
rect -140 -10012 -120 -9948
rect -5492 -10028 -120 -10012
rect -5492 -10092 -204 -10028
rect -140 -10092 -120 -10028
rect -5492 -10108 -120 -10092
rect -5492 -10172 -204 -10108
rect -140 -10172 -120 -10108
rect -5492 -10188 -120 -10172
rect -5492 -10252 -204 -10188
rect -140 -10252 -120 -10188
rect -5492 -10268 -120 -10252
rect -5492 -10332 -204 -10268
rect -140 -10332 -120 -10268
rect -5492 -10348 -120 -10332
rect -5492 -10412 -204 -10348
rect -140 -10412 -120 -10348
rect -5492 -10428 -120 -10412
rect -5492 -10492 -204 -10428
rect -140 -10492 -120 -10428
rect -5492 -10520 -120 -10492
rect 120 -5468 5492 -5440
rect 120 -5532 5408 -5468
rect 5472 -5532 5492 -5468
rect 120 -5548 5492 -5532
rect 120 -5612 5408 -5548
rect 5472 -5612 5492 -5548
rect 120 -5628 5492 -5612
rect 120 -5692 5408 -5628
rect 5472 -5692 5492 -5628
rect 120 -5708 5492 -5692
rect 120 -5772 5408 -5708
rect 5472 -5772 5492 -5708
rect 120 -5788 5492 -5772
rect 120 -5852 5408 -5788
rect 5472 -5852 5492 -5788
rect 120 -5868 5492 -5852
rect 120 -5932 5408 -5868
rect 5472 -5932 5492 -5868
rect 120 -5948 5492 -5932
rect 120 -6012 5408 -5948
rect 5472 -6012 5492 -5948
rect 120 -6028 5492 -6012
rect 120 -6092 5408 -6028
rect 5472 -6092 5492 -6028
rect 120 -6108 5492 -6092
rect 120 -6172 5408 -6108
rect 5472 -6172 5492 -6108
rect 120 -6188 5492 -6172
rect 120 -6252 5408 -6188
rect 5472 -6252 5492 -6188
rect 120 -6268 5492 -6252
rect 120 -6332 5408 -6268
rect 5472 -6332 5492 -6268
rect 120 -6348 5492 -6332
rect 120 -6412 5408 -6348
rect 5472 -6412 5492 -6348
rect 120 -6428 5492 -6412
rect 120 -6492 5408 -6428
rect 5472 -6492 5492 -6428
rect 120 -6508 5492 -6492
rect 120 -6572 5408 -6508
rect 5472 -6572 5492 -6508
rect 120 -6588 5492 -6572
rect 120 -6652 5408 -6588
rect 5472 -6652 5492 -6588
rect 120 -6668 5492 -6652
rect 120 -6732 5408 -6668
rect 5472 -6732 5492 -6668
rect 120 -6748 5492 -6732
rect 120 -6812 5408 -6748
rect 5472 -6812 5492 -6748
rect 120 -6828 5492 -6812
rect 120 -6892 5408 -6828
rect 5472 -6892 5492 -6828
rect 120 -6908 5492 -6892
rect 120 -6972 5408 -6908
rect 5472 -6972 5492 -6908
rect 120 -6988 5492 -6972
rect 120 -7052 5408 -6988
rect 5472 -7052 5492 -6988
rect 120 -7068 5492 -7052
rect 120 -7132 5408 -7068
rect 5472 -7132 5492 -7068
rect 120 -7148 5492 -7132
rect 120 -7212 5408 -7148
rect 5472 -7212 5492 -7148
rect 120 -7228 5492 -7212
rect 120 -7292 5408 -7228
rect 5472 -7292 5492 -7228
rect 120 -7308 5492 -7292
rect 120 -7372 5408 -7308
rect 5472 -7372 5492 -7308
rect 120 -7388 5492 -7372
rect 120 -7452 5408 -7388
rect 5472 -7452 5492 -7388
rect 120 -7468 5492 -7452
rect 120 -7532 5408 -7468
rect 5472 -7532 5492 -7468
rect 120 -7548 5492 -7532
rect 120 -7612 5408 -7548
rect 5472 -7612 5492 -7548
rect 120 -7628 5492 -7612
rect 120 -7692 5408 -7628
rect 5472 -7692 5492 -7628
rect 120 -7708 5492 -7692
rect 120 -7772 5408 -7708
rect 5472 -7772 5492 -7708
rect 120 -7788 5492 -7772
rect 120 -7852 5408 -7788
rect 5472 -7852 5492 -7788
rect 120 -7868 5492 -7852
rect 120 -7932 5408 -7868
rect 5472 -7932 5492 -7868
rect 120 -7948 5492 -7932
rect 120 -8012 5408 -7948
rect 5472 -8012 5492 -7948
rect 120 -8028 5492 -8012
rect 120 -8092 5408 -8028
rect 5472 -8092 5492 -8028
rect 120 -8108 5492 -8092
rect 120 -8172 5408 -8108
rect 5472 -8172 5492 -8108
rect 120 -8188 5492 -8172
rect 120 -8252 5408 -8188
rect 5472 -8252 5492 -8188
rect 120 -8268 5492 -8252
rect 120 -8332 5408 -8268
rect 5472 -8332 5492 -8268
rect 120 -8348 5492 -8332
rect 120 -8412 5408 -8348
rect 5472 -8412 5492 -8348
rect 120 -8428 5492 -8412
rect 120 -8492 5408 -8428
rect 5472 -8492 5492 -8428
rect 120 -8508 5492 -8492
rect 120 -8572 5408 -8508
rect 5472 -8572 5492 -8508
rect 120 -8588 5492 -8572
rect 120 -8652 5408 -8588
rect 5472 -8652 5492 -8588
rect 120 -8668 5492 -8652
rect 120 -8732 5408 -8668
rect 5472 -8732 5492 -8668
rect 120 -8748 5492 -8732
rect 120 -8812 5408 -8748
rect 5472 -8812 5492 -8748
rect 120 -8828 5492 -8812
rect 120 -8892 5408 -8828
rect 5472 -8892 5492 -8828
rect 120 -8908 5492 -8892
rect 120 -8972 5408 -8908
rect 5472 -8972 5492 -8908
rect 120 -8988 5492 -8972
rect 120 -9052 5408 -8988
rect 5472 -9052 5492 -8988
rect 120 -9068 5492 -9052
rect 120 -9132 5408 -9068
rect 5472 -9132 5492 -9068
rect 120 -9148 5492 -9132
rect 120 -9212 5408 -9148
rect 5472 -9212 5492 -9148
rect 120 -9228 5492 -9212
rect 120 -9292 5408 -9228
rect 5472 -9292 5492 -9228
rect 120 -9308 5492 -9292
rect 120 -9372 5408 -9308
rect 5472 -9372 5492 -9308
rect 120 -9388 5492 -9372
rect 120 -9452 5408 -9388
rect 5472 -9452 5492 -9388
rect 120 -9468 5492 -9452
rect 120 -9532 5408 -9468
rect 5472 -9532 5492 -9468
rect 120 -9548 5492 -9532
rect 120 -9612 5408 -9548
rect 5472 -9612 5492 -9548
rect 120 -9628 5492 -9612
rect 120 -9692 5408 -9628
rect 5472 -9692 5492 -9628
rect 120 -9708 5492 -9692
rect 120 -9772 5408 -9708
rect 5472 -9772 5492 -9708
rect 120 -9788 5492 -9772
rect 120 -9852 5408 -9788
rect 5472 -9852 5492 -9788
rect 120 -9868 5492 -9852
rect 120 -9932 5408 -9868
rect 5472 -9932 5492 -9868
rect 120 -9948 5492 -9932
rect 120 -10012 5408 -9948
rect 5472 -10012 5492 -9948
rect 120 -10028 5492 -10012
rect 120 -10092 5408 -10028
rect 5472 -10092 5492 -10028
rect 120 -10108 5492 -10092
rect 120 -10172 5408 -10108
rect 5472 -10172 5492 -10108
rect 120 -10188 5492 -10172
rect 120 -10252 5408 -10188
rect 5472 -10252 5492 -10188
rect 120 -10268 5492 -10252
rect 120 -10332 5408 -10268
rect 5472 -10332 5492 -10268
rect 120 -10348 5492 -10332
rect 120 -10412 5408 -10348
rect 5472 -10412 5492 -10348
rect 120 -10428 5492 -10412
rect 120 -10492 5408 -10428
rect 5472 -10492 5492 -10428
rect 120 -10520 5492 -10492
rect 5732 -5468 11104 -5440
rect 5732 -5532 11020 -5468
rect 11084 -5532 11104 -5468
rect 5732 -5548 11104 -5532
rect 5732 -5612 11020 -5548
rect 11084 -5612 11104 -5548
rect 5732 -5628 11104 -5612
rect 5732 -5692 11020 -5628
rect 11084 -5692 11104 -5628
rect 5732 -5708 11104 -5692
rect 5732 -5772 11020 -5708
rect 11084 -5772 11104 -5708
rect 5732 -5788 11104 -5772
rect 5732 -5852 11020 -5788
rect 11084 -5852 11104 -5788
rect 5732 -5868 11104 -5852
rect 5732 -5932 11020 -5868
rect 11084 -5932 11104 -5868
rect 5732 -5948 11104 -5932
rect 5732 -6012 11020 -5948
rect 11084 -6012 11104 -5948
rect 5732 -6028 11104 -6012
rect 5732 -6092 11020 -6028
rect 11084 -6092 11104 -6028
rect 5732 -6108 11104 -6092
rect 5732 -6172 11020 -6108
rect 11084 -6172 11104 -6108
rect 5732 -6188 11104 -6172
rect 5732 -6252 11020 -6188
rect 11084 -6252 11104 -6188
rect 5732 -6268 11104 -6252
rect 5732 -6332 11020 -6268
rect 11084 -6332 11104 -6268
rect 5732 -6348 11104 -6332
rect 5732 -6412 11020 -6348
rect 11084 -6412 11104 -6348
rect 5732 -6428 11104 -6412
rect 5732 -6492 11020 -6428
rect 11084 -6492 11104 -6428
rect 5732 -6508 11104 -6492
rect 5732 -6572 11020 -6508
rect 11084 -6572 11104 -6508
rect 5732 -6588 11104 -6572
rect 5732 -6652 11020 -6588
rect 11084 -6652 11104 -6588
rect 5732 -6668 11104 -6652
rect 5732 -6732 11020 -6668
rect 11084 -6732 11104 -6668
rect 5732 -6748 11104 -6732
rect 5732 -6812 11020 -6748
rect 11084 -6812 11104 -6748
rect 5732 -6828 11104 -6812
rect 5732 -6892 11020 -6828
rect 11084 -6892 11104 -6828
rect 5732 -6908 11104 -6892
rect 5732 -6972 11020 -6908
rect 11084 -6972 11104 -6908
rect 5732 -6988 11104 -6972
rect 5732 -7052 11020 -6988
rect 11084 -7052 11104 -6988
rect 5732 -7068 11104 -7052
rect 5732 -7132 11020 -7068
rect 11084 -7132 11104 -7068
rect 5732 -7148 11104 -7132
rect 5732 -7212 11020 -7148
rect 11084 -7212 11104 -7148
rect 5732 -7228 11104 -7212
rect 5732 -7292 11020 -7228
rect 11084 -7292 11104 -7228
rect 5732 -7308 11104 -7292
rect 5732 -7372 11020 -7308
rect 11084 -7372 11104 -7308
rect 5732 -7388 11104 -7372
rect 5732 -7452 11020 -7388
rect 11084 -7452 11104 -7388
rect 5732 -7468 11104 -7452
rect 5732 -7532 11020 -7468
rect 11084 -7532 11104 -7468
rect 5732 -7548 11104 -7532
rect 5732 -7612 11020 -7548
rect 11084 -7612 11104 -7548
rect 5732 -7628 11104 -7612
rect 5732 -7692 11020 -7628
rect 11084 -7692 11104 -7628
rect 5732 -7708 11104 -7692
rect 5732 -7772 11020 -7708
rect 11084 -7772 11104 -7708
rect 5732 -7788 11104 -7772
rect 5732 -7852 11020 -7788
rect 11084 -7852 11104 -7788
rect 5732 -7868 11104 -7852
rect 5732 -7932 11020 -7868
rect 11084 -7932 11104 -7868
rect 5732 -7948 11104 -7932
rect 5732 -8012 11020 -7948
rect 11084 -8012 11104 -7948
rect 5732 -8028 11104 -8012
rect 5732 -8092 11020 -8028
rect 11084 -8092 11104 -8028
rect 5732 -8108 11104 -8092
rect 5732 -8172 11020 -8108
rect 11084 -8172 11104 -8108
rect 5732 -8188 11104 -8172
rect 5732 -8252 11020 -8188
rect 11084 -8252 11104 -8188
rect 5732 -8268 11104 -8252
rect 5732 -8332 11020 -8268
rect 11084 -8332 11104 -8268
rect 5732 -8348 11104 -8332
rect 5732 -8412 11020 -8348
rect 11084 -8412 11104 -8348
rect 5732 -8428 11104 -8412
rect 5732 -8492 11020 -8428
rect 11084 -8492 11104 -8428
rect 5732 -8508 11104 -8492
rect 5732 -8572 11020 -8508
rect 11084 -8572 11104 -8508
rect 5732 -8588 11104 -8572
rect 5732 -8652 11020 -8588
rect 11084 -8652 11104 -8588
rect 5732 -8668 11104 -8652
rect 5732 -8732 11020 -8668
rect 11084 -8732 11104 -8668
rect 5732 -8748 11104 -8732
rect 5732 -8812 11020 -8748
rect 11084 -8812 11104 -8748
rect 5732 -8828 11104 -8812
rect 5732 -8892 11020 -8828
rect 11084 -8892 11104 -8828
rect 5732 -8908 11104 -8892
rect 5732 -8972 11020 -8908
rect 11084 -8972 11104 -8908
rect 5732 -8988 11104 -8972
rect 5732 -9052 11020 -8988
rect 11084 -9052 11104 -8988
rect 5732 -9068 11104 -9052
rect 5732 -9132 11020 -9068
rect 11084 -9132 11104 -9068
rect 5732 -9148 11104 -9132
rect 5732 -9212 11020 -9148
rect 11084 -9212 11104 -9148
rect 5732 -9228 11104 -9212
rect 5732 -9292 11020 -9228
rect 11084 -9292 11104 -9228
rect 5732 -9308 11104 -9292
rect 5732 -9372 11020 -9308
rect 11084 -9372 11104 -9308
rect 5732 -9388 11104 -9372
rect 5732 -9452 11020 -9388
rect 11084 -9452 11104 -9388
rect 5732 -9468 11104 -9452
rect 5732 -9532 11020 -9468
rect 11084 -9532 11104 -9468
rect 5732 -9548 11104 -9532
rect 5732 -9612 11020 -9548
rect 11084 -9612 11104 -9548
rect 5732 -9628 11104 -9612
rect 5732 -9692 11020 -9628
rect 11084 -9692 11104 -9628
rect 5732 -9708 11104 -9692
rect 5732 -9772 11020 -9708
rect 11084 -9772 11104 -9708
rect 5732 -9788 11104 -9772
rect 5732 -9852 11020 -9788
rect 11084 -9852 11104 -9788
rect 5732 -9868 11104 -9852
rect 5732 -9932 11020 -9868
rect 11084 -9932 11104 -9868
rect 5732 -9948 11104 -9932
rect 5732 -10012 11020 -9948
rect 11084 -10012 11104 -9948
rect 5732 -10028 11104 -10012
rect 5732 -10092 11020 -10028
rect 11084 -10092 11104 -10028
rect 5732 -10108 11104 -10092
rect 5732 -10172 11020 -10108
rect 11084 -10172 11104 -10108
rect 5732 -10188 11104 -10172
rect 5732 -10252 11020 -10188
rect 11084 -10252 11104 -10188
rect 5732 -10268 11104 -10252
rect 5732 -10332 11020 -10268
rect 11084 -10332 11104 -10268
rect 5732 -10348 11104 -10332
rect 5732 -10412 11020 -10348
rect 11084 -10412 11104 -10348
rect 5732 -10428 11104 -10412
rect 5732 -10492 11020 -10428
rect 11084 -10492 11104 -10428
rect 5732 -10520 11104 -10492
rect 11344 -5468 16716 -5440
rect 11344 -5532 16632 -5468
rect 16696 -5532 16716 -5468
rect 11344 -5548 16716 -5532
rect 11344 -5612 16632 -5548
rect 16696 -5612 16716 -5548
rect 11344 -5628 16716 -5612
rect 11344 -5692 16632 -5628
rect 16696 -5692 16716 -5628
rect 11344 -5708 16716 -5692
rect 11344 -5772 16632 -5708
rect 16696 -5772 16716 -5708
rect 11344 -5788 16716 -5772
rect 11344 -5852 16632 -5788
rect 16696 -5852 16716 -5788
rect 11344 -5868 16716 -5852
rect 11344 -5932 16632 -5868
rect 16696 -5932 16716 -5868
rect 11344 -5948 16716 -5932
rect 11344 -6012 16632 -5948
rect 16696 -6012 16716 -5948
rect 11344 -6028 16716 -6012
rect 11344 -6092 16632 -6028
rect 16696 -6092 16716 -6028
rect 11344 -6108 16716 -6092
rect 11344 -6172 16632 -6108
rect 16696 -6172 16716 -6108
rect 11344 -6188 16716 -6172
rect 11344 -6252 16632 -6188
rect 16696 -6252 16716 -6188
rect 11344 -6268 16716 -6252
rect 11344 -6332 16632 -6268
rect 16696 -6332 16716 -6268
rect 11344 -6348 16716 -6332
rect 11344 -6412 16632 -6348
rect 16696 -6412 16716 -6348
rect 11344 -6428 16716 -6412
rect 11344 -6492 16632 -6428
rect 16696 -6492 16716 -6428
rect 11344 -6508 16716 -6492
rect 11344 -6572 16632 -6508
rect 16696 -6572 16716 -6508
rect 11344 -6588 16716 -6572
rect 11344 -6652 16632 -6588
rect 16696 -6652 16716 -6588
rect 11344 -6668 16716 -6652
rect 11344 -6732 16632 -6668
rect 16696 -6732 16716 -6668
rect 11344 -6748 16716 -6732
rect 11344 -6812 16632 -6748
rect 16696 -6812 16716 -6748
rect 11344 -6828 16716 -6812
rect 11344 -6892 16632 -6828
rect 16696 -6892 16716 -6828
rect 11344 -6908 16716 -6892
rect 11344 -6972 16632 -6908
rect 16696 -6972 16716 -6908
rect 11344 -6988 16716 -6972
rect 11344 -7052 16632 -6988
rect 16696 -7052 16716 -6988
rect 11344 -7068 16716 -7052
rect 11344 -7132 16632 -7068
rect 16696 -7132 16716 -7068
rect 11344 -7148 16716 -7132
rect 11344 -7212 16632 -7148
rect 16696 -7212 16716 -7148
rect 11344 -7228 16716 -7212
rect 11344 -7292 16632 -7228
rect 16696 -7292 16716 -7228
rect 11344 -7308 16716 -7292
rect 11344 -7372 16632 -7308
rect 16696 -7372 16716 -7308
rect 11344 -7388 16716 -7372
rect 11344 -7452 16632 -7388
rect 16696 -7452 16716 -7388
rect 11344 -7468 16716 -7452
rect 11344 -7532 16632 -7468
rect 16696 -7532 16716 -7468
rect 11344 -7548 16716 -7532
rect 11344 -7612 16632 -7548
rect 16696 -7612 16716 -7548
rect 11344 -7628 16716 -7612
rect 11344 -7692 16632 -7628
rect 16696 -7692 16716 -7628
rect 11344 -7708 16716 -7692
rect 11344 -7772 16632 -7708
rect 16696 -7772 16716 -7708
rect 11344 -7788 16716 -7772
rect 11344 -7852 16632 -7788
rect 16696 -7852 16716 -7788
rect 11344 -7868 16716 -7852
rect 11344 -7932 16632 -7868
rect 16696 -7932 16716 -7868
rect 11344 -7948 16716 -7932
rect 11344 -8012 16632 -7948
rect 16696 -8012 16716 -7948
rect 11344 -8028 16716 -8012
rect 11344 -8092 16632 -8028
rect 16696 -8092 16716 -8028
rect 11344 -8108 16716 -8092
rect 11344 -8172 16632 -8108
rect 16696 -8172 16716 -8108
rect 11344 -8188 16716 -8172
rect 11344 -8252 16632 -8188
rect 16696 -8252 16716 -8188
rect 11344 -8268 16716 -8252
rect 11344 -8332 16632 -8268
rect 16696 -8332 16716 -8268
rect 11344 -8348 16716 -8332
rect 11344 -8412 16632 -8348
rect 16696 -8412 16716 -8348
rect 11344 -8428 16716 -8412
rect 11344 -8492 16632 -8428
rect 16696 -8492 16716 -8428
rect 11344 -8508 16716 -8492
rect 11344 -8572 16632 -8508
rect 16696 -8572 16716 -8508
rect 11344 -8588 16716 -8572
rect 11344 -8652 16632 -8588
rect 16696 -8652 16716 -8588
rect 11344 -8668 16716 -8652
rect 11344 -8732 16632 -8668
rect 16696 -8732 16716 -8668
rect 11344 -8748 16716 -8732
rect 11344 -8812 16632 -8748
rect 16696 -8812 16716 -8748
rect 11344 -8828 16716 -8812
rect 11344 -8892 16632 -8828
rect 16696 -8892 16716 -8828
rect 11344 -8908 16716 -8892
rect 11344 -8972 16632 -8908
rect 16696 -8972 16716 -8908
rect 11344 -8988 16716 -8972
rect 11344 -9052 16632 -8988
rect 16696 -9052 16716 -8988
rect 11344 -9068 16716 -9052
rect 11344 -9132 16632 -9068
rect 16696 -9132 16716 -9068
rect 11344 -9148 16716 -9132
rect 11344 -9212 16632 -9148
rect 16696 -9212 16716 -9148
rect 11344 -9228 16716 -9212
rect 11344 -9292 16632 -9228
rect 16696 -9292 16716 -9228
rect 11344 -9308 16716 -9292
rect 11344 -9372 16632 -9308
rect 16696 -9372 16716 -9308
rect 11344 -9388 16716 -9372
rect 11344 -9452 16632 -9388
rect 16696 -9452 16716 -9388
rect 11344 -9468 16716 -9452
rect 11344 -9532 16632 -9468
rect 16696 -9532 16716 -9468
rect 11344 -9548 16716 -9532
rect 11344 -9612 16632 -9548
rect 16696 -9612 16716 -9548
rect 11344 -9628 16716 -9612
rect 11344 -9692 16632 -9628
rect 16696 -9692 16716 -9628
rect 11344 -9708 16716 -9692
rect 11344 -9772 16632 -9708
rect 16696 -9772 16716 -9708
rect 11344 -9788 16716 -9772
rect 11344 -9852 16632 -9788
rect 16696 -9852 16716 -9788
rect 11344 -9868 16716 -9852
rect 11344 -9932 16632 -9868
rect 16696 -9932 16716 -9868
rect 11344 -9948 16716 -9932
rect 11344 -10012 16632 -9948
rect 16696 -10012 16716 -9948
rect 11344 -10028 16716 -10012
rect 11344 -10092 16632 -10028
rect 16696 -10092 16716 -10028
rect 11344 -10108 16716 -10092
rect 11344 -10172 16632 -10108
rect 16696 -10172 16716 -10108
rect 11344 -10188 16716 -10172
rect 11344 -10252 16632 -10188
rect 16696 -10252 16716 -10188
rect 11344 -10268 16716 -10252
rect 11344 -10332 16632 -10268
rect 16696 -10332 16716 -10268
rect 11344 -10348 16716 -10332
rect 11344 -10412 16632 -10348
rect 16696 -10412 16716 -10348
rect 11344 -10428 16716 -10412
rect 11344 -10492 16632 -10428
rect 16696 -10492 16716 -10428
rect 11344 -10520 16716 -10492
rect 16956 -5468 22328 -5440
rect 16956 -5532 22244 -5468
rect 22308 -5532 22328 -5468
rect 16956 -5548 22328 -5532
rect 16956 -5612 22244 -5548
rect 22308 -5612 22328 -5548
rect 16956 -5628 22328 -5612
rect 16956 -5692 22244 -5628
rect 22308 -5692 22328 -5628
rect 16956 -5708 22328 -5692
rect 16956 -5772 22244 -5708
rect 22308 -5772 22328 -5708
rect 16956 -5788 22328 -5772
rect 16956 -5852 22244 -5788
rect 22308 -5852 22328 -5788
rect 16956 -5868 22328 -5852
rect 16956 -5932 22244 -5868
rect 22308 -5932 22328 -5868
rect 16956 -5948 22328 -5932
rect 16956 -6012 22244 -5948
rect 22308 -6012 22328 -5948
rect 16956 -6028 22328 -6012
rect 16956 -6092 22244 -6028
rect 22308 -6092 22328 -6028
rect 16956 -6108 22328 -6092
rect 16956 -6172 22244 -6108
rect 22308 -6172 22328 -6108
rect 16956 -6188 22328 -6172
rect 16956 -6252 22244 -6188
rect 22308 -6252 22328 -6188
rect 16956 -6268 22328 -6252
rect 16956 -6332 22244 -6268
rect 22308 -6332 22328 -6268
rect 16956 -6348 22328 -6332
rect 16956 -6412 22244 -6348
rect 22308 -6412 22328 -6348
rect 16956 -6428 22328 -6412
rect 16956 -6492 22244 -6428
rect 22308 -6492 22328 -6428
rect 16956 -6508 22328 -6492
rect 16956 -6572 22244 -6508
rect 22308 -6572 22328 -6508
rect 16956 -6588 22328 -6572
rect 16956 -6652 22244 -6588
rect 22308 -6652 22328 -6588
rect 16956 -6668 22328 -6652
rect 16956 -6732 22244 -6668
rect 22308 -6732 22328 -6668
rect 16956 -6748 22328 -6732
rect 16956 -6812 22244 -6748
rect 22308 -6812 22328 -6748
rect 16956 -6828 22328 -6812
rect 16956 -6892 22244 -6828
rect 22308 -6892 22328 -6828
rect 16956 -6908 22328 -6892
rect 16956 -6972 22244 -6908
rect 22308 -6972 22328 -6908
rect 16956 -6988 22328 -6972
rect 16956 -7052 22244 -6988
rect 22308 -7052 22328 -6988
rect 16956 -7068 22328 -7052
rect 16956 -7132 22244 -7068
rect 22308 -7132 22328 -7068
rect 16956 -7148 22328 -7132
rect 16956 -7212 22244 -7148
rect 22308 -7212 22328 -7148
rect 16956 -7228 22328 -7212
rect 16956 -7292 22244 -7228
rect 22308 -7292 22328 -7228
rect 16956 -7308 22328 -7292
rect 16956 -7372 22244 -7308
rect 22308 -7372 22328 -7308
rect 16956 -7388 22328 -7372
rect 16956 -7452 22244 -7388
rect 22308 -7452 22328 -7388
rect 16956 -7468 22328 -7452
rect 16956 -7532 22244 -7468
rect 22308 -7532 22328 -7468
rect 16956 -7548 22328 -7532
rect 16956 -7612 22244 -7548
rect 22308 -7612 22328 -7548
rect 16956 -7628 22328 -7612
rect 16956 -7692 22244 -7628
rect 22308 -7692 22328 -7628
rect 16956 -7708 22328 -7692
rect 16956 -7772 22244 -7708
rect 22308 -7772 22328 -7708
rect 16956 -7788 22328 -7772
rect 16956 -7852 22244 -7788
rect 22308 -7852 22328 -7788
rect 16956 -7868 22328 -7852
rect 16956 -7932 22244 -7868
rect 22308 -7932 22328 -7868
rect 16956 -7948 22328 -7932
rect 16956 -8012 22244 -7948
rect 22308 -8012 22328 -7948
rect 16956 -8028 22328 -8012
rect 16956 -8092 22244 -8028
rect 22308 -8092 22328 -8028
rect 16956 -8108 22328 -8092
rect 16956 -8172 22244 -8108
rect 22308 -8172 22328 -8108
rect 16956 -8188 22328 -8172
rect 16956 -8252 22244 -8188
rect 22308 -8252 22328 -8188
rect 16956 -8268 22328 -8252
rect 16956 -8332 22244 -8268
rect 22308 -8332 22328 -8268
rect 16956 -8348 22328 -8332
rect 16956 -8412 22244 -8348
rect 22308 -8412 22328 -8348
rect 16956 -8428 22328 -8412
rect 16956 -8492 22244 -8428
rect 22308 -8492 22328 -8428
rect 16956 -8508 22328 -8492
rect 16956 -8572 22244 -8508
rect 22308 -8572 22328 -8508
rect 16956 -8588 22328 -8572
rect 16956 -8652 22244 -8588
rect 22308 -8652 22328 -8588
rect 16956 -8668 22328 -8652
rect 16956 -8732 22244 -8668
rect 22308 -8732 22328 -8668
rect 16956 -8748 22328 -8732
rect 16956 -8812 22244 -8748
rect 22308 -8812 22328 -8748
rect 16956 -8828 22328 -8812
rect 16956 -8892 22244 -8828
rect 22308 -8892 22328 -8828
rect 16956 -8908 22328 -8892
rect 16956 -8972 22244 -8908
rect 22308 -8972 22328 -8908
rect 16956 -8988 22328 -8972
rect 16956 -9052 22244 -8988
rect 22308 -9052 22328 -8988
rect 16956 -9068 22328 -9052
rect 16956 -9132 22244 -9068
rect 22308 -9132 22328 -9068
rect 16956 -9148 22328 -9132
rect 16956 -9212 22244 -9148
rect 22308 -9212 22328 -9148
rect 16956 -9228 22328 -9212
rect 16956 -9292 22244 -9228
rect 22308 -9292 22328 -9228
rect 16956 -9308 22328 -9292
rect 16956 -9372 22244 -9308
rect 22308 -9372 22328 -9308
rect 16956 -9388 22328 -9372
rect 16956 -9452 22244 -9388
rect 22308 -9452 22328 -9388
rect 16956 -9468 22328 -9452
rect 16956 -9532 22244 -9468
rect 22308 -9532 22328 -9468
rect 16956 -9548 22328 -9532
rect 16956 -9612 22244 -9548
rect 22308 -9612 22328 -9548
rect 16956 -9628 22328 -9612
rect 16956 -9692 22244 -9628
rect 22308 -9692 22328 -9628
rect 16956 -9708 22328 -9692
rect 16956 -9772 22244 -9708
rect 22308 -9772 22328 -9708
rect 16956 -9788 22328 -9772
rect 16956 -9852 22244 -9788
rect 22308 -9852 22328 -9788
rect 16956 -9868 22328 -9852
rect 16956 -9932 22244 -9868
rect 22308 -9932 22328 -9868
rect 16956 -9948 22328 -9932
rect 16956 -10012 22244 -9948
rect 22308 -10012 22328 -9948
rect 16956 -10028 22328 -10012
rect 16956 -10092 22244 -10028
rect 22308 -10092 22328 -10028
rect 16956 -10108 22328 -10092
rect 16956 -10172 22244 -10108
rect 22308 -10172 22328 -10108
rect 16956 -10188 22328 -10172
rect 16956 -10252 22244 -10188
rect 22308 -10252 22328 -10188
rect 16956 -10268 22328 -10252
rect 16956 -10332 22244 -10268
rect 22308 -10332 22328 -10268
rect 16956 -10348 22328 -10332
rect 16956 -10412 22244 -10348
rect 22308 -10412 22328 -10348
rect 16956 -10428 22328 -10412
rect 16956 -10492 22244 -10428
rect 22308 -10492 22328 -10428
rect 16956 -10520 22328 -10492
rect 22568 -5468 27940 -5440
rect 22568 -5532 27856 -5468
rect 27920 -5532 27940 -5468
rect 22568 -5548 27940 -5532
rect 22568 -5612 27856 -5548
rect 27920 -5612 27940 -5548
rect 22568 -5628 27940 -5612
rect 22568 -5692 27856 -5628
rect 27920 -5692 27940 -5628
rect 22568 -5708 27940 -5692
rect 22568 -5772 27856 -5708
rect 27920 -5772 27940 -5708
rect 22568 -5788 27940 -5772
rect 22568 -5852 27856 -5788
rect 27920 -5852 27940 -5788
rect 22568 -5868 27940 -5852
rect 22568 -5932 27856 -5868
rect 27920 -5932 27940 -5868
rect 22568 -5948 27940 -5932
rect 22568 -6012 27856 -5948
rect 27920 -6012 27940 -5948
rect 22568 -6028 27940 -6012
rect 22568 -6092 27856 -6028
rect 27920 -6092 27940 -6028
rect 22568 -6108 27940 -6092
rect 22568 -6172 27856 -6108
rect 27920 -6172 27940 -6108
rect 22568 -6188 27940 -6172
rect 22568 -6252 27856 -6188
rect 27920 -6252 27940 -6188
rect 22568 -6268 27940 -6252
rect 22568 -6332 27856 -6268
rect 27920 -6332 27940 -6268
rect 22568 -6348 27940 -6332
rect 22568 -6412 27856 -6348
rect 27920 -6412 27940 -6348
rect 22568 -6428 27940 -6412
rect 22568 -6492 27856 -6428
rect 27920 -6492 27940 -6428
rect 22568 -6508 27940 -6492
rect 22568 -6572 27856 -6508
rect 27920 -6572 27940 -6508
rect 22568 -6588 27940 -6572
rect 22568 -6652 27856 -6588
rect 27920 -6652 27940 -6588
rect 22568 -6668 27940 -6652
rect 22568 -6732 27856 -6668
rect 27920 -6732 27940 -6668
rect 22568 -6748 27940 -6732
rect 22568 -6812 27856 -6748
rect 27920 -6812 27940 -6748
rect 22568 -6828 27940 -6812
rect 22568 -6892 27856 -6828
rect 27920 -6892 27940 -6828
rect 22568 -6908 27940 -6892
rect 22568 -6972 27856 -6908
rect 27920 -6972 27940 -6908
rect 22568 -6988 27940 -6972
rect 22568 -7052 27856 -6988
rect 27920 -7052 27940 -6988
rect 22568 -7068 27940 -7052
rect 22568 -7132 27856 -7068
rect 27920 -7132 27940 -7068
rect 22568 -7148 27940 -7132
rect 22568 -7212 27856 -7148
rect 27920 -7212 27940 -7148
rect 22568 -7228 27940 -7212
rect 22568 -7292 27856 -7228
rect 27920 -7292 27940 -7228
rect 22568 -7308 27940 -7292
rect 22568 -7372 27856 -7308
rect 27920 -7372 27940 -7308
rect 22568 -7388 27940 -7372
rect 22568 -7452 27856 -7388
rect 27920 -7452 27940 -7388
rect 22568 -7468 27940 -7452
rect 22568 -7532 27856 -7468
rect 27920 -7532 27940 -7468
rect 22568 -7548 27940 -7532
rect 22568 -7612 27856 -7548
rect 27920 -7612 27940 -7548
rect 22568 -7628 27940 -7612
rect 22568 -7692 27856 -7628
rect 27920 -7692 27940 -7628
rect 22568 -7708 27940 -7692
rect 22568 -7772 27856 -7708
rect 27920 -7772 27940 -7708
rect 22568 -7788 27940 -7772
rect 22568 -7852 27856 -7788
rect 27920 -7852 27940 -7788
rect 22568 -7868 27940 -7852
rect 22568 -7932 27856 -7868
rect 27920 -7932 27940 -7868
rect 22568 -7948 27940 -7932
rect 22568 -8012 27856 -7948
rect 27920 -8012 27940 -7948
rect 22568 -8028 27940 -8012
rect 22568 -8092 27856 -8028
rect 27920 -8092 27940 -8028
rect 22568 -8108 27940 -8092
rect 22568 -8172 27856 -8108
rect 27920 -8172 27940 -8108
rect 22568 -8188 27940 -8172
rect 22568 -8252 27856 -8188
rect 27920 -8252 27940 -8188
rect 22568 -8268 27940 -8252
rect 22568 -8332 27856 -8268
rect 27920 -8332 27940 -8268
rect 22568 -8348 27940 -8332
rect 22568 -8412 27856 -8348
rect 27920 -8412 27940 -8348
rect 22568 -8428 27940 -8412
rect 22568 -8492 27856 -8428
rect 27920 -8492 27940 -8428
rect 22568 -8508 27940 -8492
rect 22568 -8572 27856 -8508
rect 27920 -8572 27940 -8508
rect 22568 -8588 27940 -8572
rect 22568 -8652 27856 -8588
rect 27920 -8652 27940 -8588
rect 22568 -8668 27940 -8652
rect 22568 -8732 27856 -8668
rect 27920 -8732 27940 -8668
rect 22568 -8748 27940 -8732
rect 22568 -8812 27856 -8748
rect 27920 -8812 27940 -8748
rect 22568 -8828 27940 -8812
rect 22568 -8892 27856 -8828
rect 27920 -8892 27940 -8828
rect 22568 -8908 27940 -8892
rect 22568 -8972 27856 -8908
rect 27920 -8972 27940 -8908
rect 22568 -8988 27940 -8972
rect 22568 -9052 27856 -8988
rect 27920 -9052 27940 -8988
rect 22568 -9068 27940 -9052
rect 22568 -9132 27856 -9068
rect 27920 -9132 27940 -9068
rect 22568 -9148 27940 -9132
rect 22568 -9212 27856 -9148
rect 27920 -9212 27940 -9148
rect 22568 -9228 27940 -9212
rect 22568 -9292 27856 -9228
rect 27920 -9292 27940 -9228
rect 22568 -9308 27940 -9292
rect 22568 -9372 27856 -9308
rect 27920 -9372 27940 -9308
rect 22568 -9388 27940 -9372
rect 22568 -9452 27856 -9388
rect 27920 -9452 27940 -9388
rect 22568 -9468 27940 -9452
rect 22568 -9532 27856 -9468
rect 27920 -9532 27940 -9468
rect 22568 -9548 27940 -9532
rect 22568 -9612 27856 -9548
rect 27920 -9612 27940 -9548
rect 22568 -9628 27940 -9612
rect 22568 -9692 27856 -9628
rect 27920 -9692 27940 -9628
rect 22568 -9708 27940 -9692
rect 22568 -9772 27856 -9708
rect 27920 -9772 27940 -9708
rect 22568 -9788 27940 -9772
rect 22568 -9852 27856 -9788
rect 27920 -9852 27940 -9788
rect 22568 -9868 27940 -9852
rect 22568 -9932 27856 -9868
rect 27920 -9932 27940 -9868
rect 22568 -9948 27940 -9932
rect 22568 -10012 27856 -9948
rect 27920 -10012 27940 -9948
rect 22568 -10028 27940 -10012
rect 22568 -10092 27856 -10028
rect 27920 -10092 27940 -10028
rect 22568 -10108 27940 -10092
rect 22568 -10172 27856 -10108
rect 27920 -10172 27940 -10108
rect 22568 -10188 27940 -10172
rect 22568 -10252 27856 -10188
rect 27920 -10252 27940 -10188
rect 22568 -10268 27940 -10252
rect 22568 -10332 27856 -10268
rect 27920 -10332 27940 -10268
rect 22568 -10348 27940 -10332
rect 22568 -10412 27856 -10348
rect 27920 -10412 27940 -10348
rect 22568 -10428 27940 -10412
rect 22568 -10492 27856 -10428
rect 27920 -10492 27940 -10428
rect 22568 -10520 27940 -10492
rect 28180 -5468 33552 -5440
rect 28180 -5532 33468 -5468
rect 33532 -5532 33552 -5468
rect 28180 -5548 33552 -5532
rect 28180 -5612 33468 -5548
rect 33532 -5612 33552 -5548
rect 28180 -5628 33552 -5612
rect 28180 -5692 33468 -5628
rect 33532 -5692 33552 -5628
rect 28180 -5708 33552 -5692
rect 28180 -5772 33468 -5708
rect 33532 -5772 33552 -5708
rect 28180 -5788 33552 -5772
rect 28180 -5852 33468 -5788
rect 33532 -5852 33552 -5788
rect 28180 -5868 33552 -5852
rect 28180 -5932 33468 -5868
rect 33532 -5932 33552 -5868
rect 28180 -5948 33552 -5932
rect 28180 -6012 33468 -5948
rect 33532 -6012 33552 -5948
rect 28180 -6028 33552 -6012
rect 28180 -6092 33468 -6028
rect 33532 -6092 33552 -6028
rect 28180 -6108 33552 -6092
rect 28180 -6172 33468 -6108
rect 33532 -6172 33552 -6108
rect 28180 -6188 33552 -6172
rect 28180 -6252 33468 -6188
rect 33532 -6252 33552 -6188
rect 28180 -6268 33552 -6252
rect 28180 -6332 33468 -6268
rect 33532 -6332 33552 -6268
rect 28180 -6348 33552 -6332
rect 28180 -6412 33468 -6348
rect 33532 -6412 33552 -6348
rect 28180 -6428 33552 -6412
rect 28180 -6492 33468 -6428
rect 33532 -6492 33552 -6428
rect 28180 -6508 33552 -6492
rect 28180 -6572 33468 -6508
rect 33532 -6572 33552 -6508
rect 28180 -6588 33552 -6572
rect 28180 -6652 33468 -6588
rect 33532 -6652 33552 -6588
rect 28180 -6668 33552 -6652
rect 28180 -6732 33468 -6668
rect 33532 -6732 33552 -6668
rect 28180 -6748 33552 -6732
rect 28180 -6812 33468 -6748
rect 33532 -6812 33552 -6748
rect 28180 -6828 33552 -6812
rect 28180 -6892 33468 -6828
rect 33532 -6892 33552 -6828
rect 28180 -6908 33552 -6892
rect 28180 -6972 33468 -6908
rect 33532 -6972 33552 -6908
rect 28180 -6988 33552 -6972
rect 28180 -7052 33468 -6988
rect 33532 -7052 33552 -6988
rect 28180 -7068 33552 -7052
rect 28180 -7132 33468 -7068
rect 33532 -7132 33552 -7068
rect 28180 -7148 33552 -7132
rect 28180 -7212 33468 -7148
rect 33532 -7212 33552 -7148
rect 28180 -7228 33552 -7212
rect 28180 -7292 33468 -7228
rect 33532 -7292 33552 -7228
rect 28180 -7308 33552 -7292
rect 28180 -7372 33468 -7308
rect 33532 -7372 33552 -7308
rect 28180 -7388 33552 -7372
rect 28180 -7452 33468 -7388
rect 33532 -7452 33552 -7388
rect 28180 -7468 33552 -7452
rect 28180 -7532 33468 -7468
rect 33532 -7532 33552 -7468
rect 28180 -7548 33552 -7532
rect 28180 -7612 33468 -7548
rect 33532 -7612 33552 -7548
rect 28180 -7628 33552 -7612
rect 28180 -7692 33468 -7628
rect 33532 -7692 33552 -7628
rect 28180 -7708 33552 -7692
rect 28180 -7772 33468 -7708
rect 33532 -7772 33552 -7708
rect 28180 -7788 33552 -7772
rect 28180 -7852 33468 -7788
rect 33532 -7852 33552 -7788
rect 28180 -7868 33552 -7852
rect 28180 -7932 33468 -7868
rect 33532 -7932 33552 -7868
rect 28180 -7948 33552 -7932
rect 28180 -8012 33468 -7948
rect 33532 -8012 33552 -7948
rect 28180 -8028 33552 -8012
rect 28180 -8092 33468 -8028
rect 33532 -8092 33552 -8028
rect 28180 -8108 33552 -8092
rect 28180 -8172 33468 -8108
rect 33532 -8172 33552 -8108
rect 28180 -8188 33552 -8172
rect 28180 -8252 33468 -8188
rect 33532 -8252 33552 -8188
rect 28180 -8268 33552 -8252
rect 28180 -8332 33468 -8268
rect 33532 -8332 33552 -8268
rect 28180 -8348 33552 -8332
rect 28180 -8412 33468 -8348
rect 33532 -8412 33552 -8348
rect 28180 -8428 33552 -8412
rect 28180 -8492 33468 -8428
rect 33532 -8492 33552 -8428
rect 28180 -8508 33552 -8492
rect 28180 -8572 33468 -8508
rect 33532 -8572 33552 -8508
rect 28180 -8588 33552 -8572
rect 28180 -8652 33468 -8588
rect 33532 -8652 33552 -8588
rect 28180 -8668 33552 -8652
rect 28180 -8732 33468 -8668
rect 33532 -8732 33552 -8668
rect 28180 -8748 33552 -8732
rect 28180 -8812 33468 -8748
rect 33532 -8812 33552 -8748
rect 28180 -8828 33552 -8812
rect 28180 -8892 33468 -8828
rect 33532 -8892 33552 -8828
rect 28180 -8908 33552 -8892
rect 28180 -8972 33468 -8908
rect 33532 -8972 33552 -8908
rect 28180 -8988 33552 -8972
rect 28180 -9052 33468 -8988
rect 33532 -9052 33552 -8988
rect 28180 -9068 33552 -9052
rect 28180 -9132 33468 -9068
rect 33532 -9132 33552 -9068
rect 28180 -9148 33552 -9132
rect 28180 -9212 33468 -9148
rect 33532 -9212 33552 -9148
rect 28180 -9228 33552 -9212
rect 28180 -9292 33468 -9228
rect 33532 -9292 33552 -9228
rect 28180 -9308 33552 -9292
rect 28180 -9372 33468 -9308
rect 33532 -9372 33552 -9308
rect 28180 -9388 33552 -9372
rect 28180 -9452 33468 -9388
rect 33532 -9452 33552 -9388
rect 28180 -9468 33552 -9452
rect 28180 -9532 33468 -9468
rect 33532 -9532 33552 -9468
rect 28180 -9548 33552 -9532
rect 28180 -9612 33468 -9548
rect 33532 -9612 33552 -9548
rect 28180 -9628 33552 -9612
rect 28180 -9692 33468 -9628
rect 33532 -9692 33552 -9628
rect 28180 -9708 33552 -9692
rect 28180 -9772 33468 -9708
rect 33532 -9772 33552 -9708
rect 28180 -9788 33552 -9772
rect 28180 -9852 33468 -9788
rect 33532 -9852 33552 -9788
rect 28180 -9868 33552 -9852
rect 28180 -9932 33468 -9868
rect 33532 -9932 33552 -9868
rect 28180 -9948 33552 -9932
rect 28180 -10012 33468 -9948
rect 33532 -10012 33552 -9948
rect 28180 -10028 33552 -10012
rect 28180 -10092 33468 -10028
rect 33532 -10092 33552 -10028
rect 28180 -10108 33552 -10092
rect 28180 -10172 33468 -10108
rect 33532 -10172 33552 -10108
rect 28180 -10188 33552 -10172
rect 28180 -10252 33468 -10188
rect 33532 -10252 33552 -10188
rect 28180 -10268 33552 -10252
rect 28180 -10332 33468 -10268
rect 33532 -10332 33552 -10268
rect 28180 -10348 33552 -10332
rect 28180 -10412 33468 -10348
rect 33532 -10412 33552 -10348
rect 28180 -10428 33552 -10412
rect 28180 -10492 33468 -10428
rect 33532 -10492 33552 -10428
rect 28180 -10520 33552 -10492
rect 33792 -5468 39164 -5440
rect 33792 -5532 39080 -5468
rect 39144 -5532 39164 -5468
rect 33792 -5548 39164 -5532
rect 33792 -5612 39080 -5548
rect 39144 -5612 39164 -5548
rect 33792 -5628 39164 -5612
rect 33792 -5692 39080 -5628
rect 39144 -5692 39164 -5628
rect 33792 -5708 39164 -5692
rect 33792 -5772 39080 -5708
rect 39144 -5772 39164 -5708
rect 33792 -5788 39164 -5772
rect 33792 -5852 39080 -5788
rect 39144 -5852 39164 -5788
rect 33792 -5868 39164 -5852
rect 33792 -5932 39080 -5868
rect 39144 -5932 39164 -5868
rect 33792 -5948 39164 -5932
rect 33792 -6012 39080 -5948
rect 39144 -6012 39164 -5948
rect 33792 -6028 39164 -6012
rect 33792 -6092 39080 -6028
rect 39144 -6092 39164 -6028
rect 33792 -6108 39164 -6092
rect 33792 -6172 39080 -6108
rect 39144 -6172 39164 -6108
rect 33792 -6188 39164 -6172
rect 33792 -6252 39080 -6188
rect 39144 -6252 39164 -6188
rect 33792 -6268 39164 -6252
rect 33792 -6332 39080 -6268
rect 39144 -6332 39164 -6268
rect 33792 -6348 39164 -6332
rect 33792 -6412 39080 -6348
rect 39144 -6412 39164 -6348
rect 33792 -6428 39164 -6412
rect 33792 -6492 39080 -6428
rect 39144 -6492 39164 -6428
rect 33792 -6508 39164 -6492
rect 33792 -6572 39080 -6508
rect 39144 -6572 39164 -6508
rect 33792 -6588 39164 -6572
rect 33792 -6652 39080 -6588
rect 39144 -6652 39164 -6588
rect 33792 -6668 39164 -6652
rect 33792 -6732 39080 -6668
rect 39144 -6732 39164 -6668
rect 33792 -6748 39164 -6732
rect 33792 -6812 39080 -6748
rect 39144 -6812 39164 -6748
rect 33792 -6828 39164 -6812
rect 33792 -6892 39080 -6828
rect 39144 -6892 39164 -6828
rect 33792 -6908 39164 -6892
rect 33792 -6972 39080 -6908
rect 39144 -6972 39164 -6908
rect 33792 -6988 39164 -6972
rect 33792 -7052 39080 -6988
rect 39144 -7052 39164 -6988
rect 33792 -7068 39164 -7052
rect 33792 -7132 39080 -7068
rect 39144 -7132 39164 -7068
rect 33792 -7148 39164 -7132
rect 33792 -7212 39080 -7148
rect 39144 -7212 39164 -7148
rect 33792 -7228 39164 -7212
rect 33792 -7292 39080 -7228
rect 39144 -7292 39164 -7228
rect 33792 -7308 39164 -7292
rect 33792 -7372 39080 -7308
rect 39144 -7372 39164 -7308
rect 33792 -7388 39164 -7372
rect 33792 -7452 39080 -7388
rect 39144 -7452 39164 -7388
rect 33792 -7468 39164 -7452
rect 33792 -7532 39080 -7468
rect 39144 -7532 39164 -7468
rect 33792 -7548 39164 -7532
rect 33792 -7612 39080 -7548
rect 39144 -7612 39164 -7548
rect 33792 -7628 39164 -7612
rect 33792 -7692 39080 -7628
rect 39144 -7692 39164 -7628
rect 33792 -7708 39164 -7692
rect 33792 -7772 39080 -7708
rect 39144 -7772 39164 -7708
rect 33792 -7788 39164 -7772
rect 33792 -7852 39080 -7788
rect 39144 -7852 39164 -7788
rect 33792 -7868 39164 -7852
rect 33792 -7932 39080 -7868
rect 39144 -7932 39164 -7868
rect 33792 -7948 39164 -7932
rect 33792 -8012 39080 -7948
rect 39144 -8012 39164 -7948
rect 33792 -8028 39164 -8012
rect 33792 -8092 39080 -8028
rect 39144 -8092 39164 -8028
rect 33792 -8108 39164 -8092
rect 33792 -8172 39080 -8108
rect 39144 -8172 39164 -8108
rect 33792 -8188 39164 -8172
rect 33792 -8252 39080 -8188
rect 39144 -8252 39164 -8188
rect 33792 -8268 39164 -8252
rect 33792 -8332 39080 -8268
rect 39144 -8332 39164 -8268
rect 33792 -8348 39164 -8332
rect 33792 -8412 39080 -8348
rect 39144 -8412 39164 -8348
rect 33792 -8428 39164 -8412
rect 33792 -8492 39080 -8428
rect 39144 -8492 39164 -8428
rect 33792 -8508 39164 -8492
rect 33792 -8572 39080 -8508
rect 39144 -8572 39164 -8508
rect 33792 -8588 39164 -8572
rect 33792 -8652 39080 -8588
rect 39144 -8652 39164 -8588
rect 33792 -8668 39164 -8652
rect 33792 -8732 39080 -8668
rect 39144 -8732 39164 -8668
rect 33792 -8748 39164 -8732
rect 33792 -8812 39080 -8748
rect 39144 -8812 39164 -8748
rect 33792 -8828 39164 -8812
rect 33792 -8892 39080 -8828
rect 39144 -8892 39164 -8828
rect 33792 -8908 39164 -8892
rect 33792 -8972 39080 -8908
rect 39144 -8972 39164 -8908
rect 33792 -8988 39164 -8972
rect 33792 -9052 39080 -8988
rect 39144 -9052 39164 -8988
rect 33792 -9068 39164 -9052
rect 33792 -9132 39080 -9068
rect 39144 -9132 39164 -9068
rect 33792 -9148 39164 -9132
rect 33792 -9212 39080 -9148
rect 39144 -9212 39164 -9148
rect 33792 -9228 39164 -9212
rect 33792 -9292 39080 -9228
rect 39144 -9292 39164 -9228
rect 33792 -9308 39164 -9292
rect 33792 -9372 39080 -9308
rect 39144 -9372 39164 -9308
rect 33792 -9388 39164 -9372
rect 33792 -9452 39080 -9388
rect 39144 -9452 39164 -9388
rect 33792 -9468 39164 -9452
rect 33792 -9532 39080 -9468
rect 39144 -9532 39164 -9468
rect 33792 -9548 39164 -9532
rect 33792 -9612 39080 -9548
rect 39144 -9612 39164 -9548
rect 33792 -9628 39164 -9612
rect 33792 -9692 39080 -9628
rect 39144 -9692 39164 -9628
rect 33792 -9708 39164 -9692
rect 33792 -9772 39080 -9708
rect 39144 -9772 39164 -9708
rect 33792 -9788 39164 -9772
rect 33792 -9852 39080 -9788
rect 39144 -9852 39164 -9788
rect 33792 -9868 39164 -9852
rect 33792 -9932 39080 -9868
rect 39144 -9932 39164 -9868
rect 33792 -9948 39164 -9932
rect 33792 -10012 39080 -9948
rect 39144 -10012 39164 -9948
rect 33792 -10028 39164 -10012
rect 33792 -10092 39080 -10028
rect 39144 -10092 39164 -10028
rect 33792 -10108 39164 -10092
rect 33792 -10172 39080 -10108
rect 39144 -10172 39164 -10108
rect 33792 -10188 39164 -10172
rect 33792 -10252 39080 -10188
rect 39144 -10252 39164 -10188
rect 33792 -10268 39164 -10252
rect 33792 -10332 39080 -10268
rect 39144 -10332 39164 -10268
rect 33792 -10348 39164 -10332
rect 33792 -10412 39080 -10348
rect 39144 -10412 39164 -10348
rect 33792 -10428 39164 -10412
rect 33792 -10492 39080 -10428
rect 39144 -10492 39164 -10428
rect 33792 -10520 39164 -10492
rect -39164 -10788 -33792 -10760
rect -39164 -10852 -33876 -10788
rect -33812 -10852 -33792 -10788
rect -39164 -10868 -33792 -10852
rect -39164 -10932 -33876 -10868
rect -33812 -10932 -33792 -10868
rect -39164 -10948 -33792 -10932
rect -39164 -11012 -33876 -10948
rect -33812 -11012 -33792 -10948
rect -39164 -11028 -33792 -11012
rect -39164 -11092 -33876 -11028
rect -33812 -11092 -33792 -11028
rect -39164 -11108 -33792 -11092
rect -39164 -11172 -33876 -11108
rect -33812 -11172 -33792 -11108
rect -39164 -11188 -33792 -11172
rect -39164 -11252 -33876 -11188
rect -33812 -11252 -33792 -11188
rect -39164 -11268 -33792 -11252
rect -39164 -11332 -33876 -11268
rect -33812 -11332 -33792 -11268
rect -39164 -11348 -33792 -11332
rect -39164 -11412 -33876 -11348
rect -33812 -11412 -33792 -11348
rect -39164 -11428 -33792 -11412
rect -39164 -11492 -33876 -11428
rect -33812 -11492 -33792 -11428
rect -39164 -11508 -33792 -11492
rect -39164 -11572 -33876 -11508
rect -33812 -11572 -33792 -11508
rect -39164 -11588 -33792 -11572
rect -39164 -11652 -33876 -11588
rect -33812 -11652 -33792 -11588
rect -39164 -11668 -33792 -11652
rect -39164 -11732 -33876 -11668
rect -33812 -11732 -33792 -11668
rect -39164 -11748 -33792 -11732
rect -39164 -11812 -33876 -11748
rect -33812 -11812 -33792 -11748
rect -39164 -11828 -33792 -11812
rect -39164 -11892 -33876 -11828
rect -33812 -11892 -33792 -11828
rect -39164 -11908 -33792 -11892
rect -39164 -11972 -33876 -11908
rect -33812 -11972 -33792 -11908
rect -39164 -11988 -33792 -11972
rect -39164 -12052 -33876 -11988
rect -33812 -12052 -33792 -11988
rect -39164 -12068 -33792 -12052
rect -39164 -12132 -33876 -12068
rect -33812 -12132 -33792 -12068
rect -39164 -12148 -33792 -12132
rect -39164 -12212 -33876 -12148
rect -33812 -12212 -33792 -12148
rect -39164 -12228 -33792 -12212
rect -39164 -12292 -33876 -12228
rect -33812 -12292 -33792 -12228
rect -39164 -12308 -33792 -12292
rect -39164 -12372 -33876 -12308
rect -33812 -12372 -33792 -12308
rect -39164 -12388 -33792 -12372
rect -39164 -12452 -33876 -12388
rect -33812 -12452 -33792 -12388
rect -39164 -12468 -33792 -12452
rect -39164 -12532 -33876 -12468
rect -33812 -12532 -33792 -12468
rect -39164 -12548 -33792 -12532
rect -39164 -12612 -33876 -12548
rect -33812 -12612 -33792 -12548
rect -39164 -12628 -33792 -12612
rect -39164 -12692 -33876 -12628
rect -33812 -12692 -33792 -12628
rect -39164 -12708 -33792 -12692
rect -39164 -12772 -33876 -12708
rect -33812 -12772 -33792 -12708
rect -39164 -12788 -33792 -12772
rect -39164 -12852 -33876 -12788
rect -33812 -12852 -33792 -12788
rect -39164 -12868 -33792 -12852
rect -39164 -12932 -33876 -12868
rect -33812 -12932 -33792 -12868
rect -39164 -12948 -33792 -12932
rect -39164 -13012 -33876 -12948
rect -33812 -13012 -33792 -12948
rect -39164 -13028 -33792 -13012
rect -39164 -13092 -33876 -13028
rect -33812 -13092 -33792 -13028
rect -39164 -13108 -33792 -13092
rect -39164 -13172 -33876 -13108
rect -33812 -13172 -33792 -13108
rect -39164 -13188 -33792 -13172
rect -39164 -13252 -33876 -13188
rect -33812 -13252 -33792 -13188
rect -39164 -13268 -33792 -13252
rect -39164 -13332 -33876 -13268
rect -33812 -13332 -33792 -13268
rect -39164 -13348 -33792 -13332
rect -39164 -13412 -33876 -13348
rect -33812 -13412 -33792 -13348
rect -39164 -13428 -33792 -13412
rect -39164 -13492 -33876 -13428
rect -33812 -13492 -33792 -13428
rect -39164 -13508 -33792 -13492
rect -39164 -13572 -33876 -13508
rect -33812 -13572 -33792 -13508
rect -39164 -13588 -33792 -13572
rect -39164 -13652 -33876 -13588
rect -33812 -13652 -33792 -13588
rect -39164 -13668 -33792 -13652
rect -39164 -13732 -33876 -13668
rect -33812 -13732 -33792 -13668
rect -39164 -13748 -33792 -13732
rect -39164 -13812 -33876 -13748
rect -33812 -13812 -33792 -13748
rect -39164 -13828 -33792 -13812
rect -39164 -13892 -33876 -13828
rect -33812 -13892 -33792 -13828
rect -39164 -13908 -33792 -13892
rect -39164 -13972 -33876 -13908
rect -33812 -13972 -33792 -13908
rect -39164 -13988 -33792 -13972
rect -39164 -14052 -33876 -13988
rect -33812 -14052 -33792 -13988
rect -39164 -14068 -33792 -14052
rect -39164 -14132 -33876 -14068
rect -33812 -14132 -33792 -14068
rect -39164 -14148 -33792 -14132
rect -39164 -14212 -33876 -14148
rect -33812 -14212 -33792 -14148
rect -39164 -14228 -33792 -14212
rect -39164 -14292 -33876 -14228
rect -33812 -14292 -33792 -14228
rect -39164 -14308 -33792 -14292
rect -39164 -14372 -33876 -14308
rect -33812 -14372 -33792 -14308
rect -39164 -14388 -33792 -14372
rect -39164 -14452 -33876 -14388
rect -33812 -14452 -33792 -14388
rect -39164 -14468 -33792 -14452
rect -39164 -14532 -33876 -14468
rect -33812 -14532 -33792 -14468
rect -39164 -14548 -33792 -14532
rect -39164 -14612 -33876 -14548
rect -33812 -14612 -33792 -14548
rect -39164 -14628 -33792 -14612
rect -39164 -14692 -33876 -14628
rect -33812 -14692 -33792 -14628
rect -39164 -14708 -33792 -14692
rect -39164 -14772 -33876 -14708
rect -33812 -14772 -33792 -14708
rect -39164 -14788 -33792 -14772
rect -39164 -14852 -33876 -14788
rect -33812 -14852 -33792 -14788
rect -39164 -14868 -33792 -14852
rect -39164 -14932 -33876 -14868
rect -33812 -14932 -33792 -14868
rect -39164 -14948 -33792 -14932
rect -39164 -15012 -33876 -14948
rect -33812 -15012 -33792 -14948
rect -39164 -15028 -33792 -15012
rect -39164 -15092 -33876 -15028
rect -33812 -15092 -33792 -15028
rect -39164 -15108 -33792 -15092
rect -39164 -15172 -33876 -15108
rect -33812 -15172 -33792 -15108
rect -39164 -15188 -33792 -15172
rect -39164 -15252 -33876 -15188
rect -33812 -15252 -33792 -15188
rect -39164 -15268 -33792 -15252
rect -39164 -15332 -33876 -15268
rect -33812 -15332 -33792 -15268
rect -39164 -15348 -33792 -15332
rect -39164 -15412 -33876 -15348
rect -33812 -15412 -33792 -15348
rect -39164 -15428 -33792 -15412
rect -39164 -15492 -33876 -15428
rect -33812 -15492 -33792 -15428
rect -39164 -15508 -33792 -15492
rect -39164 -15572 -33876 -15508
rect -33812 -15572 -33792 -15508
rect -39164 -15588 -33792 -15572
rect -39164 -15652 -33876 -15588
rect -33812 -15652 -33792 -15588
rect -39164 -15668 -33792 -15652
rect -39164 -15732 -33876 -15668
rect -33812 -15732 -33792 -15668
rect -39164 -15748 -33792 -15732
rect -39164 -15812 -33876 -15748
rect -33812 -15812 -33792 -15748
rect -39164 -15840 -33792 -15812
rect -33552 -10788 -28180 -10760
rect -33552 -10852 -28264 -10788
rect -28200 -10852 -28180 -10788
rect -33552 -10868 -28180 -10852
rect -33552 -10932 -28264 -10868
rect -28200 -10932 -28180 -10868
rect -33552 -10948 -28180 -10932
rect -33552 -11012 -28264 -10948
rect -28200 -11012 -28180 -10948
rect -33552 -11028 -28180 -11012
rect -33552 -11092 -28264 -11028
rect -28200 -11092 -28180 -11028
rect -33552 -11108 -28180 -11092
rect -33552 -11172 -28264 -11108
rect -28200 -11172 -28180 -11108
rect -33552 -11188 -28180 -11172
rect -33552 -11252 -28264 -11188
rect -28200 -11252 -28180 -11188
rect -33552 -11268 -28180 -11252
rect -33552 -11332 -28264 -11268
rect -28200 -11332 -28180 -11268
rect -33552 -11348 -28180 -11332
rect -33552 -11412 -28264 -11348
rect -28200 -11412 -28180 -11348
rect -33552 -11428 -28180 -11412
rect -33552 -11492 -28264 -11428
rect -28200 -11492 -28180 -11428
rect -33552 -11508 -28180 -11492
rect -33552 -11572 -28264 -11508
rect -28200 -11572 -28180 -11508
rect -33552 -11588 -28180 -11572
rect -33552 -11652 -28264 -11588
rect -28200 -11652 -28180 -11588
rect -33552 -11668 -28180 -11652
rect -33552 -11732 -28264 -11668
rect -28200 -11732 -28180 -11668
rect -33552 -11748 -28180 -11732
rect -33552 -11812 -28264 -11748
rect -28200 -11812 -28180 -11748
rect -33552 -11828 -28180 -11812
rect -33552 -11892 -28264 -11828
rect -28200 -11892 -28180 -11828
rect -33552 -11908 -28180 -11892
rect -33552 -11972 -28264 -11908
rect -28200 -11972 -28180 -11908
rect -33552 -11988 -28180 -11972
rect -33552 -12052 -28264 -11988
rect -28200 -12052 -28180 -11988
rect -33552 -12068 -28180 -12052
rect -33552 -12132 -28264 -12068
rect -28200 -12132 -28180 -12068
rect -33552 -12148 -28180 -12132
rect -33552 -12212 -28264 -12148
rect -28200 -12212 -28180 -12148
rect -33552 -12228 -28180 -12212
rect -33552 -12292 -28264 -12228
rect -28200 -12292 -28180 -12228
rect -33552 -12308 -28180 -12292
rect -33552 -12372 -28264 -12308
rect -28200 -12372 -28180 -12308
rect -33552 -12388 -28180 -12372
rect -33552 -12452 -28264 -12388
rect -28200 -12452 -28180 -12388
rect -33552 -12468 -28180 -12452
rect -33552 -12532 -28264 -12468
rect -28200 -12532 -28180 -12468
rect -33552 -12548 -28180 -12532
rect -33552 -12612 -28264 -12548
rect -28200 -12612 -28180 -12548
rect -33552 -12628 -28180 -12612
rect -33552 -12692 -28264 -12628
rect -28200 -12692 -28180 -12628
rect -33552 -12708 -28180 -12692
rect -33552 -12772 -28264 -12708
rect -28200 -12772 -28180 -12708
rect -33552 -12788 -28180 -12772
rect -33552 -12852 -28264 -12788
rect -28200 -12852 -28180 -12788
rect -33552 -12868 -28180 -12852
rect -33552 -12932 -28264 -12868
rect -28200 -12932 -28180 -12868
rect -33552 -12948 -28180 -12932
rect -33552 -13012 -28264 -12948
rect -28200 -13012 -28180 -12948
rect -33552 -13028 -28180 -13012
rect -33552 -13092 -28264 -13028
rect -28200 -13092 -28180 -13028
rect -33552 -13108 -28180 -13092
rect -33552 -13172 -28264 -13108
rect -28200 -13172 -28180 -13108
rect -33552 -13188 -28180 -13172
rect -33552 -13252 -28264 -13188
rect -28200 -13252 -28180 -13188
rect -33552 -13268 -28180 -13252
rect -33552 -13332 -28264 -13268
rect -28200 -13332 -28180 -13268
rect -33552 -13348 -28180 -13332
rect -33552 -13412 -28264 -13348
rect -28200 -13412 -28180 -13348
rect -33552 -13428 -28180 -13412
rect -33552 -13492 -28264 -13428
rect -28200 -13492 -28180 -13428
rect -33552 -13508 -28180 -13492
rect -33552 -13572 -28264 -13508
rect -28200 -13572 -28180 -13508
rect -33552 -13588 -28180 -13572
rect -33552 -13652 -28264 -13588
rect -28200 -13652 -28180 -13588
rect -33552 -13668 -28180 -13652
rect -33552 -13732 -28264 -13668
rect -28200 -13732 -28180 -13668
rect -33552 -13748 -28180 -13732
rect -33552 -13812 -28264 -13748
rect -28200 -13812 -28180 -13748
rect -33552 -13828 -28180 -13812
rect -33552 -13892 -28264 -13828
rect -28200 -13892 -28180 -13828
rect -33552 -13908 -28180 -13892
rect -33552 -13972 -28264 -13908
rect -28200 -13972 -28180 -13908
rect -33552 -13988 -28180 -13972
rect -33552 -14052 -28264 -13988
rect -28200 -14052 -28180 -13988
rect -33552 -14068 -28180 -14052
rect -33552 -14132 -28264 -14068
rect -28200 -14132 -28180 -14068
rect -33552 -14148 -28180 -14132
rect -33552 -14212 -28264 -14148
rect -28200 -14212 -28180 -14148
rect -33552 -14228 -28180 -14212
rect -33552 -14292 -28264 -14228
rect -28200 -14292 -28180 -14228
rect -33552 -14308 -28180 -14292
rect -33552 -14372 -28264 -14308
rect -28200 -14372 -28180 -14308
rect -33552 -14388 -28180 -14372
rect -33552 -14452 -28264 -14388
rect -28200 -14452 -28180 -14388
rect -33552 -14468 -28180 -14452
rect -33552 -14532 -28264 -14468
rect -28200 -14532 -28180 -14468
rect -33552 -14548 -28180 -14532
rect -33552 -14612 -28264 -14548
rect -28200 -14612 -28180 -14548
rect -33552 -14628 -28180 -14612
rect -33552 -14692 -28264 -14628
rect -28200 -14692 -28180 -14628
rect -33552 -14708 -28180 -14692
rect -33552 -14772 -28264 -14708
rect -28200 -14772 -28180 -14708
rect -33552 -14788 -28180 -14772
rect -33552 -14852 -28264 -14788
rect -28200 -14852 -28180 -14788
rect -33552 -14868 -28180 -14852
rect -33552 -14932 -28264 -14868
rect -28200 -14932 -28180 -14868
rect -33552 -14948 -28180 -14932
rect -33552 -15012 -28264 -14948
rect -28200 -15012 -28180 -14948
rect -33552 -15028 -28180 -15012
rect -33552 -15092 -28264 -15028
rect -28200 -15092 -28180 -15028
rect -33552 -15108 -28180 -15092
rect -33552 -15172 -28264 -15108
rect -28200 -15172 -28180 -15108
rect -33552 -15188 -28180 -15172
rect -33552 -15252 -28264 -15188
rect -28200 -15252 -28180 -15188
rect -33552 -15268 -28180 -15252
rect -33552 -15332 -28264 -15268
rect -28200 -15332 -28180 -15268
rect -33552 -15348 -28180 -15332
rect -33552 -15412 -28264 -15348
rect -28200 -15412 -28180 -15348
rect -33552 -15428 -28180 -15412
rect -33552 -15492 -28264 -15428
rect -28200 -15492 -28180 -15428
rect -33552 -15508 -28180 -15492
rect -33552 -15572 -28264 -15508
rect -28200 -15572 -28180 -15508
rect -33552 -15588 -28180 -15572
rect -33552 -15652 -28264 -15588
rect -28200 -15652 -28180 -15588
rect -33552 -15668 -28180 -15652
rect -33552 -15732 -28264 -15668
rect -28200 -15732 -28180 -15668
rect -33552 -15748 -28180 -15732
rect -33552 -15812 -28264 -15748
rect -28200 -15812 -28180 -15748
rect -33552 -15840 -28180 -15812
rect -27940 -10788 -22568 -10760
rect -27940 -10852 -22652 -10788
rect -22588 -10852 -22568 -10788
rect -27940 -10868 -22568 -10852
rect -27940 -10932 -22652 -10868
rect -22588 -10932 -22568 -10868
rect -27940 -10948 -22568 -10932
rect -27940 -11012 -22652 -10948
rect -22588 -11012 -22568 -10948
rect -27940 -11028 -22568 -11012
rect -27940 -11092 -22652 -11028
rect -22588 -11092 -22568 -11028
rect -27940 -11108 -22568 -11092
rect -27940 -11172 -22652 -11108
rect -22588 -11172 -22568 -11108
rect -27940 -11188 -22568 -11172
rect -27940 -11252 -22652 -11188
rect -22588 -11252 -22568 -11188
rect -27940 -11268 -22568 -11252
rect -27940 -11332 -22652 -11268
rect -22588 -11332 -22568 -11268
rect -27940 -11348 -22568 -11332
rect -27940 -11412 -22652 -11348
rect -22588 -11412 -22568 -11348
rect -27940 -11428 -22568 -11412
rect -27940 -11492 -22652 -11428
rect -22588 -11492 -22568 -11428
rect -27940 -11508 -22568 -11492
rect -27940 -11572 -22652 -11508
rect -22588 -11572 -22568 -11508
rect -27940 -11588 -22568 -11572
rect -27940 -11652 -22652 -11588
rect -22588 -11652 -22568 -11588
rect -27940 -11668 -22568 -11652
rect -27940 -11732 -22652 -11668
rect -22588 -11732 -22568 -11668
rect -27940 -11748 -22568 -11732
rect -27940 -11812 -22652 -11748
rect -22588 -11812 -22568 -11748
rect -27940 -11828 -22568 -11812
rect -27940 -11892 -22652 -11828
rect -22588 -11892 -22568 -11828
rect -27940 -11908 -22568 -11892
rect -27940 -11972 -22652 -11908
rect -22588 -11972 -22568 -11908
rect -27940 -11988 -22568 -11972
rect -27940 -12052 -22652 -11988
rect -22588 -12052 -22568 -11988
rect -27940 -12068 -22568 -12052
rect -27940 -12132 -22652 -12068
rect -22588 -12132 -22568 -12068
rect -27940 -12148 -22568 -12132
rect -27940 -12212 -22652 -12148
rect -22588 -12212 -22568 -12148
rect -27940 -12228 -22568 -12212
rect -27940 -12292 -22652 -12228
rect -22588 -12292 -22568 -12228
rect -27940 -12308 -22568 -12292
rect -27940 -12372 -22652 -12308
rect -22588 -12372 -22568 -12308
rect -27940 -12388 -22568 -12372
rect -27940 -12452 -22652 -12388
rect -22588 -12452 -22568 -12388
rect -27940 -12468 -22568 -12452
rect -27940 -12532 -22652 -12468
rect -22588 -12532 -22568 -12468
rect -27940 -12548 -22568 -12532
rect -27940 -12612 -22652 -12548
rect -22588 -12612 -22568 -12548
rect -27940 -12628 -22568 -12612
rect -27940 -12692 -22652 -12628
rect -22588 -12692 -22568 -12628
rect -27940 -12708 -22568 -12692
rect -27940 -12772 -22652 -12708
rect -22588 -12772 -22568 -12708
rect -27940 -12788 -22568 -12772
rect -27940 -12852 -22652 -12788
rect -22588 -12852 -22568 -12788
rect -27940 -12868 -22568 -12852
rect -27940 -12932 -22652 -12868
rect -22588 -12932 -22568 -12868
rect -27940 -12948 -22568 -12932
rect -27940 -13012 -22652 -12948
rect -22588 -13012 -22568 -12948
rect -27940 -13028 -22568 -13012
rect -27940 -13092 -22652 -13028
rect -22588 -13092 -22568 -13028
rect -27940 -13108 -22568 -13092
rect -27940 -13172 -22652 -13108
rect -22588 -13172 -22568 -13108
rect -27940 -13188 -22568 -13172
rect -27940 -13252 -22652 -13188
rect -22588 -13252 -22568 -13188
rect -27940 -13268 -22568 -13252
rect -27940 -13332 -22652 -13268
rect -22588 -13332 -22568 -13268
rect -27940 -13348 -22568 -13332
rect -27940 -13412 -22652 -13348
rect -22588 -13412 -22568 -13348
rect -27940 -13428 -22568 -13412
rect -27940 -13492 -22652 -13428
rect -22588 -13492 -22568 -13428
rect -27940 -13508 -22568 -13492
rect -27940 -13572 -22652 -13508
rect -22588 -13572 -22568 -13508
rect -27940 -13588 -22568 -13572
rect -27940 -13652 -22652 -13588
rect -22588 -13652 -22568 -13588
rect -27940 -13668 -22568 -13652
rect -27940 -13732 -22652 -13668
rect -22588 -13732 -22568 -13668
rect -27940 -13748 -22568 -13732
rect -27940 -13812 -22652 -13748
rect -22588 -13812 -22568 -13748
rect -27940 -13828 -22568 -13812
rect -27940 -13892 -22652 -13828
rect -22588 -13892 -22568 -13828
rect -27940 -13908 -22568 -13892
rect -27940 -13972 -22652 -13908
rect -22588 -13972 -22568 -13908
rect -27940 -13988 -22568 -13972
rect -27940 -14052 -22652 -13988
rect -22588 -14052 -22568 -13988
rect -27940 -14068 -22568 -14052
rect -27940 -14132 -22652 -14068
rect -22588 -14132 -22568 -14068
rect -27940 -14148 -22568 -14132
rect -27940 -14212 -22652 -14148
rect -22588 -14212 -22568 -14148
rect -27940 -14228 -22568 -14212
rect -27940 -14292 -22652 -14228
rect -22588 -14292 -22568 -14228
rect -27940 -14308 -22568 -14292
rect -27940 -14372 -22652 -14308
rect -22588 -14372 -22568 -14308
rect -27940 -14388 -22568 -14372
rect -27940 -14452 -22652 -14388
rect -22588 -14452 -22568 -14388
rect -27940 -14468 -22568 -14452
rect -27940 -14532 -22652 -14468
rect -22588 -14532 -22568 -14468
rect -27940 -14548 -22568 -14532
rect -27940 -14612 -22652 -14548
rect -22588 -14612 -22568 -14548
rect -27940 -14628 -22568 -14612
rect -27940 -14692 -22652 -14628
rect -22588 -14692 -22568 -14628
rect -27940 -14708 -22568 -14692
rect -27940 -14772 -22652 -14708
rect -22588 -14772 -22568 -14708
rect -27940 -14788 -22568 -14772
rect -27940 -14852 -22652 -14788
rect -22588 -14852 -22568 -14788
rect -27940 -14868 -22568 -14852
rect -27940 -14932 -22652 -14868
rect -22588 -14932 -22568 -14868
rect -27940 -14948 -22568 -14932
rect -27940 -15012 -22652 -14948
rect -22588 -15012 -22568 -14948
rect -27940 -15028 -22568 -15012
rect -27940 -15092 -22652 -15028
rect -22588 -15092 -22568 -15028
rect -27940 -15108 -22568 -15092
rect -27940 -15172 -22652 -15108
rect -22588 -15172 -22568 -15108
rect -27940 -15188 -22568 -15172
rect -27940 -15252 -22652 -15188
rect -22588 -15252 -22568 -15188
rect -27940 -15268 -22568 -15252
rect -27940 -15332 -22652 -15268
rect -22588 -15332 -22568 -15268
rect -27940 -15348 -22568 -15332
rect -27940 -15412 -22652 -15348
rect -22588 -15412 -22568 -15348
rect -27940 -15428 -22568 -15412
rect -27940 -15492 -22652 -15428
rect -22588 -15492 -22568 -15428
rect -27940 -15508 -22568 -15492
rect -27940 -15572 -22652 -15508
rect -22588 -15572 -22568 -15508
rect -27940 -15588 -22568 -15572
rect -27940 -15652 -22652 -15588
rect -22588 -15652 -22568 -15588
rect -27940 -15668 -22568 -15652
rect -27940 -15732 -22652 -15668
rect -22588 -15732 -22568 -15668
rect -27940 -15748 -22568 -15732
rect -27940 -15812 -22652 -15748
rect -22588 -15812 -22568 -15748
rect -27940 -15840 -22568 -15812
rect -22328 -10788 -16956 -10760
rect -22328 -10852 -17040 -10788
rect -16976 -10852 -16956 -10788
rect -22328 -10868 -16956 -10852
rect -22328 -10932 -17040 -10868
rect -16976 -10932 -16956 -10868
rect -22328 -10948 -16956 -10932
rect -22328 -11012 -17040 -10948
rect -16976 -11012 -16956 -10948
rect -22328 -11028 -16956 -11012
rect -22328 -11092 -17040 -11028
rect -16976 -11092 -16956 -11028
rect -22328 -11108 -16956 -11092
rect -22328 -11172 -17040 -11108
rect -16976 -11172 -16956 -11108
rect -22328 -11188 -16956 -11172
rect -22328 -11252 -17040 -11188
rect -16976 -11252 -16956 -11188
rect -22328 -11268 -16956 -11252
rect -22328 -11332 -17040 -11268
rect -16976 -11332 -16956 -11268
rect -22328 -11348 -16956 -11332
rect -22328 -11412 -17040 -11348
rect -16976 -11412 -16956 -11348
rect -22328 -11428 -16956 -11412
rect -22328 -11492 -17040 -11428
rect -16976 -11492 -16956 -11428
rect -22328 -11508 -16956 -11492
rect -22328 -11572 -17040 -11508
rect -16976 -11572 -16956 -11508
rect -22328 -11588 -16956 -11572
rect -22328 -11652 -17040 -11588
rect -16976 -11652 -16956 -11588
rect -22328 -11668 -16956 -11652
rect -22328 -11732 -17040 -11668
rect -16976 -11732 -16956 -11668
rect -22328 -11748 -16956 -11732
rect -22328 -11812 -17040 -11748
rect -16976 -11812 -16956 -11748
rect -22328 -11828 -16956 -11812
rect -22328 -11892 -17040 -11828
rect -16976 -11892 -16956 -11828
rect -22328 -11908 -16956 -11892
rect -22328 -11972 -17040 -11908
rect -16976 -11972 -16956 -11908
rect -22328 -11988 -16956 -11972
rect -22328 -12052 -17040 -11988
rect -16976 -12052 -16956 -11988
rect -22328 -12068 -16956 -12052
rect -22328 -12132 -17040 -12068
rect -16976 -12132 -16956 -12068
rect -22328 -12148 -16956 -12132
rect -22328 -12212 -17040 -12148
rect -16976 -12212 -16956 -12148
rect -22328 -12228 -16956 -12212
rect -22328 -12292 -17040 -12228
rect -16976 -12292 -16956 -12228
rect -22328 -12308 -16956 -12292
rect -22328 -12372 -17040 -12308
rect -16976 -12372 -16956 -12308
rect -22328 -12388 -16956 -12372
rect -22328 -12452 -17040 -12388
rect -16976 -12452 -16956 -12388
rect -22328 -12468 -16956 -12452
rect -22328 -12532 -17040 -12468
rect -16976 -12532 -16956 -12468
rect -22328 -12548 -16956 -12532
rect -22328 -12612 -17040 -12548
rect -16976 -12612 -16956 -12548
rect -22328 -12628 -16956 -12612
rect -22328 -12692 -17040 -12628
rect -16976 -12692 -16956 -12628
rect -22328 -12708 -16956 -12692
rect -22328 -12772 -17040 -12708
rect -16976 -12772 -16956 -12708
rect -22328 -12788 -16956 -12772
rect -22328 -12852 -17040 -12788
rect -16976 -12852 -16956 -12788
rect -22328 -12868 -16956 -12852
rect -22328 -12932 -17040 -12868
rect -16976 -12932 -16956 -12868
rect -22328 -12948 -16956 -12932
rect -22328 -13012 -17040 -12948
rect -16976 -13012 -16956 -12948
rect -22328 -13028 -16956 -13012
rect -22328 -13092 -17040 -13028
rect -16976 -13092 -16956 -13028
rect -22328 -13108 -16956 -13092
rect -22328 -13172 -17040 -13108
rect -16976 -13172 -16956 -13108
rect -22328 -13188 -16956 -13172
rect -22328 -13252 -17040 -13188
rect -16976 -13252 -16956 -13188
rect -22328 -13268 -16956 -13252
rect -22328 -13332 -17040 -13268
rect -16976 -13332 -16956 -13268
rect -22328 -13348 -16956 -13332
rect -22328 -13412 -17040 -13348
rect -16976 -13412 -16956 -13348
rect -22328 -13428 -16956 -13412
rect -22328 -13492 -17040 -13428
rect -16976 -13492 -16956 -13428
rect -22328 -13508 -16956 -13492
rect -22328 -13572 -17040 -13508
rect -16976 -13572 -16956 -13508
rect -22328 -13588 -16956 -13572
rect -22328 -13652 -17040 -13588
rect -16976 -13652 -16956 -13588
rect -22328 -13668 -16956 -13652
rect -22328 -13732 -17040 -13668
rect -16976 -13732 -16956 -13668
rect -22328 -13748 -16956 -13732
rect -22328 -13812 -17040 -13748
rect -16976 -13812 -16956 -13748
rect -22328 -13828 -16956 -13812
rect -22328 -13892 -17040 -13828
rect -16976 -13892 -16956 -13828
rect -22328 -13908 -16956 -13892
rect -22328 -13972 -17040 -13908
rect -16976 -13972 -16956 -13908
rect -22328 -13988 -16956 -13972
rect -22328 -14052 -17040 -13988
rect -16976 -14052 -16956 -13988
rect -22328 -14068 -16956 -14052
rect -22328 -14132 -17040 -14068
rect -16976 -14132 -16956 -14068
rect -22328 -14148 -16956 -14132
rect -22328 -14212 -17040 -14148
rect -16976 -14212 -16956 -14148
rect -22328 -14228 -16956 -14212
rect -22328 -14292 -17040 -14228
rect -16976 -14292 -16956 -14228
rect -22328 -14308 -16956 -14292
rect -22328 -14372 -17040 -14308
rect -16976 -14372 -16956 -14308
rect -22328 -14388 -16956 -14372
rect -22328 -14452 -17040 -14388
rect -16976 -14452 -16956 -14388
rect -22328 -14468 -16956 -14452
rect -22328 -14532 -17040 -14468
rect -16976 -14532 -16956 -14468
rect -22328 -14548 -16956 -14532
rect -22328 -14612 -17040 -14548
rect -16976 -14612 -16956 -14548
rect -22328 -14628 -16956 -14612
rect -22328 -14692 -17040 -14628
rect -16976 -14692 -16956 -14628
rect -22328 -14708 -16956 -14692
rect -22328 -14772 -17040 -14708
rect -16976 -14772 -16956 -14708
rect -22328 -14788 -16956 -14772
rect -22328 -14852 -17040 -14788
rect -16976 -14852 -16956 -14788
rect -22328 -14868 -16956 -14852
rect -22328 -14932 -17040 -14868
rect -16976 -14932 -16956 -14868
rect -22328 -14948 -16956 -14932
rect -22328 -15012 -17040 -14948
rect -16976 -15012 -16956 -14948
rect -22328 -15028 -16956 -15012
rect -22328 -15092 -17040 -15028
rect -16976 -15092 -16956 -15028
rect -22328 -15108 -16956 -15092
rect -22328 -15172 -17040 -15108
rect -16976 -15172 -16956 -15108
rect -22328 -15188 -16956 -15172
rect -22328 -15252 -17040 -15188
rect -16976 -15252 -16956 -15188
rect -22328 -15268 -16956 -15252
rect -22328 -15332 -17040 -15268
rect -16976 -15332 -16956 -15268
rect -22328 -15348 -16956 -15332
rect -22328 -15412 -17040 -15348
rect -16976 -15412 -16956 -15348
rect -22328 -15428 -16956 -15412
rect -22328 -15492 -17040 -15428
rect -16976 -15492 -16956 -15428
rect -22328 -15508 -16956 -15492
rect -22328 -15572 -17040 -15508
rect -16976 -15572 -16956 -15508
rect -22328 -15588 -16956 -15572
rect -22328 -15652 -17040 -15588
rect -16976 -15652 -16956 -15588
rect -22328 -15668 -16956 -15652
rect -22328 -15732 -17040 -15668
rect -16976 -15732 -16956 -15668
rect -22328 -15748 -16956 -15732
rect -22328 -15812 -17040 -15748
rect -16976 -15812 -16956 -15748
rect -22328 -15840 -16956 -15812
rect -16716 -10788 -11344 -10760
rect -16716 -10852 -11428 -10788
rect -11364 -10852 -11344 -10788
rect -16716 -10868 -11344 -10852
rect -16716 -10932 -11428 -10868
rect -11364 -10932 -11344 -10868
rect -16716 -10948 -11344 -10932
rect -16716 -11012 -11428 -10948
rect -11364 -11012 -11344 -10948
rect -16716 -11028 -11344 -11012
rect -16716 -11092 -11428 -11028
rect -11364 -11092 -11344 -11028
rect -16716 -11108 -11344 -11092
rect -16716 -11172 -11428 -11108
rect -11364 -11172 -11344 -11108
rect -16716 -11188 -11344 -11172
rect -16716 -11252 -11428 -11188
rect -11364 -11252 -11344 -11188
rect -16716 -11268 -11344 -11252
rect -16716 -11332 -11428 -11268
rect -11364 -11332 -11344 -11268
rect -16716 -11348 -11344 -11332
rect -16716 -11412 -11428 -11348
rect -11364 -11412 -11344 -11348
rect -16716 -11428 -11344 -11412
rect -16716 -11492 -11428 -11428
rect -11364 -11492 -11344 -11428
rect -16716 -11508 -11344 -11492
rect -16716 -11572 -11428 -11508
rect -11364 -11572 -11344 -11508
rect -16716 -11588 -11344 -11572
rect -16716 -11652 -11428 -11588
rect -11364 -11652 -11344 -11588
rect -16716 -11668 -11344 -11652
rect -16716 -11732 -11428 -11668
rect -11364 -11732 -11344 -11668
rect -16716 -11748 -11344 -11732
rect -16716 -11812 -11428 -11748
rect -11364 -11812 -11344 -11748
rect -16716 -11828 -11344 -11812
rect -16716 -11892 -11428 -11828
rect -11364 -11892 -11344 -11828
rect -16716 -11908 -11344 -11892
rect -16716 -11972 -11428 -11908
rect -11364 -11972 -11344 -11908
rect -16716 -11988 -11344 -11972
rect -16716 -12052 -11428 -11988
rect -11364 -12052 -11344 -11988
rect -16716 -12068 -11344 -12052
rect -16716 -12132 -11428 -12068
rect -11364 -12132 -11344 -12068
rect -16716 -12148 -11344 -12132
rect -16716 -12212 -11428 -12148
rect -11364 -12212 -11344 -12148
rect -16716 -12228 -11344 -12212
rect -16716 -12292 -11428 -12228
rect -11364 -12292 -11344 -12228
rect -16716 -12308 -11344 -12292
rect -16716 -12372 -11428 -12308
rect -11364 -12372 -11344 -12308
rect -16716 -12388 -11344 -12372
rect -16716 -12452 -11428 -12388
rect -11364 -12452 -11344 -12388
rect -16716 -12468 -11344 -12452
rect -16716 -12532 -11428 -12468
rect -11364 -12532 -11344 -12468
rect -16716 -12548 -11344 -12532
rect -16716 -12612 -11428 -12548
rect -11364 -12612 -11344 -12548
rect -16716 -12628 -11344 -12612
rect -16716 -12692 -11428 -12628
rect -11364 -12692 -11344 -12628
rect -16716 -12708 -11344 -12692
rect -16716 -12772 -11428 -12708
rect -11364 -12772 -11344 -12708
rect -16716 -12788 -11344 -12772
rect -16716 -12852 -11428 -12788
rect -11364 -12852 -11344 -12788
rect -16716 -12868 -11344 -12852
rect -16716 -12932 -11428 -12868
rect -11364 -12932 -11344 -12868
rect -16716 -12948 -11344 -12932
rect -16716 -13012 -11428 -12948
rect -11364 -13012 -11344 -12948
rect -16716 -13028 -11344 -13012
rect -16716 -13092 -11428 -13028
rect -11364 -13092 -11344 -13028
rect -16716 -13108 -11344 -13092
rect -16716 -13172 -11428 -13108
rect -11364 -13172 -11344 -13108
rect -16716 -13188 -11344 -13172
rect -16716 -13252 -11428 -13188
rect -11364 -13252 -11344 -13188
rect -16716 -13268 -11344 -13252
rect -16716 -13332 -11428 -13268
rect -11364 -13332 -11344 -13268
rect -16716 -13348 -11344 -13332
rect -16716 -13412 -11428 -13348
rect -11364 -13412 -11344 -13348
rect -16716 -13428 -11344 -13412
rect -16716 -13492 -11428 -13428
rect -11364 -13492 -11344 -13428
rect -16716 -13508 -11344 -13492
rect -16716 -13572 -11428 -13508
rect -11364 -13572 -11344 -13508
rect -16716 -13588 -11344 -13572
rect -16716 -13652 -11428 -13588
rect -11364 -13652 -11344 -13588
rect -16716 -13668 -11344 -13652
rect -16716 -13732 -11428 -13668
rect -11364 -13732 -11344 -13668
rect -16716 -13748 -11344 -13732
rect -16716 -13812 -11428 -13748
rect -11364 -13812 -11344 -13748
rect -16716 -13828 -11344 -13812
rect -16716 -13892 -11428 -13828
rect -11364 -13892 -11344 -13828
rect -16716 -13908 -11344 -13892
rect -16716 -13972 -11428 -13908
rect -11364 -13972 -11344 -13908
rect -16716 -13988 -11344 -13972
rect -16716 -14052 -11428 -13988
rect -11364 -14052 -11344 -13988
rect -16716 -14068 -11344 -14052
rect -16716 -14132 -11428 -14068
rect -11364 -14132 -11344 -14068
rect -16716 -14148 -11344 -14132
rect -16716 -14212 -11428 -14148
rect -11364 -14212 -11344 -14148
rect -16716 -14228 -11344 -14212
rect -16716 -14292 -11428 -14228
rect -11364 -14292 -11344 -14228
rect -16716 -14308 -11344 -14292
rect -16716 -14372 -11428 -14308
rect -11364 -14372 -11344 -14308
rect -16716 -14388 -11344 -14372
rect -16716 -14452 -11428 -14388
rect -11364 -14452 -11344 -14388
rect -16716 -14468 -11344 -14452
rect -16716 -14532 -11428 -14468
rect -11364 -14532 -11344 -14468
rect -16716 -14548 -11344 -14532
rect -16716 -14612 -11428 -14548
rect -11364 -14612 -11344 -14548
rect -16716 -14628 -11344 -14612
rect -16716 -14692 -11428 -14628
rect -11364 -14692 -11344 -14628
rect -16716 -14708 -11344 -14692
rect -16716 -14772 -11428 -14708
rect -11364 -14772 -11344 -14708
rect -16716 -14788 -11344 -14772
rect -16716 -14852 -11428 -14788
rect -11364 -14852 -11344 -14788
rect -16716 -14868 -11344 -14852
rect -16716 -14932 -11428 -14868
rect -11364 -14932 -11344 -14868
rect -16716 -14948 -11344 -14932
rect -16716 -15012 -11428 -14948
rect -11364 -15012 -11344 -14948
rect -16716 -15028 -11344 -15012
rect -16716 -15092 -11428 -15028
rect -11364 -15092 -11344 -15028
rect -16716 -15108 -11344 -15092
rect -16716 -15172 -11428 -15108
rect -11364 -15172 -11344 -15108
rect -16716 -15188 -11344 -15172
rect -16716 -15252 -11428 -15188
rect -11364 -15252 -11344 -15188
rect -16716 -15268 -11344 -15252
rect -16716 -15332 -11428 -15268
rect -11364 -15332 -11344 -15268
rect -16716 -15348 -11344 -15332
rect -16716 -15412 -11428 -15348
rect -11364 -15412 -11344 -15348
rect -16716 -15428 -11344 -15412
rect -16716 -15492 -11428 -15428
rect -11364 -15492 -11344 -15428
rect -16716 -15508 -11344 -15492
rect -16716 -15572 -11428 -15508
rect -11364 -15572 -11344 -15508
rect -16716 -15588 -11344 -15572
rect -16716 -15652 -11428 -15588
rect -11364 -15652 -11344 -15588
rect -16716 -15668 -11344 -15652
rect -16716 -15732 -11428 -15668
rect -11364 -15732 -11344 -15668
rect -16716 -15748 -11344 -15732
rect -16716 -15812 -11428 -15748
rect -11364 -15812 -11344 -15748
rect -16716 -15840 -11344 -15812
rect -11104 -10788 -5732 -10760
rect -11104 -10852 -5816 -10788
rect -5752 -10852 -5732 -10788
rect -11104 -10868 -5732 -10852
rect -11104 -10932 -5816 -10868
rect -5752 -10932 -5732 -10868
rect -11104 -10948 -5732 -10932
rect -11104 -11012 -5816 -10948
rect -5752 -11012 -5732 -10948
rect -11104 -11028 -5732 -11012
rect -11104 -11092 -5816 -11028
rect -5752 -11092 -5732 -11028
rect -11104 -11108 -5732 -11092
rect -11104 -11172 -5816 -11108
rect -5752 -11172 -5732 -11108
rect -11104 -11188 -5732 -11172
rect -11104 -11252 -5816 -11188
rect -5752 -11252 -5732 -11188
rect -11104 -11268 -5732 -11252
rect -11104 -11332 -5816 -11268
rect -5752 -11332 -5732 -11268
rect -11104 -11348 -5732 -11332
rect -11104 -11412 -5816 -11348
rect -5752 -11412 -5732 -11348
rect -11104 -11428 -5732 -11412
rect -11104 -11492 -5816 -11428
rect -5752 -11492 -5732 -11428
rect -11104 -11508 -5732 -11492
rect -11104 -11572 -5816 -11508
rect -5752 -11572 -5732 -11508
rect -11104 -11588 -5732 -11572
rect -11104 -11652 -5816 -11588
rect -5752 -11652 -5732 -11588
rect -11104 -11668 -5732 -11652
rect -11104 -11732 -5816 -11668
rect -5752 -11732 -5732 -11668
rect -11104 -11748 -5732 -11732
rect -11104 -11812 -5816 -11748
rect -5752 -11812 -5732 -11748
rect -11104 -11828 -5732 -11812
rect -11104 -11892 -5816 -11828
rect -5752 -11892 -5732 -11828
rect -11104 -11908 -5732 -11892
rect -11104 -11972 -5816 -11908
rect -5752 -11972 -5732 -11908
rect -11104 -11988 -5732 -11972
rect -11104 -12052 -5816 -11988
rect -5752 -12052 -5732 -11988
rect -11104 -12068 -5732 -12052
rect -11104 -12132 -5816 -12068
rect -5752 -12132 -5732 -12068
rect -11104 -12148 -5732 -12132
rect -11104 -12212 -5816 -12148
rect -5752 -12212 -5732 -12148
rect -11104 -12228 -5732 -12212
rect -11104 -12292 -5816 -12228
rect -5752 -12292 -5732 -12228
rect -11104 -12308 -5732 -12292
rect -11104 -12372 -5816 -12308
rect -5752 -12372 -5732 -12308
rect -11104 -12388 -5732 -12372
rect -11104 -12452 -5816 -12388
rect -5752 -12452 -5732 -12388
rect -11104 -12468 -5732 -12452
rect -11104 -12532 -5816 -12468
rect -5752 -12532 -5732 -12468
rect -11104 -12548 -5732 -12532
rect -11104 -12612 -5816 -12548
rect -5752 -12612 -5732 -12548
rect -11104 -12628 -5732 -12612
rect -11104 -12692 -5816 -12628
rect -5752 -12692 -5732 -12628
rect -11104 -12708 -5732 -12692
rect -11104 -12772 -5816 -12708
rect -5752 -12772 -5732 -12708
rect -11104 -12788 -5732 -12772
rect -11104 -12852 -5816 -12788
rect -5752 -12852 -5732 -12788
rect -11104 -12868 -5732 -12852
rect -11104 -12932 -5816 -12868
rect -5752 -12932 -5732 -12868
rect -11104 -12948 -5732 -12932
rect -11104 -13012 -5816 -12948
rect -5752 -13012 -5732 -12948
rect -11104 -13028 -5732 -13012
rect -11104 -13092 -5816 -13028
rect -5752 -13092 -5732 -13028
rect -11104 -13108 -5732 -13092
rect -11104 -13172 -5816 -13108
rect -5752 -13172 -5732 -13108
rect -11104 -13188 -5732 -13172
rect -11104 -13252 -5816 -13188
rect -5752 -13252 -5732 -13188
rect -11104 -13268 -5732 -13252
rect -11104 -13332 -5816 -13268
rect -5752 -13332 -5732 -13268
rect -11104 -13348 -5732 -13332
rect -11104 -13412 -5816 -13348
rect -5752 -13412 -5732 -13348
rect -11104 -13428 -5732 -13412
rect -11104 -13492 -5816 -13428
rect -5752 -13492 -5732 -13428
rect -11104 -13508 -5732 -13492
rect -11104 -13572 -5816 -13508
rect -5752 -13572 -5732 -13508
rect -11104 -13588 -5732 -13572
rect -11104 -13652 -5816 -13588
rect -5752 -13652 -5732 -13588
rect -11104 -13668 -5732 -13652
rect -11104 -13732 -5816 -13668
rect -5752 -13732 -5732 -13668
rect -11104 -13748 -5732 -13732
rect -11104 -13812 -5816 -13748
rect -5752 -13812 -5732 -13748
rect -11104 -13828 -5732 -13812
rect -11104 -13892 -5816 -13828
rect -5752 -13892 -5732 -13828
rect -11104 -13908 -5732 -13892
rect -11104 -13972 -5816 -13908
rect -5752 -13972 -5732 -13908
rect -11104 -13988 -5732 -13972
rect -11104 -14052 -5816 -13988
rect -5752 -14052 -5732 -13988
rect -11104 -14068 -5732 -14052
rect -11104 -14132 -5816 -14068
rect -5752 -14132 -5732 -14068
rect -11104 -14148 -5732 -14132
rect -11104 -14212 -5816 -14148
rect -5752 -14212 -5732 -14148
rect -11104 -14228 -5732 -14212
rect -11104 -14292 -5816 -14228
rect -5752 -14292 -5732 -14228
rect -11104 -14308 -5732 -14292
rect -11104 -14372 -5816 -14308
rect -5752 -14372 -5732 -14308
rect -11104 -14388 -5732 -14372
rect -11104 -14452 -5816 -14388
rect -5752 -14452 -5732 -14388
rect -11104 -14468 -5732 -14452
rect -11104 -14532 -5816 -14468
rect -5752 -14532 -5732 -14468
rect -11104 -14548 -5732 -14532
rect -11104 -14612 -5816 -14548
rect -5752 -14612 -5732 -14548
rect -11104 -14628 -5732 -14612
rect -11104 -14692 -5816 -14628
rect -5752 -14692 -5732 -14628
rect -11104 -14708 -5732 -14692
rect -11104 -14772 -5816 -14708
rect -5752 -14772 -5732 -14708
rect -11104 -14788 -5732 -14772
rect -11104 -14852 -5816 -14788
rect -5752 -14852 -5732 -14788
rect -11104 -14868 -5732 -14852
rect -11104 -14932 -5816 -14868
rect -5752 -14932 -5732 -14868
rect -11104 -14948 -5732 -14932
rect -11104 -15012 -5816 -14948
rect -5752 -15012 -5732 -14948
rect -11104 -15028 -5732 -15012
rect -11104 -15092 -5816 -15028
rect -5752 -15092 -5732 -15028
rect -11104 -15108 -5732 -15092
rect -11104 -15172 -5816 -15108
rect -5752 -15172 -5732 -15108
rect -11104 -15188 -5732 -15172
rect -11104 -15252 -5816 -15188
rect -5752 -15252 -5732 -15188
rect -11104 -15268 -5732 -15252
rect -11104 -15332 -5816 -15268
rect -5752 -15332 -5732 -15268
rect -11104 -15348 -5732 -15332
rect -11104 -15412 -5816 -15348
rect -5752 -15412 -5732 -15348
rect -11104 -15428 -5732 -15412
rect -11104 -15492 -5816 -15428
rect -5752 -15492 -5732 -15428
rect -11104 -15508 -5732 -15492
rect -11104 -15572 -5816 -15508
rect -5752 -15572 -5732 -15508
rect -11104 -15588 -5732 -15572
rect -11104 -15652 -5816 -15588
rect -5752 -15652 -5732 -15588
rect -11104 -15668 -5732 -15652
rect -11104 -15732 -5816 -15668
rect -5752 -15732 -5732 -15668
rect -11104 -15748 -5732 -15732
rect -11104 -15812 -5816 -15748
rect -5752 -15812 -5732 -15748
rect -11104 -15840 -5732 -15812
rect -5492 -10788 -120 -10760
rect -5492 -10852 -204 -10788
rect -140 -10852 -120 -10788
rect -5492 -10868 -120 -10852
rect -5492 -10932 -204 -10868
rect -140 -10932 -120 -10868
rect -5492 -10948 -120 -10932
rect -5492 -11012 -204 -10948
rect -140 -11012 -120 -10948
rect -5492 -11028 -120 -11012
rect -5492 -11092 -204 -11028
rect -140 -11092 -120 -11028
rect -5492 -11108 -120 -11092
rect -5492 -11172 -204 -11108
rect -140 -11172 -120 -11108
rect -5492 -11188 -120 -11172
rect -5492 -11252 -204 -11188
rect -140 -11252 -120 -11188
rect -5492 -11268 -120 -11252
rect -5492 -11332 -204 -11268
rect -140 -11332 -120 -11268
rect -5492 -11348 -120 -11332
rect -5492 -11412 -204 -11348
rect -140 -11412 -120 -11348
rect -5492 -11428 -120 -11412
rect -5492 -11492 -204 -11428
rect -140 -11492 -120 -11428
rect -5492 -11508 -120 -11492
rect -5492 -11572 -204 -11508
rect -140 -11572 -120 -11508
rect -5492 -11588 -120 -11572
rect -5492 -11652 -204 -11588
rect -140 -11652 -120 -11588
rect -5492 -11668 -120 -11652
rect -5492 -11732 -204 -11668
rect -140 -11732 -120 -11668
rect -5492 -11748 -120 -11732
rect -5492 -11812 -204 -11748
rect -140 -11812 -120 -11748
rect -5492 -11828 -120 -11812
rect -5492 -11892 -204 -11828
rect -140 -11892 -120 -11828
rect -5492 -11908 -120 -11892
rect -5492 -11972 -204 -11908
rect -140 -11972 -120 -11908
rect -5492 -11988 -120 -11972
rect -5492 -12052 -204 -11988
rect -140 -12052 -120 -11988
rect -5492 -12068 -120 -12052
rect -5492 -12132 -204 -12068
rect -140 -12132 -120 -12068
rect -5492 -12148 -120 -12132
rect -5492 -12212 -204 -12148
rect -140 -12212 -120 -12148
rect -5492 -12228 -120 -12212
rect -5492 -12292 -204 -12228
rect -140 -12292 -120 -12228
rect -5492 -12308 -120 -12292
rect -5492 -12372 -204 -12308
rect -140 -12372 -120 -12308
rect -5492 -12388 -120 -12372
rect -5492 -12452 -204 -12388
rect -140 -12452 -120 -12388
rect -5492 -12468 -120 -12452
rect -5492 -12532 -204 -12468
rect -140 -12532 -120 -12468
rect -5492 -12548 -120 -12532
rect -5492 -12612 -204 -12548
rect -140 -12612 -120 -12548
rect -5492 -12628 -120 -12612
rect -5492 -12692 -204 -12628
rect -140 -12692 -120 -12628
rect -5492 -12708 -120 -12692
rect -5492 -12772 -204 -12708
rect -140 -12772 -120 -12708
rect -5492 -12788 -120 -12772
rect -5492 -12852 -204 -12788
rect -140 -12852 -120 -12788
rect -5492 -12868 -120 -12852
rect -5492 -12932 -204 -12868
rect -140 -12932 -120 -12868
rect -5492 -12948 -120 -12932
rect -5492 -13012 -204 -12948
rect -140 -13012 -120 -12948
rect -5492 -13028 -120 -13012
rect -5492 -13092 -204 -13028
rect -140 -13092 -120 -13028
rect -5492 -13108 -120 -13092
rect -5492 -13172 -204 -13108
rect -140 -13172 -120 -13108
rect -5492 -13188 -120 -13172
rect -5492 -13252 -204 -13188
rect -140 -13252 -120 -13188
rect -5492 -13268 -120 -13252
rect -5492 -13332 -204 -13268
rect -140 -13332 -120 -13268
rect -5492 -13348 -120 -13332
rect -5492 -13412 -204 -13348
rect -140 -13412 -120 -13348
rect -5492 -13428 -120 -13412
rect -5492 -13492 -204 -13428
rect -140 -13492 -120 -13428
rect -5492 -13508 -120 -13492
rect -5492 -13572 -204 -13508
rect -140 -13572 -120 -13508
rect -5492 -13588 -120 -13572
rect -5492 -13652 -204 -13588
rect -140 -13652 -120 -13588
rect -5492 -13668 -120 -13652
rect -5492 -13732 -204 -13668
rect -140 -13732 -120 -13668
rect -5492 -13748 -120 -13732
rect -5492 -13812 -204 -13748
rect -140 -13812 -120 -13748
rect -5492 -13828 -120 -13812
rect -5492 -13892 -204 -13828
rect -140 -13892 -120 -13828
rect -5492 -13908 -120 -13892
rect -5492 -13972 -204 -13908
rect -140 -13972 -120 -13908
rect -5492 -13988 -120 -13972
rect -5492 -14052 -204 -13988
rect -140 -14052 -120 -13988
rect -5492 -14068 -120 -14052
rect -5492 -14132 -204 -14068
rect -140 -14132 -120 -14068
rect -5492 -14148 -120 -14132
rect -5492 -14212 -204 -14148
rect -140 -14212 -120 -14148
rect -5492 -14228 -120 -14212
rect -5492 -14292 -204 -14228
rect -140 -14292 -120 -14228
rect -5492 -14308 -120 -14292
rect -5492 -14372 -204 -14308
rect -140 -14372 -120 -14308
rect -5492 -14388 -120 -14372
rect -5492 -14452 -204 -14388
rect -140 -14452 -120 -14388
rect -5492 -14468 -120 -14452
rect -5492 -14532 -204 -14468
rect -140 -14532 -120 -14468
rect -5492 -14548 -120 -14532
rect -5492 -14612 -204 -14548
rect -140 -14612 -120 -14548
rect -5492 -14628 -120 -14612
rect -5492 -14692 -204 -14628
rect -140 -14692 -120 -14628
rect -5492 -14708 -120 -14692
rect -5492 -14772 -204 -14708
rect -140 -14772 -120 -14708
rect -5492 -14788 -120 -14772
rect -5492 -14852 -204 -14788
rect -140 -14852 -120 -14788
rect -5492 -14868 -120 -14852
rect -5492 -14932 -204 -14868
rect -140 -14932 -120 -14868
rect -5492 -14948 -120 -14932
rect -5492 -15012 -204 -14948
rect -140 -15012 -120 -14948
rect -5492 -15028 -120 -15012
rect -5492 -15092 -204 -15028
rect -140 -15092 -120 -15028
rect -5492 -15108 -120 -15092
rect -5492 -15172 -204 -15108
rect -140 -15172 -120 -15108
rect -5492 -15188 -120 -15172
rect -5492 -15252 -204 -15188
rect -140 -15252 -120 -15188
rect -5492 -15268 -120 -15252
rect -5492 -15332 -204 -15268
rect -140 -15332 -120 -15268
rect -5492 -15348 -120 -15332
rect -5492 -15412 -204 -15348
rect -140 -15412 -120 -15348
rect -5492 -15428 -120 -15412
rect -5492 -15492 -204 -15428
rect -140 -15492 -120 -15428
rect -5492 -15508 -120 -15492
rect -5492 -15572 -204 -15508
rect -140 -15572 -120 -15508
rect -5492 -15588 -120 -15572
rect -5492 -15652 -204 -15588
rect -140 -15652 -120 -15588
rect -5492 -15668 -120 -15652
rect -5492 -15732 -204 -15668
rect -140 -15732 -120 -15668
rect -5492 -15748 -120 -15732
rect -5492 -15812 -204 -15748
rect -140 -15812 -120 -15748
rect -5492 -15840 -120 -15812
rect 120 -10788 5492 -10760
rect 120 -10852 5408 -10788
rect 5472 -10852 5492 -10788
rect 120 -10868 5492 -10852
rect 120 -10932 5408 -10868
rect 5472 -10932 5492 -10868
rect 120 -10948 5492 -10932
rect 120 -11012 5408 -10948
rect 5472 -11012 5492 -10948
rect 120 -11028 5492 -11012
rect 120 -11092 5408 -11028
rect 5472 -11092 5492 -11028
rect 120 -11108 5492 -11092
rect 120 -11172 5408 -11108
rect 5472 -11172 5492 -11108
rect 120 -11188 5492 -11172
rect 120 -11252 5408 -11188
rect 5472 -11252 5492 -11188
rect 120 -11268 5492 -11252
rect 120 -11332 5408 -11268
rect 5472 -11332 5492 -11268
rect 120 -11348 5492 -11332
rect 120 -11412 5408 -11348
rect 5472 -11412 5492 -11348
rect 120 -11428 5492 -11412
rect 120 -11492 5408 -11428
rect 5472 -11492 5492 -11428
rect 120 -11508 5492 -11492
rect 120 -11572 5408 -11508
rect 5472 -11572 5492 -11508
rect 120 -11588 5492 -11572
rect 120 -11652 5408 -11588
rect 5472 -11652 5492 -11588
rect 120 -11668 5492 -11652
rect 120 -11732 5408 -11668
rect 5472 -11732 5492 -11668
rect 120 -11748 5492 -11732
rect 120 -11812 5408 -11748
rect 5472 -11812 5492 -11748
rect 120 -11828 5492 -11812
rect 120 -11892 5408 -11828
rect 5472 -11892 5492 -11828
rect 120 -11908 5492 -11892
rect 120 -11972 5408 -11908
rect 5472 -11972 5492 -11908
rect 120 -11988 5492 -11972
rect 120 -12052 5408 -11988
rect 5472 -12052 5492 -11988
rect 120 -12068 5492 -12052
rect 120 -12132 5408 -12068
rect 5472 -12132 5492 -12068
rect 120 -12148 5492 -12132
rect 120 -12212 5408 -12148
rect 5472 -12212 5492 -12148
rect 120 -12228 5492 -12212
rect 120 -12292 5408 -12228
rect 5472 -12292 5492 -12228
rect 120 -12308 5492 -12292
rect 120 -12372 5408 -12308
rect 5472 -12372 5492 -12308
rect 120 -12388 5492 -12372
rect 120 -12452 5408 -12388
rect 5472 -12452 5492 -12388
rect 120 -12468 5492 -12452
rect 120 -12532 5408 -12468
rect 5472 -12532 5492 -12468
rect 120 -12548 5492 -12532
rect 120 -12612 5408 -12548
rect 5472 -12612 5492 -12548
rect 120 -12628 5492 -12612
rect 120 -12692 5408 -12628
rect 5472 -12692 5492 -12628
rect 120 -12708 5492 -12692
rect 120 -12772 5408 -12708
rect 5472 -12772 5492 -12708
rect 120 -12788 5492 -12772
rect 120 -12852 5408 -12788
rect 5472 -12852 5492 -12788
rect 120 -12868 5492 -12852
rect 120 -12932 5408 -12868
rect 5472 -12932 5492 -12868
rect 120 -12948 5492 -12932
rect 120 -13012 5408 -12948
rect 5472 -13012 5492 -12948
rect 120 -13028 5492 -13012
rect 120 -13092 5408 -13028
rect 5472 -13092 5492 -13028
rect 120 -13108 5492 -13092
rect 120 -13172 5408 -13108
rect 5472 -13172 5492 -13108
rect 120 -13188 5492 -13172
rect 120 -13252 5408 -13188
rect 5472 -13252 5492 -13188
rect 120 -13268 5492 -13252
rect 120 -13332 5408 -13268
rect 5472 -13332 5492 -13268
rect 120 -13348 5492 -13332
rect 120 -13412 5408 -13348
rect 5472 -13412 5492 -13348
rect 120 -13428 5492 -13412
rect 120 -13492 5408 -13428
rect 5472 -13492 5492 -13428
rect 120 -13508 5492 -13492
rect 120 -13572 5408 -13508
rect 5472 -13572 5492 -13508
rect 120 -13588 5492 -13572
rect 120 -13652 5408 -13588
rect 5472 -13652 5492 -13588
rect 120 -13668 5492 -13652
rect 120 -13732 5408 -13668
rect 5472 -13732 5492 -13668
rect 120 -13748 5492 -13732
rect 120 -13812 5408 -13748
rect 5472 -13812 5492 -13748
rect 120 -13828 5492 -13812
rect 120 -13892 5408 -13828
rect 5472 -13892 5492 -13828
rect 120 -13908 5492 -13892
rect 120 -13972 5408 -13908
rect 5472 -13972 5492 -13908
rect 120 -13988 5492 -13972
rect 120 -14052 5408 -13988
rect 5472 -14052 5492 -13988
rect 120 -14068 5492 -14052
rect 120 -14132 5408 -14068
rect 5472 -14132 5492 -14068
rect 120 -14148 5492 -14132
rect 120 -14212 5408 -14148
rect 5472 -14212 5492 -14148
rect 120 -14228 5492 -14212
rect 120 -14292 5408 -14228
rect 5472 -14292 5492 -14228
rect 120 -14308 5492 -14292
rect 120 -14372 5408 -14308
rect 5472 -14372 5492 -14308
rect 120 -14388 5492 -14372
rect 120 -14452 5408 -14388
rect 5472 -14452 5492 -14388
rect 120 -14468 5492 -14452
rect 120 -14532 5408 -14468
rect 5472 -14532 5492 -14468
rect 120 -14548 5492 -14532
rect 120 -14612 5408 -14548
rect 5472 -14612 5492 -14548
rect 120 -14628 5492 -14612
rect 120 -14692 5408 -14628
rect 5472 -14692 5492 -14628
rect 120 -14708 5492 -14692
rect 120 -14772 5408 -14708
rect 5472 -14772 5492 -14708
rect 120 -14788 5492 -14772
rect 120 -14852 5408 -14788
rect 5472 -14852 5492 -14788
rect 120 -14868 5492 -14852
rect 120 -14932 5408 -14868
rect 5472 -14932 5492 -14868
rect 120 -14948 5492 -14932
rect 120 -15012 5408 -14948
rect 5472 -15012 5492 -14948
rect 120 -15028 5492 -15012
rect 120 -15092 5408 -15028
rect 5472 -15092 5492 -15028
rect 120 -15108 5492 -15092
rect 120 -15172 5408 -15108
rect 5472 -15172 5492 -15108
rect 120 -15188 5492 -15172
rect 120 -15252 5408 -15188
rect 5472 -15252 5492 -15188
rect 120 -15268 5492 -15252
rect 120 -15332 5408 -15268
rect 5472 -15332 5492 -15268
rect 120 -15348 5492 -15332
rect 120 -15412 5408 -15348
rect 5472 -15412 5492 -15348
rect 120 -15428 5492 -15412
rect 120 -15492 5408 -15428
rect 5472 -15492 5492 -15428
rect 120 -15508 5492 -15492
rect 120 -15572 5408 -15508
rect 5472 -15572 5492 -15508
rect 120 -15588 5492 -15572
rect 120 -15652 5408 -15588
rect 5472 -15652 5492 -15588
rect 120 -15668 5492 -15652
rect 120 -15732 5408 -15668
rect 5472 -15732 5492 -15668
rect 120 -15748 5492 -15732
rect 120 -15812 5408 -15748
rect 5472 -15812 5492 -15748
rect 120 -15840 5492 -15812
rect 5732 -10788 11104 -10760
rect 5732 -10852 11020 -10788
rect 11084 -10852 11104 -10788
rect 5732 -10868 11104 -10852
rect 5732 -10932 11020 -10868
rect 11084 -10932 11104 -10868
rect 5732 -10948 11104 -10932
rect 5732 -11012 11020 -10948
rect 11084 -11012 11104 -10948
rect 5732 -11028 11104 -11012
rect 5732 -11092 11020 -11028
rect 11084 -11092 11104 -11028
rect 5732 -11108 11104 -11092
rect 5732 -11172 11020 -11108
rect 11084 -11172 11104 -11108
rect 5732 -11188 11104 -11172
rect 5732 -11252 11020 -11188
rect 11084 -11252 11104 -11188
rect 5732 -11268 11104 -11252
rect 5732 -11332 11020 -11268
rect 11084 -11332 11104 -11268
rect 5732 -11348 11104 -11332
rect 5732 -11412 11020 -11348
rect 11084 -11412 11104 -11348
rect 5732 -11428 11104 -11412
rect 5732 -11492 11020 -11428
rect 11084 -11492 11104 -11428
rect 5732 -11508 11104 -11492
rect 5732 -11572 11020 -11508
rect 11084 -11572 11104 -11508
rect 5732 -11588 11104 -11572
rect 5732 -11652 11020 -11588
rect 11084 -11652 11104 -11588
rect 5732 -11668 11104 -11652
rect 5732 -11732 11020 -11668
rect 11084 -11732 11104 -11668
rect 5732 -11748 11104 -11732
rect 5732 -11812 11020 -11748
rect 11084 -11812 11104 -11748
rect 5732 -11828 11104 -11812
rect 5732 -11892 11020 -11828
rect 11084 -11892 11104 -11828
rect 5732 -11908 11104 -11892
rect 5732 -11972 11020 -11908
rect 11084 -11972 11104 -11908
rect 5732 -11988 11104 -11972
rect 5732 -12052 11020 -11988
rect 11084 -12052 11104 -11988
rect 5732 -12068 11104 -12052
rect 5732 -12132 11020 -12068
rect 11084 -12132 11104 -12068
rect 5732 -12148 11104 -12132
rect 5732 -12212 11020 -12148
rect 11084 -12212 11104 -12148
rect 5732 -12228 11104 -12212
rect 5732 -12292 11020 -12228
rect 11084 -12292 11104 -12228
rect 5732 -12308 11104 -12292
rect 5732 -12372 11020 -12308
rect 11084 -12372 11104 -12308
rect 5732 -12388 11104 -12372
rect 5732 -12452 11020 -12388
rect 11084 -12452 11104 -12388
rect 5732 -12468 11104 -12452
rect 5732 -12532 11020 -12468
rect 11084 -12532 11104 -12468
rect 5732 -12548 11104 -12532
rect 5732 -12612 11020 -12548
rect 11084 -12612 11104 -12548
rect 5732 -12628 11104 -12612
rect 5732 -12692 11020 -12628
rect 11084 -12692 11104 -12628
rect 5732 -12708 11104 -12692
rect 5732 -12772 11020 -12708
rect 11084 -12772 11104 -12708
rect 5732 -12788 11104 -12772
rect 5732 -12852 11020 -12788
rect 11084 -12852 11104 -12788
rect 5732 -12868 11104 -12852
rect 5732 -12932 11020 -12868
rect 11084 -12932 11104 -12868
rect 5732 -12948 11104 -12932
rect 5732 -13012 11020 -12948
rect 11084 -13012 11104 -12948
rect 5732 -13028 11104 -13012
rect 5732 -13092 11020 -13028
rect 11084 -13092 11104 -13028
rect 5732 -13108 11104 -13092
rect 5732 -13172 11020 -13108
rect 11084 -13172 11104 -13108
rect 5732 -13188 11104 -13172
rect 5732 -13252 11020 -13188
rect 11084 -13252 11104 -13188
rect 5732 -13268 11104 -13252
rect 5732 -13332 11020 -13268
rect 11084 -13332 11104 -13268
rect 5732 -13348 11104 -13332
rect 5732 -13412 11020 -13348
rect 11084 -13412 11104 -13348
rect 5732 -13428 11104 -13412
rect 5732 -13492 11020 -13428
rect 11084 -13492 11104 -13428
rect 5732 -13508 11104 -13492
rect 5732 -13572 11020 -13508
rect 11084 -13572 11104 -13508
rect 5732 -13588 11104 -13572
rect 5732 -13652 11020 -13588
rect 11084 -13652 11104 -13588
rect 5732 -13668 11104 -13652
rect 5732 -13732 11020 -13668
rect 11084 -13732 11104 -13668
rect 5732 -13748 11104 -13732
rect 5732 -13812 11020 -13748
rect 11084 -13812 11104 -13748
rect 5732 -13828 11104 -13812
rect 5732 -13892 11020 -13828
rect 11084 -13892 11104 -13828
rect 5732 -13908 11104 -13892
rect 5732 -13972 11020 -13908
rect 11084 -13972 11104 -13908
rect 5732 -13988 11104 -13972
rect 5732 -14052 11020 -13988
rect 11084 -14052 11104 -13988
rect 5732 -14068 11104 -14052
rect 5732 -14132 11020 -14068
rect 11084 -14132 11104 -14068
rect 5732 -14148 11104 -14132
rect 5732 -14212 11020 -14148
rect 11084 -14212 11104 -14148
rect 5732 -14228 11104 -14212
rect 5732 -14292 11020 -14228
rect 11084 -14292 11104 -14228
rect 5732 -14308 11104 -14292
rect 5732 -14372 11020 -14308
rect 11084 -14372 11104 -14308
rect 5732 -14388 11104 -14372
rect 5732 -14452 11020 -14388
rect 11084 -14452 11104 -14388
rect 5732 -14468 11104 -14452
rect 5732 -14532 11020 -14468
rect 11084 -14532 11104 -14468
rect 5732 -14548 11104 -14532
rect 5732 -14612 11020 -14548
rect 11084 -14612 11104 -14548
rect 5732 -14628 11104 -14612
rect 5732 -14692 11020 -14628
rect 11084 -14692 11104 -14628
rect 5732 -14708 11104 -14692
rect 5732 -14772 11020 -14708
rect 11084 -14772 11104 -14708
rect 5732 -14788 11104 -14772
rect 5732 -14852 11020 -14788
rect 11084 -14852 11104 -14788
rect 5732 -14868 11104 -14852
rect 5732 -14932 11020 -14868
rect 11084 -14932 11104 -14868
rect 5732 -14948 11104 -14932
rect 5732 -15012 11020 -14948
rect 11084 -15012 11104 -14948
rect 5732 -15028 11104 -15012
rect 5732 -15092 11020 -15028
rect 11084 -15092 11104 -15028
rect 5732 -15108 11104 -15092
rect 5732 -15172 11020 -15108
rect 11084 -15172 11104 -15108
rect 5732 -15188 11104 -15172
rect 5732 -15252 11020 -15188
rect 11084 -15252 11104 -15188
rect 5732 -15268 11104 -15252
rect 5732 -15332 11020 -15268
rect 11084 -15332 11104 -15268
rect 5732 -15348 11104 -15332
rect 5732 -15412 11020 -15348
rect 11084 -15412 11104 -15348
rect 5732 -15428 11104 -15412
rect 5732 -15492 11020 -15428
rect 11084 -15492 11104 -15428
rect 5732 -15508 11104 -15492
rect 5732 -15572 11020 -15508
rect 11084 -15572 11104 -15508
rect 5732 -15588 11104 -15572
rect 5732 -15652 11020 -15588
rect 11084 -15652 11104 -15588
rect 5732 -15668 11104 -15652
rect 5732 -15732 11020 -15668
rect 11084 -15732 11104 -15668
rect 5732 -15748 11104 -15732
rect 5732 -15812 11020 -15748
rect 11084 -15812 11104 -15748
rect 5732 -15840 11104 -15812
rect 11344 -10788 16716 -10760
rect 11344 -10852 16632 -10788
rect 16696 -10852 16716 -10788
rect 11344 -10868 16716 -10852
rect 11344 -10932 16632 -10868
rect 16696 -10932 16716 -10868
rect 11344 -10948 16716 -10932
rect 11344 -11012 16632 -10948
rect 16696 -11012 16716 -10948
rect 11344 -11028 16716 -11012
rect 11344 -11092 16632 -11028
rect 16696 -11092 16716 -11028
rect 11344 -11108 16716 -11092
rect 11344 -11172 16632 -11108
rect 16696 -11172 16716 -11108
rect 11344 -11188 16716 -11172
rect 11344 -11252 16632 -11188
rect 16696 -11252 16716 -11188
rect 11344 -11268 16716 -11252
rect 11344 -11332 16632 -11268
rect 16696 -11332 16716 -11268
rect 11344 -11348 16716 -11332
rect 11344 -11412 16632 -11348
rect 16696 -11412 16716 -11348
rect 11344 -11428 16716 -11412
rect 11344 -11492 16632 -11428
rect 16696 -11492 16716 -11428
rect 11344 -11508 16716 -11492
rect 11344 -11572 16632 -11508
rect 16696 -11572 16716 -11508
rect 11344 -11588 16716 -11572
rect 11344 -11652 16632 -11588
rect 16696 -11652 16716 -11588
rect 11344 -11668 16716 -11652
rect 11344 -11732 16632 -11668
rect 16696 -11732 16716 -11668
rect 11344 -11748 16716 -11732
rect 11344 -11812 16632 -11748
rect 16696 -11812 16716 -11748
rect 11344 -11828 16716 -11812
rect 11344 -11892 16632 -11828
rect 16696 -11892 16716 -11828
rect 11344 -11908 16716 -11892
rect 11344 -11972 16632 -11908
rect 16696 -11972 16716 -11908
rect 11344 -11988 16716 -11972
rect 11344 -12052 16632 -11988
rect 16696 -12052 16716 -11988
rect 11344 -12068 16716 -12052
rect 11344 -12132 16632 -12068
rect 16696 -12132 16716 -12068
rect 11344 -12148 16716 -12132
rect 11344 -12212 16632 -12148
rect 16696 -12212 16716 -12148
rect 11344 -12228 16716 -12212
rect 11344 -12292 16632 -12228
rect 16696 -12292 16716 -12228
rect 11344 -12308 16716 -12292
rect 11344 -12372 16632 -12308
rect 16696 -12372 16716 -12308
rect 11344 -12388 16716 -12372
rect 11344 -12452 16632 -12388
rect 16696 -12452 16716 -12388
rect 11344 -12468 16716 -12452
rect 11344 -12532 16632 -12468
rect 16696 -12532 16716 -12468
rect 11344 -12548 16716 -12532
rect 11344 -12612 16632 -12548
rect 16696 -12612 16716 -12548
rect 11344 -12628 16716 -12612
rect 11344 -12692 16632 -12628
rect 16696 -12692 16716 -12628
rect 11344 -12708 16716 -12692
rect 11344 -12772 16632 -12708
rect 16696 -12772 16716 -12708
rect 11344 -12788 16716 -12772
rect 11344 -12852 16632 -12788
rect 16696 -12852 16716 -12788
rect 11344 -12868 16716 -12852
rect 11344 -12932 16632 -12868
rect 16696 -12932 16716 -12868
rect 11344 -12948 16716 -12932
rect 11344 -13012 16632 -12948
rect 16696 -13012 16716 -12948
rect 11344 -13028 16716 -13012
rect 11344 -13092 16632 -13028
rect 16696 -13092 16716 -13028
rect 11344 -13108 16716 -13092
rect 11344 -13172 16632 -13108
rect 16696 -13172 16716 -13108
rect 11344 -13188 16716 -13172
rect 11344 -13252 16632 -13188
rect 16696 -13252 16716 -13188
rect 11344 -13268 16716 -13252
rect 11344 -13332 16632 -13268
rect 16696 -13332 16716 -13268
rect 11344 -13348 16716 -13332
rect 11344 -13412 16632 -13348
rect 16696 -13412 16716 -13348
rect 11344 -13428 16716 -13412
rect 11344 -13492 16632 -13428
rect 16696 -13492 16716 -13428
rect 11344 -13508 16716 -13492
rect 11344 -13572 16632 -13508
rect 16696 -13572 16716 -13508
rect 11344 -13588 16716 -13572
rect 11344 -13652 16632 -13588
rect 16696 -13652 16716 -13588
rect 11344 -13668 16716 -13652
rect 11344 -13732 16632 -13668
rect 16696 -13732 16716 -13668
rect 11344 -13748 16716 -13732
rect 11344 -13812 16632 -13748
rect 16696 -13812 16716 -13748
rect 11344 -13828 16716 -13812
rect 11344 -13892 16632 -13828
rect 16696 -13892 16716 -13828
rect 11344 -13908 16716 -13892
rect 11344 -13972 16632 -13908
rect 16696 -13972 16716 -13908
rect 11344 -13988 16716 -13972
rect 11344 -14052 16632 -13988
rect 16696 -14052 16716 -13988
rect 11344 -14068 16716 -14052
rect 11344 -14132 16632 -14068
rect 16696 -14132 16716 -14068
rect 11344 -14148 16716 -14132
rect 11344 -14212 16632 -14148
rect 16696 -14212 16716 -14148
rect 11344 -14228 16716 -14212
rect 11344 -14292 16632 -14228
rect 16696 -14292 16716 -14228
rect 11344 -14308 16716 -14292
rect 11344 -14372 16632 -14308
rect 16696 -14372 16716 -14308
rect 11344 -14388 16716 -14372
rect 11344 -14452 16632 -14388
rect 16696 -14452 16716 -14388
rect 11344 -14468 16716 -14452
rect 11344 -14532 16632 -14468
rect 16696 -14532 16716 -14468
rect 11344 -14548 16716 -14532
rect 11344 -14612 16632 -14548
rect 16696 -14612 16716 -14548
rect 11344 -14628 16716 -14612
rect 11344 -14692 16632 -14628
rect 16696 -14692 16716 -14628
rect 11344 -14708 16716 -14692
rect 11344 -14772 16632 -14708
rect 16696 -14772 16716 -14708
rect 11344 -14788 16716 -14772
rect 11344 -14852 16632 -14788
rect 16696 -14852 16716 -14788
rect 11344 -14868 16716 -14852
rect 11344 -14932 16632 -14868
rect 16696 -14932 16716 -14868
rect 11344 -14948 16716 -14932
rect 11344 -15012 16632 -14948
rect 16696 -15012 16716 -14948
rect 11344 -15028 16716 -15012
rect 11344 -15092 16632 -15028
rect 16696 -15092 16716 -15028
rect 11344 -15108 16716 -15092
rect 11344 -15172 16632 -15108
rect 16696 -15172 16716 -15108
rect 11344 -15188 16716 -15172
rect 11344 -15252 16632 -15188
rect 16696 -15252 16716 -15188
rect 11344 -15268 16716 -15252
rect 11344 -15332 16632 -15268
rect 16696 -15332 16716 -15268
rect 11344 -15348 16716 -15332
rect 11344 -15412 16632 -15348
rect 16696 -15412 16716 -15348
rect 11344 -15428 16716 -15412
rect 11344 -15492 16632 -15428
rect 16696 -15492 16716 -15428
rect 11344 -15508 16716 -15492
rect 11344 -15572 16632 -15508
rect 16696 -15572 16716 -15508
rect 11344 -15588 16716 -15572
rect 11344 -15652 16632 -15588
rect 16696 -15652 16716 -15588
rect 11344 -15668 16716 -15652
rect 11344 -15732 16632 -15668
rect 16696 -15732 16716 -15668
rect 11344 -15748 16716 -15732
rect 11344 -15812 16632 -15748
rect 16696 -15812 16716 -15748
rect 11344 -15840 16716 -15812
rect 16956 -10788 22328 -10760
rect 16956 -10852 22244 -10788
rect 22308 -10852 22328 -10788
rect 16956 -10868 22328 -10852
rect 16956 -10932 22244 -10868
rect 22308 -10932 22328 -10868
rect 16956 -10948 22328 -10932
rect 16956 -11012 22244 -10948
rect 22308 -11012 22328 -10948
rect 16956 -11028 22328 -11012
rect 16956 -11092 22244 -11028
rect 22308 -11092 22328 -11028
rect 16956 -11108 22328 -11092
rect 16956 -11172 22244 -11108
rect 22308 -11172 22328 -11108
rect 16956 -11188 22328 -11172
rect 16956 -11252 22244 -11188
rect 22308 -11252 22328 -11188
rect 16956 -11268 22328 -11252
rect 16956 -11332 22244 -11268
rect 22308 -11332 22328 -11268
rect 16956 -11348 22328 -11332
rect 16956 -11412 22244 -11348
rect 22308 -11412 22328 -11348
rect 16956 -11428 22328 -11412
rect 16956 -11492 22244 -11428
rect 22308 -11492 22328 -11428
rect 16956 -11508 22328 -11492
rect 16956 -11572 22244 -11508
rect 22308 -11572 22328 -11508
rect 16956 -11588 22328 -11572
rect 16956 -11652 22244 -11588
rect 22308 -11652 22328 -11588
rect 16956 -11668 22328 -11652
rect 16956 -11732 22244 -11668
rect 22308 -11732 22328 -11668
rect 16956 -11748 22328 -11732
rect 16956 -11812 22244 -11748
rect 22308 -11812 22328 -11748
rect 16956 -11828 22328 -11812
rect 16956 -11892 22244 -11828
rect 22308 -11892 22328 -11828
rect 16956 -11908 22328 -11892
rect 16956 -11972 22244 -11908
rect 22308 -11972 22328 -11908
rect 16956 -11988 22328 -11972
rect 16956 -12052 22244 -11988
rect 22308 -12052 22328 -11988
rect 16956 -12068 22328 -12052
rect 16956 -12132 22244 -12068
rect 22308 -12132 22328 -12068
rect 16956 -12148 22328 -12132
rect 16956 -12212 22244 -12148
rect 22308 -12212 22328 -12148
rect 16956 -12228 22328 -12212
rect 16956 -12292 22244 -12228
rect 22308 -12292 22328 -12228
rect 16956 -12308 22328 -12292
rect 16956 -12372 22244 -12308
rect 22308 -12372 22328 -12308
rect 16956 -12388 22328 -12372
rect 16956 -12452 22244 -12388
rect 22308 -12452 22328 -12388
rect 16956 -12468 22328 -12452
rect 16956 -12532 22244 -12468
rect 22308 -12532 22328 -12468
rect 16956 -12548 22328 -12532
rect 16956 -12612 22244 -12548
rect 22308 -12612 22328 -12548
rect 16956 -12628 22328 -12612
rect 16956 -12692 22244 -12628
rect 22308 -12692 22328 -12628
rect 16956 -12708 22328 -12692
rect 16956 -12772 22244 -12708
rect 22308 -12772 22328 -12708
rect 16956 -12788 22328 -12772
rect 16956 -12852 22244 -12788
rect 22308 -12852 22328 -12788
rect 16956 -12868 22328 -12852
rect 16956 -12932 22244 -12868
rect 22308 -12932 22328 -12868
rect 16956 -12948 22328 -12932
rect 16956 -13012 22244 -12948
rect 22308 -13012 22328 -12948
rect 16956 -13028 22328 -13012
rect 16956 -13092 22244 -13028
rect 22308 -13092 22328 -13028
rect 16956 -13108 22328 -13092
rect 16956 -13172 22244 -13108
rect 22308 -13172 22328 -13108
rect 16956 -13188 22328 -13172
rect 16956 -13252 22244 -13188
rect 22308 -13252 22328 -13188
rect 16956 -13268 22328 -13252
rect 16956 -13332 22244 -13268
rect 22308 -13332 22328 -13268
rect 16956 -13348 22328 -13332
rect 16956 -13412 22244 -13348
rect 22308 -13412 22328 -13348
rect 16956 -13428 22328 -13412
rect 16956 -13492 22244 -13428
rect 22308 -13492 22328 -13428
rect 16956 -13508 22328 -13492
rect 16956 -13572 22244 -13508
rect 22308 -13572 22328 -13508
rect 16956 -13588 22328 -13572
rect 16956 -13652 22244 -13588
rect 22308 -13652 22328 -13588
rect 16956 -13668 22328 -13652
rect 16956 -13732 22244 -13668
rect 22308 -13732 22328 -13668
rect 16956 -13748 22328 -13732
rect 16956 -13812 22244 -13748
rect 22308 -13812 22328 -13748
rect 16956 -13828 22328 -13812
rect 16956 -13892 22244 -13828
rect 22308 -13892 22328 -13828
rect 16956 -13908 22328 -13892
rect 16956 -13972 22244 -13908
rect 22308 -13972 22328 -13908
rect 16956 -13988 22328 -13972
rect 16956 -14052 22244 -13988
rect 22308 -14052 22328 -13988
rect 16956 -14068 22328 -14052
rect 16956 -14132 22244 -14068
rect 22308 -14132 22328 -14068
rect 16956 -14148 22328 -14132
rect 16956 -14212 22244 -14148
rect 22308 -14212 22328 -14148
rect 16956 -14228 22328 -14212
rect 16956 -14292 22244 -14228
rect 22308 -14292 22328 -14228
rect 16956 -14308 22328 -14292
rect 16956 -14372 22244 -14308
rect 22308 -14372 22328 -14308
rect 16956 -14388 22328 -14372
rect 16956 -14452 22244 -14388
rect 22308 -14452 22328 -14388
rect 16956 -14468 22328 -14452
rect 16956 -14532 22244 -14468
rect 22308 -14532 22328 -14468
rect 16956 -14548 22328 -14532
rect 16956 -14612 22244 -14548
rect 22308 -14612 22328 -14548
rect 16956 -14628 22328 -14612
rect 16956 -14692 22244 -14628
rect 22308 -14692 22328 -14628
rect 16956 -14708 22328 -14692
rect 16956 -14772 22244 -14708
rect 22308 -14772 22328 -14708
rect 16956 -14788 22328 -14772
rect 16956 -14852 22244 -14788
rect 22308 -14852 22328 -14788
rect 16956 -14868 22328 -14852
rect 16956 -14932 22244 -14868
rect 22308 -14932 22328 -14868
rect 16956 -14948 22328 -14932
rect 16956 -15012 22244 -14948
rect 22308 -15012 22328 -14948
rect 16956 -15028 22328 -15012
rect 16956 -15092 22244 -15028
rect 22308 -15092 22328 -15028
rect 16956 -15108 22328 -15092
rect 16956 -15172 22244 -15108
rect 22308 -15172 22328 -15108
rect 16956 -15188 22328 -15172
rect 16956 -15252 22244 -15188
rect 22308 -15252 22328 -15188
rect 16956 -15268 22328 -15252
rect 16956 -15332 22244 -15268
rect 22308 -15332 22328 -15268
rect 16956 -15348 22328 -15332
rect 16956 -15412 22244 -15348
rect 22308 -15412 22328 -15348
rect 16956 -15428 22328 -15412
rect 16956 -15492 22244 -15428
rect 22308 -15492 22328 -15428
rect 16956 -15508 22328 -15492
rect 16956 -15572 22244 -15508
rect 22308 -15572 22328 -15508
rect 16956 -15588 22328 -15572
rect 16956 -15652 22244 -15588
rect 22308 -15652 22328 -15588
rect 16956 -15668 22328 -15652
rect 16956 -15732 22244 -15668
rect 22308 -15732 22328 -15668
rect 16956 -15748 22328 -15732
rect 16956 -15812 22244 -15748
rect 22308 -15812 22328 -15748
rect 16956 -15840 22328 -15812
rect 22568 -10788 27940 -10760
rect 22568 -10852 27856 -10788
rect 27920 -10852 27940 -10788
rect 22568 -10868 27940 -10852
rect 22568 -10932 27856 -10868
rect 27920 -10932 27940 -10868
rect 22568 -10948 27940 -10932
rect 22568 -11012 27856 -10948
rect 27920 -11012 27940 -10948
rect 22568 -11028 27940 -11012
rect 22568 -11092 27856 -11028
rect 27920 -11092 27940 -11028
rect 22568 -11108 27940 -11092
rect 22568 -11172 27856 -11108
rect 27920 -11172 27940 -11108
rect 22568 -11188 27940 -11172
rect 22568 -11252 27856 -11188
rect 27920 -11252 27940 -11188
rect 22568 -11268 27940 -11252
rect 22568 -11332 27856 -11268
rect 27920 -11332 27940 -11268
rect 22568 -11348 27940 -11332
rect 22568 -11412 27856 -11348
rect 27920 -11412 27940 -11348
rect 22568 -11428 27940 -11412
rect 22568 -11492 27856 -11428
rect 27920 -11492 27940 -11428
rect 22568 -11508 27940 -11492
rect 22568 -11572 27856 -11508
rect 27920 -11572 27940 -11508
rect 22568 -11588 27940 -11572
rect 22568 -11652 27856 -11588
rect 27920 -11652 27940 -11588
rect 22568 -11668 27940 -11652
rect 22568 -11732 27856 -11668
rect 27920 -11732 27940 -11668
rect 22568 -11748 27940 -11732
rect 22568 -11812 27856 -11748
rect 27920 -11812 27940 -11748
rect 22568 -11828 27940 -11812
rect 22568 -11892 27856 -11828
rect 27920 -11892 27940 -11828
rect 22568 -11908 27940 -11892
rect 22568 -11972 27856 -11908
rect 27920 -11972 27940 -11908
rect 22568 -11988 27940 -11972
rect 22568 -12052 27856 -11988
rect 27920 -12052 27940 -11988
rect 22568 -12068 27940 -12052
rect 22568 -12132 27856 -12068
rect 27920 -12132 27940 -12068
rect 22568 -12148 27940 -12132
rect 22568 -12212 27856 -12148
rect 27920 -12212 27940 -12148
rect 22568 -12228 27940 -12212
rect 22568 -12292 27856 -12228
rect 27920 -12292 27940 -12228
rect 22568 -12308 27940 -12292
rect 22568 -12372 27856 -12308
rect 27920 -12372 27940 -12308
rect 22568 -12388 27940 -12372
rect 22568 -12452 27856 -12388
rect 27920 -12452 27940 -12388
rect 22568 -12468 27940 -12452
rect 22568 -12532 27856 -12468
rect 27920 -12532 27940 -12468
rect 22568 -12548 27940 -12532
rect 22568 -12612 27856 -12548
rect 27920 -12612 27940 -12548
rect 22568 -12628 27940 -12612
rect 22568 -12692 27856 -12628
rect 27920 -12692 27940 -12628
rect 22568 -12708 27940 -12692
rect 22568 -12772 27856 -12708
rect 27920 -12772 27940 -12708
rect 22568 -12788 27940 -12772
rect 22568 -12852 27856 -12788
rect 27920 -12852 27940 -12788
rect 22568 -12868 27940 -12852
rect 22568 -12932 27856 -12868
rect 27920 -12932 27940 -12868
rect 22568 -12948 27940 -12932
rect 22568 -13012 27856 -12948
rect 27920 -13012 27940 -12948
rect 22568 -13028 27940 -13012
rect 22568 -13092 27856 -13028
rect 27920 -13092 27940 -13028
rect 22568 -13108 27940 -13092
rect 22568 -13172 27856 -13108
rect 27920 -13172 27940 -13108
rect 22568 -13188 27940 -13172
rect 22568 -13252 27856 -13188
rect 27920 -13252 27940 -13188
rect 22568 -13268 27940 -13252
rect 22568 -13332 27856 -13268
rect 27920 -13332 27940 -13268
rect 22568 -13348 27940 -13332
rect 22568 -13412 27856 -13348
rect 27920 -13412 27940 -13348
rect 22568 -13428 27940 -13412
rect 22568 -13492 27856 -13428
rect 27920 -13492 27940 -13428
rect 22568 -13508 27940 -13492
rect 22568 -13572 27856 -13508
rect 27920 -13572 27940 -13508
rect 22568 -13588 27940 -13572
rect 22568 -13652 27856 -13588
rect 27920 -13652 27940 -13588
rect 22568 -13668 27940 -13652
rect 22568 -13732 27856 -13668
rect 27920 -13732 27940 -13668
rect 22568 -13748 27940 -13732
rect 22568 -13812 27856 -13748
rect 27920 -13812 27940 -13748
rect 22568 -13828 27940 -13812
rect 22568 -13892 27856 -13828
rect 27920 -13892 27940 -13828
rect 22568 -13908 27940 -13892
rect 22568 -13972 27856 -13908
rect 27920 -13972 27940 -13908
rect 22568 -13988 27940 -13972
rect 22568 -14052 27856 -13988
rect 27920 -14052 27940 -13988
rect 22568 -14068 27940 -14052
rect 22568 -14132 27856 -14068
rect 27920 -14132 27940 -14068
rect 22568 -14148 27940 -14132
rect 22568 -14212 27856 -14148
rect 27920 -14212 27940 -14148
rect 22568 -14228 27940 -14212
rect 22568 -14292 27856 -14228
rect 27920 -14292 27940 -14228
rect 22568 -14308 27940 -14292
rect 22568 -14372 27856 -14308
rect 27920 -14372 27940 -14308
rect 22568 -14388 27940 -14372
rect 22568 -14452 27856 -14388
rect 27920 -14452 27940 -14388
rect 22568 -14468 27940 -14452
rect 22568 -14532 27856 -14468
rect 27920 -14532 27940 -14468
rect 22568 -14548 27940 -14532
rect 22568 -14612 27856 -14548
rect 27920 -14612 27940 -14548
rect 22568 -14628 27940 -14612
rect 22568 -14692 27856 -14628
rect 27920 -14692 27940 -14628
rect 22568 -14708 27940 -14692
rect 22568 -14772 27856 -14708
rect 27920 -14772 27940 -14708
rect 22568 -14788 27940 -14772
rect 22568 -14852 27856 -14788
rect 27920 -14852 27940 -14788
rect 22568 -14868 27940 -14852
rect 22568 -14932 27856 -14868
rect 27920 -14932 27940 -14868
rect 22568 -14948 27940 -14932
rect 22568 -15012 27856 -14948
rect 27920 -15012 27940 -14948
rect 22568 -15028 27940 -15012
rect 22568 -15092 27856 -15028
rect 27920 -15092 27940 -15028
rect 22568 -15108 27940 -15092
rect 22568 -15172 27856 -15108
rect 27920 -15172 27940 -15108
rect 22568 -15188 27940 -15172
rect 22568 -15252 27856 -15188
rect 27920 -15252 27940 -15188
rect 22568 -15268 27940 -15252
rect 22568 -15332 27856 -15268
rect 27920 -15332 27940 -15268
rect 22568 -15348 27940 -15332
rect 22568 -15412 27856 -15348
rect 27920 -15412 27940 -15348
rect 22568 -15428 27940 -15412
rect 22568 -15492 27856 -15428
rect 27920 -15492 27940 -15428
rect 22568 -15508 27940 -15492
rect 22568 -15572 27856 -15508
rect 27920 -15572 27940 -15508
rect 22568 -15588 27940 -15572
rect 22568 -15652 27856 -15588
rect 27920 -15652 27940 -15588
rect 22568 -15668 27940 -15652
rect 22568 -15732 27856 -15668
rect 27920 -15732 27940 -15668
rect 22568 -15748 27940 -15732
rect 22568 -15812 27856 -15748
rect 27920 -15812 27940 -15748
rect 22568 -15840 27940 -15812
rect 28180 -10788 33552 -10760
rect 28180 -10852 33468 -10788
rect 33532 -10852 33552 -10788
rect 28180 -10868 33552 -10852
rect 28180 -10932 33468 -10868
rect 33532 -10932 33552 -10868
rect 28180 -10948 33552 -10932
rect 28180 -11012 33468 -10948
rect 33532 -11012 33552 -10948
rect 28180 -11028 33552 -11012
rect 28180 -11092 33468 -11028
rect 33532 -11092 33552 -11028
rect 28180 -11108 33552 -11092
rect 28180 -11172 33468 -11108
rect 33532 -11172 33552 -11108
rect 28180 -11188 33552 -11172
rect 28180 -11252 33468 -11188
rect 33532 -11252 33552 -11188
rect 28180 -11268 33552 -11252
rect 28180 -11332 33468 -11268
rect 33532 -11332 33552 -11268
rect 28180 -11348 33552 -11332
rect 28180 -11412 33468 -11348
rect 33532 -11412 33552 -11348
rect 28180 -11428 33552 -11412
rect 28180 -11492 33468 -11428
rect 33532 -11492 33552 -11428
rect 28180 -11508 33552 -11492
rect 28180 -11572 33468 -11508
rect 33532 -11572 33552 -11508
rect 28180 -11588 33552 -11572
rect 28180 -11652 33468 -11588
rect 33532 -11652 33552 -11588
rect 28180 -11668 33552 -11652
rect 28180 -11732 33468 -11668
rect 33532 -11732 33552 -11668
rect 28180 -11748 33552 -11732
rect 28180 -11812 33468 -11748
rect 33532 -11812 33552 -11748
rect 28180 -11828 33552 -11812
rect 28180 -11892 33468 -11828
rect 33532 -11892 33552 -11828
rect 28180 -11908 33552 -11892
rect 28180 -11972 33468 -11908
rect 33532 -11972 33552 -11908
rect 28180 -11988 33552 -11972
rect 28180 -12052 33468 -11988
rect 33532 -12052 33552 -11988
rect 28180 -12068 33552 -12052
rect 28180 -12132 33468 -12068
rect 33532 -12132 33552 -12068
rect 28180 -12148 33552 -12132
rect 28180 -12212 33468 -12148
rect 33532 -12212 33552 -12148
rect 28180 -12228 33552 -12212
rect 28180 -12292 33468 -12228
rect 33532 -12292 33552 -12228
rect 28180 -12308 33552 -12292
rect 28180 -12372 33468 -12308
rect 33532 -12372 33552 -12308
rect 28180 -12388 33552 -12372
rect 28180 -12452 33468 -12388
rect 33532 -12452 33552 -12388
rect 28180 -12468 33552 -12452
rect 28180 -12532 33468 -12468
rect 33532 -12532 33552 -12468
rect 28180 -12548 33552 -12532
rect 28180 -12612 33468 -12548
rect 33532 -12612 33552 -12548
rect 28180 -12628 33552 -12612
rect 28180 -12692 33468 -12628
rect 33532 -12692 33552 -12628
rect 28180 -12708 33552 -12692
rect 28180 -12772 33468 -12708
rect 33532 -12772 33552 -12708
rect 28180 -12788 33552 -12772
rect 28180 -12852 33468 -12788
rect 33532 -12852 33552 -12788
rect 28180 -12868 33552 -12852
rect 28180 -12932 33468 -12868
rect 33532 -12932 33552 -12868
rect 28180 -12948 33552 -12932
rect 28180 -13012 33468 -12948
rect 33532 -13012 33552 -12948
rect 28180 -13028 33552 -13012
rect 28180 -13092 33468 -13028
rect 33532 -13092 33552 -13028
rect 28180 -13108 33552 -13092
rect 28180 -13172 33468 -13108
rect 33532 -13172 33552 -13108
rect 28180 -13188 33552 -13172
rect 28180 -13252 33468 -13188
rect 33532 -13252 33552 -13188
rect 28180 -13268 33552 -13252
rect 28180 -13332 33468 -13268
rect 33532 -13332 33552 -13268
rect 28180 -13348 33552 -13332
rect 28180 -13412 33468 -13348
rect 33532 -13412 33552 -13348
rect 28180 -13428 33552 -13412
rect 28180 -13492 33468 -13428
rect 33532 -13492 33552 -13428
rect 28180 -13508 33552 -13492
rect 28180 -13572 33468 -13508
rect 33532 -13572 33552 -13508
rect 28180 -13588 33552 -13572
rect 28180 -13652 33468 -13588
rect 33532 -13652 33552 -13588
rect 28180 -13668 33552 -13652
rect 28180 -13732 33468 -13668
rect 33532 -13732 33552 -13668
rect 28180 -13748 33552 -13732
rect 28180 -13812 33468 -13748
rect 33532 -13812 33552 -13748
rect 28180 -13828 33552 -13812
rect 28180 -13892 33468 -13828
rect 33532 -13892 33552 -13828
rect 28180 -13908 33552 -13892
rect 28180 -13972 33468 -13908
rect 33532 -13972 33552 -13908
rect 28180 -13988 33552 -13972
rect 28180 -14052 33468 -13988
rect 33532 -14052 33552 -13988
rect 28180 -14068 33552 -14052
rect 28180 -14132 33468 -14068
rect 33532 -14132 33552 -14068
rect 28180 -14148 33552 -14132
rect 28180 -14212 33468 -14148
rect 33532 -14212 33552 -14148
rect 28180 -14228 33552 -14212
rect 28180 -14292 33468 -14228
rect 33532 -14292 33552 -14228
rect 28180 -14308 33552 -14292
rect 28180 -14372 33468 -14308
rect 33532 -14372 33552 -14308
rect 28180 -14388 33552 -14372
rect 28180 -14452 33468 -14388
rect 33532 -14452 33552 -14388
rect 28180 -14468 33552 -14452
rect 28180 -14532 33468 -14468
rect 33532 -14532 33552 -14468
rect 28180 -14548 33552 -14532
rect 28180 -14612 33468 -14548
rect 33532 -14612 33552 -14548
rect 28180 -14628 33552 -14612
rect 28180 -14692 33468 -14628
rect 33532 -14692 33552 -14628
rect 28180 -14708 33552 -14692
rect 28180 -14772 33468 -14708
rect 33532 -14772 33552 -14708
rect 28180 -14788 33552 -14772
rect 28180 -14852 33468 -14788
rect 33532 -14852 33552 -14788
rect 28180 -14868 33552 -14852
rect 28180 -14932 33468 -14868
rect 33532 -14932 33552 -14868
rect 28180 -14948 33552 -14932
rect 28180 -15012 33468 -14948
rect 33532 -15012 33552 -14948
rect 28180 -15028 33552 -15012
rect 28180 -15092 33468 -15028
rect 33532 -15092 33552 -15028
rect 28180 -15108 33552 -15092
rect 28180 -15172 33468 -15108
rect 33532 -15172 33552 -15108
rect 28180 -15188 33552 -15172
rect 28180 -15252 33468 -15188
rect 33532 -15252 33552 -15188
rect 28180 -15268 33552 -15252
rect 28180 -15332 33468 -15268
rect 33532 -15332 33552 -15268
rect 28180 -15348 33552 -15332
rect 28180 -15412 33468 -15348
rect 33532 -15412 33552 -15348
rect 28180 -15428 33552 -15412
rect 28180 -15492 33468 -15428
rect 33532 -15492 33552 -15428
rect 28180 -15508 33552 -15492
rect 28180 -15572 33468 -15508
rect 33532 -15572 33552 -15508
rect 28180 -15588 33552 -15572
rect 28180 -15652 33468 -15588
rect 33532 -15652 33552 -15588
rect 28180 -15668 33552 -15652
rect 28180 -15732 33468 -15668
rect 33532 -15732 33552 -15668
rect 28180 -15748 33552 -15732
rect 28180 -15812 33468 -15748
rect 33532 -15812 33552 -15748
rect 28180 -15840 33552 -15812
rect 33792 -10788 39164 -10760
rect 33792 -10852 39080 -10788
rect 39144 -10852 39164 -10788
rect 33792 -10868 39164 -10852
rect 33792 -10932 39080 -10868
rect 39144 -10932 39164 -10868
rect 33792 -10948 39164 -10932
rect 33792 -11012 39080 -10948
rect 39144 -11012 39164 -10948
rect 33792 -11028 39164 -11012
rect 33792 -11092 39080 -11028
rect 39144 -11092 39164 -11028
rect 33792 -11108 39164 -11092
rect 33792 -11172 39080 -11108
rect 39144 -11172 39164 -11108
rect 33792 -11188 39164 -11172
rect 33792 -11252 39080 -11188
rect 39144 -11252 39164 -11188
rect 33792 -11268 39164 -11252
rect 33792 -11332 39080 -11268
rect 39144 -11332 39164 -11268
rect 33792 -11348 39164 -11332
rect 33792 -11412 39080 -11348
rect 39144 -11412 39164 -11348
rect 33792 -11428 39164 -11412
rect 33792 -11492 39080 -11428
rect 39144 -11492 39164 -11428
rect 33792 -11508 39164 -11492
rect 33792 -11572 39080 -11508
rect 39144 -11572 39164 -11508
rect 33792 -11588 39164 -11572
rect 33792 -11652 39080 -11588
rect 39144 -11652 39164 -11588
rect 33792 -11668 39164 -11652
rect 33792 -11732 39080 -11668
rect 39144 -11732 39164 -11668
rect 33792 -11748 39164 -11732
rect 33792 -11812 39080 -11748
rect 39144 -11812 39164 -11748
rect 33792 -11828 39164 -11812
rect 33792 -11892 39080 -11828
rect 39144 -11892 39164 -11828
rect 33792 -11908 39164 -11892
rect 33792 -11972 39080 -11908
rect 39144 -11972 39164 -11908
rect 33792 -11988 39164 -11972
rect 33792 -12052 39080 -11988
rect 39144 -12052 39164 -11988
rect 33792 -12068 39164 -12052
rect 33792 -12132 39080 -12068
rect 39144 -12132 39164 -12068
rect 33792 -12148 39164 -12132
rect 33792 -12212 39080 -12148
rect 39144 -12212 39164 -12148
rect 33792 -12228 39164 -12212
rect 33792 -12292 39080 -12228
rect 39144 -12292 39164 -12228
rect 33792 -12308 39164 -12292
rect 33792 -12372 39080 -12308
rect 39144 -12372 39164 -12308
rect 33792 -12388 39164 -12372
rect 33792 -12452 39080 -12388
rect 39144 -12452 39164 -12388
rect 33792 -12468 39164 -12452
rect 33792 -12532 39080 -12468
rect 39144 -12532 39164 -12468
rect 33792 -12548 39164 -12532
rect 33792 -12612 39080 -12548
rect 39144 -12612 39164 -12548
rect 33792 -12628 39164 -12612
rect 33792 -12692 39080 -12628
rect 39144 -12692 39164 -12628
rect 33792 -12708 39164 -12692
rect 33792 -12772 39080 -12708
rect 39144 -12772 39164 -12708
rect 33792 -12788 39164 -12772
rect 33792 -12852 39080 -12788
rect 39144 -12852 39164 -12788
rect 33792 -12868 39164 -12852
rect 33792 -12932 39080 -12868
rect 39144 -12932 39164 -12868
rect 33792 -12948 39164 -12932
rect 33792 -13012 39080 -12948
rect 39144 -13012 39164 -12948
rect 33792 -13028 39164 -13012
rect 33792 -13092 39080 -13028
rect 39144 -13092 39164 -13028
rect 33792 -13108 39164 -13092
rect 33792 -13172 39080 -13108
rect 39144 -13172 39164 -13108
rect 33792 -13188 39164 -13172
rect 33792 -13252 39080 -13188
rect 39144 -13252 39164 -13188
rect 33792 -13268 39164 -13252
rect 33792 -13332 39080 -13268
rect 39144 -13332 39164 -13268
rect 33792 -13348 39164 -13332
rect 33792 -13412 39080 -13348
rect 39144 -13412 39164 -13348
rect 33792 -13428 39164 -13412
rect 33792 -13492 39080 -13428
rect 39144 -13492 39164 -13428
rect 33792 -13508 39164 -13492
rect 33792 -13572 39080 -13508
rect 39144 -13572 39164 -13508
rect 33792 -13588 39164 -13572
rect 33792 -13652 39080 -13588
rect 39144 -13652 39164 -13588
rect 33792 -13668 39164 -13652
rect 33792 -13732 39080 -13668
rect 39144 -13732 39164 -13668
rect 33792 -13748 39164 -13732
rect 33792 -13812 39080 -13748
rect 39144 -13812 39164 -13748
rect 33792 -13828 39164 -13812
rect 33792 -13892 39080 -13828
rect 39144 -13892 39164 -13828
rect 33792 -13908 39164 -13892
rect 33792 -13972 39080 -13908
rect 39144 -13972 39164 -13908
rect 33792 -13988 39164 -13972
rect 33792 -14052 39080 -13988
rect 39144 -14052 39164 -13988
rect 33792 -14068 39164 -14052
rect 33792 -14132 39080 -14068
rect 39144 -14132 39164 -14068
rect 33792 -14148 39164 -14132
rect 33792 -14212 39080 -14148
rect 39144 -14212 39164 -14148
rect 33792 -14228 39164 -14212
rect 33792 -14292 39080 -14228
rect 39144 -14292 39164 -14228
rect 33792 -14308 39164 -14292
rect 33792 -14372 39080 -14308
rect 39144 -14372 39164 -14308
rect 33792 -14388 39164 -14372
rect 33792 -14452 39080 -14388
rect 39144 -14452 39164 -14388
rect 33792 -14468 39164 -14452
rect 33792 -14532 39080 -14468
rect 39144 -14532 39164 -14468
rect 33792 -14548 39164 -14532
rect 33792 -14612 39080 -14548
rect 39144 -14612 39164 -14548
rect 33792 -14628 39164 -14612
rect 33792 -14692 39080 -14628
rect 39144 -14692 39164 -14628
rect 33792 -14708 39164 -14692
rect 33792 -14772 39080 -14708
rect 39144 -14772 39164 -14708
rect 33792 -14788 39164 -14772
rect 33792 -14852 39080 -14788
rect 39144 -14852 39164 -14788
rect 33792 -14868 39164 -14852
rect 33792 -14932 39080 -14868
rect 39144 -14932 39164 -14868
rect 33792 -14948 39164 -14932
rect 33792 -15012 39080 -14948
rect 39144 -15012 39164 -14948
rect 33792 -15028 39164 -15012
rect 33792 -15092 39080 -15028
rect 39144 -15092 39164 -15028
rect 33792 -15108 39164 -15092
rect 33792 -15172 39080 -15108
rect 39144 -15172 39164 -15108
rect 33792 -15188 39164 -15172
rect 33792 -15252 39080 -15188
rect 39144 -15252 39164 -15188
rect 33792 -15268 39164 -15252
rect 33792 -15332 39080 -15268
rect 39144 -15332 39164 -15268
rect 33792 -15348 39164 -15332
rect 33792 -15412 39080 -15348
rect 39144 -15412 39164 -15348
rect 33792 -15428 39164 -15412
rect 33792 -15492 39080 -15428
rect 39144 -15492 39164 -15428
rect 33792 -15508 39164 -15492
rect 33792 -15572 39080 -15508
rect 39144 -15572 39164 -15508
rect 33792 -15588 39164 -15572
rect 33792 -15652 39080 -15588
rect 39144 -15652 39164 -15588
rect 33792 -15668 39164 -15652
rect 33792 -15732 39080 -15668
rect 39144 -15732 39164 -15668
rect 33792 -15748 39164 -15732
rect 33792 -15812 39080 -15748
rect 39144 -15812 39164 -15748
rect 33792 -15840 39164 -15812
rect -39164 -16108 -33792 -16080
rect -39164 -16172 -33876 -16108
rect -33812 -16172 -33792 -16108
rect -39164 -16188 -33792 -16172
rect -39164 -16252 -33876 -16188
rect -33812 -16252 -33792 -16188
rect -39164 -16268 -33792 -16252
rect -39164 -16332 -33876 -16268
rect -33812 -16332 -33792 -16268
rect -39164 -16348 -33792 -16332
rect -39164 -16412 -33876 -16348
rect -33812 -16412 -33792 -16348
rect -39164 -16428 -33792 -16412
rect -39164 -16492 -33876 -16428
rect -33812 -16492 -33792 -16428
rect -39164 -16508 -33792 -16492
rect -39164 -16572 -33876 -16508
rect -33812 -16572 -33792 -16508
rect -39164 -16588 -33792 -16572
rect -39164 -16652 -33876 -16588
rect -33812 -16652 -33792 -16588
rect -39164 -16668 -33792 -16652
rect -39164 -16732 -33876 -16668
rect -33812 -16732 -33792 -16668
rect -39164 -16748 -33792 -16732
rect -39164 -16812 -33876 -16748
rect -33812 -16812 -33792 -16748
rect -39164 -16828 -33792 -16812
rect -39164 -16892 -33876 -16828
rect -33812 -16892 -33792 -16828
rect -39164 -16908 -33792 -16892
rect -39164 -16972 -33876 -16908
rect -33812 -16972 -33792 -16908
rect -39164 -16988 -33792 -16972
rect -39164 -17052 -33876 -16988
rect -33812 -17052 -33792 -16988
rect -39164 -17068 -33792 -17052
rect -39164 -17132 -33876 -17068
rect -33812 -17132 -33792 -17068
rect -39164 -17148 -33792 -17132
rect -39164 -17212 -33876 -17148
rect -33812 -17212 -33792 -17148
rect -39164 -17228 -33792 -17212
rect -39164 -17292 -33876 -17228
rect -33812 -17292 -33792 -17228
rect -39164 -17308 -33792 -17292
rect -39164 -17372 -33876 -17308
rect -33812 -17372 -33792 -17308
rect -39164 -17388 -33792 -17372
rect -39164 -17452 -33876 -17388
rect -33812 -17452 -33792 -17388
rect -39164 -17468 -33792 -17452
rect -39164 -17532 -33876 -17468
rect -33812 -17532 -33792 -17468
rect -39164 -17548 -33792 -17532
rect -39164 -17612 -33876 -17548
rect -33812 -17612 -33792 -17548
rect -39164 -17628 -33792 -17612
rect -39164 -17692 -33876 -17628
rect -33812 -17692 -33792 -17628
rect -39164 -17708 -33792 -17692
rect -39164 -17772 -33876 -17708
rect -33812 -17772 -33792 -17708
rect -39164 -17788 -33792 -17772
rect -39164 -17852 -33876 -17788
rect -33812 -17852 -33792 -17788
rect -39164 -17868 -33792 -17852
rect -39164 -17932 -33876 -17868
rect -33812 -17932 -33792 -17868
rect -39164 -17948 -33792 -17932
rect -39164 -18012 -33876 -17948
rect -33812 -18012 -33792 -17948
rect -39164 -18028 -33792 -18012
rect -39164 -18092 -33876 -18028
rect -33812 -18092 -33792 -18028
rect -39164 -18108 -33792 -18092
rect -39164 -18172 -33876 -18108
rect -33812 -18172 -33792 -18108
rect -39164 -18188 -33792 -18172
rect -39164 -18252 -33876 -18188
rect -33812 -18252 -33792 -18188
rect -39164 -18268 -33792 -18252
rect -39164 -18332 -33876 -18268
rect -33812 -18332 -33792 -18268
rect -39164 -18348 -33792 -18332
rect -39164 -18412 -33876 -18348
rect -33812 -18412 -33792 -18348
rect -39164 -18428 -33792 -18412
rect -39164 -18492 -33876 -18428
rect -33812 -18492 -33792 -18428
rect -39164 -18508 -33792 -18492
rect -39164 -18572 -33876 -18508
rect -33812 -18572 -33792 -18508
rect -39164 -18588 -33792 -18572
rect -39164 -18652 -33876 -18588
rect -33812 -18652 -33792 -18588
rect -39164 -18668 -33792 -18652
rect -39164 -18732 -33876 -18668
rect -33812 -18732 -33792 -18668
rect -39164 -18748 -33792 -18732
rect -39164 -18812 -33876 -18748
rect -33812 -18812 -33792 -18748
rect -39164 -18828 -33792 -18812
rect -39164 -18892 -33876 -18828
rect -33812 -18892 -33792 -18828
rect -39164 -18908 -33792 -18892
rect -39164 -18972 -33876 -18908
rect -33812 -18972 -33792 -18908
rect -39164 -18988 -33792 -18972
rect -39164 -19052 -33876 -18988
rect -33812 -19052 -33792 -18988
rect -39164 -19068 -33792 -19052
rect -39164 -19132 -33876 -19068
rect -33812 -19132 -33792 -19068
rect -39164 -19148 -33792 -19132
rect -39164 -19212 -33876 -19148
rect -33812 -19212 -33792 -19148
rect -39164 -19228 -33792 -19212
rect -39164 -19292 -33876 -19228
rect -33812 -19292 -33792 -19228
rect -39164 -19308 -33792 -19292
rect -39164 -19372 -33876 -19308
rect -33812 -19372 -33792 -19308
rect -39164 -19388 -33792 -19372
rect -39164 -19452 -33876 -19388
rect -33812 -19452 -33792 -19388
rect -39164 -19468 -33792 -19452
rect -39164 -19532 -33876 -19468
rect -33812 -19532 -33792 -19468
rect -39164 -19548 -33792 -19532
rect -39164 -19612 -33876 -19548
rect -33812 -19612 -33792 -19548
rect -39164 -19628 -33792 -19612
rect -39164 -19692 -33876 -19628
rect -33812 -19692 -33792 -19628
rect -39164 -19708 -33792 -19692
rect -39164 -19772 -33876 -19708
rect -33812 -19772 -33792 -19708
rect -39164 -19788 -33792 -19772
rect -39164 -19852 -33876 -19788
rect -33812 -19852 -33792 -19788
rect -39164 -19868 -33792 -19852
rect -39164 -19932 -33876 -19868
rect -33812 -19932 -33792 -19868
rect -39164 -19948 -33792 -19932
rect -39164 -20012 -33876 -19948
rect -33812 -20012 -33792 -19948
rect -39164 -20028 -33792 -20012
rect -39164 -20092 -33876 -20028
rect -33812 -20092 -33792 -20028
rect -39164 -20108 -33792 -20092
rect -39164 -20172 -33876 -20108
rect -33812 -20172 -33792 -20108
rect -39164 -20188 -33792 -20172
rect -39164 -20252 -33876 -20188
rect -33812 -20252 -33792 -20188
rect -39164 -20268 -33792 -20252
rect -39164 -20332 -33876 -20268
rect -33812 -20332 -33792 -20268
rect -39164 -20348 -33792 -20332
rect -39164 -20412 -33876 -20348
rect -33812 -20412 -33792 -20348
rect -39164 -20428 -33792 -20412
rect -39164 -20492 -33876 -20428
rect -33812 -20492 -33792 -20428
rect -39164 -20508 -33792 -20492
rect -39164 -20572 -33876 -20508
rect -33812 -20572 -33792 -20508
rect -39164 -20588 -33792 -20572
rect -39164 -20652 -33876 -20588
rect -33812 -20652 -33792 -20588
rect -39164 -20668 -33792 -20652
rect -39164 -20732 -33876 -20668
rect -33812 -20732 -33792 -20668
rect -39164 -20748 -33792 -20732
rect -39164 -20812 -33876 -20748
rect -33812 -20812 -33792 -20748
rect -39164 -20828 -33792 -20812
rect -39164 -20892 -33876 -20828
rect -33812 -20892 -33792 -20828
rect -39164 -20908 -33792 -20892
rect -39164 -20972 -33876 -20908
rect -33812 -20972 -33792 -20908
rect -39164 -20988 -33792 -20972
rect -39164 -21052 -33876 -20988
rect -33812 -21052 -33792 -20988
rect -39164 -21068 -33792 -21052
rect -39164 -21132 -33876 -21068
rect -33812 -21132 -33792 -21068
rect -39164 -21160 -33792 -21132
rect -33552 -16108 -28180 -16080
rect -33552 -16172 -28264 -16108
rect -28200 -16172 -28180 -16108
rect -33552 -16188 -28180 -16172
rect -33552 -16252 -28264 -16188
rect -28200 -16252 -28180 -16188
rect -33552 -16268 -28180 -16252
rect -33552 -16332 -28264 -16268
rect -28200 -16332 -28180 -16268
rect -33552 -16348 -28180 -16332
rect -33552 -16412 -28264 -16348
rect -28200 -16412 -28180 -16348
rect -33552 -16428 -28180 -16412
rect -33552 -16492 -28264 -16428
rect -28200 -16492 -28180 -16428
rect -33552 -16508 -28180 -16492
rect -33552 -16572 -28264 -16508
rect -28200 -16572 -28180 -16508
rect -33552 -16588 -28180 -16572
rect -33552 -16652 -28264 -16588
rect -28200 -16652 -28180 -16588
rect -33552 -16668 -28180 -16652
rect -33552 -16732 -28264 -16668
rect -28200 -16732 -28180 -16668
rect -33552 -16748 -28180 -16732
rect -33552 -16812 -28264 -16748
rect -28200 -16812 -28180 -16748
rect -33552 -16828 -28180 -16812
rect -33552 -16892 -28264 -16828
rect -28200 -16892 -28180 -16828
rect -33552 -16908 -28180 -16892
rect -33552 -16972 -28264 -16908
rect -28200 -16972 -28180 -16908
rect -33552 -16988 -28180 -16972
rect -33552 -17052 -28264 -16988
rect -28200 -17052 -28180 -16988
rect -33552 -17068 -28180 -17052
rect -33552 -17132 -28264 -17068
rect -28200 -17132 -28180 -17068
rect -33552 -17148 -28180 -17132
rect -33552 -17212 -28264 -17148
rect -28200 -17212 -28180 -17148
rect -33552 -17228 -28180 -17212
rect -33552 -17292 -28264 -17228
rect -28200 -17292 -28180 -17228
rect -33552 -17308 -28180 -17292
rect -33552 -17372 -28264 -17308
rect -28200 -17372 -28180 -17308
rect -33552 -17388 -28180 -17372
rect -33552 -17452 -28264 -17388
rect -28200 -17452 -28180 -17388
rect -33552 -17468 -28180 -17452
rect -33552 -17532 -28264 -17468
rect -28200 -17532 -28180 -17468
rect -33552 -17548 -28180 -17532
rect -33552 -17612 -28264 -17548
rect -28200 -17612 -28180 -17548
rect -33552 -17628 -28180 -17612
rect -33552 -17692 -28264 -17628
rect -28200 -17692 -28180 -17628
rect -33552 -17708 -28180 -17692
rect -33552 -17772 -28264 -17708
rect -28200 -17772 -28180 -17708
rect -33552 -17788 -28180 -17772
rect -33552 -17852 -28264 -17788
rect -28200 -17852 -28180 -17788
rect -33552 -17868 -28180 -17852
rect -33552 -17932 -28264 -17868
rect -28200 -17932 -28180 -17868
rect -33552 -17948 -28180 -17932
rect -33552 -18012 -28264 -17948
rect -28200 -18012 -28180 -17948
rect -33552 -18028 -28180 -18012
rect -33552 -18092 -28264 -18028
rect -28200 -18092 -28180 -18028
rect -33552 -18108 -28180 -18092
rect -33552 -18172 -28264 -18108
rect -28200 -18172 -28180 -18108
rect -33552 -18188 -28180 -18172
rect -33552 -18252 -28264 -18188
rect -28200 -18252 -28180 -18188
rect -33552 -18268 -28180 -18252
rect -33552 -18332 -28264 -18268
rect -28200 -18332 -28180 -18268
rect -33552 -18348 -28180 -18332
rect -33552 -18412 -28264 -18348
rect -28200 -18412 -28180 -18348
rect -33552 -18428 -28180 -18412
rect -33552 -18492 -28264 -18428
rect -28200 -18492 -28180 -18428
rect -33552 -18508 -28180 -18492
rect -33552 -18572 -28264 -18508
rect -28200 -18572 -28180 -18508
rect -33552 -18588 -28180 -18572
rect -33552 -18652 -28264 -18588
rect -28200 -18652 -28180 -18588
rect -33552 -18668 -28180 -18652
rect -33552 -18732 -28264 -18668
rect -28200 -18732 -28180 -18668
rect -33552 -18748 -28180 -18732
rect -33552 -18812 -28264 -18748
rect -28200 -18812 -28180 -18748
rect -33552 -18828 -28180 -18812
rect -33552 -18892 -28264 -18828
rect -28200 -18892 -28180 -18828
rect -33552 -18908 -28180 -18892
rect -33552 -18972 -28264 -18908
rect -28200 -18972 -28180 -18908
rect -33552 -18988 -28180 -18972
rect -33552 -19052 -28264 -18988
rect -28200 -19052 -28180 -18988
rect -33552 -19068 -28180 -19052
rect -33552 -19132 -28264 -19068
rect -28200 -19132 -28180 -19068
rect -33552 -19148 -28180 -19132
rect -33552 -19212 -28264 -19148
rect -28200 -19212 -28180 -19148
rect -33552 -19228 -28180 -19212
rect -33552 -19292 -28264 -19228
rect -28200 -19292 -28180 -19228
rect -33552 -19308 -28180 -19292
rect -33552 -19372 -28264 -19308
rect -28200 -19372 -28180 -19308
rect -33552 -19388 -28180 -19372
rect -33552 -19452 -28264 -19388
rect -28200 -19452 -28180 -19388
rect -33552 -19468 -28180 -19452
rect -33552 -19532 -28264 -19468
rect -28200 -19532 -28180 -19468
rect -33552 -19548 -28180 -19532
rect -33552 -19612 -28264 -19548
rect -28200 -19612 -28180 -19548
rect -33552 -19628 -28180 -19612
rect -33552 -19692 -28264 -19628
rect -28200 -19692 -28180 -19628
rect -33552 -19708 -28180 -19692
rect -33552 -19772 -28264 -19708
rect -28200 -19772 -28180 -19708
rect -33552 -19788 -28180 -19772
rect -33552 -19852 -28264 -19788
rect -28200 -19852 -28180 -19788
rect -33552 -19868 -28180 -19852
rect -33552 -19932 -28264 -19868
rect -28200 -19932 -28180 -19868
rect -33552 -19948 -28180 -19932
rect -33552 -20012 -28264 -19948
rect -28200 -20012 -28180 -19948
rect -33552 -20028 -28180 -20012
rect -33552 -20092 -28264 -20028
rect -28200 -20092 -28180 -20028
rect -33552 -20108 -28180 -20092
rect -33552 -20172 -28264 -20108
rect -28200 -20172 -28180 -20108
rect -33552 -20188 -28180 -20172
rect -33552 -20252 -28264 -20188
rect -28200 -20252 -28180 -20188
rect -33552 -20268 -28180 -20252
rect -33552 -20332 -28264 -20268
rect -28200 -20332 -28180 -20268
rect -33552 -20348 -28180 -20332
rect -33552 -20412 -28264 -20348
rect -28200 -20412 -28180 -20348
rect -33552 -20428 -28180 -20412
rect -33552 -20492 -28264 -20428
rect -28200 -20492 -28180 -20428
rect -33552 -20508 -28180 -20492
rect -33552 -20572 -28264 -20508
rect -28200 -20572 -28180 -20508
rect -33552 -20588 -28180 -20572
rect -33552 -20652 -28264 -20588
rect -28200 -20652 -28180 -20588
rect -33552 -20668 -28180 -20652
rect -33552 -20732 -28264 -20668
rect -28200 -20732 -28180 -20668
rect -33552 -20748 -28180 -20732
rect -33552 -20812 -28264 -20748
rect -28200 -20812 -28180 -20748
rect -33552 -20828 -28180 -20812
rect -33552 -20892 -28264 -20828
rect -28200 -20892 -28180 -20828
rect -33552 -20908 -28180 -20892
rect -33552 -20972 -28264 -20908
rect -28200 -20972 -28180 -20908
rect -33552 -20988 -28180 -20972
rect -33552 -21052 -28264 -20988
rect -28200 -21052 -28180 -20988
rect -33552 -21068 -28180 -21052
rect -33552 -21132 -28264 -21068
rect -28200 -21132 -28180 -21068
rect -33552 -21160 -28180 -21132
rect -27940 -16108 -22568 -16080
rect -27940 -16172 -22652 -16108
rect -22588 -16172 -22568 -16108
rect -27940 -16188 -22568 -16172
rect -27940 -16252 -22652 -16188
rect -22588 -16252 -22568 -16188
rect -27940 -16268 -22568 -16252
rect -27940 -16332 -22652 -16268
rect -22588 -16332 -22568 -16268
rect -27940 -16348 -22568 -16332
rect -27940 -16412 -22652 -16348
rect -22588 -16412 -22568 -16348
rect -27940 -16428 -22568 -16412
rect -27940 -16492 -22652 -16428
rect -22588 -16492 -22568 -16428
rect -27940 -16508 -22568 -16492
rect -27940 -16572 -22652 -16508
rect -22588 -16572 -22568 -16508
rect -27940 -16588 -22568 -16572
rect -27940 -16652 -22652 -16588
rect -22588 -16652 -22568 -16588
rect -27940 -16668 -22568 -16652
rect -27940 -16732 -22652 -16668
rect -22588 -16732 -22568 -16668
rect -27940 -16748 -22568 -16732
rect -27940 -16812 -22652 -16748
rect -22588 -16812 -22568 -16748
rect -27940 -16828 -22568 -16812
rect -27940 -16892 -22652 -16828
rect -22588 -16892 -22568 -16828
rect -27940 -16908 -22568 -16892
rect -27940 -16972 -22652 -16908
rect -22588 -16972 -22568 -16908
rect -27940 -16988 -22568 -16972
rect -27940 -17052 -22652 -16988
rect -22588 -17052 -22568 -16988
rect -27940 -17068 -22568 -17052
rect -27940 -17132 -22652 -17068
rect -22588 -17132 -22568 -17068
rect -27940 -17148 -22568 -17132
rect -27940 -17212 -22652 -17148
rect -22588 -17212 -22568 -17148
rect -27940 -17228 -22568 -17212
rect -27940 -17292 -22652 -17228
rect -22588 -17292 -22568 -17228
rect -27940 -17308 -22568 -17292
rect -27940 -17372 -22652 -17308
rect -22588 -17372 -22568 -17308
rect -27940 -17388 -22568 -17372
rect -27940 -17452 -22652 -17388
rect -22588 -17452 -22568 -17388
rect -27940 -17468 -22568 -17452
rect -27940 -17532 -22652 -17468
rect -22588 -17532 -22568 -17468
rect -27940 -17548 -22568 -17532
rect -27940 -17612 -22652 -17548
rect -22588 -17612 -22568 -17548
rect -27940 -17628 -22568 -17612
rect -27940 -17692 -22652 -17628
rect -22588 -17692 -22568 -17628
rect -27940 -17708 -22568 -17692
rect -27940 -17772 -22652 -17708
rect -22588 -17772 -22568 -17708
rect -27940 -17788 -22568 -17772
rect -27940 -17852 -22652 -17788
rect -22588 -17852 -22568 -17788
rect -27940 -17868 -22568 -17852
rect -27940 -17932 -22652 -17868
rect -22588 -17932 -22568 -17868
rect -27940 -17948 -22568 -17932
rect -27940 -18012 -22652 -17948
rect -22588 -18012 -22568 -17948
rect -27940 -18028 -22568 -18012
rect -27940 -18092 -22652 -18028
rect -22588 -18092 -22568 -18028
rect -27940 -18108 -22568 -18092
rect -27940 -18172 -22652 -18108
rect -22588 -18172 -22568 -18108
rect -27940 -18188 -22568 -18172
rect -27940 -18252 -22652 -18188
rect -22588 -18252 -22568 -18188
rect -27940 -18268 -22568 -18252
rect -27940 -18332 -22652 -18268
rect -22588 -18332 -22568 -18268
rect -27940 -18348 -22568 -18332
rect -27940 -18412 -22652 -18348
rect -22588 -18412 -22568 -18348
rect -27940 -18428 -22568 -18412
rect -27940 -18492 -22652 -18428
rect -22588 -18492 -22568 -18428
rect -27940 -18508 -22568 -18492
rect -27940 -18572 -22652 -18508
rect -22588 -18572 -22568 -18508
rect -27940 -18588 -22568 -18572
rect -27940 -18652 -22652 -18588
rect -22588 -18652 -22568 -18588
rect -27940 -18668 -22568 -18652
rect -27940 -18732 -22652 -18668
rect -22588 -18732 -22568 -18668
rect -27940 -18748 -22568 -18732
rect -27940 -18812 -22652 -18748
rect -22588 -18812 -22568 -18748
rect -27940 -18828 -22568 -18812
rect -27940 -18892 -22652 -18828
rect -22588 -18892 -22568 -18828
rect -27940 -18908 -22568 -18892
rect -27940 -18972 -22652 -18908
rect -22588 -18972 -22568 -18908
rect -27940 -18988 -22568 -18972
rect -27940 -19052 -22652 -18988
rect -22588 -19052 -22568 -18988
rect -27940 -19068 -22568 -19052
rect -27940 -19132 -22652 -19068
rect -22588 -19132 -22568 -19068
rect -27940 -19148 -22568 -19132
rect -27940 -19212 -22652 -19148
rect -22588 -19212 -22568 -19148
rect -27940 -19228 -22568 -19212
rect -27940 -19292 -22652 -19228
rect -22588 -19292 -22568 -19228
rect -27940 -19308 -22568 -19292
rect -27940 -19372 -22652 -19308
rect -22588 -19372 -22568 -19308
rect -27940 -19388 -22568 -19372
rect -27940 -19452 -22652 -19388
rect -22588 -19452 -22568 -19388
rect -27940 -19468 -22568 -19452
rect -27940 -19532 -22652 -19468
rect -22588 -19532 -22568 -19468
rect -27940 -19548 -22568 -19532
rect -27940 -19612 -22652 -19548
rect -22588 -19612 -22568 -19548
rect -27940 -19628 -22568 -19612
rect -27940 -19692 -22652 -19628
rect -22588 -19692 -22568 -19628
rect -27940 -19708 -22568 -19692
rect -27940 -19772 -22652 -19708
rect -22588 -19772 -22568 -19708
rect -27940 -19788 -22568 -19772
rect -27940 -19852 -22652 -19788
rect -22588 -19852 -22568 -19788
rect -27940 -19868 -22568 -19852
rect -27940 -19932 -22652 -19868
rect -22588 -19932 -22568 -19868
rect -27940 -19948 -22568 -19932
rect -27940 -20012 -22652 -19948
rect -22588 -20012 -22568 -19948
rect -27940 -20028 -22568 -20012
rect -27940 -20092 -22652 -20028
rect -22588 -20092 -22568 -20028
rect -27940 -20108 -22568 -20092
rect -27940 -20172 -22652 -20108
rect -22588 -20172 -22568 -20108
rect -27940 -20188 -22568 -20172
rect -27940 -20252 -22652 -20188
rect -22588 -20252 -22568 -20188
rect -27940 -20268 -22568 -20252
rect -27940 -20332 -22652 -20268
rect -22588 -20332 -22568 -20268
rect -27940 -20348 -22568 -20332
rect -27940 -20412 -22652 -20348
rect -22588 -20412 -22568 -20348
rect -27940 -20428 -22568 -20412
rect -27940 -20492 -22652 -20428
rect -22588 -20492 -22568 -20428
rect -27940 -20508 -22568 -20492
rect -27940 -20572 -22652 -20508
rect -22588 -20572 -22568 -20508
rect -27940 -20588 -22568 -20572
rect -27940 -20652 -22652 -20588
rect -22588 -20652 -22568 -20588
rect -27940 -20668 -22568 -20652
rect -27940 -20732 -22652 -20668
rect -22588 -20732 -22568 -20668
rect -27940 -20748 -22568 -20732
rect -27940 -20812 -22652 -20748
rect -22588 -20812 -22568 -20748
rect -27940 -20828 -22568 -20812
rect -27940 -20892 -22652 -20828
rect -22588 -20892 -22568 -20828
rect -27940 -20908 -22568 -20892
rect -27940 -20972 -22652 -20908
rect -22588 -20972 -22568 -20908
rect -27940 -20988 -22568 -20972
rect -27940 -21052 -22652 -20988
rect -22588 -21052 -22568 -20988
rect -27940 -21068 -22568 -21052
rect -27940 -21132 -22652 -21068
rect -22588 -21132 -22568 -21068
rect -27940 -21160 -22568 -21132
rect -22328 -16108 -16956 -16080
rect -22328 -16172 -17040 -16108
rect -16976 -16172 -16956 -16108
rect -22328 -16188 -16956 -16172
rect -22328 -16252 -17040 -16188
rect -16976 -16252 -16956 -16188
rect -22328 -16268 -16956 -16252
rect -22328 -16332 -17040 -16268
rect -16976 -16332 -16956 -16268
rect -22328 -16348 -16956 -16332
rect -22328 -16412 -17040 -16348
rect -16976 -16412 -16956 -16348
rect -22328 -16428 -16956 -16412
rect -22328 -16492 -17040 -16428
rect -16976 -16492 -16956 -16428
rect -22328 -16508 -16956 -16492
rect -22328 -16572 -17040 -16508
rect -16976 -16572 -16956 -16508
rect -22328 -16588 -16956 -16572
rect -22328 -16652 -17040 -16588
rect -16976 -16652 -16956 -16588
rect -22328 -16668 -16956 -16652
rect -22328 -16732 -17040 -16668
rect -16976 -16732 -16956 -16668
rect -22328 -16748 -16956 -16732
rect -22328 -16812 -17040 -16748
rect -16976 -16812 -16956 -16748
rect -22328 -16828 -16956 -16812
rect -22328 -16892 -17040 -16828
rect -16976 -16892 -16956 -16828
rect -22328 -16908 -16956 -16892
rect -22328 -16972 -17040 -16908
rect -16976 -16972 -16956 -16908
rect -22328 -16988 -16956 -16972
rect -22328 -17052 -17040 -16988
rect -16976 -17052 -16956 -16988
rect -22328 -17068 -16956 -17052
rect -22328 -17132 -17040 -17068
rect -16976 -17132 -16956 -17068
rect -22328 -17148 -16956 -17132
rect -22328 -17212 -17040 -17148
rect -16976 -17212 -16956 -17148
rect -22328 -17228 -16956 -17212
rect -22328 -17292 -17040 -17228
rect -16976 -17292 -16956 -17228
rect -22328 -17308 -16956 -17292
rect -22328 -17372 -17040 -17308
rect -16976 -17372 -16956 -17308
rect -22328 -17388 -16956 -17372
rect -22328 -17452 -17040 -17388
rect -16976 -17452 -16956 -17388
rect -22328 -17468 -16956 -17452
rect -22328 -17532 -17040 -17468
rect -16976 -17532 -16956 -17468
rect -22328 -17548 -16956 -17532
rect -22328 -17612 -17040 -17548
rect -16976 -17612 -16956 -17548
rect -22328 -17628 -16956 -17612
rect -22328 -17692 -17040 -17628
rect -16976 -17692 -16956 -17628
rect -22328 -17708 -16956 -17692
rect -22328 -17772 -17040 -17708
rect -16976 -17772 -16956 -17708
rect -22328 -17788 -16956 -17772
rect -22328 -17852 -17040 -17788
rect -16976 -17852 -16956 -17788
rect -22328 -17868 -16956 -17852
rect -22328 -17932 -17040 -17868
rect -16976 -17932 -16956 -17868
rect -22328 -17948 -16956 -17932
rect -22328 -18012 -17040 -17948
rect -16976 -18012 -16956 -17948
rect -22328 -18028 -16956 -18012
rect -22328 -18092 -17040 -18028
rect -16976 -18092 -16956 -18028
rect -22328 -18108 -16956 -18092
rect -22328 -18172 -17040 -18108
rect -16976 -18172 -16956 -18108
rect -22328 -18188 -16956 -18172
rect -22328 -18252 -17040 -18188
rect -16976 -18252 -16956 -18188
rect -22328 -18268 -16956 -18252
rect -22328 -18332 -17040 -18268
rect -16976 -18332 -16956 -18268
rect -22328 -18348 -16956 -18332
rect -22328 -18412 -17040 -18348
rect -16976 -18412 -16956 -18348
rect -22328 -18428 -16956 -18412
rect -22328 -18492 -17040 -18428
rect -16976 -18492 -16956 -18428
rect -22328 -18508 -16956 -18492
rect -22328 -18572 -17040 -18508
rect -16976 -18572 -16956 -18508
rect -22328 -18588 -16956 -18572
rect -22328 -18652 -17040 -18588
rect -16976 -18652 -16956 -18588
rect -22328 -18668 -16956 -18652
rect -22328 -18732 -17040 -18668
rect -16976 -18732 -16956 -18668
rect -22328 -18748 -16956 -18732
rect -22328 -18812 -17040 -18748
rect -16976 -18812 -16956 -18748
rect -22328 -18828 -16956 -18812
rect -22328 -18892 -17040 -18828
rect -16976 -18892 -16956 -18828
rect -22328 -18908 -16956 -18892
rect -22328 -18972 -17040 -18908
rect -16976 -18972 -16956 -18908
rect -22328 -18988 -16956 -18972
rect -22328 -19052 -17040 -18988
rect -16976 -19052 -16956 -18988
rect -22328 -19068 -16956 -19052
rect -22328 -19132 -17040 -19068
rect -16976 -19132 -16956 -19068
rect -22328 -19148 -16956 -19132
rect -22328 -19212 -17040 -19148
rect -16976 -19212 -16956 -19148
rect -22328 -19228 -16956 -19212
rect -22328 -19292 -17040 -19228
rect -16976 -19292 -16956 -19228
rect -22328 -19308 -16956 -19292
rect -22328 -19372 -17040 -19308
rect -16976 -19372 -16956 -19308
rect -22328 -19388 -16956 -19372
rect -22328 -19452 -17040 -19388
rect -16976 -19452 -16956 -19388
rect -22328 -19468 -16956 -19452
rect -22328 -19532 -17040 -19468
rect -16976 -19532 -16956 -19468
rect -22328 -19548 -16956 -19532
rect -22328 -19612 -17040 -19548
rect -16976 -19612 -16956 -19548
rect -22328 -19628 -16956 -19612
rect -22328 -19692 -17040 -19628
rect -16976 -19692 -16956 -19628
rect -22328 -19708 -16956 -19692
rect -22328 -19772 -17040 -19708
rect -16976 -19772 -16956 -19708
rect -22328 -19788 -16956 -19772
rect -22328 -19852 -17040 -19788
rect -16976 -19852 -16956 -19788
rect -22328 -19868 -16956 -19852
rect -22328 -19932 -17040 -19868
rect -16976 -19932 -16956 -19868
rect -22328 -19948 -16956 -19932
rect -22328 -20012 -17040 -19948
rect -16976 -20012 -16956 -19948
rect -22328 -20028 -16956 -20012
rect -22328 -20092 -17040 -20028
rect -16976 -20092 -16956 -20028
rect -22328 -20108 -16956 -20092
rect -22328 -20172 -17040 -20108
rect -16976 -20172 -16956 -20108
rect -22328 -20188 -16956 -20172
rect -22328 -20252 -17040 -20188
rect -16976 -20252 -16956 -20188
rect -22328 -20268 -16956 -20252
rect -22328 -20332 -17040 -20268
rect -16976 -20332 -16956 -20268
rect -22328 -20348 -16956 -20332
rect -22328 -20412 -17040 -20348
rect -16976 -20412 -16956 -20348
rect -22328 -20428 -16956 -20412
rect -22328 -20492 -17040 -20428
rect -16976 -20492 -16956 -20428
rect -22328 -20508 -16956 -20492
rect -22328 -20572 -17040 -20508
rect -16976 -20572 -16956 -20508
rect -22328 -20588 -16956 -20572
rect -22328 -20652 -17040 -20588
rect -16976 -20652 -16956 -20588
rect -22328 -20668 -16956 -20652
rect -22328 -20732 -17040 -20668
rect -16976 -20732 -16956 -20668
rect -22328 -20748 -16956 -20732
rect -22328 -20812 -17040 -20748
rect -16976 -20812 -16956 -20748
rect -22328 -20828 -16956 -20812
rect -22328 -20892 -17040 -20828
rect -16976 -20892 -16956 -20828
rect -22328 -20908 -16956 -20892
rect -22328 -20972 -17040 -20908
rect -16976 -20972 -16956 -20908
rect -22328 -20988 -16956 -20972
rect -22328 -21052 -17040 -20988
rect -16976 -21052 -16956 -20988
rect -22328 -21068 -16956 -21052
rect -22328 -21132 -17040 -21068
rect -16976 -21132 -16956 -21068
rect -22328 -21160 -16956 -21132
rect -16716 -16108 -11344 -16080
rect -16716 -16172 -11428 -16108
rect -11364 -16172 -11344 -16108
rect -16716 -16188 -11344 -16172
rect -16716 -16252 -11428 -16188
rect -11364 -16252 -11344 -16188
rect -16716 -16268 -11344 -16252
rect -16716 -16332 -11428 -16268
rect -11364 -16332 -11344 -16268
rect -16716 -16348 -11344 -16332
rect -16716 -16412 -11428 -16348
rect -11364 -16412 -11344 -16348
rect -16716 -16428 -11344 -16412
rect -16716 -16492 -11428 -16428
rect -11364 -16492 -11344 -16428
rect -16716 -16508 -11344 -16492
rect -16716 -16572 -11428 -16508
rect -11364 -16572 -11344 -16508
rect -16716 -16588 -11344 -16572
rect -16716 -16652 -11428 -16588
rect -11364 -16652 -11344 -16588
rect -16716 -16668 -11344 -16652
rect -16716 -16732 -11428 -16668
rect -11364 -16732 -11344 -16668
rect -16716 -16748 -11344 -16732
rect -16716 -16812 -11428 -16748
rect -11364 -16812 -11344 -16748
rect -16716 -16828 -11344 -16812
rect -16716 -16892 -11428 -16828
rect -11364 -16892 -11344 -16828
rect -16716 -16908 -11344 -16892
rect -16716 -16972 -11428 -16908
rect -11364 -16972 -11344 -16908
rect -16716 -16988 -11344 -16972
rect -16716 -17052 -11428 -16988
rect -11364 -17052 -11344 -16988
rect -16716 -17068 -11344 -17052
rect -16716 -17132 -11428 -17068
rect -11364 -17132 -11344 -17068
rect -16716 -17148 -11344 -17132
rect -16716 -17212 -11428 -17148
rect -11364 -17212 -11344 -17148
rect -16716 -17228 -11344 -17212
rect -16716 -17292 -11428 -17228
rect -11364 -17292 -11344 -17228
rect -16716 -17308 -11344 -17292
rect -16716 -17372 -11428 -17308
rect -11364 -17372 -11344 -17308
rect -16716 -17388 -11344 -17372
rect -16716 -17452 -11428 -17388
rect -11364 -17452 -11344 -17388
rect -16716 -17468 -11344 -17452
rect -16716 -17532 -11428 -17468
rect -11364 -17532 -11344 -17468
rect -16716 -17548 -11344 -17532
rect -16716 -17612 -11428 -17548
rect -11364 -17612 -11344 -17548
rect -16716 -17628 -11344 -17612
rect -16716 -17692 -11428 -17628
rect -11364 -17692 -11344 -17628
rect -16716 -17708 -11344 -17692
rect -16716 -17772 -11428 -17708
rect -11364 -17772 -11344 -17708
rect -16716 -17788 -11344 -17772
rect -16716 -17852 -11428 -17788
rect -11364 -17852 -11344 -17788
rect -16716 -17868 -11344 -17852
rect -16716 -17932 -11428 -17868
rect -11364 -17932 -11344 -17868
rect -16716 -17948 -11344 -17932
rect -16716 -18012 -11428 -17948
rect -11364 -18012 -11344 -17948
rect -16716 -18028 -11344 -18012
rect -16716 -18092 -11428 -18028
rect -11364 -18092 -11344 -18028
rect -16716 -18108 -11344 -18092
rect -16716 -18172 -11428 -18108
rect -11364 -18172 -11344 -18108
rect -16716 -18188 -11344 -18172
rect -16716 -18252 -11428 -18188
rect -11364 -18252 -11344 -18188
rect -16716 -18268 -11344 -18252
rect -16716 -18332 -11428 -18268
rect -11364 -18332 -11344 -18268
rect -16716 -18348 -11344 -18332
rect -16716 -18412 -11428 -18348
rect -11364 -18412 -11344 -18348
rect -16716 -18428 -11344 -18412
rect -16716 -18492 -11428 -18428
rect -11364 -18492 -11344 -18428
rect -16716 -18508 -11344 -18492
rect -16716 -18572 -11428 -18508
rect -11364 -18572 -11344 -18508
rect -16716 -18588 -11344 -18572
rect -16716 -18652 -11428 -18588
rect -11364 -18652 -11344 -18588
rect -16716 -18668 -11344 -18652
rect -16716 -18732 -11428 -18668
rect -11364 -18732 -11344 -18668
rect -16716 -18748 -11344 -18732
rect -16716 -18812 -11428 -18748
rect -11364 -18812 -11344 -18748
rect -16716 -18828 -11344 -18812
rect -16716 -18892 -11428 -18828
rect -11364 -18892 -11344 -18828
rect -16716 -18908 -11344 -18892
rect -16716 -18972 -11428 -18908
rect -11364 -18972 -11344 -18908
rect -16716 -18988 -11344 -18972
rect -16716 -19052 -11428 -18988
rect -11364 -19052 -11344 -18988
rect -16716 -19068 -11344 -19052
rect -16716 -19132 -11428 -19068
rect -11364 -19132 -11344 -19068
rect -16716 -19148 -11344 -19132
rect -16716 -19212 -11428 -19148
rect -11364 -19212 -11344 -19148
rect -16716 -19228 -11344 -19212
rect -16716 -19292 -11428 -19228
rect -11364 -19292 -11344 -19228
rect -16716 -19308 -11344 -19292
rect -16716 -19372 -11428 -19308
rect -11364 -19372 -11344 -19308
rect -16716 -19388 -11344 -19372
rect -16716 -19452 -11428 -19388
rect -11364 -19452 -11344 -19388
rect -16716 -19468 -11344 -19452
rect -16716 -19532 -11428 -19468
rect -11364 -19532 -11344 -19468
rect -16716 -19548 -11344 -19532
rect -16716 -19612 -11428 -19548
rect -11364 -19612 -11344 -19548
rect -16716 -19628 -11344 -19612
rect -16716 -19692 -11428 -19628
rect -11364 -19692 -11344 -19628
rect -16716 -19708 -11344 -19692
rect -16716 -19772 -11428 -19708
rect -11364 -19772 -11344 -19708
rect -16716 -19788 -11344 -19772
rect -16716 -19852 -11428 -19788
rect -11364 -19852 -11344 -19788
rect -16716 -19868 -11344 -19852
rect -16716 -19932 -11428 -19868
rect -11364 -19932 -11344 -19868
rect -16716 -19948 -11344 -19932
rect -16716 -20012 -11428 -19948
rect -11364 -20012 -11344 -19948
rect -16716 -20028 -11344 -20012
rect -16716 -20092 -11428 -20028
rect -11364 -20092 -11344 -20028
rect -16716 -20108 -11344 -20092
rect -16716 -20172 -11428 -20108
rect -11364 -20172 -11344 -20108
rect -16716 -20188 -11344 -20172
rect -16716 -20252 -11428 -20188
rect -11364 -20252 -11344 -20188
rect -16716 -20268 -11344 -20252
rect -16716 -20332 -11428 -20268
rect -11364 -20332 -11344 -20268
rect -16716 -20348 -11344 -20332
rect -16716 -20412 -11428 -20348
rect -11364 -20412 -11344 -20348
rect -16716 -20428 -11344 -20412
rect -16716 -20492 -11428 -20428
rect -11364 -20492 -11344 -20428
rect -16716 -20508 -11344 -20492
rect -16716 -20572 -11428 -20508
rect -11364 -20572 -11344 -20508
rect -16716 -20588 -11344 -20572
rect -16716 -20652 -11428 -20588
rect -11364 -20652 -11344 -20588
rect -16716 -20668 -11344 -20652
rect -16716 -20732 -11428 -20668
rect -11364 -20732 -11344 -20668
rect -16716 -20748 -11344 -20732
rect -16716 -20812 -11428 -20748
rect -11364 -20812 -11344 -20748
rect -16716 -20828 -11344 -20812
rect -16716 -20892 -11428 -20828
rect -11364 -20892 -11344 -20828
rect -16716 -20908 -11344 -20892
rect -16716 -20972 -11428 -20908
rect -11364 -20972 -11344 -20908
rect -16716 -20988 -11344 -20972
rect -16716 -21052 -11428 -20988
rect -11364 -21052 -11344 -20988
rect -16716 -21068 -11344 -21052
rect -16716 -21132 -11428 -21068
rect -11364 -21132 -11344 -21068
rect -16716 -21160 -11344 -21132
rect -11104 -16108 -5732 -16080
rect -11104 -16172 -5816 -16108
rect -5752 -16172 -5732 -16108
rect -11104 -16188 -5732 -16172
rect -11104 -16252 -5816 -16188
rect -5752 -16252 -5732 -16188
rect -11104 -16268 -5732 -16252
rect -11104 -16332 -5816 -16268
rect -5752 -16332 -5732 -16268
rect -11104 -16348 -5732 -16332
rect -11104 -16412 -5816 -16348
rect -5752 -16412 -5732 -16348
rect -11104 -16428 -5732 -16412
rect -11104 -16492 -5816 -16428
rect -5752 -16492 -5732 -16428
rect -11104 -16508 -5732 -16492
rect -11104 -16572 -5816 -16508
rect -5752 -16572 -5732 -16508
rect -11104 -16588 -5732 -16572
rect -11104 -16652 -5816 -16588
rect -5752 -16652 -5732 -16588
rect -11104 -16668 -5732 -16652
rect -11104 -16732 -5816 -16668
rect -5752 -16732 -5732 -16668
rect -11104 -16748 -5732 -16732
rect -11104 -16812 -5816 -16748
rect -5752 -16812 -5732 -16748
rect -11104 -16828 -5732 -16812
rect -11104 -16892 -5816 -16828
rect -5752 -16892 -5732 -16828
rect -11104 -16908 -5732 -16892
rect -11104 -16972 -5816 -16908
rect -5752 -16972 -5732 -16908
rect -11104 -16988 -5732 -16972
rect -11104 -17052 -5816 -16988
rect -5752 -17052 -5732 -16988
rect -11104 -17068 -5732 -17052
rect -11104 -17132 -5816 -17068
rect -5752 -17132 -5732 -17068
rect -11104 -17148 -5732 -17132
rect -11104 -17212 -5816 -17148
rect -5752 -17212 -5732 -17148
rect -11104 -17228 -5732 -17212
rect -11104 -17292 -5816 -17228
rect -5752 -17292 -5732 -17228
rect -11104 -17308 -5732 -17292
rect -11104 -17372 -5816 -17308
rect -5752 -17372 -5732 -17308
rect -11104 -17388 -5732 -17372
rect -11104 -17452 -5816 -17388
rect -5752 -17452 -5732 -17388
rect -11104 -17468 -5732 -17452
rect -11104 -17532 -5816 -17468
rect -5752 -17532 -5732 -17468
rect -11104 -17548 -5732 -17532
rect -11104 -17612 -5816 -17548
rect -5752 -17612 -5732 -17548
rect -11104 -17628 -5732 -17612
rect -11104 -17692 -5816 -17628
rect -5752 -17692 -5732 -17628
rect -11104 -17708 -5732 -17692
rect -11104 -17772 -5816 -17708
rect -5752 -17772 -5732 -17708
rect -11104 -17788 -5732 -17772
rect -11104 -17852 -5816 -17788
rect -5752 -17852 -5732 -17788
rect -11104 -17868 -5732 -17852
rect -11104 -17932 -5816 -17868
rect -5752 -17932 -5732 -17868
rect -11104 -17948 -5732 -17932
rect -11104 -18012 -5816 -17948
rect -5752 -18012 -5732 -17948
rect -11104 -18028 -5732 -18012
rect -11104 -18092 -5816 -18028
rect -5752 -18092 -5732 -18028
rect -11104 -18108 -5732 -18092
rect -11104 -18172 -5816 -18108
rect -5752 -18172 -5732 -18108
rect -11104 -18188 -5732 -18172
rect -11104 -18252 -5816 -18188
rect -5752 -18252 -5732 -18188
rect -11104 -18268 -5732 -18252
rect -11104 -18332 -5816 -18268
rect -5752 -18332 -5732 -18268
rect -11104 -18348 -5732 -18332
rect -11104 -18412 -5816 -18348
rect -5752 -18412 -5732 -18348
rect -11104 -18428 -5732 -18412
rect -11104 -18492 -5816 -18428
rect -5752 -18492 -5732 -18428
rect -11104 -18508 -5732 -18492
rect -11104 -18572 -5816 -18508
rect -5752 -18572 -5732 -18508
rect -11104 -18588 -5732 -18572
rect -11104 -18652 -5816 -18588
rect -5752 -18652 -5732 -18588
rect -11104 -18668 -5732 -18652
rect -11104 -18732 -5816 -18668
rect -5752 -18732 -5732 -18668
rect -11104 -18748 -5732 -18732
rect -11104 -18812 -5816 -18748
rect -5752 -18812 -5732 -18748
rect -11104 -18828 -5732 -18812
rect -11104 -18892 -5816 -18828
rect -5752 -18892 -5732 -18828
rect -11104 -18908 -5732 -18892
rect -11104 -18972 -5816 -18908
rect -5752 -18972 -5732 -18908
rect -11104 -18988 -5732 -18972
rect -11104 -19052 -5816 -18988
rect -5752 -19052 -5732 -18988
rect -11104 -19068 -5732 -19052
rect -11104 -19132 -5816 -19068
rect -5752 -19132 -5732 -19068
rect -11104 -19148 -5732 -19132
rect -11104 -19212 -5816 -19148
rect -5752 -19212 -5732 -19148
rect -11104 -19228 -5732 -19212
rect -11104 -19292 -5816 -19228
rect -5752 -19292 -5732 -19228
rect -11104 -19308 -5732 -19292
rect -11104 -19372 -5816 -19308
rect -5752 -19372 -5732 -19308
rect -11104 -19388 -5732 -19372
rect -11104 -19452 -5816 -19388
rect -5752 -19452 -5732 -19388
rect -11104 -19468 -5732 -19452
rect -11104 -19532 -5816 -19468
rect -5752 -19532 -5732 -19468
rect -11104 -19548 -5732 -19532
rect -11104 -19612 -5816 -19548
rect -5752 -19612 -5732 -19548
rect -11104 -19628 -5732 -19612
rect -11104 -19692 -5816 -19628
rect -5752 -19692 -5732 -19628
rect -11104 -19708 -5732 -19692
rect -11104 -19772 -5816 -19708
rect -5752 -19772 -5732 -19708
rect -11104 -19788 -5732 -19772
rect -11104 -19852 -5816 -19788
rect -5752 -19852 -5732 -19788
rect -11104 -19868 -5732 -19852
rect -11104 -19932 -5816 -19868
rect -5752 -19932 -5732 -19868
rect -11104 -19948 -5732 -19932
rect -11104 -20012 -5816 -19948
rect -5752 -20012 -5732 -19948
rect -11104 -20028 -5732 -20012
rect -11104 -20092 -5816 -20028
rect -5752 -20092 -5732 -20028
rect -11104 -20108 -5732 -20092
rect -11104 -20172 -5816 -20108
rect -5752 -20172 -5732 -20108
rect -11104 -20188 -5732 -20172
rect -11104 -20252 -5816 -20188
rect -5752 -20252 -5732 -20188
rect -11104 -20268 -5732 -20252
rect -11104 -20332 -5816 -20268
rect -5752 -20332 -5732 -20268
rect -11104 -20348 -5732 -20332
rect -11104 -20412 -5816 -20348
rect -5752 -20412 -5732 -20348
rect -11104 -20428 -5732 -20412
rect -11104 -20492 -5816 -20428
rect -5752 -20492 -5732 -20428
rect -11104 -20508 -5732 -20492
rect -11104 -20572 -5816 -20508
rect -5752 -20572 -5732 -20508
rect -11104 -20588 -5732 -20572
rect -11104 -20652 -5816 -20588
rect -5752 -20652 -5732 -20588
rect -11104 -20668 -5732 -20652
rect -11104 -20732 -5816 -20668
rect -5752 -20732 -5732 -20668
rect -11104 -20748 -5732 -20732
rect -11104 -20812 -5816 -20748
rect -5752 -20812 -5732 -20748
rect -11104 -20828 -5732 -20812
rect -11104 -20892 -5816 -20828
rect -5752 -20892 -5732 -20828
rect -11104 -20908 -5732 -20892
rect -11104 -20972 -5816 -20908
rect -5752 -20972 -5732 -20908
rect -11104 -20988 -5732 -20972
rect -11104 -21052 -5816 -20988
rect -5752 -21052 -5732 -20988
rect -11104 -21068 -5732 -21052
rect -11104 -21132 -5816 -21068
rect -5752 -21132 -5732 -21068
rect -11104 -21160 -5732 -21132
rect -5492 -16108 -120 -16080
rect -5492 -16172 -204 -16108
rect -140 -16172 -120 -16108
rect -5492 -16188 -120 -16172
rect -5492 -16252 -204 -16188
rect -140 -16252 -120 -16188
rect -5492 -16268 -120 -16252
rect -5492 -16332 -204 -16268
rect -140 -16332 -120 -16268
rect -5492 -16348 -120 -16332
rect -5492 -16412 -204 -16348
rect -140 -16412 -120 -16348
rect -5492 -16428 -120 -16412
rect -5492 -16492 -204 -16428
rect -140 -16492 -120 -16428
rect -5492 -16508 -120 -16492
rect -5492 -16572 -204 -16508
rect -140 -16572 -120 -16508
rect -5492 -16588 -120 -16572
rect -5492 -16652 -204 -16588
rect -140 -16652 -120 -16588
rect -5492 -16668 -120 -16652
rect -5492 -16732 -204 -16668
rect -140 -16732 -120 -16668
rect -5492 -16748 -120 -16732
rect -5492 -16812 -204 -16748
rect -140 -16812 -120 -16748
rect -5492 -16828 -120 -16812
rect -5492 -16892 -204 -16828
rect -140 -16892 -120 -16828
rect -5492 -16908 -120 -16892
rect -5492 -16972 -204 -16908
rect -140 -16972 -120 -16908
rect -5492 -16988 -120 -16972
rect -5492 -17052 -204 -16988
rect -140 -17052 -120 -16988
rect -5492 -17068 -120 -17052
rect -5492 -17132 -204 -17068
rect -140 -17132 -120 -17068
rect -5492 -17148 -120 -17132
rect -5492 -17212 -204 -17148
rect -140 -17212 -120 -17148
rect -5492 -17228 -120 -17212
rect -5492 -17292 -204 -17228
rect -140 -17292 -120 -17228
rect -5492 -17308 -120 -17292
rect -5492 -17372 -204 -17308
rect -140 -17372 -120 -17308
rect -5492 -17388 -120 -17372
rect -5492 -17452 -204 -17388
rect -140 -17452 -120 -17388
rect -5492 -17468 -120 -17452
rect -5492 -17532 -204 -17468
rect -140 -17532 -120 -17468
rect -5492 -17548 -120 -17532
rect -5492 -17612 -204 -17548
rect -140 -17612 -120 -17548
rect -5492 -17628 -120 -17612
rect -5492 -17692 -204 -17628
rect -140 -17692 -120 -17628
rect -5492 -17708 -120 -17692
rect -5492 -17772 -204 -17708
rect -140 -17772 -120 -17708
rect -5492 -17788 -120 -17772
rect -5492 -17852 -204 -17788
rect -140 -17852 -120 -17788
rect -5492 -17868 -120 -17852
rect -5492 -17932 -204 -17868
rect -140 -17932 -120 -17868
rect -5492 -17948 -120 -17932
rect -5492 -18012 -204 -17948
rect -140 -18012 -120 -17948
rect -5492 -18028 -120 -18012
rect -5492 -18092 -204 -18028
rect -140 -18092 -120 -18028
rect -5492 -18108 -120 -18092
rect -5492 -18172 -204 -18108
rect -140 -18172 -120 -18108
rect -5492 -18188 -120 -18172
rect -5492 -18252 -204 -18188
rect -140 -18252 -120 -18188
rect -5492 -18268 -120 -18252
rect -5492 -18332 -204 -18268
rect -140 -18332 -120 -18268
rect -5492 -18348 -120 -18332
rect -5492 -18412 -204 -18348
rect -140 -18412 -120 -18348
rect -5492 -18428 -120 -18412
rect -5492 -18492 -204 -18428
rect -140 -18492 -120 -18428
rect -5492 -18508 -120 -18492
rect -5492 -18572 -204 -18508
rect -140 -18572 -120 -18508
rect -5492 -18588 -120 -18572
rect -5492 -18652 -204 -18588
rect -140 -18652 -120 -18588
rect -5492 -18668 -120 -18652
rect -5492 -18732 -204 -18668
rect -140 -18732 -120 -18668
rect -5492 -18748 -120 -18732
rect -5492 -18812 -204 -18748
rect -140 -18812 -120 -18748
rect -5492 -18828 -120 -18812
rect -5492 -18892 -204 -18828
rect -140 -18892 -120 -18828
rect -5492 -18908 -120 -18892
rect -5492 -18972 -204 -18908
rect -140 -18972 -120 -18908
rect -5492 -18988 -120 -18972
rect -5492 -19052 -204 -18988
rect -140 -19052 -120 -18988
rect -5492 -19068 -120 -19052
rect -5492 -19132 -204 -19068
rect -140 -19132 -120 -19068
rect -5492 -19148 -120 -19132
rect -5492 -19212 -204 -19148
rect -140 -19212 -120 -19148
rect -5492 -19228 -120 -19212
rect -5492 -19292 -204 -19228
rect -140 -19292 -120 -19228
rect -5492 -19308 -120 -19292
rect -5492 -19372 -204 -19308
rect -140 -19372 -120 -19308
rect -5492 -19388 -120 -19372
rect -5492 -19452 -204 -19388
rect -140 -19452 -120 -19388
rect -5492 -19468 -120 -19452
rect -5492 -19532 -204 -19468
rect -140 -19532 -120 -19468
rect -5492 -19548 -120 -19532
rect -5492 -19612 -204 -19548
rect -140 -19612 -120 -19548
rect -5492 -19628 -120 -19612
rect -5492 -19692 -204 -19628
rect -140 -19692 -120 -19628
rect -5492 -19708 -120 -19692
rect -5492 -19772 -204 -19708
rect -140 -19772 -120 -19708
rect -5492 -19788 -120 -19772
rect -5492 -19852 -204 -19788
rect -140 -19852 -120 -19788
rect -5492 -19868 -120 -19852
rect -5492 -19932 -204 -19868
rect -140 -19932 -120 -19868
rect -5492 -19948 -120 -19932
rect -5492 -20012 -204 -19948
rect -140 -20012 -120 -19948
rect -5492 -20028 -120 -20012
rect -5492 -20092 -204 -20028
rect -140 -20092 -120 -20028
rect -5492 -20108 -120 -20092
rect -5492 -20172 -204 -20108
rect -140 -20172 -120 -20108
rect -5492 -20188 -120 -20172
rect -5492 -20252 -204 -20188
rect -140 -20252 -120 -20188
rect -5492 -20268 -120 -20252
rect -5492 -20332 -204 -20268
rect -140 -20332 -120 -20268
rect -5492 -20348 -120 -20332
rect -5492 -20412 -204 -20348
rect -140 -20412 -120 -20348
rect -5492 -20428 -120 -20412
rect -5492 -20492 -204 -20428
rect -140 -20492 -120 -20428
rect -5492 -20508 -120 -20492
rect -5492 -20572 -204 -20508
rect -140 -20572 -120 -20508
rect -5492 -20588 -120 -20572
rect -5492 -20652 -204 -20588
rect -140 -20652 -120 -20588
rect -5492 -20668 -120 -20652
rect -5492 -20732 -204 -20668
rect -140 -20732 -120 -20668
rect -5492 -20748 -120 -20732
rect -5492 -20812 -204 -20748
rect -140 -20812 -120 -20748
rect -5492 -20828 -120 -20812
rect -5492 -20892 -204 -20828
rect -140 -20892 -120 -20828
rect -5492 -20908 -120 -20892
rect -5492 -20972 -204 -20908
rect -140 -20972 -120 -20908
rect -5492 -20988 -120 -20972
rect -5492 -21052 -204 -20988
rect -140 -21052 -120 -20988
rect -5492 -21068 -120 -21052
rect -5492 -21132 -204 -21068
rect -140 -21132 -120 -21068
rect -5492 -21160 -120 -21132
rect 120 -16108 5492 -16080
rect 120 -16172 5408 -16108
rect 5472 -16172 5492 -16108
rect 120 -16188 5492 -16172
rect 120 -16252 5408 -16188
rect 5472 -16252 5492 -16188
rect 120 -16268 5492 -16252
rect 120 -16332 5408 -16268
rect 5472 -16332 5492 -16268
rect 120 -16348 5492 -16332
rect 120 -16412 5408 -16348
rect 5472 -16412 5492 -16348
rect 120 -16428 5492 -16412
rect 120 -16492 5408 -16428
rect 5472 -16492 5492 -16428
rect 120 -16508 5492 -16492
rect 120 -16572 5408 -16508
rect 5472 -16572 5492 -16508
rect 120 -16588 5492 -16572
rect 120 -16652 5408 -16588
rect 5472 -16652 5492 -16588
rect 120 -16668 5492 -16652
rect 120 -16732 5408 -16668
rect 5472 -16732 5492 -16668
rect 120 -16748 5492 -16732
rect 120 -16812 5408 -16748
rect 5472 -16812 5492 -16748
rect 120 -16828 5492 -16812
rect 120 -16892 5408 -16828
rect 5472 -16892 5492 -16828
rect 120 -16908 5492 -16892
rect 120 -16972 5408 -16908
rect 5472 -16972 5492 -16908
rect 120 -16988 5492 -16972
rect 120 -17052 5408 -16988
rect 5472 -17052 5492 -16988
rect 120 -17068 5492 -17052
rect 120 -17132 5408 -17068
rect 5472 -17132 5492 -17068
rect 120 -17148 5492 -17132
rect 120 -17212 5408 -17148
rect 5472 -17212 5492 -17148
rect 120 -17228 5492 -17212
rect 120 -17292 5408 -17228
rect 5472 -17292 5492 -17228
rect 120 -17308 5492 -17292
rect 120 -17372 5408 -17308
rect 5472 -17372 5492 -17308
rect 120 -17388 5492 -17372
rect 120 -17452 5408 -17388
rect 5472 -17452 5492 -17388
rect 120 -17468 5492 -17452
rect 120 -17532 5408 -17468
rect 5472 -17532 5492 -17468
rect 120 -17548 5492 -17532
rect 120 -17612 5408 -17548
rect 5472 -17612 5492 -17548
rect 120 -17628 5492 -17612
rect 120 -17692 5408 -17628
rect 5472 -17692 5492 -17628
rect 120 -17708 5492 -17692
rect 120 -17772 5408 -17708
rect 5472 -17772 5492 -17708
rect 120 -17788 5492 -17772
rect 120 -17852 5408 -17788
rect 5472 -17852 5492 -17788
rect 120 -17868 5492 -17852
rect 120 -17932 5408 -17868
rect 5472 -17932 5492 -17868
rect 120 -17948 5492 -17932
rect 120 -18012 5408 -17948
rect 5472 -18012 5492 -17948
rect 120 -18028 5492 -18012
rect 120 -18092 5408 -18028
rect 5472 -18092 5492 -18028
rect 120 -18108 5492 -18092
rect 120 -18172 5408 -18108
rect 5472 -18172 5492 -18108
rect 120 -18188 5492 -18172
rect 120 -18252 5408 -18188
rect 5472 -18252 5492 -18188
rect 120 -18268 5492 -18252
rect 120 -18332 5408 -18268
rect 5472 -18332 5492 -18268
rect 120 -18348 5492 -18332
rect 120 -18412 5408 -18348
rect 5472 -18412 5492 -18348
rect 120 -18428 5492 -18412
rect 120 -18492 5408 -18428
rect 5472 -18492 5492 -18428
rect 120 -18508 5492 -18492
rect 120 -18572 5408 -18508
rect 5472 -18572 5492 -18508
rect 120 -18588 5492 -18572
rect 120 -18652 5408 -18588
rect 5472 -18652 5492 -18588
rect 120 -18668 5492 -18652
rect 120 -18732 5408 -18668
rect 5472 -18732 5492 -18668
rect 120 -18748 5492 -18732
rect 120 -18812 5408 -18748
rect 5472 -18812 5492 -18748
rect 120 -18828 5492 -18812
rect 120 -18892 5408 -18828
rect 5472 -18892 5492 -18828
rect 120 -18908 5492 -18892
rect 120 -18972 5408 -18908
rect 5472 -18972 5492 -18908
rect 120 -18988 5492 -18972
rect 120 -19052 5408 -18988
rect 5472 -19052 5492 -18988
rect 120 -19068 5492 -19052
rect 120 -19132 5408 -19068
rect 5472 -19132 5492 -19068
rect 120 -19148 5492 -19132
rect 120 -19212 5408 -19148
rect 5472 -19212 5492 -19148
rect 120 -19228 5492 -19212
rect 120 -19292 5408 -19228
rect 5472 -19292 5492 -19228
rect 120 -19308 5492 -19292
rect 120 -19372 5408 -19308
rect 5472 -19372 5492 -19308
rect 120 -19388 5492 -19372
rect 120 -19452 5408 -19388
rect 5472 -19452 5492 -19388
rect 120 -19468 5492 -19452
rect 120 -19532 5408 -19468
rect 5472 -19532 5492 -19468
rect 120 -19548 5492 -19532
rect 120 -19612 5408 -19548
rect 5472 -19612 5492 -19548
rect 120 -19628 5492 -19612
rect 120 -19692 5408 -19628
rect 5472 -19692 5492 -19628
rect 120 -19708 5492 -19692
rect 120 -19772 5408 -19708
rect 5472 -19772 5492 -19708
rect 120 -19788 5492 -19772
rect 120 -19852 5408 -19788
rect 5472 -19852 5492 -19788
rect 120 -19868 5492 -19852
rect 120 -19932 5408 -19868
rect 5472 -19932 5492 -19868
rect 120 -19948 5492 -19932
rect 120 -20012 5408 -19948
rect 5472 -20012 5492 -19948
rect 120 -20028 5492 -20012
rect 120 -20092 5408 -20028
rect 5472 -20092 5492 -20028
rect 120 -20108 5492 -20092
rect 120 -20172 5408 -20108
rect 5472 -20172 5492 -20108
rect 120 -20188 5492 -20172
rect 120 -20252 5408 -20188
rect 5472 -20252 5492 -20188
rect 120 -20268 5492 -20252
rect 120 -20332 5408 -20268
rect 5472 -20332 5492 -20268
rect 120 -20348 5492 -20332
rect 120 -20412 5408 -20348
rect 5472 -20412 5492 -20348
rect 120 -20428 5492 -20412
rect 120 -20492 5408 -20428
rect 5472 -20492 5492 -20428
rect 120 -20508 5492 -20492
rect 120 -20572 5408 -20508
rect 5472 -20572 5492 -20508
rect 120 -20588 5492 -20572
rect 120 -20652 5408 -20588
rect 5472 -20652 5492 -20588
rect 120 -20668 5492 -20652
rect 120 -20732 5408 -20668
rect 5472 -20732 5492 -20668
rect 120 -20748 5492 -20732
rect 120 -20812 5408 -20748
rect 5472 -20812 5492 -20748
rect 120 -20828 5492 -20812
rect 120 -20892 5408 -20828
rect 5472 -20892 5492 -20828
rect 120 -20908 5492 -20892
rect 120 -20972 5408 -20908
rect 5472 -20972 5492 -20908
rect 120 -20988 5492 -20972
rect 120 -21052 5408 -20988
rect 5472 -21052 5492 -20988
rect 120 -21068 5492 -21052
rect 120 -21132 5408 -21068
rect 5472 -21132 5492 -21068
rect 120 -21160 5492 -21132
rect 5732 -16108 11104 -16080
rect 5732 -16172 11020 -16108
rect 11084 -16172 11104 -16108
rect 5732 -16188 11104 -16172
rect 5732 -16252 11020 -16188
rect 11084 -16252 11104 -16188
rect 5732 -16268 11104 -16252
rect 5732 -16332 11020 -16268
rect 11084 -16332 11104 -16268
rect 5732 -16348 11104 -16332
rect 5732 -16412 11020 -16348
rect 11084 -16412 11104 -16348
rect 5732 -16428 11104 -16412
rect 5732 -16492 11020 -16428
rect 11084 -16492 11104 -16428
rect 5732 -16508 11104 -16492
rect 5732 -16572 11020 -16508
rect 11084 -16572 11104 -16508
rect 5732 -16588 11104 -16572
rect 5732 -16652 11020 -16588
rect 11084 -16652 11104 -16588
rect 5732 -16668 11104 -16652
rect 5732 -16732 11020 -16668
rect 11084 -16732 11104 -16668
rect 5732 -16748 11104 -16732
rect 5732 -16812 11020 -16748
rect 11084 -16812 11104 -16748
rect 5732 -16828 11104 -16812
rect 5732 -16892 11020 -16828
rect 11084 -16892 11104 -16828
rect 5732 -16908 11104 -16892
rect 5732 -16972 11020 -16908
rect 11084 -16972 11104 -16908
rect 5732 -16988 11104 -16972
rect 5732 -17052 11020 -16988
rect 11084 -17052 11104 -16988
rect 5732 -17068 11104 -17052
rect 5732 -17132 11020 -17068
rect 11084 -17132 11104 -17068
rect 5732 -17148 11104 -17132
rect 5732 -17212 11020 -17148
rect 11084 -17212 11104 -17148
rect 5732 -17228 11104 -17212
rect 5732 -17292 11020 -17228
rect 11084 -17292 11104 -17228
rect 5732 -17308 11104 -17292
rect 5732 -17372 11020 -17308
rect 11084 -17372 11104 -17308
rect 5732 -17388 11104 -17372
rect 5732 -17452 11020 -17388
rect 11084 -17452 11104 -17388
rect 5732 -17468 11104 -17452
rect 5732 -17532 11020 -17468
rect 11084 -17532 11104 -17468
rect 5732 -17548 11104 -17532
rect 5732 -17612 11020 -17548
rect 11084 -17612 11104 -17548
rect 5732 -17628 11104 -17612
rect 5732 -17692 11020 -17628
rect 11084 -17692 11104 -17628
rect 5732 -17708 11104 -17692
rect 5732 -17772 11020 -17708
rect 11084 -17772 11104 -17708
rect 5732 -17788 11104 -17772
rect 5732 -17852 11020 -17788
rect 11084 -17852 11104 -17788
rect 5732 -17868 11104 -17852
rect 5732 -17932 11020 -17868
rect 11084 -17932 11104 -17868
rect 5732 -17948 11104 -17932
rect 5732 -18012 11020 -17948
rect 11084 -18012 11104 -17948
rect 5732 -18028 11104 -18012
rect 5732 -18092 11020 -18028
rect 11084 -18092 11104 -18028
rect 5732 -18108 11104 -18092
rect 5732 -18172 11020 -18108
rect 11084 -18172 11104 -18108
rect 5732 -18188 11104 -18172
rect 5732 -18252 11020 -18188
rect 11084 -18252 11104 -18188
rect 5732 -18268 11104 -18252
rect 5732 -18332 11020 -18268
rect 11084 -18332 11104 -18268
rect 5732 -18348 11104 -18332
rect 5732 -18412 11020 -18348
rect 11084 -18412 11104 -18348
rect 5732 -18428 11104 -18412
rect 5732 -18492 11020 -18428
rect 11084 -18492 11104 -18428
rect 5732 -18508 11104 -18492
rect 5732 -18572 11020 -18508
rect 11084 -18572 11104 -18508
rect 5732 -18588 11104 -18572
rect 5732 -18652 11020 -18588
rect 11084 -18652 11104 -18588
rect 5732 -18668 11104 -18652
rect 5732 -18732 11020 -18668
rect 11084 -18732 11104 -18668
rect 5732 -18748 11104 -18732
rect 5732 -18812 11020 -18748
rect 11084 -18812 11104 -18748
rect 5732 -18828 11104 -18812
rect 5732 -18892 11020 -18828
rect 11084 -18892 11104 -18828
rect 5732 -18908 11104 -18892
rect 5732 -18972 11020 -18908
rect 11084 -18972 11104 -18908
rect 5732 -18988 11104 -18972
rect 5732 -19052 11020 -18988
rect 11084 -19052 11104 -18988
rect 5732 -19068 11104 -19052
rect 5732 -19132 11020 -19068
rect 11084 -19132 11104 -19068
rect 5732 -19148 11104 -19132
rect 5732 -19212 11020 -19148
rect 11084 -19212 11104 -19148
rect 5732 -19228 11104 -19212
rect 5732 -19292 11020 -19228
rect 11084 -19292 11104 -19228
rect 5732 -19308 11104 -19292
rect 5732 -19372 11020 -19308
rect 11084 -19372 11104 -19308
rect 5732 -19388 11104 -19372
rect 5732 -19452 11020 -19388
rect 11084 -19452 11104 -19388
rect 5732 -19468 11104 -19452
rect 5732 -19532 11020 -19468
rect 11084 -19532 11104 -19468
rect 5732 -19548 11104 -19532
rect 5732 -19612 11020 -19548
rect 11084 -19612 11104 -19548
rect 5732 -19628 11104 -19612
rect 5732 -19692 11020 -19628
rect 11084 -19692 11104 -19628
rect 5732 -19708 11104 -19692
rect 5732 -19772 11020 -19708
rect 11084 -19772 11104 -19708
rect 5732 -19788 11104 -19772
rect 5732 -19852 11020 -19788
rect 11084 -19852 11104 -19788
rect 5732 -19868 11104 -19852
rect 5732 -19932 11020 -19868
rect 11084 -19932 11104 -19868
rect 5732 -19948 11104 -19932
rect 5732 -20012 11020 -19948
rect 11084 -20012 11104 -19948
rect 5732 -20028 11104 -20012
rect 5732 -20092 11020 -20028
rect 11084 -20092 11104 -20028
rect 5732 -20108 11104 -20092
rect 5732 -20172 11020 -20108
rect 11084 -20172 11104 -20108
rect 5732 -20188 11104 -20172
rect 5732 -20252 11020 -20188
rect 11084 -20252 11104 -20188
rect 5732 -20268 11104 -20252
rect 5732 -20332 11020 -20268
rect 11084 -20332 11104 -20268
rect 5732 -20348 11104 -20332
rect 5732 -20412 11020 -20348
rect 11084 -20412 11104 -20348
rect 5732 -20428 11104 -20412
rect 5732 -20492 11020 -20428
rect 11084 -20492 11104 -20428
rect 5732 -20508 11104 -20492
rect 5732 -20572 11020 -20508
rect 11084 -20572 11104 -20508
rect 5732 -20588 11104 -20572
rect 5732 -20652 11020 -20588
rect 11084 -20652 11104 -20588
rect 5732 -20668 11104 -20652
rect 5732 -20732 11020 -20668
rect 11084 -20732 11104 -20668
rect 5732 -20748 11104 -20732
rect 5732 -20812 11020 -20748
rect 11084 -20812 11104 -20748
rect 5732 -20828 11104 -20812
rect 5732 -20892 11020 -20828
rect 11084 -20892 11104 -20828
rect 5732 -20908 11104 -20892
rect 5732 -20972 11020 -20908
rect 11084 -20972 11104 -20908
rect 5732 -20988 11104 -20972
rect 5732 -21052 11020 -20988
rect 11084 -21052 11104 -20988
rect 5732 -21068 11104 -21052
rect 5732 -21132 11020 -21068
rect 11084 -21132 11104 -21068
rect 5732 -21160 11104 -21132
rect 11344 -16108 16716 -16080
rect 11344 -16172 16632 -16108
rect 16696 -16172 16716 -16108
rect 11344 -16188 16716 -16172
rect 11344 -16252 16632 -16188
rect 16696 -16252 16716 -16188
rect 11344 -16268 16716 -16252
rect 11344 -16332 16632 -16268
rect 16696 -16332 16716 -16268
rect 11344 -16348 16716 -16332
rect 11344 -16412 16632 -16348
rect 16696 -16412 16716 -16348
rect 11344 -16428 16716 -16412
rect 11344 -16492 16632 -16428
rect 16696 -16492 16716 -16428
rect 11344 -16508 16716 -16492
rect 11344 -16572 16632 -16508
rect 16696 -16572 16716 -16508
rect 11344 -16588 16716 -16572
rect 11344 -16652 16632 -16588
rect 16696 -16652 16716 -16588
rect 11344 -16668 16716 -16652
rect 11344 -16732 16632 -16668
rect 16696 -16732 16716 -16668
rect 11344 -16748 16716 -16732
rect 11344 -16812 16632 -16748
rect 16696 -16812 16716 -16748
rect 11344 -16828 16716 -16812
rect 11344 -16892 16632 -16828
rect 16696 -16892 16716 -16828
rect 11344 -16908 16716 -16892
rect 11344 -16972 16632 -16908
rect 16696 -16972 16716 -16908
rect 11344 -16988 16716 -16972
rect 11344 -17052 16632 -16988
rect 16696 -17052 16716 -16988
rect 11344 -17068 16716 -17052
rect 11344 -17132 16632 -17068
rect 16696 -17132 16716 -17068
rect 11344 -17148 16716 -17132
rect 11344 -17212 16632 -17148
rect 16696 -17212 16716 -17148
rect 11344 -17228 16716 -17212
rect 11344 -17292 16632 -17228
rect 16696 -17292 16716 -17228
rect 11344 -17308 16716 -17292
rect 11344 -17372 16632 -17308
rect 16696 -17372 16716 -17308
rect 11344 -17388 16716 -17372
rect 11344 -17452 16632 -17388
rect 16696 -17452 16716 -17388
rect 11344 -17468 16716 -17452
rect 11344 -17532 16632 -17468
rect 16696 -17532 16716 -17468
rect 11344 -17548 16716 -17532
rect 11344 -17612 16632 -17548
rect 16696 -17612 16716 -17548
rect 11344 -17628 16716 -17612
rect 11344 -17692 16632 -17628
rect 16696 -17692 16716 -17628
rect 11344 -17708 16716 -17692
rect 11344 -17772 16632 -17708
rect 16696 -17772 16716 -17708
rect 11344 -17788 16716 -17772
rect 11344 -17852 16632 -17788
rect 16696 -17852 16716 -17788
rect 11344 -17868 16716 -17852
rect 11344 -17932 16632 -17868
rect 16696 -17932 16716 -17868
rect 11344 -17948 16716 -17932
rect 11344 -18012 16632 -17948
rect 16696 -18012 16716 -17948
rect 11344 -18028 16716 -18012
rect 11344 -18092 16632 -18028
rect 16696 -18092 16716 -18028
rect 11344 -18108 16716 -18092
rect 11344 -18172 16632 -18108
rect 16696 -18172 16716 -18108
rect 11344 -18188 16716 -18172
rect 11344 -18252 16632 -18188
rect 16696 -18252 16716 -18188
rect 11344 -18268 16716 -18252
rect 11344 -18332 16632 -18268
rect 16696 -18332 16716 -18268
rect 11344 -18348 16716 -18332
rect 11344 -18412 16632 -18348
rect 16696 -18412 16716 -18348
rect 11344 -18428 16716 -18412
rect 11344 -18492 16632 -18428
rect 16696 -18492 16716 -18428
rect 11344 -18508 16716 -18492
rect 11344 -18572 16632 -18508
rect 16696 -18572 16716 -18508
rect 11344 -18588 16716 -18572
rect 11344 -18652 16632 -18588
rect 16696 -18652 16716 -18588
rect 11344 -18668 16716 -18652
rect 11344 -18732 16632 -18668
rect 16696 -18732 16716 -18668
rect 11344 -18748 16716 -18732
rect 11344 -18812 16632 -18748
rect 16696 -18812 16716 -18748
rect 11344 -18828 16716 -18812
rect 11344 -18892 16632 -18828
rect 16696 -18892 16716 -18828
rect 11344 -18908 16716 -18892
rect 11344 -18972 16632 -18908
rect 16696 -18972 16716 -18908
rect 11344 -18988 16716 -18972
rect 11344 -19052 16632 -18988
rect 16696 -19052 16716 -18988
rect 11344 -19068 16716 -19052
rect 11344 -19132 16632 -19068
rect 16696 -19132 16716 -19068
rect 11344 -19148 16716 -19132
rect 11344 -19212 16632 -19148
rect 16696 -19212 16716 -19148
rect 11344 -19228 16716 -19212
rect 11344 -19292 16632 -19228
rect 16696 -19292 16716 -19228
rect 11344 -19308 16716 -19292
rect 11344 -19372 16632 -19308
rect 16696 -19372 16716 -19308
rect 11344 -19388 16716 -19372
rect 11344 -19452 16632 -19388
rect 16696 -19452 16716 -19388
rect 11344 -19468 16716 -19452
rect 11344 -19532 16632 -19468
rect 16696 -19532 16716 -19468
rect 11344 -19548 16716 -19532
rect 11344 -19612 16632 -19548
rect 16696 -19612 16716 -19548
rect 11344 -19628 16716 -19612
rect 11344 -19692 16632 -19628
rect 16696 -19692 16716 -19628
rect 11344 -19708 16716 -19692
rect 11344 -19772 16632 -19708
rect 16696 -19772 16716 -19708
rect 11344 -19788 16716 -19772
rect 11344 -19852 16632 -19788
rect 16696 -19852 16716 -19788
rect 11344 -19868 16716 -19852
rect 11344 -19932 16632 -19868
rect 16696 -19932 16716 -19868
rect 11344 -19948 16716 -19932
rect 11344 -20012 16632 -19948
rect 16696 -20012 16716 -19948
rect 11344 -20028 16716 -20012
rect 11344 -20092 16632 -20028
rect 16696 -20092 16716 -20028
rect 11344 -20108 16716 -20092
rect 11344 -20172 16632 -20108
rect 16696 -20172 16716 -20108
rect 11344 -20188 16716 -20172
rect 11344 -20252 16632 -20188
rect 16696 -20252 16716 -20188
rect 11344 -20268 16716 -20252
rect 11344 -20332 16632 -20268
rect 16696 -20332 16716 -20268
rect 11344 -20348 16716 -20332
rect 11344 -20412 16632 -20348
rect 16696 -20412 16716 -20348
rect 11344 -20428 16716 -20412
rect 11344 -20492 16632 -20428
rect 16696 -20492 16716 -20428
rect 11344 -20508 16716 -20492
rect 11344 -20572 16632 -20508
rect 16696 -20572 16716 -20508
rect 11344 -20588 16716 -20572
rect 11344 -20652 16632 -20588
rect 16696 -20652 16716 -20588
rect 11344 -20668 16716 -20652
rect 11344 -20732 16632 -20668
rect 16696 -20732 16716 -20668
rect 11344 -20748 16716 -20732
rect 11344 -20812 16632 -20748
rect 16696 -20812 16716 -20748
rect 11344 -20828 16716 -20812
rect 11344 -20892 16632 -20828
rect 16696 -20892 16716 -20828
rect 11344 -20908 16716 -20892
rect 11344 -20972 16632 -20908
rect 16696 -20972 16716 -20908
rect 11344 -20988 16716 -20972
rect 11344 -21052 16632 -20988
rect 16696 -21052 16716 -20988
rect 11344 -21068 16716 -21052
rect 11344 -21132 16632 -21068
rect 16696 -21132 16716 -21068
rect 11344 -21160 16716 -21132
rect 16956 -16108 22328 -16080
rect 16956 -16172 22244 -16108
rect 22308 -16172 22328 -16108
rect 16956 -16188 22328 -16172
rect 16956 -16252 22244 -16188
rect 22308 -16252 22328 -16188
rect 16956 -16268 22328 -16252
rect 16956 -16332 22244 -16268
rect 22308 -16332 22328 -16268
rect 16956 -16348 22328 -16332
rect 16956 -16412 22244 -16348
rect 22308 -16412 22328 -16348
rect 16956 -16428 22328 -16412
rect 16956 -16492 22244 -16428
rect 22308 -16492 22328 -16428
rect 16956 -16508 22328 -16492
rect 16956 -16572 22244 -16508
rect 22308 -16572 22328 -16508
rect 16956 -16588 22328 -16572
rect 16956 -16652 22244 -16588
rect 22308 -16652 22328 -16588
rect 16956 -16668 22328 -16652
rect 16956 -16732 22244 -16668
rect 22308 -16732 22328 -16668
rect 16956 -16748 22328 -16732
rect 16956 -16812 22244 -16748
rect 22308 -16812 22328 -16748
rect 16956 -16828 22328 -16812
rect 16956 -16892 22244 -16828
rect 22308 -16892 22328 -16828
rect 16956 -16908 22328 -16892
rect 16956 -16972 22244 -16908
rect 22308 -16972 22328 -16908
rect 16956 -16988 22328 -16972
rect 16956 -17052 22244 -16988
rect 22308 -17052 22328 -16988
rect 16956 -17068 22328 -17052
rect 16956 -17132 22244 -17068
rect 22308 -17132 22328 -17068
rect 16956 -17148 22328 -17132
rect 16956 -17212 22244 -17148
rect 22308 -17212 22328 -17148
rect 16956 -17228 22328 -17212
rect 16956 -17292 22244 -17228
rect 22308 -17292 22328 -17228
rect 16956 -17308 22328 -17292
rect 16956 -17372 22244 -17308
rect 22308 -17372 22328 -17308
rect 16956 -17388 22328 -17372
rect 16956 -17452 22244 -17388
rect 22308 -17452 22328 -17388
rect 16956 -17468 22328 -17452
rect 16956 -17532 22244 -17468
rect 22308 -17532 22328 -17468
rect 16956 -17548 22328 -17532
rect 16956 -17612 22244 -17548
rect 22308 -17612 22328 -17548
rect 16956 -17628 22328 -17612
rect 16956 -17692 22244 -17628
rect 22308 -17692 22328 -17628
rect 16956 -17708 22328 -17692
rect 16956 -17772 22244 -17708
rect 22308 -17772 22328 -17708
rect 16956 -17788 22328 -17772
rect 16956 -17852 22244 -17788
rect 22308 -17852 22328 -17788
rect 16956 -17868 22328 -17852
rect 16956 -17932 22244 -17868
rect 22308 -17932 22328 -17868
rect 16956 -17948 22328 -17932
rect 16956 -18012 22244 -17948
rect 22308 -18012 22328 -17948
rect 16956 -18028 22328 -18012
rect 16956 -18092 22244 -18028
rect 22308 -18092 22328 -18028
rect 16956 -18108 22328 -18092
rect 16956 -18172 22244 -18108
rect 22308 -18172 22328 -18108
rect 16956 -18188 22328 -18172
rect 16956 -18252 22244 -18188
rect 22308 -18252 22328 -18188
rect 16956 -18268 22328 -18252
rect 16956 -18332 22244 -18268
rect 22308 -18332 22328 -18268
rect 16956 -18348 22328 -18332
rect 16956 -18412 22244 -18348
rect 22308 -18412 22328 -18348
rect 16956 -18428 22328 -18412
rect 16956 -18492 22244 -18428
rect 22308 -18492 22328 -18428
rect 16956 -18508 22328 -18492
rect 16956 -18572 22244 -18508
rect 22308 -18572 22328 -18508
rect 16956 -18588 22328 -18572
rect 16956 -18652 22244 -18588
rect 22308 -18652 22328 -18588
rect 16956 -18668 22328 -18652
rect 16956 -18732 22244 -18668
rect 22308 -18732 22328 -18668
rect 16956 -18748 22328 -18732
rect 16956 -18812 22244 -18748
rect 22308 -18812 22328 -18748
rect 16956 -18828 22328 -18812
rect 16956 -18892 22244 -18828
rect 22308 -18892 22328 -18828
rect 16956 -18908 22328 -18892
rect 16956 -18972 22244 -18908
rect 22308 -18972 22328 -18908
rect 16956 -18988 22328 -18972
rect 16956 -19052 22244 -18988
rect 22308 -19052 22328 -18988
rect 16956 -19068 22328 -19052
rect 16956 -19132 22244 -19068
rect 22308 -19132 22328 -19068
rect 16956 -19148 22328 -19132
rect 16956 -19212 22244 -19148
rect 22308 -19212 22328 -19148
rect 16956 -19228 22328 -19212
rect 16956 -19292 22244 -19228
rect 22308 -19292 22328 -19228
rect 16956 -19308 22328 -19292
rect 16956 -19372 22244 -19308
rect 22308 -19372 22328 -19308
rect 16956 -19388 22328 -19372
rect 16956 -19452 22244 -19388
rect 22308 -19452 22328 -19388
rect 16956 -19468 22328 -19452
rect 16956 -19532 22244 -19468
rect 22308 -19532 22328 -19468
rect 16956 -19548 22328 -19532
rect 16956 -19612 22244 -19548
rect 22308 -19612 22328 -19548
rect 16956 -19628 22328 -19612
rect 16956 -19692 22244 -19628
rect 22308 -19692 22328 -19628
rect 16956 -19708 22328 -19692
rect 16956 -19772 22244 -19708
rect 22308 -19772 22328 -19708
rect 16956 -19788 22328 -19772
rect 16956 -19852 22244 -19788
rect 22308 -19852 22328 -19788
rect 16956 -19868 22328 -19852
rect 16956 -19932 22244 -19868
rect 22308 -19932 22328 -19868
rect 16956 -19948 22328 -19932
rect 16956 -20012 22244 -19948
rect 22308 -20012 22328 -19948
rect 16956 -20028 22328 -20012
rect 16956 -20092 22244 -20028
rect 22308 -20092 22328 -20028
rect 16956 -20108 22328 -20092
rect 16956 -20172 22244 -20108
rect 22308 -20172 22328 -20108
rect 16956 -20188 22328 -20172
rect 16956 -20252 22244 -20188
rect 22308 -20252 22328 -20188
rect 16956 -20268 22328 -20252
rect 16956 -20332 22244 -20268
rect 22308 -20332 22328 -20268
rect 16956 -20348 22328 -20332
rect 16956 -20412 22244 -20348
rect 22308 -20412 22328 -20348
rect 16956 -20428 22328 -20412
rect 16956 -20492 22244 -20428
rect 22308 -20492 22328 -20428
rect 16956 -20508 22328 -20492
rect 16956 -20572 22244 -20508
rect 22308 -20572 22328 -20508
rect 16956 -20588 22328 -20572
rect 16956 -20652 22244 -20588
rect 22308 -20652 22328 -20588
rect 16956 -20668 22328 -20652
rect 16956 -20732 22244 -20668
rect 22308 -20732 22328 -20668
rect 16956 -20748 22328 -20732
rect 16956 -20812 22244 -20748
rect 22308 -20812 22328 -20748
rect 16956 -20828 22328 -20812
rect 16956 -20892 22244 -20828
rect 22308 -20892 22328 -20828
rect 16956 -20908 22328 -20892
rect 16956 -20972 22244 -20908
rect 22308 -20972 22328 -20908
rect 16956 -20988 22328 -20972
rect 16956 -21052 22244 -20988
rect 22308 -21052 22328 -20988
rect 16956 -21068 22328 -21052
rect 16956 -21132 22244 -21068
rect 22308 -21132 22328 -21068
rect 16956 -21160 22328 -21132
rect 22568 -16108 27940 -16080
rect 22568 -16172 27856 -16108
rect 27920 -16172 27940 -16108
rect 22568 -16188 27940 -16172
rect 22568 -16252 27856 -16188
rect 27920 -16252 27940 -16188
rect 22568 -16268 27940 -16252
rect 22568 -16332 27856 -16268
rect 27920 -16332 27940 -16268
rect 22568 -16348 27940 -16332
rect 22568 -16412 27856 -16348
rect 27920 -16412 27940 -16348
rect 22568 -16428 27940 -16412
rect 22568 -16492 27856 -16428
rect 27920 -16492 27940 -16428
rect 22568 -16508 27940 -16492
rect 22568 -16572 27856 -16508
rect 27920 -16572 27940 -16508
rect 22568 -16588 27940 -16572
rect 22568 -16652 27856 -16588
rect 27920 -16652 27940 -16588
rect 22568 -16668 27940 -16652
rect 22568 -16732 27856 -16668
rect 27920 -16732 27940 -16668
rect 22568 -16748 27940 -16732
rect 22568 -16812 27856 -16748
rect 27920 -16812 27940 -16748
rect 22568 -16828 27940 -16812
rect 22568 -16892 27856 -16828
rect 27920 -16892 27940 -16828
rect 22568 -16908 27940 -16892
rect 22568 -16972 27856 -16908
rect 27920 -16972 27940 -16908
rect 22568 -16988 27940 -16972
rect 22568 -17052 27856 -16988
rect 27920 -17052 27940 -16988
rect 22568 -17068 27940 -17052
rect 22568 -17132 27856 -17068
rect 27920 -17132 27940 -17068
rect 22568 -17148 27940 -17132
rect 22568 -17212 27856 -17148
rect 27920 -17212 27940 -17148
rect 22568 -17228 27940 -17212
rect 22568 -17292 27856 -17228
rect 27920 -17292 27940 -17228
rect 22568 -17308 27940 -17292
rect 22568 -17372 27856 -17308
rect 27920 -17372 27940 -17308
rect 22568 -17388 27940 -17372
rect 22568 -17452 27856 -17388
rect 27920 -17452 27940 -17388
rect 22568 -17468 27940 -17452
rect 22568 -17532 27856 -17468
rect 27920 -17532 27940 -17468
rect 22568 -17548 27940 -17532
rect 22568 -17612 27856 -17548
rect 27920 -17612 27940 -17548
rect 22568 -17628 27940 -17612
rect 22568 -17692 27856 -17628
rect 27920 -17692 27940 -17628
rect 22568 -17708 27940 -17692
rect 22568 -17772 27856 -17708
rect 27920 -17772 27940 -17708
rect 22568 -17788 27940 -17772
rect 22568 -17852 27856 -17788
rect 27920 -17852 27940 -17788
rect 22568 -17868 27940 -17852
rect 22568 -17932 27856 -17868
rect 27920 -17932 27940 -17868
rect 22568 -17948 27940 -17932
rect 22568 -18012 27856 -17948
rect 27920 -18012 27940 -17948
rect 22568 -18028 27940 -18012
rect 22568 -18092 27856 -18028
rect 27920 -18092 27940 -18028
rect 22568 -18108 27940 -18092
rect 22568 -18172 27856 -18108
rect 27920 -18172 27940 -18108
rect 22568 -18188 27940 -18172
rect 22568 -18252 27856 -18188
rect 27920 -18252 27940 -18188
rect 22568 -18268 27940 -18252
rect 22568 -18332 27856 -18268
rect 27920 -18332 27940 -18268
rect 22568 -18348 27940 -18332
rect 22568 -18412 27856 -18348
rect 27920 -18412 27940 -18348
rect 22568 -18428 27940 -18412
rect 22568 -18492 27856 -18428
rect 27920 -18492 27940 -18428
rect 22568 -18508 27940 -18492
rect 22568 -18572 27856 -18508
rect 27920 -18572 27940 -18508
rect 22568 -18588 27940 -18572
rect 22568 -18652 27856 -18588
rect 27920 -18652 27940 -18588
rect 22568 -18668 27940 -18652
rect 22568 -18732 27856 -18668
rect 27920 -18732 27940 -18668
rect 22568 -18748 27940 -18732
rect 22568 -18812 27856 -18748
rect 27920 -18812 27940 -18748
rect 22568 -18828 27940 -18812
rect 22568 -18892 27856 -18828
rect 27920 -18892 27940 -18828
rect 22568 -18908 27940 -18892
rect 22568 -18972 27856 -18908
rect 27920 -18972 27940 -18908
rect 22568 -18988 27940 -18972
rect 22568 -19052 27856 -18988
rect 27920 -19052 27940 -18988
rect 22568 -19068 27940 -19052
rect 22568 -19132 27856 -19068
rect 27920 -19132 27940 -19068
rect 22568 -19148 27940 -19132
rect 22568 -19212 27856 -19148
rect 27920 -19212 27940 -19148
rect 22568 -19228 27940 -19212
rect 22568 -19292 27856 -19228
rect 27920 -19292 27940 -19228
rect 22568 -19308 27940 -19292
rect 22568 -19372 27856 -19308
rect 27920 -19372 27940 -19308
rect 22568 -19388 27940 -19372
rect 22568 -19452 27856 -19388
rect 27920 -19452 27940 -19388
rect 22568 -19468 27940 -19452
rect 22568 -19532 27856 -19468
rect 27920 -19532 27940 -19468
rect 22568 -19548 27940 -19532
rect 22568 -19612 27856 -19548
rect 27920 -19612 27940 -19548
rect 22568 -19628 27940 -19612
rect 22568 -19692 27856 -19628
rect 27920 -19692 27940 -19628
rect 22568 -19708 27940 -19692
rect 22568 -19772 27856 -19708
rect 27920 -19772 27940 -19708
rect 22568 -19788 27940 -19772
rect 22568 -19852 27856 -19788
rect 27920 -19852 27940 -19788
rect 22568 -19868 27940 -19852
rect 22568 -19932 27856 -19868
rect 27920 -19932 27940 -19868
rect 22568 -19948 27940 -19932
rect 22568 -20012 27856 -19948
rect 27920 -20012 27940 -19948
rect 22568 -20028 27940 -20012
rect 22568 -20092 27856 -20028
rect 27920 -20092 27940 -20028
rect 22568 -20108 27940 -20092
rect 22568 -20172 27856 -20108
rect 27920 -20172 27940 -20108
rect 22568 -20188 27940 -20172
rect 22568 -20252 27856 -20188
rect 27920 -20252 27940 -20188
rect 22568 -20268 27940 -20252
rect 22568 -20332 27856 -20268
rect 27920 -20332 27940 -20268
rect 22568 -20348 27940 -20332
rect 22568 -20412 27856 -20348
rect 27920 -20412 27940 -20348
rect 22568 -20428 27940 -20412
rect 22568 -20492 27856 -20428
rect 27920 -20492 27940 -20428
rect 22568 -20508 27940 -20492
rect 22568 -20572 27856 -20508
rect 27920 -20572 27940 -20508
rect 22568 -20588 27940 -20572
rect 22568 -20652 27856 -20588
rect 27920 -20652 27940 -20588
rect 22568 -20668 27940 -20652
rect 22568 -20732 27856 -20668
rect 27920 -20732 27940 -20668
rect 22568 -20748 27940 -20732
rect 22568 -20812 27856 -20748
rect 27920 -20812 27940 -20748
rect 22568 -20828 27940 -20812
rect 22568 -20892 27856 -20828
rect 27920 -20892 27940 -20828
rect 22568 -20908 27940 -20892
rect 22568 -20972 27856 -20908
rect 27920 -20972 27940 -20908
rect 22568 -20988 27940 -20972
rect 22568 -21052 27856 -20988
rect 27920 -21052 27940 -20988
rect 22568 -21068 27940 -21052
rect 22568 -21132 27856 -21068
rect 27920 -21132 27940 -21068
rect 22568 -21160 27940 -21132
rect 28180 -16108 33552 -16080
rect 28180 -16172 33468 -16108
rect 33532 -16172 33552 -16108
rect 28180 -16188 33552 -16172
rect 28180 -16252 33468 -16188
rect 33532 -16252 33552 -16188
rect 28180 -16268 33552 -16252
rect 28180 -16332 33468 -16268
rect 33532 -16332 33552 -16268
rect 28180 -16348 33552 -16332
rect 28180 -16412 33468 -16348
rect 33532 -16412 33552 -16348
rect 28180 -16428 33552 -16412
rect 28180 -16492 33468 -16428
rect 33532 -16492 33552 -16428
rect 28180 -16508 33552 -16492
rect 28180 -16572 33468 -16508
rect 33532 -16572 33552 -16508
rect 28180 -16588 33552 -16572
rect 28180 -16652 33468 -16588
rect 33532 -16652 33552 -16588
rect 28180 -16668 33552 -16652
rect 28180 -16732 33468 -16668
rect 33532 -16732 33552 -16668
rect 28180 -16748 33552 -16732
rect 28180 -16812 33468 -16748
rect 33532 -16812 33552 -16748
rect 28180 -16828 33552 -16812
rect 28180 -16892 33468 -16828
rect 33532 -16892 33552 -16828
rect 28180 -16908 33552 -16892
rect 28180 -16972 33468 -16908
rect 33532 -16972 33552 -16908
rect 28180 -16988 33552 -16972
rect 28180 -17052 33468 -16988
rect 33532 -17052 33552 -16988
rect 28180 -17068 33552 -17052
rect 28180 -17132 33468 -17068
rect 33532 -17132 33552 -17068
rect 28180 -17148 33552 -17132
rect 28180 -17212 33468 -17148
rect 33532 -17212 33552 -17148
rect 28180 -17228 33552 -17212
rect 28180 -17292 33468 -17228
rect 33532 -17292 33552 -17228
rect 28180 -17308 33552 -17292
rect 28180 -17372 33468 -17308
rect 33532 -17372 33552 -17308
rect 28180 -17388 33552 -17372
rect 28180 -17452 33468 -17388
rect 33532 -17452 33552 -17388
rect 28180 -17468 33552 -17452
rect 28180 -17532 33468 -17468
rect 33532 -17532 33552 -17468
rect 28180 -17548 33552 -17532
rect 28180 -17612 33468 -17548
rect 33532 -17612 33552 -17548
rect 28180 -17628 33552 -17612
rect 28180 -17692 33468 -17628
rect 33532 -17692 33552 -17628
rect 28180 -17708 33552 -17692
rect 28180 -17772 33468 -17708
rect 33532 -17772 33552 -17708
rect 28180 -17788 33552 -17772
rect 28180 -17852 33468 -17788
rect 33532 -17852 33552 -17788
rect 28180 -17868 33552 -17852
rect 28180 -17932 33468 -17868
rect 33532 -17932 33552 -17868
rect 28180 -17948 33552 -17932
rect 28180 -18012 33468 -17948
rect 33532 -18012 33552 -17948
rect 28180 -18028 33552 -18012
rect 28180 -18092 33468 -18028
rect 33532 -18092 33552 -18028
rect 28180 -18108 33552 -18092
rect 28180 -18172 33468 -18108
rect 33532 -18172 33552 -18108
rect 28180 -18188 33552 -18172
rect 28180 -18252 33468 -18188
rect 33532 -18252 33552 -18188
rect 28180 -18268 33552 -18252
rect 28180 -18332 33468 -18268
rect 33532 -18332 33552 -18268
rect 28180 -18348 33552 -18332
rect 28180 -18412 33468 -18348
rect 33532 -18412 33552 -18348
rect 28180 -18428 33552 -18412
rect 28180 -18492 33468 -18428
rect 33532 -18492 33552 -18428
rect 28180 -18508 33552 -18492
rect 28180 -18572 33468 -18508
rect 33532 -18572 33552 -18508
rect 28180 -18588 33552 -18572
rect 28180 -18652 33468 -18588
rect 33532 -18652 33552 -18588
rect 28180 -18668 33552 -18652
rect 28180 -18732 33468 -18668
rect 33532 -18732 33552 -18668
rect 28180 -18748 33552 -18732
rect 28180 -18812 33468 -18748
rect 33532 -18812 33552 -18748
rect 28180 -18828 33552 -18812
rect 28180 -18892 33468 -18828
rect 33532 -18892 33552 -18828
rect 28180 -18908 33552 -18892
rect 28180 -18972 33468 -18908
rect 33532 -18972 33552 -18908
rect 28180 -18988 33552 -18972
rect 28180 -19052 33468 -18988
rect 33532 -19052 33552 -18988
rect 28180 -19068 33552 -19052
rect 28180 -19132 33468 -19068
rect 33532 -19132 33552 -19068
rect 28180 -19148 33552 -19132
rect 28180 -19212 33468 -19148
rect 33532 -19212 33552 -19148
rect 28180 -19228 33552 -19212
rect 28180 -19292 33468 -19228
rect 33532 -19292 33552 -19228
rect 28180 -19308 33552 -19292
rect 28180 -19372 33468 -19308
rect 33532 -19372 33552 -19308
rect 28180 -19388 33552 -19372
rect 28180 -19452 33468 -19388
rect 33532 -19452 33552 -19388
rect 28180 -19468 33552 -19452
rect 28180 -19532 33468 -19468
rect 33532 -19532 33552 -19468
rect 28180 -19548 33552 -19532
rect 28180 -19612 33468 -19548
rect 33532 -19612 33552 -19548
rect 28180 -19628 33552 -19612
rect 28180 -19692 33468 -19628
rect 33532 -19692 33552 -19628
rect 28180 -19708 33552 -19692
rect 28180 -19772 33468 -19708
rect 33532 -19772 33552 -19708
rect 28180 -19788 33552 -19772
rect 28180 -19852 33468 -19788
rect 33532 -19852 33552 -19788
rect 28180 -19868 33552 -19852
rect 28180 -19932 33468 -19868
rect 33532 -19932 33552 -19868
rect 28180 -19948 33552 -19932
rect 28180 -20012 33468 -19948
rect 33532 -20012 33552 -19948
rect 28180 -20028 33552 -20012
rect 28180 -20092 33468 -20028
rect 33532 -20092 33552 -20028
rect 28180 -20108 33552 -20092
rect 28180 -20172 33468 -20108
rect 33532 -20172 33552 -20108
rect 28180 -20188 33552 -20172
rect 28180 -20252 33468 -20188
rect 33532 -20252 33552 -20188
rect 28180 -20268 33552 -20252
rect 28180 -20332 33468 -20268
rect 33532 -20332 33552 -20268
rect 28180 -20348 33552 -20332
rect 28180 -20412 33468 -20348
rect 33532 -20412 33552 -20348
rect 28180 -20428 33552 -20412
rect 28180 -20492 33468 -20428
rect 33532 -20492 33552 -20428
rect 28180 -20508 33552 -20492
rect 28180 -20572 33468 -20508
rect 33532 -20572 33552 -20508
rect 28180 -20588 33552 -20572
rect 28180 -20652 33468 -20588
rect 33532 -20652 33552 -20588
rect 28180 -20668 33552 -20652
rect 28180 -20732 33468 -20668
rect 33532 -20732 33552 -20668
rect 28180 -20748 33552 -20732
rect 28180 -20812 33468 -20748
rect 33532 -20812 33552 -20748
rect 28180 -20828 33552 -20812
rect 28180 -20892 33468 -20828
rect 33532 -20892 33552 -20828
rect 28180 -20908 33552 -20892
rect 28180 -20972 33468 -20908
rect 33532 -20972 33552 -20908
rect 28180 -20988 33552 -20972
rect 28180 -21052 33468 -20988
rect 33532 -21052 33552 -20988
rect 28180 -21068 33552 -21052
rect 28180 -21132 33468 -21068
rect 33532 -21132 33552 -21068
rect 28180 -21160 33552 -21132
rect 33792 -16108 39164 -16080
rect 33792 -16172 39080 -16108
rect 39144 -16172 39164 -16108
rect 33792 -16188 39164 -16172
rect 33792 -16252 39080 -16188
rect 39144 -16252 39164 -16188
rect 33792 -16268 39164 -16252
rect 33792 -16332 39080 -16268
rect 39144 -16332 39164 -16268
rect 33792 -16348 39164 -16332
rect 33792 -16412 39080 -16348
rect 39144 -16412 39164 -16348
rect 33792 -16428 39164 -16412
rect 33792 -16492 39080 -16428
rect 39144 -16492 39164 -16428
rect 33792 -16508 39164 -16492
rect 33792 -16572 39080 -16508
rect 39144 -16572 39164 -16508
rect 33792 -16588 39164 -16572
rect 33792 -16652 39080 -16588
rect 39144 -16652 39164 -16588
rect 33792 -16668 39164 -16652
rect 33792 -16732 39080 -16668
rect 39144 -16732 39164 -16668
rect 33792 -16748 39164 -16732
rect 33792 -16812 39080 -16748
rect 39144 -16812 39164 -16748
rect 33792 -16828 39164 -16812
rect 33792 -16892 39080 -16828
rect 39144 -16892 39164 -16828
rect 33792 -16908 39164 -16892
rect 33792 -16972 39080 -16908
rect 39144 -16972 39164 -16908
rect 33792 -16988 39164 -16972
rect 33792 -17052 39080 -16988
rect 39144 -17052 39164 -16988
rect 33792 -17068 39164 -17052
rect 33792 -17132 39080 -17068
rect 39144 -17132 39164 -17068
rect 33792 -17148 39164 -17132
rect 33792 -17212 39080 -17148
rect 39144 -17212 39164 -17148
rect 33792 -17228 39164 -17212
rect 33792 -17292 39080 -17228
rect 39144 -17292 39164 -17228
rect 33792 -17308 39164 -17292
rect 33792 -17372 39080 -17308
rect 39144 -17372 39164 -17308
rect 33792 -17388 39164 -17372
rect 33792 -17452 39080 -17388
rect 39144 -17452 39164 -17388
rect 33792 -17468 39164 -17452
rect 33792 -17532 39080 -17468
rect 39144 -17532 39164 -17468
rect 33792 -17548 39164 -17532
rect 33792 -17612 39080 -17548
rect 39144 -17612 39164 -17548
rect 33792 -17628 39164 -17612
rect 33792 -17692 39080 -17628
rect 39144 -17692 39164 -17628
rect 33792 -17708 39164 -17692
rect 33792 -17772 39080 -17708
rect 39144 -17772 39164 -17708
rect 33792 -17788 39164 -17772
rect 33792 -17852 39080 -17788
rect 39144 -17852 39164 -17788
rect 33792 -17868 39164 -17852
rect 33792 -17932 39080 -17868
rect 39144 -17932 39164 -17868
rect 33792 -17948 39164 -17932
rect 33792 -18012 39080 -17948
rect 39144 -18012 39164 -17948
rect 33792 -18028 39164 -18012
rect 33792 -18092 39080 -18028
rect 39144 -18092 39164 -18028
rect 33792 -18108 39164 -18092
rect 33792 -18172 39080 -18108
rect 39144 -18172 39164 -18108
rect 33792 -18188 39164 -18172
rect 33792 -18252 39080 -18188
rect 39144 -18252 39164 -18188
rect 33792 -18268 39164 -18252
rect 33792 -18332 39080 -18268
rect 39144 -18332 39164 -18268
rect 33792 -18348 39164 -18332
rect 33792 -18412 39080 -18348
rect 39144 -18412 39164 -18348
rect 33792 -18428 39164 -18412
rect 33792 -18492 39080 -18428
rect 39144 -18492 39164 -18428
rect 33792 -18508 39164 -18492
rect 33792 -18572 39080 -18508
rect 39144 -18572 39164 -18508
rect 33792 -18588 39164 -18572
rect 33792 -18652 39080 -18588
rect 39144 -18652 39164 -18588
rect 33792 -18668 39164 -18652
rect 33792 -18732 39080 -18668
rect 39144 -18732 39164 -18668
rect 33792 -18748 39164 -18732
rect 33792 -18812 39080 -18748
rect 39144 -18812 39164 -18748
rect 33792 -18828 39164 -18812
rect 33792 -18892 39080 -18828
rect 39144 -18892 39164 -18828
rect 33792 -18908 39164 -18892
rect 33792 -18972 39080 -18908
rect 39144 -18972 39164 -18908
rect 33792 -18988 39164 -18972
rect 33792 -19052 39080 -18988
rect 39144 -19052 39164 -18988
rect 33792 -19068 39164 -19052
rect 33792 -19132 39080 -19068
rect 39144 -19132 39164 -19068
rect 33792 -19148 39164 -19132
rect 33792 -19212 39080 -19148
rect 39144 -19212 39164 -19148
rect 33792 -19228 39164 -19212
rect 33792 -19292 39080 -19228
rect 39144 -19292 39164 -19228
rect 33792 -19308 39164 -19292
rect 33792 -19372 39080 -19308
rect 39144 -19372 39164 -19308
rect 33792 -19388 39164 -19372
rect 33792 -19452 39080 -19388
rect 39144 -19452 39164 -19388
rect 33792 -19468 39164 -19452
rect 33792 -19532 39080 -19468
rect 39144 -19532 39164 -19468
rect 33792 -19548 39164 -19532
rect 33792 -19612 39080 -19548
rect 39144 -19612 39164 -19548
rect 33792 -19628 39164 -19612
rect 33792 -19692 39080 -19628
rect 39144 -19692 39164 -19628
rect 33792 -19708 39164 -19692
rect 33792 -19772 39080 -19708
rect 39144 -19772 39164 -19708
rect 33792 -19788 39164 -19772
rect 33792 -19852 39080 -19788
rect 39144 -19852 39164 -19788
rect 33792 -19868 39164 -19852
rect 33792 -19932 39080 -19868
rect 39144 -19932 39164 -19868
rect 33792 -19948 39164 -19932
rect 33792 -20012 39080 -19948
rect 39144 -20012 39164 -19948
rect 33792 -20028 39164 -20012
rect 33792 -20092 39080 -20028
rect 39144 -20092 39164 -20028
rect 33792 -20108 39164 -20092
rect 33792 -20172 39080 -20108
rect 39144 -20172 39164 -20108
rect 33792 -20188 39164 -20172
rect 33792 -20252 39080 -20188
rect 39144 -20252 39164 -20188
rect 33792 -20268 39164 -20252
rect 33792 -20332 39080 -20268
rect 39144 -20332 39164 -20268
rect 33792 -20348 39164 -20332
rect 33792 -20412 39080 -20348
rect 39144 -20412 39164 -20348
rect 33792 -20428 39164 -20412
rect 33792 -20492 39080 -20428
rect 39144 -20492 39164 -20428
rect 33792 -20508 39164 -20492
rect 33792 -20572 39080 -20508
rect 39144 -20572 39164 -20508
rect 33792 -20588 39164 -20572
rect 33792 -20652 39080 -20588
rect 39144 -20652 39164 -20588
rect 33792 -20668 39164 -20652
rect 33792 -20732 39080 -20668
rect 39144 -20732 39164 -20668
rect 33792 -20748 39164 -20732
rect 33792 -20812 39080 -20748
rect 39144 -20812 39164 -20748
rect 33792 -20828 39164 -20812
rect 33792 -20892 39080 -20828
rect 39144 -20892 39164 -20828
rect 33792 -20908 39164 -20892
rect 33792 -20972 39080 -20908
rect 39144 -20972 39164 -20908
rect 33792 -20988 39164 -20972
rect 33792 -21052 39080 -20988
rect 39144 -21052 39164 -20988
rect 33792 -21068 39164 -21052
rect 33792 -21132 39080 -21068
rect 39144 -21132 39164 -21068
rect 33792 -21160 39164 -21132
rect -39164 -21428 -33792 -21400
rect -39164 -21492 -33876 -21428
rect -33812 -21492 -33792 -21428
rect -39164 -21508 -33792 -21492
rect -39164 -21572 -33876 -21508
rect -33812 -21572 -33792 -21508
rect -39164 -21588 -33792 -21572
rect -39164 -21652 -33876 -21588
rect -33812 -21652 -33792 -21588
rect -39164 -21668 -33792 -21652
rect -39164 -21732 -33876 -21668
rect -33812 -21732 -33792 -21668
rect -39164 -21748 -33792 -21732
rect -39164 -21812 -33876 -21748
rect -33812 -21812 -33792 -21748
rect -39164 -21828 -33792 -21812
rect -39164 -21892 -33876 -21828
rect -33812 -21892 -33792 -21828
rect -39164 -21908 -33792 -21892
rect -39164 -21972 -33876 -21908
rect -33812 -21972 -33792 -21908
rect -39164 -21988 -33792 -21972
rect -39164 -22052 -33876 -21988
rect -33812 -22052 -33792 -21988
rect -39164 -22068 -33792 -22052
rect -39164 -22132 -33876 -22068
rect -33812 -22132 -33792 -22068
rect -39164 -22148 -33792 -22132
rect -39164 -22212 -33876 -22148
rect -33812 -22212 -33792 -22148
rect -39164 -22228 -33792 -22212
rect -39164 -22292 -33876 -22228
rect -33812 -22292 -33792 -22228
rect -39164 -22308 -33792 -22292
rect -39164 -22372 -33876 -22308
rect -33812 -22372 -33792 -22308
rect -39164 -22388 -33792 -22372
rect -39164 -22452 -33876 -22388
rect -33812 -22452 -33792 -22388
rect -39164 -22468 -33792 -22452
rect -39164 -22532 -33876 -22468
rect -33812 -22532 -33792 -22468
rect -39164 -22548 -33792 -22532
rect -39164 -22612 -33876 -22548
rect -33812 -22612 -33792 -22548
rect -39164 -22628 -33792 -22612
rect -39164 -22692 -33876 -22628
rect -33812 -22692 -33792 -22628
rect -39164 -22708 -33792 -22692
rect -39164 -22772 -33876 -22708
rect -33812 -22772 -33792 -22708
rect -39164 -22788 -33792 -22772
rect -39164 -22852 -33876 -22788
rect -33812 -22852 -33792 -22788
rect -39164 -22868 -33792 -22852
rect -39164 -22932 -33876 -22868
rect -33812 -22932 -33792 -22868
rect -39164 -22948 -33792 -22932
rect -39164 -23012 -33876 -22948
rect -33812 -23012 -33792 -22948
rect -39164 -23028 -33792 -23012
rect -39164 -23092 -33876 -23028
rect -33812 -23092 -33792 -23028
rect -39164 -23108 -33792 -23092
rect -39164 -23172 -33876 -23108
rect -33812 -23172 -33792 -23108
rect -39164 -23188 -33792 -23172
rect -39164 -23252 -33876 -23188
rect -33812 -23252 -33792 -23188
rect -39164 -23268 -33792 -23252
rect -39164 -23332 -33876 -23268
rect -33812 -23332 -33792 -23268
rect -39164 -23348 -33792 -23332
rect -39164 -23412 -33876 -23348
rect -33812 -23412 -33792 -23348
rect -39164 -23428 -33792 -23412
rect -39164 -23492 -33876 -23428
rect -33812 -23492 -33792 -23428
rect -39164 -23508 -33792 -23492
rect -39164 -23572 -33876 -23508
rect -33812 -23572 -33792 -23508
rect -39164 -23588 -33792 -23572
rect -39164 -23652 -33876 -23588
rect -33812 -23652 -33792 -23588
rect -39164 -23668 -33792 -23652
rect -39164 -23732 -33876 -23668
rect -33812 -23732 -33792 -23668
rect -39164 -23748 -33792 -23732
rect -39164 -23812 -33876 -23748
rect -33812 -23812 -33792 -23748
rect -39164 -23828 -33792 -23812
rect -39164 -23892 -33876 -23828
rect -33812 -23892 -33792 -23828
rect -39164 -23908 -33792 -23892
rect -39164 -23972 -33876 -23908
rect -33812 -23972 -33792 -23908
rect -39164 -23988 -33792 -23972
rect -39164 -24052 -33876 -23988
rect -33812 -24052 -33792 -23988
rect -39164 -24068 -33792 -24052
rect -39164 -24132 -33876 -24068
rect -33812 -24132 -33792 -24068
rect -39164 -24148 -33792 -24132
rect -39164 -24212 -33876 -24148
rect -33812 -24212 -33792 -24148
rect -39164 -24228 -33792 -24212
rect -39164 -24292 -33876 -24228
rect -33812 -24292 -33792 -24228
rect -39164 -24308 -33792 -24292
rect -39164 -24372 -33876 -24308
rect -33812 -24372 -33792 -24308
rect -39164 -24388 -33792 -24372
rect -39164 -24452 -33876 -24388
rect -33812 -24452 -33792 -24388
rect -39164 -24468 -33792 -24452
rect -39164 -24532 -33876 -24468
rect -33812 -24532 -33792 -24468
rect -39164 -24548 -33792 -24532
rect -39164 -24612 -33876 -24548
rect -33812 -24612 -33792 -24548
rect -39164 -24628 -33792 -24612
rect -39164 -24692 -33876 -24628
rect -33812 -24692 -33792 -24628
rect -39164 -24708 -33792 -24692
rect -39164 -24772 -33876 -24708
rect -33812 -24772 -33792 -24708
rect -39164 -24788 -33792 -24772
rect -39164 -24852 -33876 -24788
rect -33812 -24852 -33792 -24788
rect -39164 -24868 -33792 -24852
rect -39164 -24932 -33876 -24868
rect -33812 -24932 -33792 -24868
rect -39164 -24948 -33792 -24932
rect -39164 -25012 -33876 -24948
rect -33812 -25012 -33792 -24948
rect -39164 -25028 -33792 -25012
rect -39164 -25092 -33876 -25028
rect -33812 -25092 -33792 -25028
rect -39164 -25108 -33792 -25092
rect -39164 -25172 -33876 -25108
rect -33812 -25172 -33792 -25108
rect -39164 -25188 -33792 -25172
rect -39164 -25252 -33876 -25188
rect -33812 -25252 -33792 -25188
rect -39164 -25268 -33792 -25252
rect -39164 -25332 -33876 -25268
rect -33812 -25332 -33792 -25268
rect -39164 -25348 -33792 -25332
rect -39164 -25412 -33876 -25348
rect -33812 -25412 -33792 -25348
rect -39164 -25428 -33792 -25412
rect -39164 -25492 -33876 -25428
rect -33812 -25492 -33792 -25428
rect -39164 -25508 -33792 -25492
rect -39164 -25572 -33876 -25508
rect -33812 -25572 -33792 -25508
rect -39164 -25588 -33792 -25572
rect -39164 -25652 -33876 -25588
rect -33812 -25652 -33792 -25588
rect -39164 -25668 -33792 -25652
rect -39164 -25732 -33876 -25668
rect -33812 -25732 -33792 -25668
rect -39164 -25748 -33792 -25732
rect -39164 -25812 -33876 -25748
rect -33812 -25812 -33792 -25748
rect -39164 -25828 -33792 -25812
rect -39164 -25892 -33876 -25828
rect -33812 -25892 -33792 -25828
rect -39164 -25908 -33792 -25892
rect -39164 -25972 -33876 -25908
rect -33812 -25972 -33792 -25908
rect -39164 -25988 -33792 -25972
rect -39164 -26052 -33876 -25988
rect -33812 -26052 -33792 -25988
rect -39164 -26068 -33792 -26052
rect -39164 -26132 -33876 -26068
rect -33812 -26132 -33792 -26068
rect -39164 -26148 -33792 -26132
rect -39164 -26212 -33876 -26148
rect -33812 -26212 -33792 -26148
rect -39164 -26228 -33792 -26212
rect -39164 -26292 -33876 -26228
rect -33812 -26292 -33792 -26228
rect -39164 -26308 -33792 -26292
rect -39164 -26372 -33876 -26308
rect -33812 -26372 -33792 -26308
rect -39164 -26388 -33792 -26372
rect -39164 -26452 -33876 -26388
rect -33812 -26452 -33792 -26388
rect -39164 -26480 -33792 -26452
rect -33552 -21428 -28180 -21400
rect -33552 -21492 -28264 -21428
rect -28200 -21492 -28180 -21428
rect -33552 -21508 -28180 -21492
rect -33552 -21572 -28264 -21508
rect -28200 -21572 -28180 -21508
rect -33552 -21588 -28180 -21572
rect -33552 -21652 -28264 -21588
rect -28200 -21652 -28180 -21588
rect -33552 -21668 -28180 -21652
rect -33552 -21732 -28264 -21668
rect -28200 -21732 -28180 -21668
rect -33552 -21748 -28180 -21732
rect -33552 -21812 -28264 -21748
rect -28200 -21812 -28180 -21748
rect -33552 -21828 -28180 -21812
rect -33552 -21892 -28264 -21828
rect -28200 -21892 -28180 -21828
rect -33552 -21908 -28180 -21892
rect -33552 -21972 -28264 -21908
rect -28200 -21972 -28180 -21908
rect -33552 -21988 -28180 -21972
rect -33552 -22052 -28264 -21988
rect -28200 -22052 -28180 -21988
rect -33552 -22068 -28180 -22052
rect -33552 -22132 -28264 -22068
rect -28200 -22132 -28180 -22068
rect -33552 -22148 -28180 -22132
rect -33552 -22212 -28264 -22148
rect -28200 -22212 -28180 -22148
rect -33552 -22228 -28180 -22212
rect -33552 -22292 -28264 -22228
rect -28200 -22292 -28180 -22228
rect -33552 -22308 -28180 -22292
rect -33552 -22372 -28264 -22308
rect -28200 -22372 -28180 -22308
rect -33552 -22388 -28180 -22372
rect -33552 -22452 -28264 -22388
rect -28200 -22452 -28180 -22388
rect -33552 -22468 -28180 -22452
rect -33552 -22532 -28264 -22468
rect -28200 -22532 -28180 -22468
rect -33552 -22548 -28180 -22532
rect -33552 -22612 -28264 -22548
rect -28200 -22612 -28180 -22548
rect -33552 -22628 -28180 -22612
rect -33552 -22692 -28264 -22628
rect -28200 -22692 -28180 -22628
rect -33552 -22708 -28180 -22692
rect -33552 -22772 -28264 -22708
rect -28200 -22772 -28180 -22708
rect -33552 -22788 -28180 -22772
rect -33552 -22852 -28264 -22788
rect -28200 -22852 -28180 -22788
rect -33552 -22868 -28180 -22852
rect -33552 -22932 -28264 -22868
rect -28200 -22932 -28180 -22868
rect -33552 -22948 -28180 -22932
rect -33552 -23012 -28264 -22948
rect -28200 -23012 -28180 -22948
rect -33552 -23028 -28180 -23012
rect -33552 -23092 -28264 -23028
rect -28200 -23092 -28180 -23028
rect -33552 -23108 -28180 -23092
rect -33552 -23172 -28264 -23108
rect -28200 -23172 -28180 -23108
rect -33552 -23188 -28180 -23172
rect -33552 -23252 -28264 -23188
rect -28200 -23252 -28180 -23188
rect -33552 -23268 -28180 -23252
rect -33552 -23332 -28264 -23268
rect -28200 -23332 -28180 -23268
rect -33552 -23348 -28180 -23332
rect -33552 -23412 -28264 -23348
rect -28200 -23412 -28180 -23348
rect -33552 -23428 -28180 -23412
rect -33552 -23492 -28264 -23428
rect -28200 -23492 -28180 -23428
rect -33552 -23508 -28180 -23492
rect -33552 -23572 -28264 -23508
rect -28200 -23572 -28180 -23508
rect -33552 -23588 -28180 -23572
rect -33552 -23652 -28264 -23588
rect -28200 -23652 -28180 -23588
rect -33552 -23668 -28180 -23652
rect -33552 -23732 -28264 -23668
rect -28200 -23732 -28180 -23668
rect -33552 -23748 -28180 -23732
rect -33552 -23812 -28264 -23748
rect -28200 -23812 -28180 -23748
rect -33552 -23828 -28180 -23812
rect -33552 -23892 -28264 -23828
rect -28200 -23892 -28180 -23828
rect -33552 -23908 -28180 -23892
rect -33552 -23972 -28264 -23908
rect -28200 -23972 -28180 -23908
rect -33552 -23988 -28180 -23972
rect -33552 -24052 -28264 -23988
rect -28200 -24052 -28180 -23988
rect -33552 -24068 -28180 -24052
rect -33552 -24132 -28264 -24068
rect -28200 -24132 -28180 -24068
rect -33552 -24148 -28180 -24132
rect -33552 -24212 -28264 -24148
rect -28200 -24212 -28180 -24148
rect -33552 -24228 -28180 -24212
rect -33552 -24292 -28264 -24228
rect -28200 -24292 -28180 -24228
rect -33552 -24308 -28180 -24292
rect -33552 -24372 -28264 -24308
rect -28200 -24372 -28180 -24308
rect -33552 -24388 -28180 -24372
rect -33552 -24452 -28264 -24388
rect -28200 -24452 -28180 -24388
rect -33552 -24468 -28180 -24452
rect -33552 -24532 -28264 -24468
rect -28200 -24532 -28180 -24468
rect -33552 -24548 -28180 -24532
rect -33552 -24612 -28264 -24548
rect -28200 -24612 -28180 -24548
rect -33552 -24628 -28180 -24612
rect -33552 -24692 -28264 -24628
rect -28200 -24692 -28180 -24628
rect -33552 -24708 -28180 -24692
rect -33552 -24772 -28264 -24708
rect -28200 -24772 -28180 -24708
rect -33552 -24788 -28180 -24772
rect -33552 -24852 -28264 -24788
rect -28200 -24852 -28180 -24788
rect -33552 -24868 -28180 -24852
rect -33552 -24932 -28264 -24868
rect -28200 -24932 -28180 -24868
rect -33552 -24948 -28180 -24932
rect -33552 -25012 -28264 -24948
rect -28200 -25012 -28180 -24948
rect -33552 -25028 -28180 -25012
rect -33552 -25092 -28264 -25028
rect -28200 -25092 -28180 -25028
rect -33552 -25108 -28180 -25092
rect -33552 -25172 -28264 -25108
rect -28200 -25172 -28180 -25108
rect -33552 -25188 -28180 -25172
rect -33552 -25252 -28264 -25188
rect -28200 -25252 -28180 -25188
rect -33552 -25268 -28180 -25252
rect -33552 -25332 -28264 -25268
rect -28200 -25332 -28180 -25268
rect -33552 -25348 -28180 -25332
rect -33552 -25412 -28264 -25348
rect -28200 -25412 -28180 -25348
rect -33552 -25428 -28180 -25412
rect -33552 -25492 -28264 -25428
rect -28200 -25492 -28180 -25428
rect -33552 -25508 -28180 -25492
rect -33552 -25572 -28264 -25508
rect -28200 -25572 -28180 -25508
rect -33552 -25588 -28180 -25572
rect -33552 -25652 -28264 -25588
rect -28200 -25652 -28180 -25588
rect -33552 -25668 -28180 -25652
rect -33552 -25732 -28264 -25668
rect -28200 -25732 -28180 -25668
rect -33552 -25748 -28180 -25732
rect -33552 -25812 -28264 -25748
rect -28200 -25812 -28180 -25748
rect -33552 -25828 -28180 -25812
rect -33552 -25892 -28264 -25828
rect -28200 -25892 -28180 -25828
rect -33552 -25908 -28180 -25892
rect -33552 -25972 -28264 -25908
rect -28200 -25972 -28180 -25908
rect -33552 -25988 -28180 -25972
rect -33552 -26052 -28264 -25988
rect -28200 -26052 -28180 -25988
rect -33552 -26068 -28180 -26052
rect -33552 -26132 -28264 -26068
rect -28200 -26132 -28180 -26068
rect -33552 -26148 -28180 -26132
rect -33552 -26212 -28264 -26148
rect -28200 -26212 -28180 -26148
rect -33552 -26228 -28180 -26212
rect -33552 -26292 -28264 -26228
rect -28200 -26292 -28180 -26228
rect -33552 -26308 -28180 -26292
rect -33552 -26372 -28264 -26308
rect -28200 -26372 -28180 -26308
rect -33552 -26388 -28180 -26372
rect -33552 -26452 -28264 -26388
rect -28200 -26452 -28180 -26388
rect -33552 -26480 -28180 -26452
rect -27940 -21428 -22568 -21400
rect -27940 -21492 -22652 -21428
rect -22588 -21492 -22568 -21428
rect -27940 -21508 -22568 -21492
rect -27940 -21572 -22652 -21508
rect -22588 -21572 -22568 -21508
rect -27940 -21588 -22568 -21572
rect -27940 -21652 -22652 -21588
rect -22588 -21652 -22568 -21588
rect -27940 -21668 -22568 -21652
rect -27940 -21732 -22652 -21668
rect -22588 -21732 -22568 -21668
rect -27940 -21748 -22568 -21732
rect -27940 -21812 -22652 -21748
rect -22588 -21812 -22568 -21748
rect -27940 -21828 -22568 -21812
rect -27940 -21892 -22652 -21828
rect -22588 -21892 -22568 -21828
rect -27940 -21908 -22568 -21892
rect -27940 -21972 -22652 -21908
rect -22588 -21972 -22568 -21908
rect -27940 -21988 -22568 -21972
rect -27940 -22052 -22652 -21988
rect -22588 -22052 -22568 -21988
rect -27940 -22068 -22568 -22052
rect -27940 -22132 -22652 -22068
rect -22588 -22132 -22568 -22068
rect -27940 -22148 -22568 -22132
rect -27940 -22212 -22652 -22148
rect -22588 -22212 -22568 -22148
rect -27940 -22228 -22568 -22212
rect -27940 -22292 -22652 -22228
rect -22588 -22292 -22568 -22228
rect -27940 -22308 -22568 -22292
rect -27940 -22372 -22652 -22308
rect -22588 -22372 -22568 -22308
rect -27940 -22388 -22568 -22372
rect -27940 -22452 -22652 -22388
rect -22588 -22452 -22568 -22388
rect -27940 -22468 -22568 -22452
rect -27940 -22532 -22652 -22468
rect -22588 -22532 -22568 -22468
rect -27940 -22548 -22568 -22532
rect -27940 -22612 -22652 -22548
rect -22588 -22612 -22568 -22548
rect -27940 -22628 -22568 -22612
rect -27940 -22692 -22652 -22628
rect -22588 -22692 -22568 -22628
rect -27940 -22708 -22568 -22692
rect -27940 -22772 -22652 -22708
rect -22588 -22772 -22568 -22708
rect -27940 -22788 -22568 -22772
rect -27940 -22852 -22652 -22788
rect -22588 -22852 -22568 -22788
rect -27940 -22868 -22568 -22852
rect -27940 -22932 -22652 -22868
rect -22588 -22932 -22568 -22868
rect -27940 -22948 -22568 -22932
rect -27940 -23012 -22652 -22948
rect -22588 -23012 -22568 -22948
rect -27940 -23028 -22568 -23012
rect -27940 -23092 -22652 -23028
rect -22588 -23092 -22568 -23028
rect -27940 -23108 -22568 -23092
rect -27940 -23172 -22652 -23108
rect -22588 -23172 -22568 -23108
rect -27940 -23188 -22568 -23172
rect -27940 -23252 -22652 -23188
rect -22588 -23252 -22568 -23188
rect -27940 -23268 -22568 -23252
rect -27940 -23332 -22652 -23268
rect -22588 -23332 -22568 -23268
rect -27940 -23348 -22568 -23332
rect -27940 -23412 -22652 -23348
rect -22588 -23412 -22568 -23348
rect -27940 -23428 -22568 -23412
rect -27940 -23492 -22652 -23428
rect -22588 -23492 -22568 -23428
rect -27940 -23508 -22568 -23492
rect -27940 -23572 -22652 -23508
rect -22588 -23572 -22568 -23508
rect -27940 -23588 -22568 -23572
rect -27940 -23652 -22652 -23588
rect -22588 -23652 -22568 -23588
rect -27940 -23668 -22568 -23652
rect -27940 -23732 -22652 -23668
rect -22588 -23732 -22568 -23668
rect -27940 -23748 -22568 -23732
rect -27940 -23812 -22652 -23748
rect -22588 -23812 -22568 -23748
rect -27940 -23828 -22568 -23812
rect -27940 -23892 -22652 -23828
rect -22588 -23892 -22568 -23828
rect -27940 -23908 -22568 -23892
rect -27940 -23972 -22652 -23908
rect -22588 -23972 -22568 -23908
rect -27940 -23988 -22568 -23972
rect -27940 -24052 -22652 -23988
rect -22588 -24052 -22568 -23988
rect -27940 -24068 -22568 -24052
rect -27940 -24132 -22652 -24068
rect -22588 -24132 -22568 -24068
rect -27940 -24148 -22568 -24132
rect -27940 -24212 -22652 -24148
rect -22588 -24212 -22568 -24148
rect -27940 -24228 -22568 -24212
rect -27940 -24292 -22652 -24228
rect -22588 -24292 -22568 -24228
rect -27940 -24308 -22568 -24292
rect -27940 -24372 -22652 -24308
rect -22588 -24372 -22568 -24308
rect -27940 -24388 -22568 -24372
rect -27940 -24452 -22652 -24388
rect -22588 -24452 -22568 -24388
rect -27940 -24468 -22568 -24452
rect -27940 -24532 -22652 -24468
rect -22588 -24532 -22568 -24468
rect -27940 -24548 -22568 -24532
rect -27940 -24612 -22652 -24548
rect -22588 -24612 -22568 -24548
rect -27940 -24628 -22568 -24612
rect -27940 -24692 -22652 -24628
rect -22588 -24692 -22568 -24628
rect -27940 -24708 -22568 -24692
rect -27940 -24772 -22652 -24708
rect -22588 -24772 -22568 -24708
rect -27940 -24788 -22568 -24772
rect -27940 -24852 -22652 -24788
rect -22588 -24852 -22568 -24788
rect -27940 -24868 -22568 -24852
rect -27940 -24932 -22652 -24868
rect -22588 -24932 -22568 -24868
rect -27940 -24948 -22568 -24932
rect -27940 -25012 -22652 -24948
rect -22588 -25012 -22568 -24948
rect -27940 -25028 -22568 -25012
rect -27940 -25092 -22652 -25028
rect -22588 -25092 -22568 -25028
rect -27940 -25108 -22568 -25092
rect -27940 -25172 -22652 -25108
rect -22588 -25172 -22568 -25108
rect -27940 -25188 -22568 -25172
rect -27940 -25252 -22652 -25188
rect -22588 -25252 -22568 -25188
rect -27940 -25268 -22568 -25252
rect -27940 -25332 -22652 -25268
rect -22588 -25332 -22568 -25268
rect -27940 -25348 -22568 -25332
rect -27940 -25412 -22652 -25348
rect -22588 -25412 -22568 -25348
rect -27940 -25428 -22568 -25412
rect -27940 -25492 -22652 -25428
rect -22588 -25492 -22568 -25428
rect -27940 -25508 -22568 -25492
rect -27940 -25572 -22652 -25508
rect -22588 -25572 -22568 -25508
rect -27940 -25588 -22568 -25572
rect -27940 -25652 -22652 -25588
rect -22588 -25652 -22568 -25588
rect -27940 -25668 -22568 -25652
rect -27940 -25732 -22652 -25668
rect -22588 -25732 -22568 -25668
rect -27940 -25748 -22568 -25732
rect -27940 -25812 -22652 -25748
rect -22588 -25812 -22568 -25748
rect -27940 -25828 -22568 -25812
rect -27940 -25892 -22652 -25828
rect -22588 -25892 -22568 -25828
rect -27940 -25908 -22568 -25892
rect -27940 -25972 -22652 -25908
rect -22588 -25972 -22568 -25908
rect -27940 -25988 -22568 -25972
rect -27940 -26052 -22652 -25988
rect -22588 -26052 -22568 -25988
rect -27940 -26068 -22568 -26052
rect -27940 -26132 -22652 -26068
rect -22588 -26132 -22568 -26068
rect -27940 -26148 -22568 -26132
rect -27940 -26212 -22652 -26148
rect -22588 -26212 -22568 -26148
rect -27940 -26228 -22568 -26212
rect -27940 -26292 -22652 -26228
rect -22588 -26292 -22568 -26228
rect -27940 -26308 -22568 -26292
rect -27940 -26372 -22652 -26308
rect -22588 -26372 -22568 -26308
rect -27940 -26388 -22568 -26372
rect -27940 -26452 -22652 -26388
rect -22588 -26452 -22568 -26388
rect -27940 -26480 -22568 -26452
rect -22328 -21428 -16956 -21400
rect -22328 -21492 -17040 -21428
rect -16976 -21492 -16956 -21428
rect -22328 -21508 -16956 -21492
rect -22328 -21572 -17040 -21508
rect -16976 -21572 -16956 -21508
rect -22328 -21588 -16956 -21572
rect -22328 -21652 -17040 -21588
rect -16976 -21652 -16956 -21588
rect -22328 -21668 -16956 -21652
rect -22328 -21732 -17040 -21668
rect -16976 -21732 -16956 -21668
rect -22328 -21748 -16956 -21732
rect -22328 -21812 -17040 -21748
rect -16976 -21812 -16956 -21748
rect -22328 -21828 -16956 -21812
rect -22328 -21892 -17040 -21828
rect -16976 -21892 -16956 -21828
rect -22328 -21908 -16956 -21892
rect -22328 -21972 -17040 -21908
rect -16976 -21972 -16956 -21908
rect -22328 -21988 -16956 -21972
rect -22328 -22052 -17040 -21988
rect -16976 -22052 -16956 -21988
rect -22328 -22068 -16956 -22052
rect -22328 -22132 -17040 -22068
rect -16976 -22132 -16956 -22068
rect -22328 -22148 -16956 -22132
rect -22328 -22212 -17040 -22148
rect -16976 -22212 -16956 -22148
rect -22328 -22228 -16956 -22212
rect -22328 -22292 -17040 -22228
rect -16976 -22292 -16956 -22228
rect -22328 -22308 -16956 -22292
rect -22328 -22372 -17040 -22308
rect -16976 -22372 -16956 -22308
rect -22328 -22388 -16956 -22372
rect -22328 -22452 -17040 -22388
rect -16976 -22452 -16956 -22388
rect -22328 -22468 -16956 -22452
rect -22328 -22532 -17040 -22468
rect -16976 -22532 -16956 -22468
rect -22328 -22548 -16956 -22532
rect -22328 -22612 -17040 -22548
rect -16976 -22612 -16956 -22548
rect -22328 -22628 -16956 -22612
rect -22328 -22692 -17040 -22628
rect -16976 -22692 -16956 -22628
rect -22328 -22708 -16956 -22692
rect -22328 -22772 -17040 -22708
rect -16976 -22772 -16956 -22708
rect -22328 -22788 -16956 -22772
rect -22328 -22852 -17040 -22788
rect -16976 -22852 -16956 -22788
rect -22328 -22868 -16956 -22852
rect -22328 -22932 -17040 -22868
rect -16976 -22932 -16956 -22868
rect -22328 -22948 -16956 -22932
rect -22328 -23012 -17040 -22948
rect -16976 -23012 -16956 -22948
rect -22328 -23028 -16956 -23012
rect -22328 -23092 -17040 -23028
rect -16976 -23092 -16956 -23028
rect -22328 -23108 -16956 -23092
rect -22328 -23172 -17040 -23108
rect -16976 -23172 -16956 -23108
rect -22328 -23188 -16956 -23172
rect -22328 -23252 -17040 -23188
rect -16976 -23252 -16956 -23188
rect -22328 -23268 -16956 -23252
rect -22328 -23332 -17040 -23268
rect -16976 -23332 -16956 -23268
rect -22328 -23348 -16956 -23332
rect -22328 -23412 -17040 -23348
rect -16976 -23412 -16956 -23348
rect -22328 -23428 -16956 -23412
rect -22328 -23492 -17040 -23428
rect -16976 -23492 -16956 -23428
rect -22328 -23508 -16956 -23492
rect -22328 -23572 -17040 -23508
rect -16976 -23572 -16956 -23508
rect -22328 -23588 -16956 -23572
rect -22328 -23652 -17040 -23588
rect -16976 -23652 -16956 -23588
rect -22328 -23668 -16956 -23652
rect -22328 -23732 -17040 -23668
rect -16976 -23732 -16956 -23668
rect -22328 -23748 -16956 -23732
rect -22328 -23812 -17040 -23748
rect -16976 -23812 -16956 -23748
rect -22328 -23828 -16956 -23812
rect -22328 -23892 -17040 -23828
rect -16976 -23892 -16956 -23828
rect -22328 -23908 -16956 -23892
rect -22328 -23972 -17040 -23908
rect -16976 -23972 -16956 -23908
rect -22328 -23988 -16956 -23972
rect -22328 -24052 -17040 -23988
rect -16976 -24052 -16956 -23988
rect -22328 -24068 -16956 -24052
rect -22328 -24132 -17040 -24068
rect -16976 -24132 -16956 -24068
rect -22328 -24148 -16956 -24132
rect -22328 -24212 -17040 -24148
rect -16976 -24212 -16956 -24148
rect -22328 -24228 -16956 -24212
rect -22328 -24292 -17040 -24228
rect -16976 -24292 -16956 -24228
rect -22328 -24308 -16956 -24292
rect -22328 -24372 -17040 -24308
rect -16976 -24372 -16956 -24308
rect -22328 -24388 -16956 -24372
rect -22328 -24452 -17040 -24388
rect -16976 -24452 -16956 -24388
rect -22328 -24468 -16956 -24452
rect -22328 -24532 -17040 -24468
rect -16976 -24532 -16956 -24468
rect -22328 -24548 -16956 -24532
rect -22328 -24612 -17040 -24548
rect -16976 -24612 -16956 -24548
rect -22328 -24628 -16956 -24612
rect -22328 -24692 -17040 -24628
rect -16976 -24692 -16956 -24628
rect -22328 -24708 -16956 -24692
rect -22328 -24772 -17040 -24708
rect -16976 -24772 -16956 -24708
rect -22328 -24788 -16956 -24772
rect -22328 -24852 -17040 -24788
rect -16976 -24852 -16956 -24788
rect -22328 -24868 -16956 -24852
rect -22328 -24932 -17040 -24868
rect -16976 -24932 -16956 -24868
rect -22328 -24948 -16956 -24932
rect -22328 -25012 -17040 -24948
rect -16976 -25012 -16956 -24948
rect -22328 -25028 -16956 -25012
rect -22328 -25092 -17040 -25028
rect -16976 -25092 -16956 -25028
rect -22328 -25108 -16956 -25092
rect -22328 -25172 -17040 -25108
rect -16976 -25172 -16956 -25108
rect -22328 -25188 -16956 -25172
rect -22328 -25252 -17040 -25188
rect -16976 -25252 -16956 -25188
rect -22328 -25268 -16956 -25252
rect -22328 -25332 -17040 -25268
rect -16976 -25332 -16956 -25268
rect -22328 -25348 -16956 -25332
rect -22328 -25412 -17040 -25348
rect -16976 -25412 -16956 -25348
rect -22328 -25428 -16956 -25412
rect -22328 -25492 -17040 -25428
rect -16976 -25492 -16956 -25428
rect -22328 -25508 -16956 -25492
rect -22328 -25572 -17040 -25508
rect -16976 -25572 -16956 -25508
rect -22328 -25588 -16956 -25572
rect -22328 -25652 -17040 -25588
rect -16976 -25652 -16956 -25588
rect -22328 -25668 -16956 -25652
rect -22328 -25732 -17040 -25668
rect -16976 -25732 -16956 -25668
rect -22328 -25748 -16956 -25732
rect -22328 -25812 -17040 -25748
rect -16976 -25812 -16956 -25748
rect -22328 -25828 -16956 -25812
rect -22328 -25892 -17040 -25828
rect -16976 -25892 -16956 -25828
rect -22328 -25908 -16956 -25892
rect -22328 -25972 -17040 -25908
rect -16976 -25972 -16956 -25908
rect -22328 -25988 -16956 -25972
rect -22328 -26052 -17040 -25988
rect -16976 -26052 -16956 -25988
rect -22328 -26068 -16956 -26052
rect -22328 -26132 -17040 -26068
rect -16976 -26132 -16956 -26068
rect -22328 -26148 -16956 -26132
rect -22328 -26212 -17040 -26148
rect -16976 -26212 -16956 -26148
rect -22328 -26228 -16956 -26212
rect -22328 -26292 -17040 -26228
rect -16976 -26292 -16956 -26228
rect -22328 -26308 -16956 -26292
rect -22328 -26372 -17040 -26308
rect -16976 -26372 -16956 -26308
rect -22328 -26388 -16956 -26372
rect -22328 -26452 -17040 -26388
rect -16976 -26452 -16956 -26388
rect -22328 -26480 -16956 -26452
rect -16716 -21428 -11344 -21400
rect -16716 -21492 -11428 -21428
rect -11364 -21492 -11344 -21428
rect -16716 -21508 -11344 -21492
rect -16716 -21572 -11428 -21508
rect -11364 -21572 -11344 -21508
rect -16716 -21588 -11344 -21572
rect -16716 -21652 -11428 -21588
rect -11364 -21652 -11344 -21588
rect -16716 -21668 -11344 -21652
rect -16716 -21732 -11428 -21668
rect -11364 -21732 -11344 -21668
rect -16716 -21748 -11344 -21732
rect -16716 -21812 -11428 -21748
rect -11364 -21812 -11344 -21748
rect -16716 -21828 -11344 -21812
rect -16716 -21892 -11428 -21828
rect -11364 -21892 -11344 -21828
rect -16716 -21908 -11344 -21892
rect -16716 -21972 -11428 -21908
rect -11364 -21972 -11344 -21908
rect -16716 -21988 -11344 -21972
rect -16716 -22052 -11428 -21988
rect -11364 -22052 -11344 -21988
rect -16716 -22068 -11344 -22052
rect -16716 -22132 -11428 -22068
rect -11364 -22132 -11344 -22068
rect -16716 -22148 -11344 -22132
rect -16716 -22212 -11428 -22148
rect -11364 -22212 -11344 -22148
rect -16716 -22228 -11344 -22212
rect -16716 -22292 -11428 -22228
rect -11364 -22292 -11344 -22228
rect -16716 -22308 -11344 -22292
rect -16716 -22372 -11428 -22308
rect -11364 -22372 -11344 -22308
rect -16716 -22388 -11344 -22372
rect -16716 -22452 -11428 -22388
rect -11364 -22452 -11344 -22388
rect -16716 -22468 -11344 -22452
rect -16716 -22532 -11428 -22468
rect -11364 -22532 -11344 -22468
rect -16716 -22548 -11344 -22532
rect -16716 -22612 -11428 -22548
rect -11364 -22612 -11344 -22548
rect -16716 -22628 -11344 -22612
rect -16716 -22692 -11428 -22628
rect -11364 -22692 -11344 -22628
rect -16716 -22708 -11344 -22692
rect -16716 -22772 -11428 -22708
rect -11364 -22772 -11344 -22708
rect -16716 -22788 -11344 -22772
rect -16716 -22852 -11428 -22788
rect -11364 -22852 -11344 -22788
rect -16716 -22868 -11344 -22852
rect -16716 -22932 -11428 -22868
rect -11364 -22932 -11344 -22868
rect -16716 -22948 -11344 -22932
rect -16716 -23012 -11428 -22948
rect -11364 -23012 -11344 -22948
rect -16716 -23028 -11344 -23012
rect -16716 -23092 -11428 -23028
rect -11364 -23092 -11344 -23028
rect -16716 -23108 -11344 -23092
rect -16716 -23172 -11428 -23108
rect -11364 -23172 -11344 -23108
rect -16716 -23188 -11344 -23172
rect -16716 -23252 -11428 -23188
rect -11364 -23252 -11344 -23188
rect -16716 -23268 -11344 -23252
rect -16716 -23332 -11428 -23268
rect -11364 -23332 -11344 -23268
rect -16716 -23348 -11344 -23332
rect -16716 -23412 -11428 -23348
rect -11364 -23412 -11344 -23348
rect -16716 -23428 -11344 -23412
rect -16716 -23492 -11428 -23428
rect -11364 -23492 -11344 -23428
rect -16716 -23508 -11344 -23492
rect -16716 -23572 -11428 -23508
rect -11364 -23572 -11344 -23508
rect -16716 -23588 -11344 -23572
rect -16716 -23652 -11428 -23588
rect -11364 -23652 -11344 -23588
rect -16716 -23668 -11344 -23652
rect -16716 -23732 -11428 -23668
rect -11364 -23732 -11344 -23668
rect -16716 -23748 -11344 -23732
rect -16716 -23812 -11428 -23748
rect -11364 -23812 -11344 -23748
rect -16716 -23828 -11344 -23812
rect -16716 -23892 -11428 -23828
rect -11364 -23892 -11344 -23828
rect -16716 -23908 -11344 -23892
rect -16716 -23972 -11428 -23908
rect -11364 -23972 -11344 -23908
rect -16716 -23988 -11344 -23972
rect -16716 -24052 -11428 -23988
rect -11364 -24052 -11344 -23988
rect -16716 -24068 -11344 -24052
rect -16716 -24132 -11428 -24068
rect -11364 -24132 -11344 -24068
rect -16716 -24148 -11344 -24132
rect -16716 -24212 -11428 -24148
rect -11364 -24212 -11344 -24148
rect -16716 -24228 -11344 -24212
rect -16716 -24292 -11428 -24228
rect -11364 -24292 -11344 -24228
rect -16716 -24308 -11344 -24292
rect -16716 -24372 -11428 -24308
rect -11364 -24372 -11344 -24308
rect -16716 -24388 -11344 -24372
rect -16716 -24452 -11428 -24388
rect -11364 -24452 -11344 -24388
rect -16716 -24468 -11344 -24452
rect -16716 -24532 -11428 -24468
rect -11364 -24532 -11344 -24468
rect -16716 -24548 -11344 -24532
rect -16716 -24612 -11428 -24548
rect -11364 -24612 -11344 -24548
rect -16716 -24628 -11344 -24612
rect -16716 -24692 -11428 -24628
rect -11364 -24692 -11344 -24628
rect -16716 -24708 -11344 -24692
rect -16716 -24772 -11428 -24708
rect -11364 -24772 -11344 -24708
rect -16716 -24788 -11344 -24772
rect -16716 -24852 -11428 -24788
rect -11364 -24852 -11344 -24788
rect -16716 -24868 -11344 -24852
rect -16716 -24932 -11428 -24868
rect -11364 -24932 -11344 -24868
rect -16716 -24948 -11344 -24932
rect -16716 -25012 -11428 -24948
rect -11364 -25012 -11344 -24948
rect -16716 -25028 -11344 -25012
rect -16716 -25092 -11428 -25028
rect -11364 -25092 -11344 -25028
rect -16716 -25108 -11344 -25092
rect -16716 -25172 -11428 -25108
rect -11364 -25172 -11344 -25108
rect -16716 -25188 -11344 -25172
rect -16716 -25252 -11428 -25188
rect -11364 -25252 -11344 -25188
rect -16716 -25268 -11344 -25252
rect -16716 -25332 -11428 -25268
rect -11364 -25332 -11344 -25268
rect -16716 -25348 -11344 -25332
rect -16716 -25412 -11428 -25348
rect -11364 -25412 -11344 -25348
rect -16716 -25428 -11344 -25412
rect -16716 -25492 -11428 -25428
rect -11364 -25492 -11344 -25428
rect -16716 -25508 -11344 -25492
rect -16716 -25572 -11428 -25508
rect -11364 -25572 -11344 -25508
rect -16716 -25588 -11344 -25572
rect -16716 -25652 -11428 -25588
rect -11364 -25652 -11344 -25588
rect -16716 -25668 -11344 -25652
rect -16716 -25732 -11428 -25668
rect -11364 -25732 -11344 -25668
rect -16716 -25748 -11344 -25732
rect -16716 -25812 -11428 -25748
rect -11364 -25812 -11344 -25748
rect -16716 -25828 -11344 -25812
rect -16716 -25892 -11428 -25828
rect -11364 -25892 -11344 -25828
rect -16716 -25908 -11344 -25892
rect -16716 -25972 -11428 -25908
rect -11364 -25972 -11344 -25908
rect -16716 -25988 -11344 -25972
rect -16716 -26052 -11428 -25988
rect -11364 -26052 -11344 -25988
rect -16716 -26068 -11344 -26052
rect -16716 -26132 -11428 -26068
rect -11364 -26132 -11344 -26068
rect -16716 -26148 -11344 -26132
rect -16716 -26212 -11428 -26148
rect -11364 -26212 -11344 -26148
rect -16716 -26228 -11344 -26212
rect -16716 -26292 -11428 -26228
rect -11364 -26292 -11344 -26228
rect -16716 -26308 -11344 -26292
rect -16716 -26372 -11428 -26308
rect -11364 -26372 -11344 -26308
rect -16716 -26388 -11344 -26372
rect -16716 -26452 -11428 -26388
rect -11364 -26452 -11344 -26388
rect -16716 -26480 -11344 -26452
rect -11104 -21428 -5732 -21400
rect -11104 -21492 -5816 -21428
rect -5752 -21492 -5732 -21428
rect -11104 -21508 -5732 -21492
rect -11104 -21572 -5816 -21508
rect -5752 -21572 -5732 -21508
rect -11104 -21588 -5732 -21572
rect -11104 -21652 -5816 -21588
rect -5752 -21652 -5732 -21588
rect -11104 -21668 -5732 -21652
rect -11104 -21732 -5816 -21668
rect -5752 -21732 -5732 -21668
rect -11104 -21748 -5732 -21732
rect -11104 -21812 -5816 -21748
rect -5752 -21812 -5732 -21748
rect -11104 -21828 -5732 -21812
rect -11104 -21892 -5816 -21828
rect -5752 -21892 -5732 -21828
rect -11104 -21908 -5732 -21892
rect -11104 -21972 -5816 -21908
rect -5752 -21972 -5732 -21908
rect -11104 -21988 -5732 -21972
rect -11104 -22052 -5816 -21988
rect -5752 -22052 -5732 -21988
rect -11104 -22068 -5732 -22052
rect -11104 -22132 -5816 -22068
rect -5752 -22132 -5732 -22068
rect -11104 -22148 -5732 -22132
rect -11104 -22212 -5816 -22148
rect -5752 -22212 -5732 -22148
rect -11104 -22228 -5732 -22212
rect -11104 -22292 -5816 -22228
rect -5752 -22292 -5732 -22228
rect -11104 -22308 -5732 -22292
rect -11104 -22372 -5816 -22308
rect -5752 -22372 -5732 -22308
rect -11104 -22388 -5732 -22372
rect -11104 -22452 -5816 -22388
rect -5752 -22452 -5732 -22388
rect -11104 -22468 -5732 -22452
rect -11104 -22532 -5816 -22468
rect -5752 -22532 -5732 -22468
rect -11104 -22548 -5732 -22532
rect -11104 -22612 -5816 -22548
rect -5752 -22612 -5732 -22548
rect -11104 -22628 -5732 -22612
rect -11104 -22692 -5816 -22628
rect -5752 -22692 -5732 -22628
rect -11104 -22708 -5732 -22692
rect -11104 -22772 -5816 -22708
rect -5752 -22772 -5732 -22708
rect -11104 -22788 -5732 -22772
rect -11104 -22852 -5816 -22788
rect -5752 -22852 -5732 -22788
rect -11104 -22868 -5732 -22852
rect -11104 -22932 -5816 -22868
rect -5752 -22932 -5732 -22868
rect -11104 -22948 -5732 -22932
rect -11104 -23012 -5816 -22948
rect -5752 -23012 -5732 -22948
rect -11104 -23028 -5732 -23012
rect -11104 -23092 -5816 -23028
rect -5752 -23092 -5732 -23028
rect -11104 -23108 -5732 -23092
rect -11104 -23172 -5816 -23108
rect -5752 -23172 -5732 -23108
rect -11104 -23188 -5732 -23172
rect -11104 -23252 -5816 -23188
rect -5752 -23252 -5732 -23188
rect -11104 -23268 -5732 -23252
rect -11104 -23332 -5816 -23268
rect -5752 -23332 -5732 -23268
rect -11104 -23348 -5732 -23332
rect -11104 -23412 -5816 -23348
rect -5752 -23412 -5732 -23348
rect -11104 -23428 -5732 -23412
rect -11104 -23492 -5816 -23428
rect -5752 -23492 -5732 -23428
rect -11104 -23508 -5732 -23492
rect -11104 -23572 -5816 -23508
rect -5752 -23572 -5732 -23508
rect -11104 -23588 -5732 -23572
rect -11104 -23652 -5816 -23588
rect -5752 -23652 -5732 -23588
rect -11104 -23668 -5732 -23652
rect -11104 -23732 -5816 -23668
rect -5752 -23732 -5732 -23668
rect -11104 -23748 -5732 -23732
rect -11104 -23812 -5816 -23748
rect -5752 -23812 -5732 -23748
rect -11104 -23828 -5732 -23812
rect -11104 -23892 -5816 -23828
rect -5752 -23892 -5732 -23828
rect -11104 -23908 -5732 -23892
rect -11104 -23972 -5816 -23908
rect -5752 -23972 -5732 -23908
rect -11104 -23988 -5732 -23972
rect -11104 -24052 -5816 -23988
rect -5752 -24052 -5732 -23988
rect -11104 -24068 -5732 -24052
rect -11104 -24132 -5816 -24068
rect -5752 -24132 -5732 -24068
rect -11104 -24148 -5732 -24132
rect -11104 -24212 -5816 -24148
rect -5752 -24212 -5732 -24148
rect -11104 -24228 -5732 -24212
rect -11104 -24292 -5816 -24228
rect -5752 -24292 -5732 -24228
rect -11104 -24308 -5732 -24292
rect -11104 -24372 -5816 -24308
rect -5752 -24372 -5732 -24308
rect -11104 -24388 -5732 -24372
rect -11104 -24452 -5816 -24388
rect -5752 -24452 -5732 -24388
rect -11104 -24468 -5732 -24452
rect -11104 -24532 -5816 -24468
rect -5752 -24532 -5732 -24468
rect -11104 -24548 -5732 -24532
rect -11104 -24612 -5816 -24548
rect -5752 -24612 -5732 -24548
rect -11104 -24628 -5732 -24612
rect -11104 -24692 -5816 -24628
rect -5752 -24692 -5732 -24628
rect -11104 -24708 -5732 -24692
rect -11104 -24772 -5816 -24708
rect -5752 -24772 -5732 -24708
rect -11104 -24788 -5732 -24772
rect -11104 -24852 -5816 -24788
rect -5752 -24852 -5732 -24788
rect -11104 -24868 -5732 -24852
rect -11104 -24932 -5816 -24868
rect -5752 -24932 -5732 -24868
rect -11104 -24948 -5732 -24932
rect -11104 -25012 -5816 -24948
rect -5752 -25012 -5732 -24948
rect -11104 -25028 -5732 -25012
rect -11104 -25092 -5816 -25028
rect -5752 -25092 -5732 -25028
rect -11104 -25108 -5732 -25092
rect -11104 -25172 -5816 -25108
rect -5752 -25172 -5732 -25108
rect -11104 -25188 -5732 -25172
rect -11104 -25252 -5816 -25188
rect -5752 -25252 -5732 -25188
rect -11104 -25268 -5732 -25252
rect -11104 -25332 -5816 -25268
rect -5752 -25332 -5732 -25268
rect -11104 -25348 -5732 -25332
rect -11104 -25412 -5816 -25348
rect -5752 -25412 -5732 -25348
rect -11104 -25428 -5732 -25412
rect -11104 -25492 -5816 -25428
rect -5752 -25492 -5732 -25428
rect -11104 -25508 -5732 -25492
rect -11104 -25572 -5816 -25508
rect -5752 -25572 -5732 -25508
rect -11104 -25588 -5732 -25572
rect -11104 -25652 -5816 -25588
rect -5752 -25652 -5732 -25588
rect -11104 -25668 -5732 -25652
rect -11104 -25732 -5816 -25668
rect -5752 -25732 -5732 -25668
rect -11104 -25748 -5732 -25732
rect -11104 -25812 -5816 -25748
rect -5752 -25812 -5732 -25748
rect -11104 -25828 -5732 -25812
rect -11104 -25892 -5816 -25828
rect -5752 -25892 -5732 -25828
rect -11104 -25908 -5732 -25892
rect -11104 -25972 -5816 -25908
rect -5752 -25972 -5732 -25908
rect -11104 -25988 -5732 -25972
rect -11104 -26052 -5816 -25988
rect -5752 -26052 -5732 -25988
rect -11104 -26068 -5732 -26052
rect -11104 -26132 -5816 -26068
rect -5752 -26132 -5732 -26068
rect -11104 -26148 -5732 -26132
rect -11104 -26212 -5816 -26148
rect -5752 -26212 -5732 -26148
rect -11104 -26228 -5732 -26212
rect -11104 -26292 -5816 -26228
rect -5752 -26292 -5732 -26228
rect -11104 -26308 -5732 -26292
rect -11104 -26372 -5816 -26308
rect -5752 -26372 -5732 -26308
rect -11104 -26388 -5732 -26372
rect -11104 -26452 -5816 -26388
rect -5752 -26452 -5732 -26388
rect -11104 -26480 -5732 -26452
rect -5492 -21428 -120 -21400
rect -5492 -21492 -204 -21428
rect -140 -21492 -120 -21428
rect -5492 -21508 -120 -21492
rect -5492 -21572 -204 -21508
rect -140 -21572 -120 -21508
rect -5492 -21588 -120 -21572
rect -5492 -21652 -204 -21588
rect -140 -21652 -120 -21588
rect -5492 -21668 -120 -21652
rect -5492 -21732 -204 -21668
rect -140 -21732 -120 -21668
rect -5492 -21748 -120 -21732
rect -5492 -21812 -204 -21748
rect -140 -21812 -120 -21748
rect -5492 -21828 -120 -21812
rect -5492 -21892 -204 -21828
rect -140 -21892 -120 -21828
rect -5492 -21908 -120 -21892
rect -5492 -21972 -204 -21908
rect -140 -21972 -120 -21908
rect -5492 -21988 -120 -21972
rect -5492 -22052 -204 -21988
rect -140 -22052 -120 -21988
rect -5492 -22068 -120 -22052
rect -5492 -22132 -204 -22068
rect -140 -22132 -120 -22068
rect -5492 -22148 -120 -22132
rect -5492 -22212 -204 -22148
rect -140 -22212 -120 -22148
rect -5492 -22228 -120 -22212
rect -5492 -22292 -204 -22228
rect -140 -22292 -120 -22228
rect -5492 -22308 -120 -22292
rect -5492 -22372 -204 -22308
rect -140 -22372 -120 -22308
rect -5492 -22388 -120 -22372
rect -5492 -22452 -204 -22388
rect -140 -22452 -120 -22388
rect -5492 -22468 -120 -22452
rect -5492 -22532 -204 -22468
rect -140 -22532 -120 -22468
rect -5492 -22548 -120 -22532
rect -5492 -22612 -204 -22548
rect -140 -22612 -120 -22548
rect -5492 -22628 -120 -22612
rect -5492 -22692 -204 -22628
rect -140 -22692 -120 -22628
rect -5492 -22708 -120 -22692
rect -5492 -22772 -204 -22708
rect -140 -22772 -120 -22708
rect -5492 -22788 -120 -22772
rect -5492 -22852 -204 -22788
rect -140 -22852 -120 -22788
rect -5492 -22868 -120 -22852
rect -5492 -22932 -204 -22868
rect -140 -22932 -120 -22868
rect -5492 -22948 -120 -22932
rect -5492 -23012 -204 -22948
rect -140 -23012 -120 -22948
rect -5492 -23028 -120 -23012
rect -5492 -23092 -204 -23028
rect -140 -23092 -120 -23028
rect -5492 -23108 -120 -23092
rect -5492 -23172 -204 -23108
rect -140 -23172 -120 -23108
rect -5492 -23188 -120 -23172
rect -5492 -23252 -204 -23188
rect -140 -23252 -120 -23188
rect -5492 -23268 -120 -23252
rect -5492 -23332 -204 -23268
rect -140 -23332 -120 -23268
rect -5492 -23348 -120 -23332
rect -5492 -23412 -204 -23348
rect -140 -23412 -120 -23348
rect -5492 -23428 -120 -23412
rect -5492 -23492 -204 -23428
rect -140 -23492 -120 -23428
rect -5492 -23508 -120 -23492
rect -5492 -23572 -204 -23508
rect -140 -23572 -120 -23508
rect -5492 -23588 -120 -23572
rect -5492 -23652 -204 -23588
rect -140 -23652 -120 -23588
rect -5492 -23668 -120 -23652
rect -5492 -23732 -204 -23668
rect -140 -23732 -120 -23668
rect -5492 -23748 -120 -23732
rect -5492 -23812 -204 -23748
rect -140 -23812 -120 -23748
rect -5492 -23828 -120 -23812
rect -5492 -23892 -204 -23828
rect -140 -23892 -120 -23828
rect -5492 -23908 -120 -23892
rect -5492 -23972 -204 -23908
rect -140 -23972 -120 -23908
rect -5492 -23988 -120 -23972
rect -5492 -24052 -204 -23988
rect -140 -24052 -120 -23988
rect -5492 -24068 -120 -24052
rect -5492 -24132 -204 -24068
rect -140 -24132 -120 -24068
rect -5492 -24148 -120 -24132
rect -5492 -24212 -204 -24148
rect -140 -24212 -120 -24148
rect -5492 -24228 -120 -24212
rect -5492 -24292 -204 -24228
rect -140 -24292 -120 -24228
rect -5492 -24308 -120 -24292
rect -5492 -24372 -204 -24308
rect -140 -24372 -120 -24308
rect -5492 -24388 -120 -24372
rect -5492 -24452 -204 -24388
rect -140 -24452 -120 -24388
rect -5492 -24468 -120 -24452
rect -5492 -24532 -204 -24468
rect -140 -24532 -120 -24468
rect -5492 -24548 -120 -24532
rect -5492 -24612 -204 -24548
rect -140 -24612 -120 -24548
rect -5492 -24628 -120 -24612
rect -5492 -24692 -204 -24628
rect -140 -24692 -120 -24628
rect -5492 -24708 -120 -24692
rect -5492 -24772 -204 -24708
rect -140 -24772 -120 -24708
rect -5492 -24788 -120 -24772
rect -5492 -24852 -204 -24788
rect -140 -24852 -120 -24788
rect -5492 -24868 -120 -24852
rect -5492 -24932 -204 -24868
rect -140 -24932 -120 -24868
rect -5492 -24948 -120 -24932
rect -5492 -25012 -204 -24948
rect -140 -25012 -120 -24948
rect -5492 -25028 -120 -25012
rect -5492 -25092 -204 -25028
rect -140 -25092 -120 -25028
rect -5492 -25108 -120 -25092
rect -5492 -25172 -204 -25108
rect -140 -25172 -120 -25108
rect -5492 -25188 -120 -25172
rect -5492 -25252 -204 -25188
rect -140 -25252 -120 -25188
rect -5492 -25268 -120 -25252
rect -5492 -25332 -204 -25268
rect -140 -25332 -120 -25268
rect -5492 -25348 -120 -25332
rect -5492 -25412 -204 -25348
rect -140 -25412 -120 -25348
rect -5492 -25428 -120 -25412
rect -5492 -25492 -204 -25428
rect -140 -25492 -120 -25428
rect -5492 -25508 -120 -25492
rect -5492 -25572 -204 -25508
rect -140 -25572 -120 -25508
rect -5492 -25588 -120 -25572
rect -5492 -25652 -204 -25588
rect -140 -25652 -120 -25588
rect -5492 -25668 -120 -25652
rect -5492 -25732 -204 -25668
rect -140 -25732 -120 -25668
rect -5492 -25748 -120 -25732
rect -5492 -25812 -204 -25748
rect -140 -25812 -120 -25748
rect -5492 -25828 -120 -25812
rect -5492 -25892 -204 -25828
rect -140 -25892 -120 -25828
rect -5492 -25908 -120 -25892
rect -5492 -25972 -204 -25908
rect -140 -25972 -120 -25908
rect -5492 -25988 -120 -25972
rect -5492 -26052 -204 -25988
rect -140 -26052 -120 -25988
rect -5492 -26068 -120 -26052
rect -5492 -26132 -204 -26068
rect -140 -26132 -120 -26068
rect -5492 -26148 -120 -26132
rect -5492 -26212 -204 -26148
rect -140 -26212 -120 -26148
rect -5492 -26228 -120 -26212
rect -5492 -26292 -204 -26228
rect -140 -26292 -120 -26228
rect -5492 -26308 -120 -26292
rect -5492 -26372 -204 -26308
rect -140 -26372 -120 -26308
rect -5492 -26388 -120 -26372
rect -5492 -26452 -204 -26388
rect -140 -26452 -120 -26388
rect -5492 -26480 -120 -26452
rect 120 -21428 5492 -21400
rect 120 -21492 5408 -21428
rect 5472 -21492 5492 -21428
rect 120 -21508 5492 -21492
rect 120 -21572 5408 -21508
rect 5472 -21572 5492 -21508
rect 120 -21588 5492 -21572
rect 120 -21652 5408 -21588
rect 5472 -21652 5492 -21588
rect 120 -21668 5492 -21652
rect 120 -21732 5408 -21668
rect 5472 -21732 5492 -21668
rect 120 -21748 5492 -21732
rect 120 -21812 5408 -21748
rect 5472 -21812 5492 -21748
rect 120 -21828 5492 -21812
rect 120 -21892 5408 -21828
rect 5472 -21892 5492 -21828
rect 120 -21908 5492 -21892
rect 120 -21972 5408 -21908
rect 5472 -21972 5492 -21908
rect 120 -21988 5492 -21972
rect 120 -22052 5408 -21988
rect 5472 -22052 5492 -21988
rect 120 -22068 5492 -22052
rect 120 -22132 5408 -22068
rect 5472 -22132 5492 -22068
rect 120 -22148 5492 -22132
rect 120 -22212 5408 -22148
rect 5472 -22212 5492 -22148
rect 120 -22228 5492 -22212
rect 120 -22292 5408 -22228
rect 5472 -22292 5492 -22228
rect 120 -22308 5492 -22292
rect 120 -22372 5408 -22308
rect 5472 -22372 5492 -22308
rect 120 -22388 5492 -22372
rect 120 -22452 5408 -22388
rect 5472 -22452 5492 -22388
rect 120 -22468 5492 -22452
rect 120 -22532 5408 -22468
rect 5472 -22532 5492 -22468
rect 120 -22548 5492 -22532
rect 120 -22612 5408 -22548
rect 5472 -22612 5492 -22548
rect 120 -22628 5492 -22612
rect 120 -22692 5408 -22628
rect 5472 -22692 5492 -22628
rect 120 -22708 5492 -22692
rect 120 -22772 5408 -22708
rect 5472 -22772 5492 -22708
rect 120 -22788 5492 -22772
rect 120 -22852 5408 -22788
rect 5472 -22852 5492 -22788
rect 120 -22868 5492 -22852
rect 120 -22932 5408 -22868
rect 5472 -22932 5492 -22868
rect 120 -22948 5492 -22932
rect 120 -23012 5408 -22948
rect 5472 -23012 5492 -22948
rect 120 -23028 5492 -23012
rect 120 -23092 5408 -23028
rect 5472 -23092 5492 -23028
rect 120 -23108 5492 -23092
rect 120 -23172 5408 -23108
rect 5472 -23172 5492 -23108
rect 120 -23188 5492 -23172
rect 120 -23252 5408 -23188
rect 5472 -23252 5492 -23188
rect 120 -23268 5492 -23252
rect 120 -23332 5408 -23268
rect 5472 -23332 5492 -23268
rect 120 -23348 5492 -23332
rect 120 -23412 5408 -23348
rect 5472 -23412 5492 -23348
rect 120 -23428 5492 -23412
rect 120 -23492 5408 -23428
rect 5472 -23492 5492 -23428
rect 120 -23508 5492 -23492
rect 120 -23572 5408 -23508
rect 5472 -23572 5492 -23508
rect 120 -23588 5492 -23572
rect 120 -23652 5408 -23588
rect 5472 -23652 5492 -23588
rect 120 -23668 5492 -23652
rect 120 -23732 5408 -23668
rect 5472 -23732 5492 -23668
rect 120 -23748 5492 -23732
rect 120 -23812 5408 -23748
rect 5472 -23812 5492 -23748
rect 120 -23828 5492 -23812
rect 120 -23892 5408 -23828
rect 5472 -23892 5492 -23828
rect 120 -23908 5492 -23892
rect 120 -23972 5408 -23908
rect 5472 -23972 5492 -23908
rect 120 -23988 5492 -23972
rect 120 -24052 5408 -23988
rect 5472 -24052 5492 -23988
rect 120 -24068 5492 -24052
rect 120 -24132 5408 -24068
rect 5472 -24132 5492 -24068
rect 120 -24148 5492 -24132
rect 120 -24212 5408 -24148
rect 5472 -24212 5492 -24148
rect 120 -24228 5492 -24212
rect 120 -24292 5408 -24228
rect 5472 -24292 5492 -24228
rect 120 -24308 5492 -24292
rect 120 -24372 5408 -24308
rect 5472 -24372 5492 -24308
rect 120 -24388 5492 -24372
rect 120 -24452 5408 -24388
rect 5472 -24452 5492 -24388
rect 120 -24468 5492 -24452
rect 120 -24532 5408 -24468
rect 5472 -24532 5492 -24468
rect 120 -24548 5492 -24532
rect 120 -24612 5408 -24548
rect 5472 -24612 5492 -24548
rect 120 -24628 5492 -24612
rect 120 -24692 5408 -24628
rect 5472 -24692 5492 -24628
rect 120 -24708 5492 -24692
rect 120 -24772 5408 -24708
rect 5472 -24772 5492 -24708
rect 120 -24788 5492 -24772
rect 120 -24852 5408 -24788
rect 5472 -24852 5492 -24788
rect 120 -24868 5492 -24852
rect 120 -24932 5408 -24868
rect 5472 -24932 5492 -24868
rect 120 -24948 5492 -24932
rect 120 -25012 5408 -24948
rect 5472 -25012 5492 -24948
rect 120 -25028 5492 -25012
rect 120 -25092 5408 -25028
rect 5472 -25092 5492 -25028
rect 120 -25108 5492 -25092
rect 120 -25172 5408 -25108
rect 5472 -25172 5492 -25108
rect 120 -25188 5492 -25172
rect 120 -25252 5408 -25188
rect 5472 -25252 5492 -25188
rect 120 -25268 5492 -25252
rect 120 -25332 5408 -25268
rect 5472 -25332 5492 -25268
rect 120 -25348 5492 -25332
rect 120 -25412 5408 -25348
rect 5472 -25412 5492 -25348
rect 120 -25428 5492 -25412
rect 120 -25492 5408 -25428
rect 5472 -25492 5492 -25428
rect 120 -25508 5492 -25492
rect 120 -25572 5408 -25508
rect 5472 -25572 5492 -25508
rect 120 -25588 5492 -25572
rect 120 -25652 5408 -25588
rect 5472 -25652 5492 -25588
rect 120 -25668 5492 -25652
rect 120 -25732 5408 -25668
rect 5472 -25732 5492 -25668
rect 120 -25748 5492 -25732
rect 120 -25812 5408 -25748
rect 5472 -25812 5492 -25748
rect 120 -25828 5492 -25812
rect 120 -25892 5408 -25828
rect 5472 -25892 5492 -25828
rect 120 -25908 5492 -25892
rect 120 -25972 5408 -25908
rect 5472 -25972 5492 -25908
rect 120 -25988 5492 -25972
rect 120 -26052 5408 -25988
rect 5472 -26052 5492 -25988
rect 120 -26068 5492 -26052
rect 120 -26132 5408 -26068
rect 5472 -26132 5492 -26068
rect 120 -26148 5492 -26132
rect 120 -26212 5408 -26148
rect 5472 -26212 5492 -26148
rect 120 -26228 5492 -26212
rect 120 -26292 5408 -26228
rect 5472 -26292 5492 -26228
rect 120 -26308 5492 -26292
rect 120 -26372 5408 -26308
rect 5472 -26372 5492 -26308
rect 120 -26388 5492 -26372
rect 120 -26452 5408 -26388
rect 5472 -26452 5492 -26388
rect 120 -26480 5492 -26452
rect 5732 -21428 11104 -21400
rect 5732 -21492 11020 -21428
rect 11084 -21492 11104 -21428
rect 5732 -21508 11104 -21492
rect 5732 -21572 11020 -21508
rect 11084 -21572 11104 -21508
rect 5732 -21588 11104 -21572
rect 5732 -21652 11020 -21588
rect 11084 -21652 11104 -21588
rect 5732 -21668 11104 -21652
rect 5732 -21732 11020 -21668
rect 11084 -21732 11104 -21668
rect 5732 -21748 11104 -21732
rect 5732 -21812 11020 -21748
rect 11084 -21812 11104 -21748
rect 5732 -21828 11104 -21812
rect 5732 -21892 11020 -21828
rect 11084 -21892 11104 -21828
rect 5732 -21908 11104 -21892
rect 5732 -21972 11020 -21908
rect 11084 -21972 11104 -21908
rect 5732 -21988 11104 -21972
rect 5732 -22052 11020 -21988
rect 11084 -22052 11104 -21988
rect 5732 -22068 11104 -22052
rect 5732 -22132 11020 -22068
rect 11084 -22132 11104 -22068
rect 5732 -22148 11104 -22132
rect 5732 -22212 11020 -22148
rect 11084 -22212 11104 -22148
rect 5732 -22228 11104 -22212
rect 5732 -22292 11020 -22228
rect 11084 -22292 11104 -22228
rect 5732 -22308 11104 -22292
rect 5732 -22372 11020 -22308
rect 11084 -22372 11104 -22308
rect 5732 -22388 11104 -22372
rect 5732 -22452 11020 -22388
rect 11084 -22452 11104 -22388
rect 5732 -22468 11104 -22452
rect 5732 -22532 11020 -22468
rect 11084 -22532 11104 -22468
rect 5732 -22548 11104 -22532
rect 5732 -22612 11020 -22548
rect 11084 -22612 11104 -22548
rect 5732 -22628 11104 -22612
rect 5732 -22692 11020 -22628
rect 11084 -22692 11104 -22628
rect 5732 -22708 11104 -22692
rect 5732 -22772 11020 -22708
rect 11084 -22772 11104 -22708
rect 5732 -22788 11104 -22772
rect 5732 -22852 11020 -22788
rect 11084 -22852 11104 -22788
rect 5732 -22868 11104 -22852
rect 5732 -22932 11020 -22868
rect 11084 -22932 11104 -22868
rect 5732 -22948 11104 -22932
rect 5732 -23012 11020 -22948
rect 11084 -23012 11104 -22948
rect 5732 -23028 11104 -23012
rect 5732 -23092 11020 -23028
rect 11084 -23092 11104 -23028
rect 5732 -23108 11104 -23092
rect 5732 -23172 11020 -23108
rect 11084 -23172 11104 -23108
rect 5732 -23188 11104 -23172
rect 5732 -23252 11020 -23188
rect 11084 -23252 11104 -23188
rect 5732 -23268 11104 -23252
rect 5732 -23332 11020 -23268
rect 11084 -23332 11104 -23268
rect 5732 -23348 11104 -23332
rect 5732 -23412 11020 -23348
rect 11084 -23412 11104 -23348
rect 5732 -23428 11104 -23412
rect 5732 -23492 11020 -23428
rect 11084 -23492 11104 -23428
rect 5732 -23508 11104 -23492
rect 5732 -23572 11020 -23508
rect 11084 -23572 11104 -23508
rect 5732 -23588 11104 -23572
rect 5732 -23652 11020 -23588
rect 11084 -23652 11104 -23588
rect 5732 -23668 11104 -23652
rect 5732 -23732 11020 -23668
rect 11084 -23732 11104 -23668
rect 5732 -23748 11104 -23732
rect 5732 -23812 11020 -23748
rect 11084 -23812 11104 -23748
rect 5732 -23828 11104 -23812
rect 5732 -23892 11020 -23828
rect 11084 -23892 11104 -23828
rect 5732 -23908 11104 -23892
rect 5732 -23972 11020 -23908
rect 11084 -23972 11104 -23908
rect 5732 -23988 11104 -23972
rect 5732 -24052 11020 -23988
rect 11084 -24052 11104 -23988
rect 5732 -24068 11104 -24052
rect 5732 -24132 11020 -24068
rect 11084 -24132 11104 -24068
rect 5732 -24148 11104 -24132
rect 5732 -24212 11020 -24148
rect 11084 -24212 11104 -24148
rect 5732 -24228 11104 -24212
rect 5732 -24292 11020 -24228
rect 11084 -24292 11104 -24228
rect 5732 -24308 11104 -24292
rect 5732 -24372 11020 -24308
rect 11084 -24372 11104 -24308
rect 5732 -24388 11104 -24372
rect 5732 -24452 11020 -24388
rect 11084 -24452 11104 -24388
rect 5732 -24468 11104 -24452
rect 5732 -24532 11020 -24468
rect 11084 -24532 11104 -24468
rect 5732 -24548 11104 -24532
rect 5732 -24612 11020 -24548
rect 11084 -24612 11104 -24548
rect 5732 -24628 11104 -24612
rect 5732 -24692 11020 -24628
rect 11084 -24692 11104 -24628
rect 5732 -24708 11104 -24692
rect 5732 -24772 11020 -24708
rect 11084 -24772 11104 -24708
rect 5732 -24788 11104 -24772
rect 5732 -24852 11020 -24788
rect 11084 -24852 11104 -24788
rect 5732 -24868 11104 -24852
rect 5732 -24932 11020 -24868
rect 11084 -24932 11104 -24868
rect 5732 -24948 11104 -24932
rect 5732 -25012 11020 -24948
rect 11084 -25012 11104 -24948
rect 5732 -25028 11104 -25012
rect 5732 -25092 11020 -25028
rect 11084 -25092 11104 -25028
rect 5732 -25108 11104 -25092
rect 5732 -25172 11020 -25108
rect 11084 -25172 11104 -25108
rect 5732 -25188 11104 -25172
rect 5732 -25252 11020 -25188
rect 11084 -25252 11104 -25188
rect 5732 -25268 11104 -25252
rect 5732 -25332 11020 -25268
rect 11084 -25332 11104 -25268
rect 5732 -25348 11104 -25332
rect 5732 -25412 11020 -25348
rect 11084 -25412 11104 -25348
rect 5732 -25428 11104 -25412
rect 5732 -25492 11020 -25428
rect 11084 -25492 11104 -25428
rect 5732 -25508 11104 -25492
rect 5732 -25572 11020 -25508
rect 11084 -25572 11104 -25508
rect 5732 -25588 11104 -25572
rect 5732 -25652 11020 -25588
rect 11084 -25652 11104 -25588
rect 5732 -25668 11104 -25652
rect 5732 -25732 11020 -25668
rect 11084 -25732 11104 -25668
rect 5732 -25748 11104 -25732
rect 5732 -25812 11020 -25748
rect 11084 -25812 11104 -25748
rect 5732 -25828 11104 -25812
rect 5732 -25892 11020 -25828
rect 11084 -25892 11104 -25828
rect 5732 -25908 11104 -25892
rect 5732 -25972 11020 -25908
rect 11084 -25972 11104 -25908
rect 5732 -25988 11104 -25972
rect 5732 -26052 11020 -25988
rect 11084 -26052 11104 -25988
rect 5732 -26068 11104 -26052
rect 5732 -26132 11020 -26068
rect 11084 -26132 11104 -26068
rect 5732 -26148 11104 -26132
rect 5732 -26212 11020 -26148
rect 11084 -26212 11104 -26148
rect 5732 -26228 11104 -26212
rect 5732 -26292 11020 -26228
rect 11084 -26292 11104 -26228
rect 5732 -26308 11104 -26292
rect 5732 -26372 11020 -26308
rect 11084 -26372 11104 -26308
rect 5732 -26388 11104 -26372
rect 5732 -26452 11020 -26388
rect 11084 -26452 11104 -26388
rect 5732 -26480 11104 -26452
rect 11344 -21428 16716 -21400
rect 11344 -21492 16632 -21428
rect 16696 -21492 16716 -21428
rect 11344 -21508 16716 -21492
rect 11344 -21572 16632 -21508
rect 16696 -21572 16716 -21508
rect 11344 -21588 16716 -21572
rect 11344 -21652 16632 -21588
rect 16696 -21652 16716 -21588
rect 11344 -21668 16716 -21652
rect 11344 -21732 16632 -21668
rect 16696 -21732 16716 -21668
rect 11344 -21748 16716 -21732
rect 11344 -21812 16632 -21748
rect 16696 -21812 16716 -21748
rect 11344 -21828 16716 -21812
rect 11344 -21892 16632 -21828
rect 16696 -21892 16716 -21828
rect 11344 -21908 16716 -21892
rect 11344 -21972 16632 -21908
rect 16696 -21972 16716 -21908
rect 11344 -21988 16716 -21972
rect 11344 -22052 16632 -21988
rect 16696 -22052 16716 -21988
rect 11344 -22068 16716 -22052
rect 11344 -22132 16632 -22068
rect 16696 -22132 16716 -22068
rect 11344 -22148 16716 -22132
rect 11344 -22212 16632 -22148
rect 16696 -22212 16716 -22148
rect 11344 -22228 16716 -22212
rect 11344 -22292 16632 -22228
rect 16696 -22292 16716 -22228
rect 11344 -22308 16716 -22292
rect 11344 -22372 16632 -22308
rect 16696 -22372 16716 -22308
rect 11344 -22388 16716 -22372
rect 11344 -22452 16632 -22388
rect 16696 -22452 16716 -22388
rect 11344 -22468 16716 -22452
rect 11344 -22532 16632 -22468
rect 16696 -22532 16716 -22468
rect 11344 -22548 16716 -22532
rect 11344 -22612 16632 -22548
rect 16696 -22612 16716 -22548
rect 11344 -22628 16716 -22612
rect 11344 -22692 16632 -22628
rect 16696 -22692 16716 -22628
rect 11344 -22708 16716 -22692
rect 11344 -22772 16632 -22708
rect 16696 -22772 16716 -22708
rect 11344 -22788 16716 -22772
rect 11344 -22852 16632 -22788
rect 16696 -22852 16716 -22788
rect 11344 -22868 16716 -22852
rect 11344 -22932 16632 -22868
rect 16696 -22932 16716 -22868
rect 11344 -22948 16716 -22932
rect 11344 -23012 16632 -22948
rect 16696 -23012 16716 -22948
rect 11344 -23028 16716 -23012
rect 11344 -23092 16632 -23028
rect 16696 -23092 16716 -23028
rect 11344 -23108 16716 -23092
rect 11344 -23172 16632 -23108
rect 16696 -23172 16716 -23108
rect 11344 -23188 16716 -23172
rect 11344 -23252 16632 -23188
rect 16696 -23252 16716 -23188
rect 11344 -23268 16716 -23252
rect 11344 -23332 16632 -23268
rect 16696 -23332 16716 -23268
rect 11344 -23348 16716 -23332
rect 11344 -23412 16632 -23348
rect 16696 -23412 16716 -23348
rect 11344 -23428 16716 -23412
rect 11344 -23492 16632 -23428
rect 16696 -23492 16716 -23428
rect 11344 -23508 16716 -23492
rect 11344 -23572 16632 -23508
rect 16696 -23572 16716 -23508
rect 11344 -23588 16716 -23572
rect 11344 -23652 16632 -23588
rect 16696 -23652 16716 -23588
rect 11344 -23668 16716 -23652
rect 11344 -23732 16632 -23668
rect 16696 -23732 16716 -23668
rect 11344 -23748 16716 -23732
rect 11344 -23812 16632 -23748
rect 16696 -23812 16716 -23748
rect 11344 -23828 16716 -23812
rect 11344 -23892 16632 -23828
rect 16696 -23892 16716 -23828
rect 11344 -23908 16716 -23892
rect 11344 -23972 16632 -23908
rect 16696 -23972 16716 -23908
rect 11344 -23988 16716 -23972
rect 11344 -24052 16632 -23988
rect 16696 -24052 16716 -23988
rect 11344 -24068 16716 -24052
rect 11344 -24132 16632 -24068
rect 16696 -24132 16716 -24068
rect 11344 -24148 16716 -24132
rect 11344 -24212 16632 -24148
rect 16696 -24212 16716 -24148
rect 11344 -24228 16716 -24212
rect 11344 -24292 16632 -24228
rect 16696 -24292 16716 -24228
rect 11344 -24308 16716 -24292
rect 11344 -24372 16632 -24308
rect 16696 -24372 16716 -24308
rect 11344 -24388 16716 -24372
rect 11344 -24452 16632 -24388
rect 16696 -24452 16716 -24388
rect 11344 -24468 16716 -24452
rect 11344 -24532 16632 -24468
rect 16696 -24532 16716 -24468
rect 11344 -24548 16716 -24532
rect 11344 -24612 16632 -24548
rect 16696 -24612 16716 -24548
rect 11344 -24628 16716 -24612
rect 11344 -24692 16632 -24628
rect 16696 -24692 16716 -24628
rect 11344 -24708 16716 -24692
rect 11344 -24772 16632 -24708
rect 16696 -24772 16716 -24708
rect 11344 -24788 16716 -24772
rect 11344 -24852 16632 -24788
rect 16696 -24852 16716 -24788
rect 11344 -24868 16716 -24852
rect 11344 -24932 16632 -24868
rect 16696 -24932 16716 -24868
rect 11344 -24948 16716 -24932
rect 11344 -25012 16632 -24948
rect 16696 -25012 16716 -24948
rect 11344 -25028 16716 -25012
rect 11344 -25092 16632 -25028
rect 16696 -25092 16716 -25028
rect 11344 -25108 16716 -25092
rect 11344 -25172 16632 -25108
rect 16696 -25172 16716 -25108
rect 11344 -25188 16716 -25172
rect 11344 -25252 16632 -25188
rect 16696 -25252 16716 -25188
rect 11344 -25268 16716 -25252
rect 11344 -25332 16632 -25268
rect 16696 -25332 16716 -25268
rect 11344 -25348 16716 -25332
rect 11344 -25412 16632 -25348
rect 16696 -25412 16716 -25348
rect 11344 -25428 16716 -25412
rect 11344 -25492 16632 -25428
rect 16696 -25492 16716 -25428
rect 11344 -25508 16716 -25492
rect 11344 -25572 16632 -25508
rect 16696 -25572 16716 -25508
rect 11344 -25588 16716 -25572
rect 11344 -25652 16632 -25588
rect 16696 -25652 16716 -25588
rect 11344 -25668 16716 -25652
rect 11344 -25732 16632 -25668
rect 16696 -25732 16716 -25668
rect 11344 -25748 16716 -25732
rect 11344 -25812 16632 -25748
rect 16696 -25812 16716 -25748
rect 11344 -25828 16716 -25812
rect 11344 -25892 16632 -25828
rect 16696 -25892 16716 -25828
rect 11344 -25908 16716 -25892
rect 11344 -25972 16632 -25908
rect 16696 -25972 16716 -25908
rect 11344 -25988 16716 -25972
rect 11344 -26052 16632 -25988
rect 16696 -26052 16716 -25988
rect 11344 -26068 16716 -26052
rect 11344 -26132 16632 -26068
rect 16696 -26132 16716 -26068
rect 11344 -26148 16716 -26132
rect 11344 -26212 16632 -26148
rect 16696 -26212 16716 -26148
rect 11344 -26228 16716 -26212
rect 11344 -26292 16632 -26228
rect 16696 -26292 16716 -26228
rect 11344 -26308 16716 -26292
rect 11344 -26372 16632 -26308
rect 16696 -26372 16716 -26308
rect 11344 -26388 16716 -26372
rect 11344 -26452 16632 -26388
rect 16696 -26452 16716 -26388
rect 11344 -26480 16716 -26452
rect 16956 -21428 22328 -21400
rect 16956 -21492 22244 -21428
rect 22308 -21492 22328 -21428
rect 16956 -21508 22328 -21492
rect 16956 -21572 22244 -21508
rect 22308 -21572 22328 -21508
rect 16956 -21588 22328 -21572
rect 16956 -21652 22244 -21588
rect 22308 -21652 22328 -21588
rect 16956 -21668 22328 -21652
rect 16956 -21732 22244 -21668
rect 22308 -21732 22328 -21668
rect 16956 -21748 22328 -21732
rect 16956 -21812 22244 -21748
rect 22308 -21812 22328 -21748
rect 16956 -21828 22328 -21812
rect 16956 -21892 22244 -21828
rect 22308 -21892 22328 -21828
rect 16956 -21908 22328 -21892
rect 16956 -21972 22244 -21908
rect 22308 -21972 22328 -21908
rect 16956 -21988 22328 -21972
rect 16956 -22052 22244 -21988
rect 22308 -22052 22328 -21988
rect 16956 -22068 22328 -22052
rect 16956 -22132 22244 -22068
rect 22308 -22132 22328 -22068
rect 16956 -22148 22328 -22132
rect 16956 -22212 22244 -22148
rect 22308 -22212 22328 -22148
rect 16956 -22228 22328 -22212
rect 16956 -22292 22244 -22228
rect 22308 -22292 22328 -22228
rect 16956 -22308 22328 -22292
rect 16956 -22372 22244 -22308
rect 22308 -22372 22328 -22308
rect 16956 -22388 22328 -22372
rect 16956 -22452 22244 -22388
rect 22308 -22452 22328 -22388
rect 16956 -22468 22328 -22452
rect 16956 -22532 22244 -22468
rect 22308 -22532 22328 -22468
rect 16956 -22548 22328 -22532
rect 16956 -22612 22244 -22548
rect 22308 -22612 22328 -22548
rect 16956 -22628 22328 -22612
rect 16956 -22692 22244 -22628
rect 22308 -22692 22328 -22628
rect 16956 -22708 22328 -22692
rect 16956 -22772 22244 -22708
rect 22308 -22772 22328 -22708
rect 16956 -22788 22328 -22772
rect 16956 -22852 22244 -22788
rect 22308 -22852 22328 -22788
rect 16956 -22868 22328 -22852
rect 16956 -22932 22244 -22868
rect 22308 -22932 22328 -22868
rect 16956 -22948 22328 -22932
rect 16956 -23012 22244 -22948
rect 22308 -23012 22328 -22948
rect 16956 -23028 22328 -23012
rect 16956 -23092 22244 -23028
rect 22308 -23092 22328 -23028
rect 16956 -23108 22328 -23092
rect 16956 -23172 22244 -23108
rect 22308 -23172 22328 -23108
rect 16956 -23188 22328 -23172
rect 16956 -23252 22244 -23188
rect 22308 -23252 22328 -23188
rect 16956 -23268 22328 -23252
rect 16956 -23332 22244 -23268
rect 22308 -23332 22328 -23268
rect 16956 -23348 22328 -23332
rect 16956 -23412 22244 -23348
rect 22308 -23412 22328 -23348
rect 16956 -23428 22328 -23412
rect 16956 -23492 22244 -23428
rect 22308 -23492 22328 -23428
rect 16956 -23508 22328 -23492
rect 16956 -23572 22244 -23508
rect 22308 -23572 22328 -23508
rect 16956 -23588 22328 -23572
rect 16956 -23652 22244 -23588
rect 22308 -23652 22328 -23588
rect 16956 -23668 22328 -23652
rect 16956 -23732 22244 -23668
rect 22308 -23732 22328 -23668
rect 16956 -23748 22328 -23732
rect 16956 -23812 22244 -23748
rect 22308 -23812 22328 -23748
rect 16956 -23828 22328 -23812
rect 16956 -23892 22244 -23828
rect 22308 -23892 22328 -23828
rect 16956 -23908 22328 -23892
rect 16956 -23972 22244 -23908
rect 22308 -23972 22328 -23908
rect 16956 -23988 22328 -23972
rect 16956 -24052 22244 -23988
rect 22308 -24052 22328 -23988
rect 16956 -24068 22328 -24052
rect 16956 -24132 22244 -24068
rect 22308 -24132 22328 -24068
rect 16956 -24148 22328 -24132
rect 16956 -24212 22244 -24148
rect 22308 -24212 22328 -24148
rect 16956 -24228 22328 -24212
rect 16956 -24292 22244 -24228
rect 22308 -24292 22328 -24228
rect 16956 -24308 22328 -24292
rect 16956 -24372 22244 -24308
rect 22308 -24372 22328 -24308
rect 16956 -24388 22328 -24372
rect 16956 -24452 22244 -24388
rect 22308 -24452 22328 -24388
rect 16956 -24468 22328 -24452
rect 16956 -24532 22244 -24468
rect 22308 -24532 22328 -24468
rect 16956 -24548 22328 -24532
rect 16956 -24612 22244 -24548
rect 22308 -24612 22328 -24548
rect 16956 -24628 22328 -24612
rect 16956 -24692 22244 -24628
rect 22308 -24692 22328 -24628
rect 16956 -24708 22328 -24692
rect 16956 -24772 22244 -24708
rect 22308 -24772 22328 -24708
rect 16956 -24788 22328 -24772
rect 16956 -24852 22244 -24788
rect 22308 -24852 22328 -24788
rect 16956 -24868 22328 -24852
rect 16956 -24932 22244 -24868
rect 22308 -24932 22328 -24868
rect 16956 -24948 22328 -24932
rect 16956 -25012 22244 -24948
rect 22308 -25012 22328 -24948
rect 16956 -25028 22328 -25012
rect 16956 -25092 22244 -25028
rect 22308 -25092 22328 -25028
rect 16956 -25108 22328 -25092
rect 16956 -25172 22244 -25108
rect 22308 -25172 22328 -25108
rect 16956 -25188 22328 -25172
rect 16956 -25252 22244 -25188
rect 22308 -25252 22328 -25188
rect 16956 -25268 22328 -25252
rect 16956 -25332 22244 -25268
rect 22308 -25332 22328 -25268
rect 16956 -25348 22328 -25332
rect 16956 -25412 22244 -25348
rect 22308 -25412 22328 -25348
rect 16956 -25428 22328 -25412
rect 16956 -25492 22244 -25428
rect 22308 -25492 22328 -25428
rect 16956 -25508 22328 -25492
rect 16956 -25572 22244 -25508
rect 22308 -25572 22328 -25508
rect 16956 -25588 22328 -25572
rect 16956 -25652 22244 -25588
rect 22308 -25652 22328 -25588
rect 16956 -25668 22328 -25652
rect 16956 -25732 22244 -25668
rect 22308 -25732 22328 -25668
rect 16956 -25748 22328 -25732
rect 16956 -25812 22244 -25748
rect 22308 -25812 22328 -25748
rect 16956 -25828 22328 -25812
rect 16956 -25892 22244 -25828
rect 22308 -25892 22328 -25828
rect 16956 -25908 22328 -25892
rect 16956 -25972 22244 -25908
rect 22308 -25972 22328 -25908
rect 16956 -25988 22328 -25972
rect 16956 -26052 22244 -25988
rect 22308 -26052 22328 -25988
rect 16956 -26068 22328 -26052
rect 16956 -26132 22244 -26068
rect 22308 -26132 22328 -26068
rect 16956 -26148 22328 -26132
rect 16956 -26212 22244 -26148
rect 22308 -26212 22328 -26148
rect 16956 -26228 22328 -26212
rect 16956 -26292 22244 -26228
rect 22308 -26292 22328 -26228
rect 16956 -26308 22328 -26292
rect 16956 -26372 22244 -26308
rect 22308 -26372 22328 -26308
rect 16956 -26388 22328 -26372
rect 16956 -26452 22244 -26388
rect 22308 -26452 22328 -26388
rect 16956 -26480 22328 -26452
rect 22568 -21428 27940 -21400
rect 22568 -21492 27856 -21428
rect 27920 -21492 27940 -21428
rect 22568 -21508 27940 -21492
rect 22568 -21572 27856 -21508
rect 27920 -21572 27940 -21508
rect 22568 -21588 27940 -21572
rect 22568 -21652 27856 -21588
rect 27920 -21652 27940 -21588
rect 22568 -21668 27940 -21652
rect 22568 -21732 27856 -21668
rect 27920 -21732 27940 -21668
rect 22568 -21748 27940 -21732
rect 22568 -21812 27856 -21748
rect 27920 -21812 27940 -21748
rect 22568 -21828 27940 -21812
rect 22568 -21892 27856 -21828
rect 27920 -21892 27940 -21828
rect 22568 -21908 27940 -21892
rect 22568 -21972 27856 -21908
rect 27920 -21972 27940 -21908
rect 22568 -21988 27940 -21972
rect 22568 -22052 27856 -21988
rect 27920 -22052 27940 -21988
rect 22568 -22068 27940 -22052
rect 22568 -22132 27856 -22068
rect 27920 -22132 27940 -22068
rect 22568 -22148 27940 -22132
rect 22568 -22212 27856 -22148
rect 27920 -22212 27940 -22148
rect 22568 -22228 27940 -22212
rect 22568 -22292 27856 -22228
rect 27920 -22292 27940 -22228
rect 22568 -22308 27940 -22292
rect 22568 -22372 27856 -22308
rect 27920 -22372 27940 -22308
rect 22568 -22388 27940 -22372
rect 22568 -22452 27856 -22388
rect 27920 -22452 27940 -22388
rect 22568 -22468 27940 -22452
rect 22568 -22532 27856 -22468
rect 27920 -22532 27940 -22468
rect 22568 -22548 27940 -22532
rect 22568 -22612 27856 -22548
rect 27920 -22612 27940 -22548
rect 22568 -22628 27940 -22612
rect 22568 -22692 27856 -22628
rect 27920 -22692 27940 -22628
rect 22568 -22708 27940 -22692
rect 22568 -22772 27856 -22708
rect 27920 -22772 27940 -22708
rect 22568 -22788 27940 -22772
rect 22568 -22852 27856 -22788
rect 27920 -22852 27940 -22788
rect 22568 -22868 27940 -22852
rect 22568 -22932 27856 -22868
rect 27920 -22932 27940 -22868
rect 22568 -22948 27940 -22932
rect 22568 -23012 27856 -22948
rect 27920 -23012 27940 -22948
rect 22568 -23028 27940 -23012
rect 22568 -23092 27856 -23028
rect 27920 -23092 27940 -23028
rect 22568 -23108 27940 -23092
rect 22568 -23172 27856 -23108
rect 27920 -23172 27940 -23108
rect 22568 -23188 27940 -23172
rect 22568 -23252 27856 -23188
rect 27920 -23252 27940 -23188
rect 22568 -23268 27940 -23252
rect 22568 -23332 27856 -23268
rect 27920 -23332 27940 -23268
rect 22568 -23348 27940 -23332
rect 22568 -23412 27856 -23348
rect 27920 -23412 27940 -23348
rect 22568 -23428 27940 -23412
rect 22568 -23492 27856 -23428
rect 27920 -23492 27940 -23428
rect 22568 -23508 27940 -23492
rect 22568 -23572 27856 -23508
rect 27920 -23572 27940 -23508
rect 22568 -23588 27940 -23572
rect 22568 -23652 27856 -23588
rect 27920 -23652 27940 -23588
rect 22568 -23668 27940 -23652
rect 22568 -23732 27856 -23668
rect 27920 -23732 27940 -23668
rect 22568 -23748 27940 -23732
rect 22568 -23812 27856 -23748
rect 27920 -23812 27940 -23748
rect 22568 -23828 27940 -23812
rect 22568 -23892 27856 -23828
rect 27920 -23892 27940 -23828
rect 22568 -23908 27940 -23892
rect 22568 -23972 27856 -23908
rect 27920 -23972 27940 -23908
rect 22568 -23988 27940 -23972
rect 22568 -24052 27856 -23988
rect 27920 -24052 27940 -23988
rect 22568 -24068 27940 -24052
rect 22568 -24132 27856 -24068
rect 27920 -24132 27940 -24068
rect 22568 -24148 27940 -24132
rect 22568 -24212 27856 -24148
rect 27920 -24212 27940 -24148
rect 22568 -24228 27940 -24212
rect 22568 -24292 27856 -24228
rect 27920 -24292 27940 -24228
rect 22568 -24308 27940 -24292
rect 22568 -24372 27856 -24308
rect 27920 -24372 27940 -24308
rect 22568 -24388 27940 -24372
rect 22568 -24452 27856 -24388
rect 27920 -24452 27940 -24388
rect 22568 -24468 27940 -24452
rect 22568 -24532 27856 -24468
rect 27920 -24532 27940 -24468
rect 22568 -24548 27940 -24532
rect 22568 -24612 27856 -24548
rect 27920 -24612 27940 -24548
rect 22568 -24628 27940 -24612
rect 22568 -24692 27856 -24628
rect 27920 -24692 27940 -24628
rect 22568 -24708 27940 -24692
rect 22568 -24772 27856 -24708
rect 27920 -24772 27940 -24708
rect 22568 -24788 27940 -24772
rect 22568 -24852 27856 -24788
rect 27920 -24852 27940 -24788
rect 22568 -24868 27940 -24852
rect 22568 -24932 27856 -24868
rect 27920 -24932 27940 -24868
rect 22568 -24948 27940 -24932
rect 22568 -25012 27856 -24948
rect 27920 -25012 27940 -24948
rect 22568 -25028 27940 -25012
rect 22568 -25092 27856 -25028
rect 27920 -25092 27940 -25028
rect 22568 -25108 27940 -25092
rect 22568 -25172 27856 -25108
rect 27920 -25172 27940 -25108
rect 22568 -25188 27940 -25172
rect 22568 -25252 27856 -25188
rect 27920 -25252 27940 -25188
rect 22568 -25268 27940 -25252
rect 22568 -25332 27856 -25268
rect 27920 -25332 27940 -25268
rect 22568 -25348 27940 -25332
rect 22568 -25412 27856 -25348
rect 27920 -25412 27940 -25348
rect 22568 -25428 27940 -25412
rect 22568 -25492 27856 -25428
rect 27920 -25492 27940 -25428
rect 22568 -25508 27940 -25492
rect 22568 -25572 27856 -25508
rect 27920 -25572 27940 -25508
rect 22568 -25588 27940 -25572
rect 22568 -25652 27856 -25588
rect 27920 -25652 27940 -25588
rect 22568 -25668 27940 -25652
rect 22568 -25732 27856 -25668
rect 27920 -25732 27940 -25668
rect 22568 -25748 27940 -25732
rect 22568 -25812 27856 -25748
rect 27920 -25812 27940 -25748
rect 22568 -25828 27940 -25812
rect 22568 -25892 27856 -25828
rect 27920 -25892 27940 -25828
rect 22568 -25908 27940 -25892
rect 22568 -25972 27856 -25908
rect 27920 -25972 27940 -25908
rect 22568 -25988 27940 -25972
rect 22568 -26052 27856 -25988
rect 27920 -26052 27940 -25988
rect 22568 -26068 27940 -26052
rect 22568 -26132 27856 -26068
rect 27920 -26132 27940 -26068
rect 22568 -26148 27940 -26132
rect 22568 -26212 27856 -26148
rect 27920 -26212 27940 -26148
rect 22568 -26228 27940 -26212
rect 22568 -26292 27856 -26228
rect 27920 -26292 27940 -26228
rect 22568 -26308 27940 -26292
rect 22568 -26372 27856 -26308
rect 27920 -26372 27940 -26308
rect 22568 -26388 27940 -26372
rect 22568 -26452 27856 -26388
rect 27920 -26452 27940 -26388
rect 22568 -26480 27940 -26452
rect 28180 -21428 33552 -21400
rect 28180 -21492 33468 -21428
rect 33532 -21492 33552 -21428
rect 28180 -21508 33552 -21492
rect 28180 -21572 33468 -21508
rect 33532 -21572 33552 -21508
rect 28180 -21588 33552 -21572
rect 28180 -21652 33468 -21588
rect 33532 -21652 33552 -21588
rect 28180 -21668 33552 -21652
rect 28180 -21732 33468 -21668
rect 33532 -21732 33552 -21668
rect 28180 -21748 33552 -21732
rect 28180 -21812 33468 -21748
rect 33532 -21812 33552 -21748
rect 28180 -21828 33552 -21812
rect 28180 -21892 33468 -21828
rect 33532 -21892 33552 -21828
rect 28180 -21908 33552 -21892
rect 28180 -21972 33468 -21908
rect 33532 -21972 33552 -21908
rect 28180 -21988 33552 -21972
rect 28180 -22052 33468 -21988
rect 33532 -22052 33552 -21988
rect 28180 -22068 33552 -22052
rect 28180 -22132 33468 -22068
rect 33532 -22132 33552 -22068
rect 28180 -22148 33552 -22132
rect 28180 -22212 33468 -22148
rect 33532 -22212 33552 -22148
rect 28180 -22228 33552 -22212
rect 28180 -22292 33468 -22228
rect 33532 -22292 33552 -22228
rect 28180 -22308 33552 -22292
rect 28180 -22372 33468 -22308
rect 33532 -22372 33552 -22308
rect 28180 -22388 33552 -22372
rect 28180 -22452 33468 -22388
rect 33532 -22452 33552 -22388
rect 28180 -22468 33552 -22452
rect 28180 -22532 33468 -22468
rect 33532 -22532 33552 -22468
rect 28180 -22548 33552 -22532
rect 28180 -22612 33468 -22548
rect 33532 -22612 33552 -22548
rect 28180 -22628 33552 -22612
rect 28180 -22692 33468 -22628
rect 33532 -22692 33552 -22628
rect 28180 -22708 33552 -22692
rect 28180 -22772 33468 -22708
rect 33532 -22772 33552 -22708
rect 28180 -22788 33552 -22772
rect 28180 -22852 33468 -22788
rect 33532 -22852 33552 -22788
rect 28180 -22868 33552 -22852
rect 28180 -22932 33468 -22868
rect 33532 -22932 33552 -22868
rect 28180 -22948 33552 -22932
rect 28180 -23012 33468 -22948
rect 33532 -23012 33552 -22948
rect 28180 -23028 33552 -23012
rect 28180 -23092 33468 -23028
rect 33532 -23092 33552 -23028
rect 28180 -23108 33552 -23092
rect 28180 -23172 33468 -23108
rect 33532 -23172 33552 -23108
rect 28180 -23188 33552 -23172
rect 28180 -23252 33468 -23188
rect 33532 -23252 33552 -23188
rect 28180 -23268 33552 -23252
rect 28180 -23332 33468 -23268
rect 33532 -23332 33552 -23268
rect 28180 -23348 33552 -23332
rect 28180 -23412 33468 -23348
rect 33532 -23412 33552 -23348
rect 28180 -23428 33552 -23412
rect 28180 -23492 33468 -23428
rect 33532 -23492 33552 -23428
rect 28180 -23508 33552 -23492
rect 28180 -23572 33468 -23508
rect 33532 -23572 33552 -23508
rect 28180 -23588 33552 -23572
rect 28180 -23652 33468 -23588
rect 33532 -23652 33552 -23588
rect 28180 -23668 33552 -23652
rect 28180 -23732 33468 -23668
rect 33532 -23732 33552 -23668
rect 28180 -23748 33552 -23732
rect 28180 -23812 33468 -23748
rect 33532 -23812 33552 -23748
rect 28180 -23828 33552 -23812
rect 28180 -23892 33468 -23828
rect 33532 -23892 33552 -23828
rect 28180 -23908 33552 -23892
rect 28180 -23972 33468 -23908
rect 33532 -23972 33552 -23908
rect 28180 -23988 33552 -23972
rect 28180 -24052 33468 -23988
rect 33532 -24052 33552 -23988
rect 28180 -24068 33552 -24052
rect 28180 -24132 33468 -24068
rect 33532 -24132 33552 -24068
rect 28180 -24148 33552 -24132
rect 28180 -24212 33468 -24148
rect 33532 -24212 33552 -24148
rect 28180 -24228 33552 -24212
rect 28180 -24292 33468 -24228
rect 33532 -24292 33552 -24228
rect 28180 -24308 33552 -24292
rect 28180 -24372 33468 -24308
rect 33532 -24372 33552 -24308
rect 28180 -24388 33552 -24372
rect 28180 -24452 33468 -24388
rect 33532 -24452 33552 -24388
rect 28180 -24468 33552 -24452
rect 28180 -24532 33468 -24468
rect 33532 -24532 33552 -24468
rect 28180 -24548 33552 -24532
rect 28180 -24612 33468 -24548
rect 33532 -24612 33552 -24548
rect 28180 -24628 33552 -24612
rect 28180 -24692 33468 -24628
rect 33532 -24692 33552 -24628
rect 28180 -24708 33552 -24692
rect 28180 -24772 33468 -24708
rect 33532 -24772 33552 -24708
rect 28180 -24788 33552 -24772
rect 28180 -24852 33468 -24788
rect 33532 -24852 33552 -24788
rect 28180 -24868 33552 -24852
rect 28180 -24932 33468 -24868
rect 33532 -24932 33552 -24868
rect 28180 -24948 33552 -24932
rect 28180 -25012 33468 -24948
rect 33532 -25012 33552 -24948
rect 28180 -25028 33552 -25012
rect 28180 -25092 33468 -25028
rect 33532 -25092 33552 -25028
rect 28180 -25108 33552 -25092
rect 28180 -25172 33468 -25108
rect 33532 -25172 33552 -25108
rect 28180 -25188 33552 -25172
rect 28180 -25252 33468 -25188
rect 33532 -25252 33552 -25188
rect 28180 -25268 33552 -25252
rect 28180 -25332 33468 -25268
rect 33532 -25332 33552 -25268
rect 28180 -25348 33552 -25332
rect 28180 -25412 33468 -25348
rect 33532 -25412 33552 -25348
rect 28180 -25428 33552 -25412
rect 28180 -25492 33468 -25428
rect 33532 -25492 33552 -25428
rect 28180 -25508 33552 -25492
rect 28180 -25572 33468 -25508
rect 33532 -25572 33552 -25508
rect 28180 -25588 33552 -25572
rect 28180 -25652 33468 -25588
rect 33532 -25652 33552 -25588
rect 28180 -25668 33552 -25652
rect 28180 -25732 33468 -25668
rect 33532 -25732 33552 -25668
rect 28180 -25748 33552 -25732
rect 28180 -25812 33468 -25748
rect 33532 -25812 33552 -25748
rect 28180 -25828 33552 -25812
rect 28180 -25892 33468 -25828
rect 33532 -25892 33552 -25828
rect 28180 -25908 33552 -25892
rect 28180 -25972 33468 -25908
rect 33532 -25972 33552 -25908
rect 28180 -25988 33552 -25972
rect 28180 -26052 33468 -25988
rect 33532 -26052 33552 -25988
rect 28180 -26068 33552 -26052
rect 28180 -26132 33468 -26068
rect 33532 -26132 33552 -26068
rect 28180 -26148 33552 -26132
rect 28180 -26212 33468 -26148
rect 33532 -26212 33552 -26148
rect 28180 -26228 33552 -26212
rect 28180 -26292 33468 -26228
rect 33532 -26292 33552 -26228
rect 28180 -26308 33552 -26292
rect 28180 -26372 33468 -26308
rect 33532 -26372 33552 -26308
rect 28180 -26388 33552 -26372
rect 28180 -26452 33468 -26388
rect 33532 -26452 33552 -26388
rect 28180 -26480 33552 -26452
rect 33792 -21428 39164 -21400
rect 33792 -21492 39080 -21428
rect 39144 -21492 39164 -21428
rect 33792 -21508 39164 -21492
rect 33792 -21572 39080 -21508
rect 39144 -21572 39164 -21508
rect 33792 -21588 39164 -21572
rect 33792 -21652 39080 -21588
rect 39144 -21652 39164 -21588
rect 33792 -21668 39164 -21652
rect 33792 -21732 39080 -21668
rect 39144 -21732 39164 -21668
rect 33792 -21748 39164 -21732
rect 33792 -21812 39080 -21748
rect 39144 -21812 39164 -21748
rect 33792 -21828 39164 -21812
rect 33792 -21892 39080 -21828
rect 39144 -21892 39164 -21828
rect 33792 -21908 39164 -21892
rect 33792 -21972 39080 -21908
rect 39144 -21972 39164 -21908
rect 33792 -21988 39164 -21972
rect 33792 -22052 39080 -21988
rect 39144 -22052 39164 -21988
rect 33792 -22068 39164 -22052
rect 33792 -22132 39080 -22068
rect 39144 -22132 39164 -22068
rect 33792 -22148 39164 -22132
rect 33792 -22212 39080 -22148
rect 39144 -22212 39164 -22148
rect 33792 -22228 39164 -22212
rect 33792 -22292 39080 -22228
rect 39144 -22292 39164 -22228
rect 33792 -22308 39164 -22292
rect 33792 -22372 39080 -22308
rect 39144 -22372 39164 -22308
rect 33792 -22388 39164 -22372
rect 33792 -22452 39080 -22388
rect 39144 -22452 39164 -22388
rect 33792 -22468 39164 -22452
rect 33792 -22532 39080 -22468
rect 39144 -22532 39164 -22468
rect 33792 -22548 39164 -22532
rect 33792 -22612 39080 -22548
rect 39144 -22612 39164 -22548
rect 33792 -22628 39164 -22612
rect 33792 -22692 39080 -22628
rect 39144 -22692 39164 -22628
rect 33792 -22708 39164 -22692
rect 33792 -22772 39080 -22708
rect 39144 -22772 39164 -22708
rect 33792 -22788 39164 -22772
rect 33792 -22852 39080 -22788
rect 39144 -22852 39164 -22788
rect 33792 -22868 39164 -22852
rect 33792 -22932 39080 -22868
rect 39144 -22932 39164 -22868
rect 33792 -22948 39164 -22932
rect 33792 -23012 39080 -22948
rect 39144 -23012 39164 -22948
rect 33792 -23028 39164 -23012
rect 33792 -23092 39080 -23028
rect 39144 -23092 39164 -23028
rect 33792 -23108 39164 -23092
rect 33792 -23172 39080 -23108
rect 39144 -23172 39164 -23108
rect 33792 -23188 39164 -23172
rect 33792 -23252 39080 -23188
rect 39144 -23252 39164 -23188
rect 33792 -23268 39164 -23252
rect 33792 -23332 39080 -23268
rect 39144 -23332 39164 -23268
rect 33792 -23348 39164 -23332
rect 33792 -23412 39080 -23348
rect 39144 -23412 39164 -23348
rect 33792 -23428 39164 -23412
rect 33792 -23492 39080 -23428
rect 39144 -23492 39164 -23428
rect 33792 -23508 39164 -23492
rect 33792 -23572 39080 -23508
rect 39144 -23572 39164 -23508
rect 33792 -23588 39164 -23572
rect 33792 -23652 39080 -23588
rect 39144 -23652 39164 -23588
rect 33792 -23668 39164 -23652
rect 33792 -23732 39080 -23668
rect 39144 -23732 39164 -23668
rect 33792 -23748 39164 -23732
rect 33792 -23812 39080 -23748
rect 39144 -23812 39164 -23748
rect 33792 -23828 39164 -23812
rect 33792 -23892 39080 -23828
rect 39144 -23892 39164 -23828
rect 33792 -23908 39164 -23892
rect 33792 -23972 39080 -23908
rect 39144 -23972 39164 -23908
rect 33792 -23988 39164 -23972
rect 33792 -24052 39080 -23988
rect 39144 -24052 39164 -23988
rect 33792 -24068 39164 -24052
rect 33792 -24132 39080 -24068
rect 39144 -24132 39164 -24068
rect 33792 -24148 39164 -24132
rect 33792 -24212 39080 -24148
rect 39144 -24212 39164 -24148
rect 33792 -24228 39164 -24212
rect 33792 -24292 39080 -24228
rect 39144 -24292 39164 -24228
rect 33792 -24308 39164 -24292
rect 33792 -24372 39080 -24308
rect 39144 -24372 39164 -24308
rect 33792 -24388 39164 -24372
rect 33792 -24452 39080 -24388
rect 39144 -24452 39164 -24388
rect 33792 -24468 39164 -24452
rect 33792 -24532 39080 -24468
rect 39144 -24532 39164 -24468
rect 33792 -24548 39164 -24532
rect 33792 -24612 39080 -24548
rect 39144 -24612 39164 -24548
rect 33792 -24628 39164 -24612
rect 33792 -24692 39080 -24628
rect 39144 -24692 39164 -24628
rect 33792 -24708 39164 -24692
rect 33792 -24772 39080 -24708
rect 39144 -24772 39164 -24708
rect 33792 -24788 39164 -24772
rect 33792 -24852 39080 -24788
rect 39144 -24852 39164 -24788
rect 33792 -24868 39164 -24852
rect 33792 -24932 39080 -24868
rect 39144 -24932 39164 -24868
rect 33792 -24948 39164 -24932
rect 33792 -25012 39080 -24948
rect 39144 -25012 39164 -24948
rect 33792 -25028 39164 -25012
rect 33792 -25092 39080 -25028
rect 39144 -25092 39164 -25028
rect 33792 -25108 39164 -25092
rect 33792 -25172 39080 -25108
rect 39144 -25172 39164 -25108
rect 33792 -25188 39164 -25172
rect 33792 -25252 39080 -25188
rect 39144 -25252 39164 -25188
rect 33792 -25268 39164 -25252
rect 33792 -25332 39080 -25268
rect 39144 -25332 39164 -25268
rect 33792 -25348 39164 -25332
rect 33792 -25412 39080 -25348
rect 39144 -25412 39164 -25348
rect 33792 -25428 39164 -25412
rect 33792 -25492 39080 -25428
rect 39144 -25492 39164 -25428
rect 33792 -25508 39164 -25492
rect 33792 -25572 39080 -25508
rect 39144 -25572 39164 -25508
rect 33792 -25588 39164 -25572
rect 33792 -25652 39080 -25588
rect 39144 -25652 39164 -25588
rect 33792 -25668 39164 -25652
rect 33792 -25732 39080 -25668
rect 39144 -25732 39164 -25668
rect 33792 -25748 39164 -25732
rect 33792 -25812 39080 -25748
rect 39144 -25812 39164 -25748
rect 33792 -25828 39164 -25812
rect 33792 -25892 39080 -25828
rect 39144 -25892 39164 -25828
rect 33792 -25908 39164 -25892
rect 33792 -25972 39080 -25908
rect 39144 -25972 39164 -25908
rect 33792 -25988 39164 -25972
rect 33792 -26052 39080 -25988
rect 39144 -26052 39164 -25988
rect 33792 -26068 39164 -26052
rect 33792 -26132 39080 -26068
rect 39144 -26132 39164 -26068
rect 33792 -26148 39164 -26132
rect 33792 -26212 39080 -26148
rect 39144 -26212 39164 -26148
rect 33792 -26228 39164 -26212
rect 33792 -26292 39080 -26228
rect 39144 -26292 39164 -26228
rect 33792 -26308 39164 -26292
rect 33792 -26372 39080 -26308
rect 39144 -26372 39164 -26308
rect 33792 -26388 39164 -26372
rect 33792 -26452 39080 -26388
rect 39144 -26452 39164 -26388
rect 33792 -26480 39164 -26452
rect -39164 -26748 -33792 -26720
rect -39164 -26812 -33876 -26748
rect -33812 -26812 -33792 -26748
rect -39164 -26828 -33792 -26812
rect -39164 -26892 -33876 -26828
rect -33812 -26892 -33792 -26828
rect -39164 -26908 -33792 -26892
rect -39164 -26972 -33876 -26908
rect -33812 -26972 -33792 -26908
rect -39164 -26988 -33792 -26972
rect -39164 -27052 -33876 -26988
rect -33812 -27052 -33792 -26988
rect -39164 -27068 -33792 -27052
rect -39164 -27132 -33876 -27068
rect -33812 -27132 -33792 -27068
rect -39164 -27148 -33792 -27132
rect -39164 -27212 -33876 -27148
rect -33812 -27212 -33792 -27148
rect -39164 -27228 -33792 -27212
rect -39164 -27292 -33876 -27228
rect -33812 -27292 -33792 -27228
rect -39164 -27308 -33792 -27292
rect -39164 -27372 -33876 -27308
rect -33812 -27372 -33792 -27308
rect -39164 -27388 -33792 -27372
rect -39164 -27452 -33876 -27388
rect -33812 -27452 -33792 -27388
rect -39164 -27468 -33792 -27452
rect -39164 -27532 -33876 -27468
rect -33812 -27532 -33792 -27468
rect -39164 -27548 -33792 -27532
rect -39164 -27612 -33876 -27548
rect -33812 -27612 -33792 -27548
rect -39164 -27628 -33792 -27612
rect -39164 -27692 -33876 -27628
rect -33812 -27692 -33792 -27628
rect -39164 -27708 -33792 -27692
rect -39164 -27772 -33876 -27708
rect -33812 -27772 -33792 -27708
rect -39164 -27788 -33792 -27772
rect -39164 -27852 -33876 -27788
rect -33812 -27852 -33792 -27788
rect -39164 -27868 -33792 -27852
rect -39164 -27932 -33876 -27868
rect -33812 -27932 -33792 -27868
rect -39164 -27948 -33792 -27932
rect -39164 -28012 -33876 -27948
rect -33812 -28012 -33792 -27948
rect -39164 -28028 -33792 -28012
rect -39164 -28092 -33876 -28028
rect -33812 -28092 -33792 -28028
rect -39164 -28108 -33792 -28092
rect -39164 -28172 -33876 -28108
rect -33812 -28172 -33792 -28108
rect -39164 -28188 -33792 -28172
rect -39164 -28252 -33876 -28188
rect -33812 -28252 -33792 -28188
rect -39164 -28268 -33792 -28252
rect -39164 -28332 -33876 -28268
rect -33812 -28332 -33792 -28268
rect -39164 -28348 -33792 -28332
rect -39164 -28412 -33876 -28348
rect -33812 -28412 -33792 -28348
rect -39164 -28428 -33792 -28412
rect -39164 -28492 -33876 -28428
rect -33812 -28492 -33792 -28428
rect -39164 -28508 -33792 -28492
rect -39164 -28572 -33876 -28508
rect -33812 -28572 -33792 -28508
rect -39164 -28588 -33792 -28572
rect -39164 -28652 -33876 -28588
rect -33812 -28652 -33792 -28588
rect -39164 -28668 -33792 -28652
rect -39164 -28732 -33876 -28668
rect -33812 -28732 -33792 -28668
rect -39164 -28748 -33792 -28732
rect -39164 -28812 -33876 -28748
rect -33812 -28812 -33792 -28748
rect -39164 -28828 -33792 -28812
rect -39164 -28892 -33876 -28828
rect -33812 -28892 -33792 -28828
rect -39164 -28908 -33792 -28892
rect -39164 -28972 -33876 -28908
rect -33812 -28972 -33792 -28908
rect -39164 -28988 -33792 -28972
rect -39164 -29052 -33876 -28988
rect -33812 -29052 -33792 -28988
rect -39164 -29068 -33792 -29052
rect -39164 -29132 -33876 -29068
rect -33812 -29132 -33792 -29068
rect -39164 -29148 -33792 -29132
rect -39164 -29212 -33876 -29148
rect -33812 -29212 -33792 -29148
rect -39164 -29228 -33792 -29212
rect -39164 -29292 -33876 -29228
rect -33812 -29292 -33792 -29228
rect -39164 -29308 -33792 -29292
rect -39164 -29372 -33876 -29308
rect -33812 -29372 -33792 -29308
rect -39164 -29388 -33792 -29372
rect -39164 -29452 -33876 -29388
rect -33812 -29452 -33792 -29388
rect -39164 -29468 -33792 -29452
rect -39164 -29532 -33876 -29468
rect -33812 -29532 -33792 -29468
rect -39164 -29548 -33792 -29532
rect -39164 -29612 -33876 -29548
rect -33812 -29612 -33792 -29548
rect -39164 -29628 -33792 -29612
rect -39164 -29692 -33876 -29628
rect -33812 -29692 -33792 -29628
rect -39164 -29708 -33792 -29692
rect -39164 -29772 -33876 -29708
rect -33812 -29772 -33792 -29708
rect -39164 -29788 -33792 -29772
rect -39164 -29852 -33876 -29788
rect -33812 -29852 -33792 -29788
rect -39164 -29868 -33792 -29852
rect -39164 -29932 -33876 -29868
rect -33812 -29932 -33792 -29868
rect -39164 -29948 -33792 -29932
rect -39164 -30012 -33876 -29948
rect -33812 -30012 -33792 -29948
rect -39164 -30028 -33792 -30012
rect -39164 -30092 -33876 -30028
rect -33812 -30092 -33792 -30028
rect -39164 -30108 -33792 -30092
rect -39164 -30172 -33876 -30108
rect -33812 -30172 -33792 -30108
rect -39164 -30188 -33792 -30172
rect -39164 -30252 -33876 -30188
rect -33812 -30252 -33792 -30188
rect -39164 -30268 -33792 -30252
rect -39164 -30332 -33876 -30268
rect -33812 -30332 -33792 -30268
rect -39164 -30348 -33792 -30332
rect -39164 -30412 -33876 -30348
rect -33812 -30412 -33792 -30348
rect -39164 -30428 -33792 -30412
rect -39164 -30492 -33876 -30428
rect -33812 -30492 -33792 -30428
rect -39164 -30508 -33792 -30492
rect -39164 -30572 -33876 -30508
rect -33812 -30572 -33792 -30508
rect -39164 -30588 -33792 -30572
rect -39164 -30652 -33876 -30588
rect -33812 -30652 -33792 -30588
rect -39164 -30668 -33792 -30652
rect -39164 -30732 -33876 -30668
rect -33812 -30732 -33792 -30668
rect -39164 -30748 -33792 -30732
rect -39164 -30812 -33876 -30748
rect -33812 -30812 -33792 -30748
rect -39164 -30828 -33792 -30812
rect -39164 -30892 -33876 -30828
rect -33812 -30892 -33792 -30828
rect -39164 -30908 -33792 -30892
rect -39164 -30972 -33876 -30908
rect -33812 -30972 -33792 -30908
rect -39164 -30988 -33792 -30972
rect -39164 -31052 -33876 -30988
rect -33812 -31052 -33792 -30988
rect -39164 -31068 -33792 -31052
rect -39164 -31132 -33876 -31068
rect -33812 -31132 -33792 -31068
rect -39164 -31148 -33792 -31132
rect -39164 -31212 -33876 -31148
rect -33812 -31212 -33792 -31148
rect -39164 -31228 -33792 -31212
rect -39164 -31292 -33876 -31228
rect -33812 -31292 -33792 -31228
rect -39164 -31308 -33792 -31292
rect -39164 -31372 -33876 -31308
rect -33812 -31372 -33792 -31308
rect -39164 -31388 -33792 -31372
rect -39164 -31452 -33876 -31388
rect -33812 -31452 -33792 -31388
rect -39164 -31468 -33792 -31452
rect -39164 -31532 -33876 -31468
rect -33812 -31532 -33792 -31468
rect -39164 -31548 -33792 -31532
rect -39164 -31612 -33876 -31548
rect -33812 -31612 -33792 -31548
rect -39164 -31628 -33792 -31612
rect -39164 -31692 -33876 -31628
rect -33812 -31692 -33792 -31628
rect -39164 -31708 -33792 -31692
rect -39164 -31772 -33876 -31708
rect -33812 -31772 -33792 -31708
rect -39164 -31800 -33792 -31772
rect -33552 -26748 -28180 -26720
rect -33552 -26812 -28264 -26748
rect -28200 -26812 -28180 -26748
rect -33552 -26828 -28180 -26812
rect -33552 -26892 -28264 -26828
rect -28200 -26892 -28180 -26828
rect -33552 -26908 -28180 -26892
rect -33552 -26972 -28264 -26908
rect -28200 -26972 -28180 -26908
rect -33552 -26988 -28180 -26972
rect -33552 -27052 -28264 -26988
rect -28200 -27052 -28180 -26988
rect -33552 -27068 -28180 -27052
rect -33552 -27132 -28264 -27068
rect -28200 -27132 -28180 -27068
rect -33552 -27148 -28180 -27132
rect -33552 -27212 -28264 -27148
rect -28200 -27212 -28180 -27148
rect -33552 -27228 -28180 -27212
rect -33552 -27292 -28264 -27228
rect -28200 -27292 -28180 -27228
rect -33552 -27308 -28180 -27292
rect -33552 -27372 -28264 -27308
rect -28200 -27372 -28180 -27308
rect -33552 -27388 -28180 -27372
rect -33552 -27452 -28264 -27388
rect -28200 -27452 -28180 -27388
rect -33552 -27468 -28180 -27452
rect -33552 -27532 -28264 -27468
rect -28200 -27532 -28180 -27468
rect -33552 -27548 -28180 -27532
rect -33552 -27612 -28264 -27548
rect -28200 -27612 -28180 -27548
rect -33552 -27628 -28180 -27612
rect -33552 -27692 -28264 -27628
rect -28200 -27692 -28180 -27628
rect -33552 -27708 -28180 -27692
rect -33552 -27772 -28264 -27708
rect -28200 -27772 -28180 -27708
rect -33552 -27788 -28180 -27772
rect -33552 -27852 -28264 -27788
rect -28200 -27852 -28180 -27788
rect -33552 -27868 -28180 -27852
rect -33552 -27932 -28264 -27868
rect -28200 -27932 -28180 -27868
rect -33552 -27948 -28180 -27932
rect -33552 -28012 -28264 -27948
rect -28200 -28012 -28180 -27948
rect -33552 -28028 -28180 -28012
rect -33552 -28092 -28264 -28028
rect -28200 -28092 -28180 -28028
rect -33552 -28108 -28180 -28092
rect -33552 -28172 -28264 -28108
rect -28200 -28172 -28180 -28108
rect -33552 -28188 -28180 -28172
rect -33552 -28252 -28264 -28188
rect -28200 -28252 -28180 -28188
rect -33552 -28268 -28180 -28252
rect -33552 -28332 -28264 -28268
rect -28200 -28332 -28180 -28268
rect -33552 -28348 -28180 -28332
rect -33552 -28412 -28264 -28348
rect -28200 -28412 -28180 -28348
rect -33552 -28428 -28180 -28412
rect -33552 -28492 -28264 -28428
rect -28200 -28492 -28180 -28428
rect -33552 -28508 -28180 -28492
rect -33552 -28572 -28264 -28508
rect -28200 -28572 -28180 -28508
rect -33552 -28588 -28180 -28572
rect -33552 -28652 -28264 -28588
rect -28200 -28652 -28180 -28588
rect -33552 -28668 -28180 -28652
rect -33552 -28732 -28264 -28668
rect -28200 -28732 -28180 -28668
rect -33552 -28748 -28180 -28732
rect -33552 -28812 -28264 -28748
rect -28200 -28812 -28180 -28748
rect -33552 -28828 -28180 -28812
rect -33552 -28892 -28264 -28828
rect -28200 -28892 -28180 -28828
rect -33552 -28908 -28180 -28892
rect -33552 -28972 -28264 -28908
rect -28200 -28972 -28180 -28908
rect -33552 -28988 -28180 -28972
rect -33552 -29052 -28264 -28988
rect -28200 -29052 -28180 -28988
rect -33552 -29068 -28180 -29052
rect -33552 -29132 -28264 -29068
rect -28200 -29132 -28180 -29068
rect -33552 -29148 -28180 -29132
rect -33552 -29212 -28264 -29148
rect -28200 -29212 -28180 -29148
rect -33552 -29228 -28180 -29212
rect -33552 -29292 -28264 -29228
rect -28200 -29292 -28180 -29228
rect -33552 -29308 -28180 -29292
rect -33552 -29372 -28264 -29308
rect -28200 -29372 -28180 -29308
rect -33552 -29388 -28180 -29372
rect -33552 -29452 -28264 -29388
rect -28200 -29452 -28180 -29388
rect -33552 -29468 -28180 -29452
rect -33552 -29532 -28264 -29468
rect -28200 -29532 -28180 -29468
rect -33552 -29548 -28180 -29532
rect -33552 -29612 -28264 -29548
rect -28200 -29612 -28180 -29548
rect -33552 -29628 -28180 -29612
rect -33552 -29692 -28264 -29628
rect -28200 -29692 -28180 -29628
rect -33552 -29708 -28180 -29692
rect -33552 -29772 -28264 -29708
rect -28200 -29772 -28180 -29708
rect -33552 -29788 -28180 -29772
rect -33552 -29852 -28264 -29788
rect -28200 -29852 -28180 -29788
rect -33552 -29868 -28180 -29852
rect -33552 -29932 -28264 -29868
rect -28200 -29932 -28180 -29868
rect -33552 -29948 -28180 -29932
rect -33552 -30012 -28264 -29948
rect -28200 -30012 -28180 -29948
rect -33552 -30028 -28180 -30012
rect -33552 -30092 -28264 -30028
rect -28200 -30092 -28180 -30028
rect -33552 -30108 -28180 -30092
rect -33552 -30172 -28264 -30108
rect -28200 -30172 -28180 -30108
rect -33552 -30188 -28180 -30172
rect -33552 -30252 -28264 -30188
rect -28200 -30252 -28180 -30188
rect -33552 -30268 -28180 -30252
rect -33552 -30332 -28264 -30268
rect -28200 -30332 -28180 -30268
rect -33552 -30348 -28180 -30332
rect -33552 -30412 -28264 -30348
rect -28200 -30412 -28180 -30348
rect -33552 -30428 -28180 -30412
rect -33552 -30492 -28264 -30428
rect -28200 -30492 -28180 -30428
rect -33552 -30508 -28180 -30492
rect -33552 -30572 -28264 -30508
rect -28200 -30572 -28180 -30508
rect -33552 -30588 -28180 -30572
rect -33552 -30652 -28264 -30588
rect -28200 -30652 -28180 -30588
rect -33552 -30668 -28180 -30652
rect -33552 -30732 -28264 -30668
rect -28200 -30732 -28180 -30668
rect -33552 -30748 -28180 -30732
rect -33552 -30812 -28264 -30748
rect -28200 -30812 -28180 -30748
rect -33552 -30828 -28180 -30812
rect -33552 -30892 -28264 -30828
rect -28200 -30892 -28180 -30828
rect -33552 -30908 -28180 -30892
rect -33552 -30972 -28264 -30908
rect -28200 -30972 -28180 -30908
rect -33552 -30988 -28180 -30972
rect -33552 -31052 -28264 -30988
rect -28200 -31052 -28180 -30988
rect -33552 -31068 -28180 -31052
rect -33552 -31132 -28264 -31068
rect -28200 -31132 -28180 -31068
rect -33552 -31148 -28180 -31132
rect -33552 -31212 -28264 -31148
rect -28200 -31212 -28180 -31148
rect -33552 -31228 -28180 -31212
rect -33552 -31292 -28264 -31228
rect -28200 -31292 -28180 -31228
rect -33552 -31308 -28180 -31292
rect -33552 -31372 -28264 -31308
rect -28200 -31372 -28180 -31308
rect -33552 -31388 -28180 -31372
rect -33552 -31452 -28264 -31388
rect -28200 -31452 -28180 -31388
rect -33552 -31468 -28180 -31452
rect -33552 -31532 -28264 -31468
rect -28200 -31532 -28180 -31468
rect -33552 -31548 -28180 -31532
rect -33552 -31612 -28264 -31548
rect -28200 -31612 -28180 -31548
rect -33552 -31628 -28180 -31612
rect -33552 -31692 -28264 -31628
rect -28200 -31692 -28180 -31628
rect -33552 -31708 -28180 -31692
rect -33552 -31772 -28264 -31708
rect -28200 -31772 -28180 -31708
rect -33552 -31800 -28180 -31772
rect -27940 -26748 -22568 -26720
rect -27940 -26812 -22652 -26748
rect -22588 -26812 -22568 -26748
rect -27940 -26828 -22568 -26812
rect -27940 -26892 -22652 -26828
rect -22588 -26892 -22568 -26828
rect -27940 -26908 -22568 -26892
rect -27940 -26972 -22652 -26908
rect -22588 -26972 -22568 -26908
rect -27940 -26988 -22568 -26972
rect -27940 -27052 -22652 -26988
rect -22588 -27052 -22568 -26988
rect -27940 -27068 -22568 -27052
rect -27940 -27132 -22652 -27068
rect -22588 -27132 -22568 -27068
rect -27940 -27148 -22568 -27132
rect -27940 -27212 -22652 -27148
rect -22588 -27212 -22568 -27148
rect -27940 -27228 -22568 -27212
rect -27940 -27292 -22652 -27228
rect -22588 -27292 -22568 -27228
rect -27940 -27308 -22568 -27292
rect -27940 -27372 -22652 -27308
rect -22588 -27372 -22568 -27308
rect -27940 -27388 -22568 -27372
rect -27940 -27452 -22652 -27388
rect -22588 -27452 -22568 -27388
rect -27940 -27468 -22568 -27452
rect -27940 -27532 -22652 -27468
rect -22588 -27532 -22568 -27468
rect -27940 -27548 -22568 -27532
rect -27940 -27612 -22652 -27548
rect -22588 -27612 -22568 -27548
rect -27940 -27628 -22568 -27612
rect -27940 -27692 -22652 -27628
rect -22588 -27692 -22568 -27628
rect -27940 -27708 -22568 -27692
rect -27940 -27772 -22652 -27708
rect -22588 -27772 -22568 -27708
rect -27940 -27788 -22568 -27772
rect -27940 -27852 -22652 -27788
rect -22588 -27852 -22568 -27788
rect -27940 -27868 -22568 -27852
rect -27940 -27932 -22652 -27868
rect -22588 -27932 -22568 -27868
rect -27940 -27948 -22568 -27932
rect -27940 -28012 -22652 -27948
rect -22588 -28012 -22568 -27948
rect -27940 -28028 -22568 -28012
rect -27940 -28092 -22652 -28028
rect -22588 -28092 -22568 -28028
rect -27940 -28108 -22568 -28092
rect -27940 -28172 -22652 -28108
rect -22588 -28172 -22568 -28108
rect -27940 -28188 -22568 -28172
rect -27940 -28252 -22652 -28188
rect -22588 -28252 -22568 -28188
rect -27940 -28268 -22568 -28252
rect -27940 -28332 -22652 -28268
rect -22588 -28332 -22568 -28268
rect -27940 -28348 -22568 -28332
rect -27940 -28412 -22652 -28348
rect -22588 -28412 -22568 -28348
rect -27940 -28428 -22568 -28412
rect -27940 -28492 -22652 -28428
rect -22588 -28492 -22568 -28428
rect -27940 -28508 -22568 -28492
rect -27940 -28572 -22652 -28508
rect -22588 -28572 -22568 -28508
rect -27940 -28588 -22568 -28572
rect -27940 -28652 -22652 -28588
rect -22588 -28652 -22568 -28588
rect -27940 -28668 -22568 -28652
rect -27940 -28732 -22652 -28668
rect -22588 -28732 -22568 -28668
rect -27940 -28748 -22568 -28732
rect -27940 -28812 -22652 -28748
rect -22588 -28812 -22568 -28748
rect -27940 -28828 -22568 -28812
rect -27940 -28892 -22652 -28828
rect -22588 -28892 -22568 -28828
rect -27940 -28908 -22568 -28892
rect -27940 -28972 -22652 -28908
rect -22588 -28972 -22568 -28908
rect -27940 -28988 -22568 -28972
rect -27940 -29052 -22652 -28988
rect -22588 -29052 -22568 -28988
rect -27940 -29068 -22568 -29052
rect -27940 -29132 -22652 -29068
rect -22588 -29132 -22568 -29068
rect -27940 -29148 -22568 -29132
rect -27940 -29212 -22652 -29148
rect -22588 -29212 -22568 -29148
rect -27940 -29228 -22568 -29212
rect -27940 -29292 -22652 -29228
rect -22588 -29292 -22568 -29228
rect -27940 -29308 -22568 -29292
rect -27940 -29372 -22652 -29308
rect -22588 -29372 -22568 -29308
rect -27940 -29388 -22568 -29372
rect -27940 -29452 -22652 -29388
rect -22588 -29452 -22568 -29388
rect -27940 -29468 -22568 -29452
rect -27940 -29532 -22652 -29468
rect -22588 -29532 -22568 -29468
rect -27940 -29548 -22568 -29532
rect -27940 -29612 -22652 -29548
rect -22588 -29612 -22568 -29548
rect -27940 -29628 -22568 -29612
rect -27940 -29692 -22652 -29628
rect -22588 -29692 -22568 -29628
rect -27940 -29708 -22568 -29692
rect -27940 -29772 -22652 -29708
rect -22588 -29772 -22568 -29708
rect -27940 -29788 -22568 -29772
rect -27940 -29852 -22652 -29788
rect -22588 -29852 -22568 -29788
rect -27940 -29868 -22568 -29852
rect -27940 -29932 -22652 -29868
rect -22588 -29932 -22568 -29868
rect -27940 -29948 -22568 -29932
rect -27940 -30012 -22652 -29948
rect -22588 -30012 -22568 -29948
rect -27940 -30028 -22568 -30012
rect -27940 -30092 -22652 -30028
rect -22588 -30092 -22568 -30028
rect -27940 -30108 -22568 -30092
rect -27940 -30172 -22652 -30108
rect -22588 -30172 -22568 -30108
rect -27940 -30188 -22568 -30172
rect -27940 -30252 -22652 -30188
rect -22588 -30252 -22568 -30188
rect -27940 -30268 -22568 -30252
rect -27940 -30332 -22652 -30268
rect -22588 -30332 -22568 -30268
rect -27940 -30348 -22568 -30332
rect -27940 -30412 -22652 -30348
rect -22588 -30412 -22568 -30348
rect -27940 -30428 -22568 -30412
rect -27940 -30492 -22652 -30428
rect -22588 -30492 -22568 -30428
rect -27940 -30508 -22568 -30492
rect -27940 -30572 -22652 -30508
rect -22588 -30572 -22568 -30508
rect -27940 -30588 -22568 -30572
rect -27940 -30652 -22652 -30588
rect -22588 -30652 -22568 -30588
rect -27940 -30668 -22568 -30652
rect -27940 -30732 -22652 -30668
rect -22588 -30732 -22568 -30668
rect -27940 -30748 -22568 -30732
rect -27940 -30812 -22652 -30748
rect -22588 -30812 -22568 -30748
rect -27940 -30828 -22568 -30812
rect -27940 -30892 -22652 -30828
rect -22588 -30892 -22568 -30828
rect -27940 -30908 -22568 -30892
rect -27940 -30972 -22652 -30908
rect -22588 -30972 -22568 -30908
rect -27940 -30988 -22568 -30972
rect -27940 -31052 -22652 -30988
rect -22588 -31052 -22568 -30988
rect -27940 -31068 -22568 -31052
rect -27940 -31132 -22652 -31068
rect -22588 -31132 -22568 -31068
rect -27940 -31148 -22568 -31132
rect -27940 -31212 -22652 -31148
rect -22588 -31212 -22568 -31148
rect -27940 -31228 -22568 -31212
rect -27940 -31292 -22652 -31228
rect -22588 -31292 -22568 -31228
rect -27940 -31308 -22568 -31292
rect -27940 -31372 -22652 -31308
rect -22588 -31372 -22568 -31308
rect -27940 -31388 -22568 -31372
rect -27940 -31452 -22652 -31388
rect -22588 -31452 -22568 -31388
rect -27940 -31468 -22568 -31452
rect -27940 -31532 -22652 -31468
rect -22588 -31532 -22568 -31468
rect -27940 -31548 -22568 -31532
rect -27940 -31612 -22652 -31548
rect -22588 -31612 -22568 -31548
rect -27940 -31628 -22568 -31612
rect -27940 -31692 -22652 -31628
rect -22588 -31692 -22568 -31628
rect -27940 -31708 -22568 -31692
rect -27940 -31772 -22652 -31708
rect -22588 -31772 -22568 -31708
rect -27940 -31800 -22568 -31772
rect -22328 -26748 -16956 -26720
rect -22328 -26812 -17040 -26748
rect -16976 -26812 -16956 -26748
rect -22328 -26828 -16956 -26812
rect -22328 -26892 -17040 -26828
rect -16976 -26892 -16956 -26828
rect -22328 -26908 -16956 -26892
rect -22328 -26972 -17040 -26908
rect -16976 -26972 -16956 -26908
rect -22328 -26988 -16956 -26972
rect -22328 -27052 -17040 -26988
rect -16976 -27052 -16956 -26988
rect -22328 -27068 -16956 -27052
rect -22328 -27132 -17040 -27068
rect -16976 -27132 -16956 -27068
rect -22328 -27148 -16956 -27132
rect -22328 -27212 -17040 -27148
rect -16976 -27212 -16956 -27148
rect -22328 -27228 -16956 -27212
rect -22328 -27292 -17040 -27228
rect -16976 -27292 -16956 -27228
rect -22328 -27308 -16956 -27292
rect -22328 -27372 -17040 -27308
rect -16976 -27372 -16956 -27308
rect -22328 -27388 -16956 -27372
rect -22328 -27452 -17040 -27388
rect -16976 -27452 -16956 -27388
rect -22328 -27468 -16956 -27452
rect -22328 -27532 -17040 -27468
rect -16976 -27532 -16956 -27468
rect -22328 -27548 -16956 -27532
rect -22328 -27612 -17040 -27548
rect -16976 -27612 -16956 -27548
rect -22328 -27628 -16956 -27612
rect -22328 -27692 -17040 -27628
rect -16976 -27692 -16956 -27628
rect -22328 -27708 -16956 -27692
rect -22328 -27772 -17040 -27708
rect -16976 -27772 -16956 -27708
rect -22328 -27788 -16956 -27772
rect -22328 -27852 -17040 -27788
rect -16976 -27852 -16956 -27788
rect -22328 -27868 -16956 -27852
rect -22328 -27932 -17040 -27868
rect -16976 -27932 -16956 -27868
rect -22328 -27948 -16956 -27932
rect -22328 -28012 -17040 -27948
rect -16976 -28012 -16956 -27948
rect -22328 -28028 -16956 -28012
rect -22328 -28092 -17040 -28028
rect -16976 -28092 -16956 -28028
rect -22328 -28108 -16956 -28092
rect -22328 -28172 -17040 -28108
rect -16976 -28172 -16956 -28108
rect -22328 -28188 -16956 -28172
rect -22328 -28252 -17040 -28188
rect -16976 -28252 -16956 -28188
rect -22328 -28268 -16956 -28252
rect -22328 -28332 -17040 -28268
rect -16976 -28332 -16956 -28268
rect -22328 -28348 -16956 -28332
rect -22328 -28412 -17040 -28348
rect -16976 -28412 -16956 -28348
rect -22328 -28428 -16956 -28412
rect -22328 -28492 -17040 -28428
rect -16976 -28492 -16956 -28428
rect -22328 -28508 -16956 -28492
rect -22328 -28572 -17040 -28508
rect -16976 -28572 -16956 -28508
rect -22328 -28588 -16956 -28572
rect -22328 -28652 -17040 -28588
rect -16976 -28652 -16956 -28588
rect -22328 -28668 -16956 -28652
rect -22328 -28732 -17040 -28668
rect -16976 -28732 -16956 -28668
rect -22328 -28748 -16956 -28732
rect -22328 -28812 -17040 -28748
rect -16976 -28812 -16956 -28748
rect -22328 -28828 -16956 -28812
rect -22328 -28892 -17040 -28828
rect -16976 -28892 -16956 -28828
rect -22328 -28908 -16956 -28892
rect -22328 -28972 -17040 -28908
rect -16976 -28972 -16956 -28908
rect -22328 -28988 -16956 -28972
rect -22328 -29052 -17040 -28988
rect -16976 -29052 -16956 -28988
rect -22328 -29068 -16956 -29052
rect -22328 -29132 -17040 -29068
rect -16976 -29132 -16956 -29068
rect -22328 -29148 -16956 -29132
rect -22328 -29212 -17040 -29148
rect -16976 -29212 -16956 -29148
rect -22328 -29228 -16956 -29212
rect -22328 -29292 -17040 -29228
rect -16976 -29292 -16956 -29228
rect -22328 -29308 -16956 -29292
rect -22328 -29372 -17040 -29308
rect -16976 -29372 -16956 -29308
rect -22328 -29388 -16956 -29372
rect -22328 -29452 -17040 -29388
rect -16976 -29452 -16956 -29388
rect -22328 -29468 -16956 -29452
rect -22328 -29532 -17040 -29468
rect -16976 -29532 -16956 -29468
rect -22328 -29548 -16956 -29532
rect -22328 -29612 -17040 -29548
rect -16976 -29612 -16956 -29548
rect -22328 -29628 -16956 -29612
rect -22328 -29692 -17040 -29628
rect -16976 -29692 -16956 -29628
rect -22328 -29708 -16956 -29692
rect -22328 -29772 -17040 -29708
rect -16976 -29772 -16956 -29708
rect -22328 -29788 -16956 -29772
rect -22328 -29852 -17040 -29788
rect -16976 -29852 -16956 -29788
rect -22328 -29868 -16956 -29852
rect -22328 -29932 -17040 -29868
rect -16976 -29932 -16956 -29868
rect -22328 -29948 -16956 -29932
rect -22328 -30012 -17040 -29948
rect -16976 -30012 -16956 -29948
rect -22328 -30028 -16956 -30012
rect -22328 -30092 -17040 -30028
rect -16976 -30092 -16956 -30028
rect -22328 -30108 -16956 -30092
rect -22328 -30172 -17040 -30108
rect -16976 -30172 -16956 -30108
rect -22328 -30188 -16956 -30172
rect -22328 -30252 -17040 -30188
rect -16976 -30252 -16956 -30188
rect -22328 -30268 -16956 -30252
rect -22328 -30332 -17040 -30268
rect -16976 -30332 -16956 -30268
rect -22328 -30348 -16956 -30332
rect -22328 -30412 -17040 -30348
rect -16976 -30412 -16956 -30348
rect -22328 -30428 -16956 -30412
rect -22328 -30492 -17040 -30428
rect -16976 -30492 -16956 -30428
rect -22328 -30508 -16956 -30492
rect -22328 -30572 -17040 -30508
rect -16976 -30572 -16956 -30508
rect -22328 -30588 -16956 -30572
rect -22328 -30652 -17040 -30588
rect -16976 -30652 -16956 -30588
rect -22328 -30668 -16956 -30652
rect -22328 -30732 -17040 -30668
rect -16976 -30732 -16956 -30668
rect -22328 -30748 -16956 -30732
rect -22328 -30812 -17040 -30748
rect -16976 -30812 -16956 -30748
rect -22328 -30828 -16956 -30812
rect -22328 -30892 -17040 -30828
rect -16976 -30892 -16956 -30828
rect -22328 -30908 -16956 -30892
rect -22328 -30972 -17040 -30908
rect -16976 -30972 -16956 -30908
rect -22328 -30988 -16956 -30972
rect -22328 -31052 -17040 -30988
rect -16976 -31052 -16956 -30988
rect -22328 -31068 -16956 -31052
rect -22328 -31132 -17040 -31068
rect -16976 -31132 -16956 -31068
rect -22328 -31148 -16956 -31132
rect -22328 -31212 -17040 -31148
rect -16976 -31212 -16956 -31148
rect -22328 -31228 -16956 -31212
rect -22328 -31292 -17040 -31228
rect -16976 -31292 -16956 -31228
rect -22328 -31308 -16956 -31292
rect -22328 -31372 -17040 -31308
rect -16976 -31372 -16956 -31308
rect -22328 -31388 -16956 -31372
rect -22328 -31452 -17040 -31388
rect -16976 -31452 -16956 -31388
rect -22328 -31468 -16956 -31452
rect -22328 -31532 -17040 -31468
rect -16976 -31532 -16956 -31468
rect -22328 -31548 -16956 -31532
rect -22328 -31612 -17040 -31548
rect -16976 -31612 -16956 -31548
rect -22328 -31628 -16956 -31612
rect -22328 -31692 -17040 -31628
rect -16976 -31692 -16956 -31628
rect -22328 -31708 -16956 -31692
rect -22328 -31772 -17040 -31708
rect -16976 -31772 -16956 -31708
rect -22328 -31800 -16956 -31772
rect -16716 -26748 -11344 -26720
rect -16716 -26812 -11428 -26748
rect -11364 -26812 -11344 -26748
rect -16716 -26828 -11344 -26812
rect -16716 -26892 -11428 -26828
rect -11364 -26892 -11344 -26828
rect -16716 -26908 -11344 -26892
rect -16716 -26972 -11428 -26908
rect -11364 -26972 -11344 -26908
rect -16716 -26988 -11344 -26972
rect -16716 -27052 -11428 -26988
rect -11364 -27052 -11344 -26988
rect -16716 -27068 -11344 -27052
rect -16716 -27132 -11428 -27068
rect -11364 -27132 -11344 -27068
rect -16716 -27148 -11344 -27132
rect -16716 -27212 -11428 -27148
rect -11364 -27212 -11344 -27148
rect -16716 -27228 -11344 -27212
rect -16716 -27292 -11428 -27228
rect -11364 -27292 -11344 -27228
rect -16716 -27308 -11344 -27292
rect -16716 -27372 -11428 -27308
rect -11364 -27372 -11344 -27308
rect -16716 -27388 -11344 -27372
rect -16716 -27452 -11428 -27388
rect -11364 -27452 -11344 -27388
rect -16716 -27468 -11344 -27452
rect -16716 -27532 -11428 -27468
rect -11364 -27532 -11344 -27468
rect -16716 -27548 -11344 -27532
rect -16716 -27612 -11428 -27548
rect -11364 -27612 -11344 -27548
rect -16716 -27628 -11344 -27612
rect -16716 -27692 -11428 -27628
rect -11364 -27692 -11344 -27628
rect -16716 -27708 -11344 -27692
rect -16716 -27772 -11428 -27708
rect -11364 -27772 -11344 -27708
rect -16716 -27788 -11344 -27772
rect -16716 -27852 -11428 -27788
rect -11364 -27852 -11344 -27788
rect -16716 -27868 -11344 -27852
rect -16716 -27932 -11428 -27868
rect -11364 -27932 -11344 -27868
rect -16716 -27948 -11344 -27932
rect -16716 -28012 -11428 -27948
rect -11364 -28012 -11344 -27948
rect -16716 -28028 -11344 -28012
rect -16716 -28092 -11428 -28028
rect -11364 -28092 -11344 -28028
rect -16716 -28108 -11344 -28092
rect -16716 -28172 -11428 -28108
rect -11364 -28172 -11344 -28108
rect -16716 -28188 -11344 -28172
rect -16716 -28252 -11428 -28188
rect -11364 -28252 -11344 -28188
rect -16716 -28268 -11344 -28252
rect -16716 -28332 -11428 -28268
rect -11364 -28332 -11344 -28268
rect -16716 -28348 -11344 -28332
rect -16716 -28412 -11428 -28348
rect -11364 -28412 -11344 -28348
rect -16716 -28428 -11344 -28412
rect -16716 -28492 -11428 -28428
rect -11364 -28492 -11344 -28428
rect -16716 -28508 -11344 -28492
rect -16716 -28572 -11428 -28508
rect -11364 -28572 -11344 -28508
rect -16716 -28588 -11344 -28572
rect -16716 -28652 -11428 -28588
rect -11364 -28652 -11344 -28588
rect -16716 -28668 -11344 -28652
rect -16716 -28732 -11428 -28668
rect -11364 -28732 -11344 -28668
rect -16716 -28748 -11344 -28732
rect -16716 -28812 -11428 -28748
rect -11364 -28812 -11344 -28748
rect -16716 -28828 -11344 -28812
rect -16716 -28892 -11428 -28828
rect -11364 -28892 -11344 -28828
rect -16716 -28908 -11344 -28892
rect -16716 -28972 -11428 -28908
rect -11364 -28972 -11344 -28908
rect -16716 -28988 -11344 -28972
rect -16716 -29052 -11428 -28988
rect -11364 -29052 -11344 -28988
rect -16716 -29068 -11344 -29052
rect -16716 -29132 -11428 -29068
rect -11364 -29132 -11344 -29068
rect -16716 -29148 -11344 -29132
rect -16716 -29212 -11428 -29148
rect -11364 -29212 -11344 -29148
rect -16716 -29228 -11344 -29212
rect -16716 -29292 -11428 -29228
rect -11364 -29292 -11344 -29228
rect -16716 -29308 -11344 -29292
rect -16716 -29372 -11428 -29308
rect -11364 -29372 -11344 -29308
rect -16716 -29388 -11344 -29372
rect -16716 -29452 -11428 -29388
rect -11364 -29452 -11344 -29388
rect -16716 -29468 -11344 -29452
rect -16716 -29532 -11428 -29468
rect -11364 -29532 -11344 -29468
rect -16716 -29548 -11344 -29532
rect -16716 -29612 -11428 -29548
rect -11364 -29612 -11344 -29548
rect -16716 -29628 -11344 -29612
rect -16716 -29692 -11428 -29628
rect -11364 -29692 -11344 -29628
rect -16716 -29708 -11344 -29692
rect -16716 -29772 -11428 -29708
rect -11364 -29772 -11344 -29708
rect -16716 -29788 -11344 -29772
rect -16716 -29852 -11428 -29788
rect -11364 -29852 -11344 -29788
rect -16716 -29868 -11344 -29852
rect -16716 -29932 -11428 -29868
rect -11364 -29932 -11344 -29868
rect -16716 -29948 -11344 -29932
rect -16716 -30012 -11428 -29948
rect -11364 -30012 -11344 -29948
rect -16716 -30028 -11344 -30012
rect -16716 -30092 -11428 -30028
rect -11364 -30092 -11344 -30028
rect -16716 -30108 -11344 -30092
rect -16716 -30172 -11428 -30108
rect -11364 -30172 -11344 -30108
rect -16716 -30188 -11344 -30172
rect -16716 -30252 -11428 -30188
rect -11364 -30252 -11344 -30188
rect -16716 -30268 -11344 -30252
rect -16716 -30332 -11428 -30268
rect -11364 -30332 -11344 -30268
rect -16716 -30348 -11344 -30332
rect -16716 -30412 -11428 -30348
rect -11364 -30412 -11344 -30348
rect -16716 -30428 -11344 -30412
rect -16716 -30492 -11428 -30428
rect -11364 -30492 -11344 -30428
rect -16716 -30508 -11344 -30492
rect -16716 -30572 -11428 -30508
rect -11364 -30572 -11344 -30508
rect -16716 -30588 -11344 -30572
rect -16716 -30652 -11428 -30588
rect -11364 -30652 -11344 -30588
rect -16716 -30668 -11344 -30652
rect -16716 -30732 -11428 -30668
rect -11364 -30732 -11344 -30668
rect -16716 -30748 -11344 -30732
rect -16716 -30812 -11428 -30748
rect -11364 -30812 -11344 -30748
rect -16716 -30828 -11344 -30812
rect -16716 -30892 -11428 -30828
rect -11364 -30892 -11344 -30828
rect -16716 -30908 -11344 -30892
rect -16716 -30972 -11428 -30908
rect -11364 -30972 -11344 -30908
rect -16716 -30988 -11344 -30972
rect -16716 -31052 -11428 -30988
rect -11364 -31052 -11344 -30988
rect -16716 -31068 -11344 -31052
rect -16716 -31132 -11428 -31068
rect -11364 -31132 -11344 -31068
rect -16716 -31148 -11344 -31132
rect -16716 -31212 -11428 -31148
rect -11364 -31212 -11344 -31148
rect -16716 -31228 -11344 -31212
rect -16716 -31292 -11428 -31228
rect -11364 -31292 -11344 -31228
rect -16716 -31308 -11344 -31292
rect -16716 -31372 -11428 -31308
rect -11364 -31372 -11344 -31308
rect -16716 -31388 -11344 -31372
rect -16716 -31452 -11428 -31388
rect -11364 -31452 -11344 -31388
rect -16716 -31468 -11344 -31452
rect -16716 -31532 -11428 -31468
rect -11364 -31532 -11344 -31468
rect -16716 -31548 -11344 -31532
rect -16716 -31612 -11428 -31548
rect -11364 -31612 -11344 -31548
rect -16716 -31628 -11344 -31612
rect -16716 -31692 -11428 -31628
rect -11364 -31692 -11344 -31628
rect -16716 -31708 -11344 -31692
rect -16716 -31772 -11428 -31708
rect -11364 -31772 -11344 -31708
rect -16716 -31800 -11344 -31772
rect -11104 -26748 -5732 -26720
rect -11104 -26812 -5816 -26748
rect -5752 -26812 -5732 -26748
rect -11104 -26828 -5732 -26812
rect -11104 -26892 -5816 -26828
rect -5752 -26892 -5732 -26828
rect -11104 -26908 -5732 -26892
rect -11104 -26972 -5816 -26908
rect -5752 -26972 -5732 -26908
rect -11104 -26988 -5732 -26972
rect -11104 -27052 -5816 -26988
rect -5752 -27052 -5732 -26988
rect -11104 -27068 -5732 -27052
rect -11104 -27132 -5816 -27068
rect -5752 -27132 -5732 -27068
rect -11104 -27148 -5732 -27132
rect -11104 -27212 -5816 -27148
rect -5752 -27212 -5732 -27148
rect -11104 -27228 -5732 -27212
rect -11104 -27292 -5816 -27228
rect -5752 -27292 -5732 -27228
rect -11104 -27308 -5732 -27292
rect -11104 -27372 -5816 -27308
rect -5752 -27372 -5732 -27308
rect -11104 -27388 -5732 -27372
rect -11104 -27452 -5816 -27388
rect -5752 -27452 -5732 -27388
rect -11104 -27468 -5732 -27452
rect -11104 -27532 -5816 -27468
rect -5752 -27532 -5732 -27468
rect -11104 -27548 -5732 -27532
rect -11104 -27612 -5816 -27548
rect -5752 -27612 -5732 -27548
rect -11104 -27628 -5732 -27612
rect -11104 -27692 -5816 -27628
rect -5752 -27692 -5732 -27628
rect -11104 -27708 -5732 -27692
rect -11104 -27772 -5816 -27708
rect -5752 -27772 -5732 -27708
rect -11104 -27788 -5732 -27772
rect -11104 -27852 -5816 -27788
rect -5752 -27852 -5732 -27788
rect -11104 -27868 -5732 -27852
rect -11104 -27932 -5816 -27868
rect -5752 -27932 -5732 -27868
rect -11104 -27948 -5732 -27932
rect -11104 -28012 -5816 -27948
rect -5752 -28012 -5732 -27948
rect -11104 -28028 -5732 -28012
rect -11104 -28092 -5816 -28028
rect -5752 -28092 -5732 -28028
rect -11104 -28108 -5732 -28092
rect -11104 -28172 -5816 -28108
rect -5752 -28172 -5732 -28108
rect -11104 -28188 -5732 -28172
rect -11104 -28252 -5816 -28188
rect -5752 -28252 -5732 -28188
rect -11104 -28268 -5732 -28252
rect -11104 -28332 -5816 -28268
rect -5752 -28332 -5732 -28268
rect -11104 -28348 -5732 -28332
rect -11104 -28412 -5816 -28348
rect -5752 -28412 -5732 -28348
rect -11104 -28428 -5732 -28412
rect -11104 -28492 -5816 -28428
rect -5752 -28492 -5732 -28428
rect -11104 -28508 -5732 -28492
rect -11104 -28572 -5816 -28508
rect -5752 -28572 -5732 -28508
rect -11104 -28588 -5732 -28572
rect -11104 -28652 -5816 -28588
rect -5752 -28652 -5732 -28588
rect -11104 -28668 -5732 -28652
rect -11104 -28732 -5816 -28668
rect -5752 -28732 -5732 -28668
rect -11104 -28748 -5732 -28732
rect -11104 -28812 -5816 -28748
rect -5752 -28812 -5732 -28748
rect -11104 -28828 -5732 -28812
rect -11104 -28892 -5816 -28828
rect -5752 -28892 -5732 -28828
rect -11104 -28908 -5732 -28892
rect -11104 -28972 -5816 -28908
rect -5752 -28972 -5732 -28908
rect -11104 -28988 -5732 -28972
rect -11104 -29052 -5816 -28988
rect -5752 -29052 -5732 -28988
rect -11104 -29068 -5732 -29052
rect -11104 -29132 -5816 -29068
rect -5752 -29132 -5732 -29068
rect -11104 -29148 -5732 -29132
rect -11104 -29212 -5816 -29148
rect -5752 -29212 -5732 -29148
rect -11104 -29228 -5732 -29212
rect -11104 -29292 -5816 -29228
rect -5752 -29292 -5732 -29228
rect -11104 -29308 -5732 -29292
rect -11104 -29372 -5816 -29308
rect -5752 -29372 -5732 -29308
rect -11104 -29388 -5732 -29372
rect -11104 -29452 -5816 -29388
rect -5752 -29452 -5732 -29388
rect -11104 -29468 -5732 -29452
rect -11104 -29532 -5816 -29468
rect -5752 -29532 -5732 -29468
rect -11104 -29548 -5732 -29532
rect -11104 -29612 -5816 -29548
rect -5752 -29612 -5732 -29548
rect -11104 -29628 -5732 -29612
rect -11104 -29692 -5816 -29628
rect -5752 -29692 -5732 -29628
rect -11104 -29708 -5732 -29692
rect -11104 -29772 -5816 -29708
rect -5752 -29772 -5732 -29708
rect -11104 -29788 -5732 -29772
rect -11104 -29852 -5816 -29788
rect -5752 -29852 -5732 -29788
rect -11104 -29868 -5732 -29852
rect -11104 -29932 -5816 -29868
rect -5752 -29932 -5732 -29868
rect -11104 -29948 -5732 -29932
rect -11104 -30012 -5816 -29948
rect -5752 -30012 -5732 -29948
rect -11104 -30028 -5732 -30012
rect -11104 -30092 -5816 -30028
rect -5752 -30092 -5732 -30028
rect -11104 -30108 -5732 -30092
rect -11104 -30172 -5816 -30108
rect -5752 -30172 -5732 -30108
rect -11104 -30188 -5732 -30172
rect -11104 -30252 -5816 -30188
rect -5752 -30252 -5732 -30188
rect -11104 -30268 -5732 -30252
rect -11104 -30332 -5816 -30268
rect -5752 -30332 -5732 -30268
rect -11104 -30348 -5732 -30332
rect -11104 -30412 -5816 -30348
rect -5752 -30412 -5732 -30348
rect -11104 -30428 -5732 -30412
rect -11104 -30492 -5816 -30428
rect -5752 -30492 -5732 -30428
rect -11104 -30508 -5732 -30492
rect -11104 -30572 -5816 -30508
rect -5752 -30572 -5732 -30508
rect -11104 -30588 -5732 -30572
rect -11104 -30652 -5816 -30588
rect -5752 -30652 -5732 -30588
rect -11104 -30668 -5732 -30652
rect -11104 -30732 -5816 -30668
rect -5752 -30732 -5732 -30668
rect -11104 -30748 -5732 -30732
rect -11104 -30812 -5816 -30748
rect -5752 -30812 -5732 -30748
rect -11104 -30828 -5732 -30812
rect -11104 -30892 -5816 -30828
rect -5752 -30892 -5732 -30828
rect -11104 -30908 -5732 -30892
rect -11104 -30972 -5816 -30908
rect -5752 -30972 -5732 -30908
rect -11104 -30988 -5732 -30972
rect -11104 -31052 -5816 -30988
rect -5752 -31052 -5732 -30988
rect -11104 -31068 -5732 -31052
rect -11104 -31132 -5816 -31068
rect -5752 -31132 -5732 -31068
rect -11104 -31148 -5732 -31132
rect -11104 -31212 -5816 -31148
rect -5752 -31212 -5732 -31148
rect -11104 -31228 -5732 -31212
rect -11104 -31292 -5816 -31228
rect -5752 -31292 -5732 -31228
rect -11104 -31308 -5732 -31292
rect -11104 -31372 -5816 -31308
rect -5752 -31372 -5732 -31308
rect -11104 -31388 -5732 -31372
rect -11104 -31452 -5816 -31388
rect -5752 -31452 -5732 -31388
rect -11104 -31468 -5732 -31452
rect -11104 -31532 -5816 -31468
rect -5752 -31532 -5732 -31468
rect -11104 -31548 -5732 -31532
rect -11104 -31612 -5816 -31548
rect -5752 -31612 -5732 -31548
rect -11104 -31628 -5732 -31612
rect -11104 -31692 -5816 -31628
rect -5752 -31692 -5732 -31628
rect -11104 -31708 -5732 -31692
rect -11104 -31772 -5816 -31708
rect -5752 -31772 -5732 -31708
rect -11104 -31800 -5732 -31772
rect -5492 -26748 -120 -26720
rect -5492 -26812 -204 -26748
rect -140 -26812 -120 -26748
rect -5492 -26828 -120 -26812
rect -5492 -26892 -204 -26828
rect -140 -26892 -120 -26828
rect -5492 -26908 -120 -26892
rect -5492 -26972 -204 -26908
rect -140 -26972 -120 -26908
rect -5492 -26988 -120 -26972
rect -5492 -27052 -204 -26988
rect -140 -27052 -120 -26988
rect -5492 -27068 -120 -27052
rect -5492 -27132 -204 -27068
rect -140 -27132 -120 -27068
rect -5492 -27148 -120 -27132
rect -5492 -27212 -204 -27148
rect -140 -27212 -120 -27148
rect -5492 -27228 -120 -27212
rect -5492 -27292 -204 -27228
rect -140 -27292 -120 -27228
rect -5492 -27308 -120 -27292
rect -5492 -27372 -204 -27308
rect -140 -27372 -120 -27308
rect -5492 -27388 -120 -27372
rect -5492 -27452 -204 -27388
rect -140 -27452 -120 -27388
rect -5492 -27468 -120 -27452
rect -5492 -27532 -204 -27468
rect -140 -27532 -120 -27468
rect -5492 -27548 -120 -27532
rect -5492 -27612 -204 -27548
rect -140 -27612 -120 -27548
rect -5492 -27628 -120 -27612
rect -5492 -27692 -204 -27628
rect -140 -27692 -120 -27628
rect -5492 -27708 -120 -27692
rect -5492 -27772 -204 -27708
rect -140 -27772 -120 -27708
rect -5492 -27788 -120 -27772
rect -5492 -27852 -204 -27788
rect -140 -27852 -120 -27788
rect -5492 -27868 -120 -27852
rect -5492 -27932 -204 -27868
rect -140 -27932 -120 -27868
rect -5492 -27948 -120 -27932
rect -5492 -28012 -204 -27948
rect -140 -28012 -120 -27948
rect -5492 -28028 -120 -28012
rect -5492 -28092 -204 -28028
rect -140 -28092 -120 -28028
rect -5492 -28108 -120 -28092
rect -5492 -28172 -204 -28108
rect -140 -28172 -120 -28108
rect -5492 -28188 -120 -28172
rect -5492 -28252 -204 -28188
rect -140 -28252 -120 -28188
rect -5492 -28268 -120 -28252
rect -5492 -28332 -204 -28268
rect -140 -28332 -120 -28268
rect -5492 -28348 -120 -28332
rect -5492 -28412 -204 -28348
rect -140 -28412 -120 -28348
rect -5492 -28428 -120 -28412
rect -5492 -28492 -204 -28428
rect -140 -28492 -120 -28428
rect -5492 -28508 -120 -28492
rect -5492 -28572 -204 -28508
rect -140 -28572 -120 -28508
rect -5492 -28588 -120 -28572
rect -5492 -28652 -204 -28588
rect -140 -28652 -120 -28588
rect -5492 -28668 -120 -28652
rect -5492 -28732 -204 -28668
rect -140 -28732 -120 -28668
rect -5492 -28748 -120 -28732
rect -5492 -28812 -204 -28748
rect -140 -28812 -120 -28748
rect -5492 -28828 -120 -28812
rect -5492 -28892 -204 -28828
rect -140 -28892 -120 -28828
rect -5492 -28908 -120 -28892
rect -5492 -28972 -204 -28908
rect -140 -28972 -120 -28908
rect -5492 -28988 -120 -28972
rect -5492 -29052 -204 -28988
rect -140 -29052 -120 -28988
rect -5492 -29068 -120 -29052
rect -5492 -29132 -204 -29068
rect -140 -29132 -120 -29068
rect -5492 -29148 -120 -29132
rect -5492 -29212 -204 -29148
rect -140 -29212 -120 -29148
rect -5492 -29228 -120 -29212
rect -5492 -29292 -204 -29228
rect -140 -29292 -120 -29228
rect -5492 -29308 -120 -29292
rect -5492 -29372 -204 -29308
rect -140 -29372 -120 -29308
rect -5492 -29388 -120 -29372
rect -5492 -29452 -204 -29388
rect -140 -29452 -120 -29388
rect -5492 -29468 -120 -29452
rect -5492 -29532 -204 -29468
rect -140 -29532 -120 -29468
rect -5492 -29548 -120 -29532
rect -5492 -29612 -204 -29548
rect -140 -29612 -120 -29548
rect -5492 -29628 -120 -29612
rect -5492 -29692 -204 -29628
rect -140 -29692 -120 -29628
rect -5492 -29708 -120 -29692
rect -5492 -29772 -204 -29708
rect -140 -29772 -120 -29708
rect -5492 -29788 -120 -29772
rect -5492 -29852 -204 -29788
rect -140 -29852 -120 -29788
rect -5492 -29868 -120 -29852
rect -5492 -29932 -204 -29868
rect -140 -29932 -120 -29868
rect -5492 -29948 -120 -29932
rect -5492 -30012 -204 -29948
rect -140 -30012 -120 -29948
rect -5492 -30028 -120 -30012
rect -5492 -30092 -204 -30028
rect -140 -30092 -120 -30028
rect -5492 -30108 -120 -30092
rect -5492 -30172 -204 -30108
rect -140 -30172 -120 -30108
rect -5492 -30188 -120 -30172
rect -5492 -30252 -204 -30188
rect -140 -30252 -120 -30188
rect -5492 -30268 -120 -30252
rect -5492 -30332 -204 -30268
rect -140 -30332 -120 -30268
rect -5492 -30348 -120 -30332
rect -5492 -30412 -204 -30348
rect -140 -30412 -120 -30348
rect -5492 -30428 -120 -30412
rect -5492 -30492 -204 -30428
rect -140 -30492 -120 -30428
rect -5492 -30508 -120 -30492
rect -5492 -30572 -204 -30508
rect -140 -30572 -120 -30508
rect -5492 -30588 -120 -30572
rect -5492 -30652 -204 -30588
rect -140 -30652 -120 -30588
rect -5492 -30668 -120 -30652
rect -5492 -30732 -204 -30668
rect -140 -30732 -120 -30668
rect -5492 -30748 -120 -30732
rect -5492 -30812 -204 -30748
rect -140 -30812 -120 -30748
rect -5492 -30828 -120 -30812
rect -5492 -30892 -204 -30828
rect -140 -30892 -120 -30828
rect -5492 -30908 -120 -30892
rect -5492 -30972 -204 -30908
rect -140 -30972 -120 -30908
rect -5492 -30988 -120 -30972
rect -5492 -31052 -204 -30988
rect -140 -31052 -120 -30988
rect -5492 -31068 -120 -31052
rect -5492 -31132 -204 -31068
rect -140 -31132 -120 -31068
rect -5492 -31148 -120 -31132
rect -5492 -31212 -204 -31148
rect -140 -31212 -120 -31148
rect -5492 -31228 -120 -31212
rect -5492 -31292 -204 -31228
rect -140 -31292 -120 -31228
rect -5492 -31308 -120 -31292
rect -5492 -31372 -204 -31308
rect -140 -31372 -120 -31308
rect -5492 -31388 -120 -31372
rect -5492 -31452 -204 -31388
rect -140 -31452 -120 -31388
rect -5492 -31468 -120 -31452
rect -5492 -31532 -204 -31468
rect -140 -31532 -120 -31468
rect -5492 -31548 -120 -31532
rect -5492 -31612 -204 -31548
rect -140 -31612 -120 -31548
rect -5492 -31628 -120 -31612
rect -5492 -31692 -204 -31628
rect -140 -31692 -120 -31628
rect -5492 -31708 -120 -31692
rect -5492 -31772 -204 -31708
rect -140 -31772 -120 -31708
rect -5492 -31800 -120 -31772
rect 120 -26748 5492 -26720
rect 120 -26812 5408 -26748
rect 5472 -26812 5492 -26748
rect 120 -26828 5492 -26812
rect 120 -26892 5408 -26828
rect 5472 -26892 5492 -26828
rect 120 -26908 5492 -26892
rect 120 -26972 5408 -26908
rect 5472 -26972 5492 -26908
rect 120 -26988 5492 -26972
rect 120 -27052 5408 -26988
rect 5472 -27052 5492 -26988
rect 120 -27068 5492 -27052
rect 120 -27132 5408 -27068
rect 5472 -27132 5492 -27068
rect 120 -27148 5492 -27132
rect 120 -27212 5408 -27148
rect 5472 -27212 5492 -27148
rect 120 -27228 5492 -27212
rect 120 -27292 5408 -27228
rect 5472 -27292 5492 -27228
rect 120 -27308 5492 -27292
rect 120 -27372 5408 -27308
rect 5472 -27372 5492 -27308
rect 120 -27388 5492 -27372
rect 120 -27452 5408 -27388
rect 5472 -27452 5492 -27388
rect 120 -27468 5492 -27452
rect 120 -27532 5408 -27468
rect 5472 -27532 5492 -27468
rect 120 -27548 5492 -27532
rect 120 -27612 5408 -27548
rect 5472 -27612 5492 -27548
rect 120 -27628 5492 -27612
rect 120 -27692 5408 -27628
rect 5472 -27692 5492 -27628
rect 120 -27708 5492 -27692
rect 120 -27772 5408 -27708
rect 5472 -27772 5492 -27708
rect 120 -27788 5492 -27772
rect 120 -27852 5408 -27788
rect 5472 -27852 5492 -27788
rect 120 -27868 5492 -27852
rect 120 -27932 5408 -27868
rect 5472 -27932 5492 -27868
rect 120 -27948 5492 -27932
rect 120 -28012 5408 -27948
rect 5472 -28012 5492 -27948
rect 120 -28028 5492 -28012
rect 120 -28092 5408 -28028
rect 5472 -28092 5492 -28028
rect 120 -28108 5492 -28092
rect 120 -28172 5408 -28108
rect 5472 -28172 5492 -28108
rect 120 -28188 5492 -28172
rect 120 -28252 5408 -28188
rect 5472 -28252 5492 -28188
rect 120 -28268 5492 -28252
rect 120 -28332 5408 -28268
rect 5472 -28332 5492 -28268
rect 120 -28348 5492 -28332
rect 120 -28412 5408 -28348
rect 5472 -28412 5492 -28348
rect 120 -28428 5492 -28412
rect 120 -28492 5408 -28428
rect 5472 -28492 5492 -28428
rect 120 -28508 5492 -28492
rect 120 -28572 5408 -28508
rect 5472 -28572 5492 -28508
rect 120 -28588 5492 -28572
rect 120 -28652 5408 -28588
rect 5472 -28652 5492 -28588
rect 120 -28668 5492 -28652
rect 120 -28732 5408 -28668
rect 5472 -28732 5492 -28668
rect 120 -28748 5492 -28732
rect 120 -28812 5408 -28748
rect 5472 -28812 5492 -28748
rect 120 -28828 5492 -28812
rect 120 -28892 5408 -28828
rect 5472 -28892 5492 -28828
rect 120 -28908 5492 -28892
rect 120 -28972 5408 -28908
rect 5472 -28972 5492 -28908
rect 120 -28988 5492 -28972
rect 120 -29052 5408 -28988
rect 5472 -29052 5492 -28988
rect 120 -29068 5492 -29052
rect 120 -29132 5408 -29068
rect 5472 -29132 5492 -29068
rect 120 -29148 5492 -29132
rect 120 -29212 5408 -29148
rect 5472 -29212 5492 -29148
rect 120 -29228 5492 -29212
rect 120 -29292 5408 -29228
rect 5472 -29292 5492 -29228
rect 120 -29308 5492 -29292
rect 120 -29372 5408 -29308
rect 5472 -29372 5492 -29308
rect 120 -29388 5492 -29372
rect 120 -29452 5408 -29388
rect 5472 -29452 5492 -29388
rect 120 -29468 5492 -29452
rect 120 -29532 5408 -29468
rect 5472 -29532 5492 -29468
rect 120 -29548 5492 -29532
rect 120 -29612 5408 -29548
rect 5472 -29612 5492 -29548
rect 120 -29628 5492 -29612
rect 120 -29692 5408 -29628
rect 5472 -29692 5492 -29628
rect 120 -29708 5492 -29692
rect 120 -29772 5408 -29708
rect 5472 -29772 5492 -29708
rect 120 -29788 5492 -29772
rect 120 -29852 5408 -29788
rect 5472 -29852 5492 -29788
rect 120 -29868 5492 -29852
rect 120 -29932 5408 -29868
rect 5472 -29932 5492 -29868
rect 120 -29948 5492 -29932
rect 120 -30012 5408 -29948
rect 5472 -30012 5492 -29948
rect 120 -30028 5492 -30012
rect 120 -30092 5408 -30028
rect 5472 -30092 5492 -30028
rect 120 -30108 5492 -30092
rect 120 -30172 5408 -30108
rect 5472 -30172 5492 -30108
rect 120 -30188 5492 -30172
rect 120 -30252 5408 -30188
rect 5472 -30252 5492 -30188
rect 120 -30268 5492 -30252
rect 120 -30332 5408 -30268
rect 5472 -30332 5492 -30268
rect 120 -30348 5492 -30332
rect 120 -30412 5408 -30348
rect 5472 -30412 5492 -30348
rect 120 -30428 5492 -30412
rect 120 -30492 5408 -30428
rect 5472 -30492 5492 -30428
rect 120 -30508 5492 -30492
rect 120 -30572 5408 -30508
rect 5472 -30572 5492 -30508
rect 120 -30588 5492 -30572
rect 120 -30652 5408 -30588
rect 5472 -30652 5492 -30588
rect 120 -30668 5492 -30652
rect 120 -30732 5408 -30668
rect 5472 -30732 5492 -30668
rect 120 -30748 5492 -30732
rect 120 -30812 5408 -30748
rect 5472 -30812 5492 -30748
rect 120 -30828 5492 -30812
rect 120 -30892 5408 -30828
rect 5472 -30892 5492 -30828
rect 120 -30908 5492 -30892
rect 120 -30972 5408 -30908
rect 5472 -30972 5492 -30908
rect 120 -30988 5492 -30972
rect 120 -31052 5408 -30988
rect 5472 -31052 5492 -30988
rect 120 -31068 5492 -31052
rect 120 -31132 5408 -31068
rect 5472 -31132 5492 -31068
rect 120 -31148 5492 -31132
rect 120 -31212 5408 -31148
rect 5472 -31212 5492 -31148
rect 120 -31228 5492 -31212
rect 120 -31292 5408 -31228
rect 5472 -31292 5492 -31228
rect 120 -31308 5492 -31292
rect 120 -31372 5408 -31308
rect 5472 -31372 5492 -31308
rect 120 -31388 5492 -31372
rect 120 -31452 5408 -31388
rect 5472 -31452 5492 -31388
rect 120 -31468 5492 -31452
rect 120 -31532 5408 -31468
rect 5472 -31532 5492 -31468
rect 120 -31548 5492 -31532
rect 120 -31612 5408 -31548
rect 5472 -31612 5492 -31548
rect 120 -31628 5492 -31612
rect 120 -31692 5408 -31628
rect 5472 -31692 5492 -31628
rect 120 -31708 5492 -31692
rect 120 -31772 5408 -31708
rect 5472 -31772 5492 -31708
rect 120 -31800 5492 -31772
rect 5732 -26748 11104 -26720
rect 5732 -26812 11020 -26748
rect 11084 -26812 11104 -26748
rect 5732 -26828 11104 -26812
rect 5732 -26892 11020 -26828
rect 11084 -26892 11104 -26828
rect 5732 -26908 11104 -26892
rect 5732 -26972 11020 -26908
rect 11084 -26972 11104 -26908
rect 5732 -26988 11104 -26972
rect 5732 -27052 11020 -26988
rect 11084 -27052 11104 -26988
rect 5732 -27068 11104 -27052
rect 5732 -27132 11020 -27068
rect 11084 -27132 11104 -27068
rect 5732 -27148 11104 -27132
rect 5732 -27212 11020 -27148
rect 11084 -27212 11104 -27148
rect 5732 -27228 11104 -27212
rect 5732 -27292 11020 -27228
rect 11084 -27292 11104 -27228
rect 5732 -27308 11104 -27292
rect 5732 -27372 11020 -27308
rect 11084 -27372 11104 -27308
rect 5732 -27388 11104 -27372
rect 5732 -27452 11020 -27388
rect 11084 -27452 11104 -27388
rect 5732 -27468 11104 -27452
rect 5732 -27532 11020 -27468
rect 11084 -27532 11104 -27468
rect 5732 -27548 11104 -27532
rect 5732 -27612 11020 -27548
rect 11084 -27612 11104 -27548
rect 5732 -27628 11104 -27612
rect 5732 -27692 11020 -27628
rect 11084 -27692 11104 -27628
rect 5732 -27708 11104 -27692
rect 5732 -27772 11020 -27708
rect 11084 -27772 11104 -27708
rect 5732 -27788 11104 -27772
rect 5732 -27852 11020 -27788
rect 11084 -27852 11104 -27788
rect 5732 -27868 11104 -27852
rect 5732 -27932 11020 -27868
rect 11084 -27932 11104 -27868
rect 5732 -27948 11104 -27932
rect 5732 -28012 11020 -27948
rect 11084 -28012 11104 -27948
rect 5732 -28028 11104 -28012
rect 5732 -28092 11020 -28028
rect 11084 -28092 11104 -28028
rect 5732 -28108 11104 -28092
rect 5732 -28172 11020 -28108
rect 11084 -28172 11104 -28108
rect 5732 -28188 11104 -28172
rect 5732 -28252 11020 -28188
rect 11084 -28252 11104 -28188
rect 5732 -28268 11104 -28252
rect 5732 -28332 11020 -28268
rect 11084 -28332 11104 -28268
rect 5732 -28348 11104 -28332
rect 5732 -28412 11020 -28348
rect 11084 -28412 11104 -28348
rect 5732 -28428 11104 -28412
rect 5732 -28492 11020 -28428
rect 11084 -28492 11104 -28428
rect 5732 -28508 11104 -28492
rect 5732 -28572 11020 -28508
rect 11084 -28572 11104 -28508
rect 5732 -28588 11104 -28572
rect 5732 -28652 11020 -28588
rect 11084 -28652 11104 -28588
rect 5732 -28668 11104 -28652
rect 5732 -28732 11020 -28668
rect 11084 -28732 11104 -28668
rect 5732 -28748 11104 -28732
rect 5732 -28812 11020 -28748
rect 11084 -28812 11104 -28748
rect 5732 -28828 11104 -28812
rect 5732 -28892 11020 -28828
rect 11084 -28892 11104 -28828
rect 5732 -28908 11104 -28892
rect 5732 -28972 11020 -28908
rect 11084 -28972 11104 -28908
rect 5732 -28988 11104 -28972
rect 5732 -29052 11020 -28988
rect 11084 -29052 11104 -28988
rect 5732 -29068 11104 -29052
rect 5732 -29132 11020 -29068
rect 11084 -29132 11104 -29068
rect 5732 -29148 11104 -29132
rect 5732 -29212 11020 -29148
rect 11084 -29212 11104 -29148
rect 5732 -29228 11104 -29212
rect 5732 -29292 11020 -29228
rect 11084 -29292 11104 -29228
rect 5732 -29308 11104 -29292
rect 5732 -29372 11020 -29308
rect 11084 -29372 11104 -29308
rect 5732 -29388 11104 -29372
rect 5732 -29452 11020 -29388
rect 11084 -29452 11104 -29388
rect 5732 -29468 11104 -29452
rect 5732 -29532 11020 -29468
rect 11084 -29532 11104 -29468
rect 5732 -29548 11104 -29532
rect 5732 -29612 11020 -29548
rect 11084 -29612 11104 -29548
rect 5732 -29628 11104 -29612
rect 5732 -29692 11020 -29628
rect 11084 -29692 11104 -29628
rect 5732 -29708 11104 -29692
rect 5732 -29772 11020 -29708
rect 11084 -29772 11104 -29708
rect 5732 -29788 11104 -29772
rect 5732 -29852 11020 -29788
rect 11084 -29852 11104 -29788
rect 5732 -29868 11104 -29852
rect 5732 -29932 11020 -29868
rect 11084 -29932 11104 -29868
rect 5732 -29948 11104 -29932
rect 5732 -30012 11020 -29948
rect 11084 -30012 11104 -29948
rect 5732 -30028 11104 -30012
rect 5732 -30092 11020 -30028
rect 11084 -30092 11104 -30028
rect 5732 -30108 11104 -30092
rect 5732 -30172 11020 -30108
rect 11084 -30172 11104 -30108
rect 5732 -30188 11104 -30172
rect 5732 -30252 11020 -30188
rect 11084 -30252 11104 -30188
rect 5732 -30268 11104 -30252
rect 5732 -30332 11020 -30268
rect 11084 -30332 11104 -30268
rect 5732 -30348 11104 -30332
rect 5732 -30412 11020 -30348
rect 11084 -30412 11104 -30348
rect 5732 -30428 11104 -30412
rect 5732 -30492 11020 -30428
rect 11084 -30492 11104 -30428
rect 5732 -30508 11104 -30492
rect 5732 -30572 11020 -30508
rect 11084 -30572 11104 -30508
rect 5732 -30588 11104 -30572
rect 5732 -30652 11020 -30588
rect 11084 -30652 11104 -30588
rect 5732 -30668 11104 -30652
rect 5732 -30732 11020 -30668
rect 11084 -30732 11104 -30668
rect 5732 -30748 11104 -30732
rect 5732 -30812 11020 -30748
rect 11084 -30812 11104 -30748
rect 5732 -30828 11104 -30812
rect 5732 -30892 11020 -30828
rect 11084 -30892 11104 -30828
rect 5732 -30908 11104 -30892
rect 5732 -30972 11020 -30908
rect 11084 -30972 11104 -30908
rect 5732 -30988 11104 -30972
rect 5732 -31052 11020 -30988
rect 11084 -31052 11104 -30988
rect 5732 -31068 11104 -31052
rect 5732 -31132 11020 -31068
rect 11084 -31132 11104 -31068
rect 5732 -31148 11104 -31132
rect 5732 -31212 11020 -31148
rect 11084 -31212 11104 -31148
rect 5732 -31228 11104 -31212
rect 5732 -31292 11020 -31228
rect 11084 -31292 11104 -31228
rect 5732 -31308 11104 -31292
rect 5732 -31372 11020 -31308
rect 11084 -31372 11104 -31308
rect 5732 -31388 11104 -31372
rect 5732 -31452 11020 -31388
rect 11084 -31452 11104 -31388
rect 5732 -31468 11104 -31452
rect 5732 -31532 11020 -31468
rect 11084 -31532 11104 -31468
rect 5732 -31548 11104 -31532
rect 5732 -31612 11020 -31548
rect 11084 -31612 11104 -31548
rect 5732 -31628 11104 -31612
rect 5732 -31692 11020 -31628
rect 11084 -31692 11104 -31628
rect 5732 -31708 11104 -31692
rect 5732 -31772 11020 -31708
rect 11084 -31772 11104 -31708
rect 5732 -31800 11104 -31772
rect 11344 -26748 16716 -26720
rect 11344 -26812 16632 -26748
rect 16696 -26812 16716 -26748
rect 11344 -26828 16716 -26812
rect 11344 -26892 16632 -26828
rect 16696 -26892 16716 -26828
rect 11344 -26908 16716 -26892
rect 11344 -26972 16632 -26908
rect 16696 -26972 16716 -26908
rect 11344 -26988 16716 -26972
rect 11344 -27052 16632 -26988
rect 16696 -27052 16716 -26988
rect 11344 -27068 16716 -27052
rect 11344 -27132 16632 -27068
rect 16696 -27132 16716 -27068
rect 11344 -27148 16716 -27132
rect 11344 -27212 16632 -27148
rect 16696 -27212 16716 -27148
rect 11344 -27228 16716 -27212
rect 11344 -27292 16632 -27228
rect 16696 -27292 16716 -27228
rect 11344 -27308 16716 -27292
rect 11344 -27372 16632 -27308
rect 16696 -27372 16716 -27308
rect 11344 -27388 16716 -27372
rect 11344 -27452 16632 -27388
rect 16696 -27452 16716 -27388
rect 11344 -27468 16716 -27452
rect 11344 -27532 16632 -27468
rect 16696 -27532 16716 -27468
rect 11344 -27548 16716 -27532
rect 11344 -27612 16632 -27548
rect 16696 -27612 16716 -27548
rect 11344 -27628 16716 -27612
rect 11344 -27692 16632 -27628
rect 16696 -27692 16716 -27628
rect 11344 -27708 16716 -27692
rect 11344 -27772 16632 -27708
rect 16696 -27772 16716 -27708
rect 11344 -27788 16716 -27772
rect 11344 -27852 16632 -27788
rect 16696 -27852 16716 -27788
rect 11344 -27868 16716 -27852
rect 11344 -27932 16632 -27868
rect 16696 -27932 16716 -27868
rect 11344 -27948 16716 -27932
rect 11344 -28012 16632 -27948
rect 16696 -28012 16716 -27948
rect 11344 -28028 16716 -28012
rect 11344 -28092 16632 -28028
rect 16696 -28092 16716 -28028
rect 11344 -28108 16716 -28092
rect 11344 -28172 16632 -28108
rect 16696 -28172 16716 -28108
rect 11344 -28188 16716 -28172
rect 11344 -28252 16632 -28188
rect 16696 -28252 16716 -28188
rect 11344 -28268 16716 -28252
rect 11344 -28332 16632 -28268
rect 16696 -28332 16716 -28268
rect 11344 -28348 16716 -28332
rect 11344 -28412 16632 -28348
rect 16696 -28412 16716 -28348
rect 11344 -28428 16716 -28412
rect 11344 -28492 16632 -28428
rect 16696 -28492 16716 -28428
rect 11344 -28508 16716 -28492
rect 11344 -28572 16632 -28508
rect 16696 -28572 16716 -28508
rect 11344 -28588 16716 -28572
rect 11344 -28652 16632 -28588
rect 16696 -28652 16716 -28588
rect 11344 -28668 16716 -28652
rect 11344 -28732 16632 -28668
rect 16696 -28732 16716 -28668
rect 11344 -28748 16716 -28732
rect 11344 -28812 16632 -28748
rect 16696 -28812 16716 -28748
rect 11344 -28828 16716 -28812
rect 11344 -28892 16632 -28828
rect 16696 -28892 16716 -28828
rect 11344 -28908 16716 -28892
rect 11344 -28972 16632 -28908
rect 16696 -28972 16716 -28908
rect 11344 -28988 16716 -28972
rect 11344 -29052 16632 -28988
rect 16696 -29052 16716 -28988
rect 11344 -29068 16716 -29052
rect 11344 -29132 16632 -29068
rect 16696 -29132 16716 -29068
rect 11344 -29148 16716 -29132
rect 11344 -29212 16632 -29148
rect 16696 -29212 16716 -29148
rect 11344 -29228 16716 -29212
rect 11344 -29292 16632 -29228
rect 16696 -29292 16716 -29228
rect 11344 -29308 16716 -29292
rect 11344 -29372 16632 -29308
rect 16696 -29372 16716 -29308
rect 11344 -29388 16716 -29372
rect 11344 -29452 16632 -29388
rect 16696 -29452 16716 -29388
rect 11344 -29468 16716 -29452
rect 11344 -29532 16632 -29468
rect 16696 -29532 16716 -29468
rect 11344 -29548 16716 -29532
rect 11344 -29612 16632 -29548
rect 16696 -29612 16716 -29548
rect 11344 -29628 16716 -29612
rect 11344 -29692 16632 -29628
rect 16696 -29692 16716 -29628
rect 11344 -29708 16716 -29692
rect 11344 -29772 16632 -29708
rect 16696 -29772 16716 -29708
rect 11344 -29788 16716 -29772
rect 11344 -29852 16632 -29788
rect 16696 -29852 16716 -29788
rect 11344 -29868 16716 -29852
rect 11344 -29932 16632 -29868
rect 16696 -29932 16716 -29868
rect 11344 -29948 16716 -29932
rect 11344 -30012 16632 -29948
rect 16696 -30012 16716 -29948
rect 11344 -30028 16716 -30012
rect 11344 -30092 16632 -30028
rect 16696 -30092 16716 -30028
rect 11344 -30108 16716 -30092
rect 11344 -30172 16632 -30108
rect 16696 -30172 16716 -30108
rect 11344 -30188 16716 -30172
rect 11344 -30252 16632 -30188
rect 16696 -30252 16716 -30188
rect 11344 -30268 16716 -30252
rect 11344 -30332 16632 -30268
rect 16696 -30332 16716 -30268
rect 11344 -30348 16716 -30332
rect 11344 -30412 16632 -30348
rect 16696 -30412 16716 -30348
rect 11344 -30428 16716 -30412
rect 11344 -30492 16632 -30428
rect 16696 -30492 16716 -30428
rect 11344 -30508 16716 -30492
rect 11344 -30572 16632 -30508
rect 16696 -30572 16716 -30508
rect 11344 -30588 16716 -30572
rect 11344 -30652 16632 -30588
rect 16696 -30652 16716 -30588
rect 11344 -30668 16716 -30652
rect 11344 -30732 16632 -30668
rect 16696 -30732 16716 -30668
rect 11344 -30748 16716 -30732
rect 11344 -30812 16632 -30748
rect 16696 -30812 16716 -30748
rect 11344 -30828 16716 -30812
rect 11344 -30892 16632 -30828
rect 16696 -30892 16716 -30828
rect 11344 -30908 16716 -30892
rect 11344 -30972 16632 -30908
rect 16696 -30972 16716 -30908
rect 11344 -30988 16716 -30972
rect 11344 -31052 16632 -30988
rect 16696 -31052 16716 -30988
rect 11344 -31068 16716 -31052
rect 11344 -31132 16632 -31068
rect 16696 -31132 16716 -31068
rect 11344 -31148 16716 -31132
rect 11344 -31212 16632 -31148
rect 16696 -31212 16716 -31148
rect 11344 -31228 16716 -31212
rect 11344 -31292 16632 -31228
rect 16696 -31292 16716 -31228
rect 11344 -31308 16716 -31292
rect 11344 -31372 16632 -31308
rect 16696 -31372 16716 -31308
rect 11344 -31388 16716 -31372
rect 11344 -31452 16632 -31388
rect 16696 -31452 16716 -31388
rect 11344 -31468 16716 -31452
rect 11344 -31532 16632 -31468
rect 16696 -31532 16716 -31468
rect 11344 -31548 16716 -31532
rect 11344 -31612 16632 -31548
rect 16696 -31612 16716 -31548
rect 11344 -31628 16716 -31612
rect 11344 -31692 16632 -31628
rect 16696 -31692 16716 -31628
rect 11344 -31708 16716 -31692
rect 11344 -31772 16632 -31708
rect 16696 -31772 16716 -31708
rect 11344 -31800 16716 -31772
rect 16956 -26748 22328 -26720
rect 16956 -26812 22244 -26748
rect 22308 -26812 22328 -26748
rect 16956 -26828 22328 -26812
rect 16956 -26892 22244 -26828
rect 22308 -26892 22328 -26828
rect 16956 -26908 22328 -26892
rect 16956 -26972 22244 -26908
rect 22308 -26972 22328 -26908
rect 16956 -26988 22328 -26972
rect 16956 -27052 22244 -26988
rect 22308 -27052 22328 -26988
rect 16956 -27068 22328 -27052
rect 16956 -27132 22244 -27068
rect 22308 -27132 22328 -27068
rect 16956 -27148 22328 -27132
rect 16956 -27212 22244 -27148
rect 22308 -27212 22328 -27148
rect 16956 -27228 22328 -27212
rect 16956 -27292 22244 -27228
rect 22308 -27292 22328 -27228
rect 16956 -27308 22328 -27292
rect 16956 -27372 22244 -27308
rect 22308 -27372 22328 -27308
rect 16956 -27388 22328 -27372
rect 16956 -27452 22244 -27388
rect 22308 -27452 22328 -27388
rect 16956 -27468 22328 -27452
rect 16956 -27532 22244 -27468
rect 22308 -27532 22328 -27468
rect 16956 -27548 22328 -27532
rect 16956 -27612 22244 -27548
rect 22308 -27612 22328 -27548
rect 16956 -27628 22328 -27612
rect 16956 -27692 22244 -27628
rect 22308 -27692 22328 -27628
rect 16956 -27708 22328 -27692
rect 16956 -27772 22244 -27708
rect 22308 -27772 22328 -27708
rect 16956 -27788 22328 -27772
rect 16956 -27852 22244 -27788
rect 22308 -27852 22328 -27788
rect 16956 -27868 22328 -27852
rect 16956 -27932 22244 -27868
rect 22308 -27932 22328 -27868
rect 16956 -27948 22328 -27932
rect 16956 -28012 22244 -27948
rect 22308 -28012 22328 -27948
rect 16956 -28028 22328 -28012
rect 16956 -28092 22244 -28028
rect 22308 -28092 22328 -28028
rect 16956 -28108 22328 -28092
rect 16956 -28172 22244 -28108
rect 22308 -28172 22328 -28108
rect 16956 -28188 22328 -28172
rect 16956 -28252 22244 -28188
rect 22308 -28252 22328 -28188
rect 16956 -28268 22328 -28252
rect 16956 -28332 22244 -28268
rect 22308 -28332 22328 -28268
rect 16956 -28348 22328 -28332
rect 16956 -28412 22244 -28348
rect 22308 -28412 22328 -28348
rect 16956 -28428 22328 -28412
rect 16956 -28492 22244 -28428
rect 22308 -28492 22328 -28428
rect 16956 -28508 22328 -28492
rect 16956 -28572 22244 -28508
rect 22308 -28572 22328 -28508
rect 16956 -28588 22328 -28572
rect 16956 -28652 22244 -28588
rect 22308 -28652 22328 -28588
rect 16956 -28668 22328 -28652
rect 16956 -28732 22244 -28668
rect 22308 -28732 22328 -28668
rect 16956 -28748 22328 -28732
rect 16956 -28812 22244 -28748
rect 22308 -28812 22328 -28748
rect 16956 -28828 22328 -28812
rect 16956 -28892 22244 -28828
rect 22308 -28892 22328 -28828
rect 16956 -28908 22328 -28892
rect 16956 -28972 22244 -28908
rect 22308 -28972 22328 -28908
rect 16956 -28988 22328 -28972
rect 16956 -29052 22244 -28988
rect 22308 -29052 22328 -28988
rect 16956 -29068 22328 -29052
rect 16956 -29132 22244 -29068
rect 22308 -29132 22328 -29068
rect 16956 -29148 22328 -29132
rect 16956 -29212 22244 -29148
rect 22308 -29212 22328 -29148
rect 16956 -29228 22328 -29212
rect 16956 -29292 22244 -29228
rect 22308 -29292 22328 -29228
rect 16956 -29308 22328 -29292
rect 16956 -29372 22244 -29308
rect 22308 -29372 22328 -29308
rect 16956 -29388 22328 -29372
rect 16956 -29452 22244 -29388
rect 22308 -29452 22328 -29388
rect 16956 -29468 22328 -29452
rect 16956 -29532 22244 -29468
rect 22308 -29532 22328 -29468
rect 16956 -29548 22328 -29532
rect 16956 -29612 22244 -29548
rect 22308 -29612 22328 -29548
rect 16956 -29628 22328 -29612
rect 16956 -29692 22244 -29628
rect 22308 -29692 22328 -29628
rect 16956 -29708 22328 -29692
rect 16956 -29772 22244 -29708
rect 22308 -29772 22328 -29708
rect 16956 -29788 22328 -29772
rect 16956 -29852 22244 -29788
rect 22308 -29852 22328 -29788
rect 16956 -29868 22328 -29852
rect 16956 -29932 22244 -29868
rect 22308 -29932 22328 -29868
rect 16956 -29948 22328 -29932
rect 16956 -30012 22244 -29948
rect 22308 -30012 22328 -29948
rect 16956 -30028 22328 -30012
rect 16956 -30092 22244 -30028
rect 22308 -30092 22328 -30028
rect 16956 -30108 22328 -30092
rect 16956 -30172 22244 -30108
rect 22308 -30172 22328 -30108
rect 16956 -30188 22328 -30172
rect 16956 -30252 22244 -30188
rect 22308 -30252 22328 -30188
rect 16956 -30268 22328 -30252
rect 16956 -30332 22244 -30268
rect 22308 -30332 22328 -30268
rect 16956 -30348 22328 -30332
rect 16956 -30412 22244 -30348
rect 22308 -30412 22328 -30348
rect 16956 -30428 22328 -30412
rect 16956 -30492 22244 -30428
rect 22308 -30492 22328 -30428
rect 16956 -30508 22328 -30492
rect 16956 -30572 22244 -30508
rect 22308 -30572 22328 -30508
rect 16956 -30588 22328 -30572
rect 16956 -30652 22244 -30588
rect 22308 -30652 22328 -30588
rect 16956 -30668 22328 -30652
rect 16956 -30732 22244 -30668
rect 22308 -30732 22328 -30668
rect 16956 -30748 22328 -30732
rect 16956 -30812 22244 -30748
rect 22308 -30812 22328 -30748
rect 16956 -30828 22328 -30812
rect 16956 -30892 22244 -30828
rect 22308 -30892 22328 -30828
rect 16956 -30908 22328 -30892
rect 16956 -30972 22244 -30908
rect 22308 -30972 22328 -30908
rect 16956 -30988 22328 -30972
rect 16956 -31052 22244 -30988
rect 22308 -31052 22328 -30988
rect 16956 -31068 22328 -31052
rect 16956 -31132 22244 -31068
rect 22308 -31132 22328 -31068
rect 16956 -31148 22328 -31132
rect 16956 -31212 22244 -31148
rect 22308 -31212 22328 -31148
rect 16956 -31228 22328 -31212
rect 16956 -31292 22244 -31228
rect 22308 -31292 22328 -31228
rect 16956 -31308 22328 -31292
rect 16956 -31372 22244 -31308
rect 22308 -31372 22328 -31308
rect 16956 -31388 22328 -31372
rect 16956 -31452 22244 -31388
rect 22308 -31452 22328 -31388
rect 16956 -31468 22328 -31452
rect 16956 -31532 22244 -31468
rect 22308 -31532 22328 -31468
rect 16956 -31548 22328 -31532
rect 16956 -31612 22244 -31548
rect 22308 -31612 22328 -31548
rect 16956 -31628 22328 -31612
rect 16956 -31692 22244 -31628
rect 22308 -31692 22328 -31628
rect 16956 -31708 22328 -31692
rect 16956 -31772 22244 -31708
rect 22308 -31772 22328 -31708
rect 16956 -31800 22328 -31772
rect 22568 -26748 27940 -26720
rect 22568 -26812 27856 -26748
rect 27920 -26812 27940 -26748
rect 22568 -26828 27940 -26812
rect 22568 -26892 27856 -26828
rect 27920 -26892 27940 -26828
rect 22568 -26908 27940 -26892
rect 22568 -26972 27856 -26908
rect 27920 -26972 27940 -26908
rect 22568 -26988 27940 -26972
rect 22568 -27052 27856 -26988
rect 27920 -27052 27940 -26988
rect 22568 -27068 27940 -27052
rect 22568 -27132 27856 -27068
rect 27920 -27132 27940 -27068
rect 22568 -27148 27940 -27132
rect 22568 -27212 27856 -27148
rect 27920 -27212 27940 -27148
rect 22568 -27228 27940 -27212
rect 22568 -27292 27856 -27228
rect 27920 -27292 27940 -27228
rect 22568 -27308 27940 -27292
rect 22568 -27372 27856 -27308
rect 27920 -27372 27940 -27308
rect 22568 -27388 27940 -27372
rect 22568 -27452 27856 -27388
rect 27920 -27452 27940 -27388
rect 22568 -27468 27940 -27452
rect 22568 -27532 27856 -27468
rect 27920 -27532 27940 -27468
rect 22568 -27548 27940 -27532
rect 22568 -27612 27856 -27548
rect 27920 -27612 27940 -27548
rect 22568 -27628 27940 -27612
rect 22568 -27692 27856 -27628
rect 27920 -27692 27940 -27628
rect 22568 -27708 27940 -27692
rect 22568 -27772 27856 -27708
rect 27920 -27772 27940 -27708
rect 22568 -27788 27940 -27772
rect 22568 -27852 27856 -27788
rect 27920 -27852 27940 -27788
rect 22568 -27868 27940 -27852
rect 22568 -27932 27856 -27868
rect 27920 -27932 27940 -27868
rect 22568 -27948 27940 -27932
rect 22568 -28012 27856 -27948
rect 27920 -28012 27940 -27948
rect 22568 -28028 27940 -28012
rect 22568 -28092 27856 -28028
rect 27920 -28092 27940 -28028
rect 22568 -28108 27940 -28092
rect 22568 -28172 27856 -28108
rect 27920 -28172 27940 -28108
rect 22568 -28188 27940 -28172
rect 22568 -28252 27856 -28188
rect 27920 -28252 27940 -28188
rect 22568 -28268 27940 -28252
rect 22568 -28332 27856 -28268
rect 27920 -28332 27940 -28268
rect 22568 -28348 27940 -28332
rect 22568 -28412 27856 -28348
rect 27920 -28412 27940 -28348
rect 22568 -28428 27940 -28412
rect 22568 -28492 27856 -28428
rect 27920 -28492 27940 -28428
rect 22568 -28508 27940 -28492
rect 22568 -28572 27856 -28508
rect 27920 -28572 27940 -28508
rect 22568 -28588 27940 -28572
rect 22568 -28652 27856 -28588
rect 27920 -28652 27940 -28588
rect 22568 -28668 27940 -28652
rect 22568 -28732 27856 -28668
rect 27920 -28732 27940 -28668
rect 22568 -28748 27940 -28732
rect 22568 -28812 27856 -28748
rect 27920 -28812 27940 -28748
rect 22568 -28828 27940 -28812
rect 22568 -28892 27856 -28828
rect 27920 -28892 27940 -28828
rect 22568 -28908 27940 -28892
rect 22568 -28972 27856 -28908
rect 27920 -28972 27940 -28908
rect 22568 -28988 27940 -28972
rect 22568 -29052 27856 -28988
rect 27920 -29052 27940 -28988
rect 22568 -29068 27940 -29052
rect 22568 -29132 27856 -29068
rect 27920 -29132 27940 -29068
rect 22568 -29148 27940 -29132
rect 22568 -29212 27856 -29148
rect 27920 -29212 27940 -29148
rect 22568 -29228 27940 -29212
rect 22568 -29292 27856 -29228
rect 27920 -29292 27940 -29228
rect 22568 -29308 27940 -29292
rect 22568 -29372 27856 -29308
rect 27920 -29372 27940 -29308
rect 22568 -29388 27940 -29372
rect 22568 -29452 27856 -29388
rect 27920 -29452 27940 -29388
rect 22568 -29468 27940 -29452
rect 22568 -29532 27856 -29468
rect 27920 -29532 27940 -29468
rect 22568 -29548 27940 -29532
rect 22568 -29612 27856 -29548
rect 27920 -29612 27940 -29548
rect 22568 -29628 27940 -29612
rect 22568 -29692 27856 -29628
rect 27920 -29692 27940 -29628
rect 22568 -29708 27940 -29692
rect 22568 -29772 27856 -29708
rect 27920 -29772 27940 -29708
rect 22568 -29788 27940 -29772
rect 22568 -29852 27856 -29788
rect 27920 -29852 27940 -29788
rect 22568 -29868 27940 -29852
rect 22568 -29932 27856 -29868
rect 27920 -29932 27940 -29868
rect 22568 -29948 27940 -29932
rect 22568 -30012 27856 -29948
rect 27920 -30012 27940 -29948
rect 22568 -30028 27940 -30012
rect 22568 -30092 27856 -30028
rect 27920 -30092 27940 -30028
rect 22568 -30108 27940 -30092
rect 22568 -30172 27856 -30108
rect 27920 -30172 27940 -30108
rect 22568 -30188 27940 -30172
rect 22568 -30252 27856 -30188
rect 27920 -30252 27940 -30188
rect 22568 -30268 27940 -30252
rect 22568 -30332 27856 -30268
rect 27920 -30332 27940 -30268
rect 22568 -30348 27940 -30332
rect 22568 -30412 27856 -30348
rect 27920 -30412 27940 -30348
rect 22568 -30428 27940 -30412
rect 22568 -30492 27856 -30428
rect 27920 -30492 27940 -30428
rect 22568 -30508 27940 -30492
rect 22568 -30572 27856 -30508
rect 27920 -30572 27940 -30508
rect 22568 -30588 27940 -30572
rect 22568 -30652 27856 -30588
rect 27920 -30652 27940 -30588
rect 22568 -30668 27940 -30652
rect 22568 -30732 27856 -30668
rect 27920 -30732 27940 -30668
rect 22568 -30748 27940 -30732
rect 22568 -30812 27856 -30748
rect 27920 -30812 27940 -30748
rect 22568 -30828 27940 -30812
rect 22568 -30892 27856 -30828
rect 27920 -30892 27940 -30828
rect 22568 -30908 27940 -30892
rect 22568 -30972 27856 -30908
rect 27920 -30972 27940 -30908
rect 22568 -30988 27940 -30972
rect 22568 -31052 27856 -30988
rect 27920 -31052 27940 -30988
rect 22568 -31068 27940 -31052
rect 22568 -31132 27856 -31068
rect 27920 -31132 27940 -31068
rect 22568 -31148 27940 -31132
rect 22568 -31212 27856 -31148
rect 27920 -31212 27940 -31148
rect 22568 -31228 27940 -31212
rect 22568 -31292 27856 -31228
rect 27920 -31292 27940 -31228
rect 22568 -31308 27940 -31292
rect 22568 -31372 27856 -31308
rect 27920 -31372 27940 -31308
rect 22568 -31388 27940 -31372
rect 22568 -31452 27856 -31388
rect 27920 -31452 27940 -31388
rect 22568 -31468 27940 -31452
rect 22568 -31532 27856 -31468
rect 27920 -31532 27940 -31468
rect 22568 -31548 27940 -31532
rect 22568 -31612 27856 -31548
rect 27920 -31612 27940 -31548
rect 22568 -31628 27940 -31612
rect 22568 -31692 27856 -31628
rect 27920 -31692 27940 -31628
rect 22568 -31708 27940 -31692
rect 22568 -31772 27856 -31708
rect 27920 -31772 27940 -31708
rect 22568 -31800 27940 -31772
rect 28180 -26748 33552 -26720
rect 28180 -26812 33468 -26748
rect 33532 -26812 33552 -26748
rect 28180 -26828 33552 -26812
rect 28180 -26892 33468 -26828
rect 33532 -26892 33552 -26828
rect 28180 -26908 33552 -26892
rect 28180 -26972 33468 -26908
rect 33532 -26972 33552 -26908
rect 28180 -26988 33552 -26972
rect 28180 -27052 33468 -26988
rect 33532 -27052 33552 -26988
rect 28180 -27068 33552 -27052
rect 28180 -27132 33468 -27068
rect 33532 -27132 33552 -27068
rect 28180 -27148 33552 -27132
rect 28180 -27212 33468 -27148
rect 33532 -27212 33552 -27148
rect 28180 -27228 33552 -27212
rect 28180 -27292 33468 -27228
rect 33532 -27292 33552 -27228
rect 28180 -27308 33552 -27292
rect 28180 -27372 33468 -27308
rect 33532 -27372 33552 -27308
rect 28180 -27388 33552 -27372
rect 28180 -27452 33468 -27388
rect 33532 -27452 33552 -27388
rect 28180 -27468 33552 -27452
rect 28180 -27532 33468 -27468
rect 33532 -27532 33552 -27468
rect 28180 -27548 33552 -27532
rect 28180 -27612 33468 -27548
rect 33532 -27612 33552 -27548
rect 28180 -27628 33552 -27612
rect 28180 -27692 33468 -27628
rect 33532 -27692 33552 -27628
rect 28180 -27708 33552 -27692
rect 28180 -27772 33468 -27708
rect 33532 -27772 33552 -27708
rect 28180 -27788 33552 -27772
rect 28180 -27852 33468 -27788
rect 33532 -27852 33552 -27788
rect 28180 -27868 33552 -27852
rect 28180 -27932 33468 -27868
rect 33532 -27932 33552 -27868
rect 28180 -27948 33552 -27932
rect 28180 -28012 33468 -27948
rect 33532 -28012 33552 -27948
rect 28180 -28028 33552 -28012
rect 28180 -28092 33468 -28028
rect 33532 -28092 33552 -28028
rect 28180 -28108 33552 -28092
rect 28180 -28172 33468 -28108
rect 33532 -28172 33552 -28108
rect 28180 -28188 33552 -28172
rect 28180 -28252 33468 -28188
rect 33532 -28252 33552 -28188
rect 28180 -28268 33552 -28252
rect 28180 -28332 33468 -28268
rect 33532 -28332 33552 -28268
rect 28180 -28348 33552 -28332
rect 28180 -28412 33468 -28348
rect 33532 -28412 33552 -28348
rect 28180 -28428 33552 -28412
rect 28180 -28492 33468 -28428
rect 33532 -28492 33552 -28428
rect 28180 -28508 33552 -28492
rect 28180 -28572 33468 -28508
rect 33532 -28572 33552 -28508
rect 28180 -28588 33552 -28572
rect 28180 -28652 33468 -28588
rect 33532 -28652 33552 -28588
rect 28180 -28668 33552 -28652
rect 28180 -28732 33468 -28668
rect 33532 -28732 33552 -28668
rect 28180 -28748 33552 -28732
rect 28180 -28812 33468 -28748
rect 33532 -28812 33552 -28748
rect 28180 -28828 33552 -28812
rect 28180 -28892 33468 -28828
rect 33532 -28892 33552 -28828
rect 28180 -28908 33552 -28892
rect 28180 -28972 33468 -28908
rect 33532 -28972 33552 -28908
rect 28180 -28988 33552 -28972
rect 28180 -29052 33468 -28988
rect 33532 -29052 33552 -28988
rect 28180 -29068 33552 -29052
rect 28180 -29132 33468 -29068
rect 33532 -29132 33552 -29068
rect 28180 -29148 33552 -29132
rect 28180 -29212 33468 -29148
rect 33532 -29212 33552 -29148
rect 28180 -29228 33552 -29212
rect 28180 -29292 33468 -29228
rect 33532 -29292 33552 -29228
rect 28180 -29308 33552 -29292
rect 28180 -29372 33468 -29308
rect 33532 -29372 33552 -29308
rect 28180 -29388 33552 -29372
rect 28180 -29452 33468 -29388
rect 33532 -29452 33552 -29388
rect 28180 -29468 33552 -29452
rect 28180 -29532 33468 -29468
rect 33532 -29532 33552 -29468
rect 28180 -29548 33552 -29532
rect 28180 -29612 33468 -29548
rect 33532 -29612 33552 -29548
rect 28180 -29628 33552 -29612
rect 28180 -29692 33468 -29628
rect 33532 -29692 33552 -29628
rect 28180 -29708 33552 -29692
rect 28180 -29772 33468 -29708
rect 33532 -29772 33552 -29708
rect 28180 -29788 33552 -29772
rect 28180 -29852 33468 -29788
rect 33532 -29852 33552 -29788
rect 28180 -29868 33552 -29852
rect 28180 -29932 33468 -29868
rect 33532 -29932 33552 -29868
rect 28180 -29948 33552 -29932
rect 28180 -30012 33468 -29948
rect 33532 -30012 33552 -29948
rect 28180 -30028 33552 -30012
rect 28180 -30092 33468 -30028
rect 33532 -30092 33552 -30028
rect 28180 -30108 33552 -30092
rect 28180 -30172 33468 -30108
rect 33532 -30172 33552 -30108
rect 28180 -30188 33552 -30172
rect 28180 -30252 33468 -30188
rect 33532 -30252 33552 -30188
rect 28180 -30268 33552 -30252
rect 28180 -30332 33468 -30268
rect 33532 -30332 33552 -30268
rect 28180 -30348 33552 -30332
rect 28180 -30412 33468 -30348
rect 33532 -30412 33552 -30348
rect 28180 -30428 33552 -30412
rect 28180 -30492 33468 -30428
rect 33532 -30492 33552 -30428
rect 28180 -30508 33552 -30492
rect 28180 -30572 33468 -30508
rect 33532 -30572 33552 -30508
rect 28180 -30588 33552 -30572
rect 28180 -30652 33468 -30588
rect 33532 -30652 33552 -30588
rect 28180 -30668 33552 -30652
rect 28180 -30732 33468 -30668
rect 33532 -30732 33552 -30668
rect 28180 -30748 33552 -30732
rect 28180 -30812 33468 -30748
rect 33532 -30812 33552 -30748
rect 28180 -30828 33552 -30812
rect 28180 -30892 33468 -30828
rect 33532 -30892 33552 -30828
rect 28180 -30908 33552 -30892
rect 28180 -30972 33468 -30908
rect 33532 -30972 33552 -30908
rect 28180 -30988 33552 -30972
rect 28180 -31052 33468 -30988
rect 33532 -31052 33552 -30988
rect 28180 -31068 33552 -31052
rect 28180 -31132 33468 -31068
rect 33532 -31132 33552 -31068
rect 28180 -31148 33552 -31132
rect 28180 -31212 33468 -31148
rect 33532 -31212 33552 -31148
rect 28180 -31228 33552 -31212
rect 28180 -31292 33468 -31228
rect 33532 -31292 33552 -31228
rect 28180 -31308 33552 -31292
rect 28180 -31372 33468 -31308
rect 33532 -31372 33552 -31308
rect 28180 -31388 33552 -31372
rect 28180 -31452 33468 -31388
rect 33532 -31452 33552 -31388
rect 28180 -31468 33552 -31452
rect 28180 -31532 33468 -31468
rect 33532 -31532 33552 -31468
rect 28180 -31548 33552 -31532
rect 28180 -31612 33468 -31548
rect 33532 -31612 33552 -31548
rect 28180 -31628 33552 -31612
rect 28180 -31692 33468 -31628
rect 33532 -31692 33552 -31628
rect 28180 -31708 33552 -31692
rect 28180 -31772 33468 -31708
rect 33532 -31772 33552 -31708
rect 28180 -31800 33552 -31772
rect 33792 -26748 39164 -26720
rect 33792 -26812 39080 -26748
rect 39144 -26812 39164 -26748
rect 33792 -26828 39164 -26812
rect 33792 -26892 39080 -26828
rect 39144 -26892 39164 -26828
rect 33792 -26908 39164 -26892
rect 33792 -26972 39080 -26908
rect 39144 -26972 39164 -26908
rect 33792 -26988 39164 -26972
rect 33792 -27052 39080 -26988
rect 39144 -27052 39164 -26988
rect 33792 -27068 39164 -27052
rect 33792 -27132 39080 -27068
rect 39144 -27132 39164 -27068
rect 33792 -27148 39164 -27132
rect 33792 -27212 39080 -27148
rect 39144 -27212 39164 -27148
rect 33792 -27228 39164 -27212
rect 33792 -27292 39080 -27228
rect 39144 -27292 39164 -27228
rect 33792 -27308 39164 -27292
rect 33792 -27372 39080 -27308
rect 39144 -27372 39164 -27308
rect 33792 -27388 39164 -27372
rect 33792 -27452 39080 -27388
rect 39144 -27452 39164 -27388
rect 33792 -27468 39164 -27452
rect 33792 -27532 39080 -27468
rect 39144 -27532 39164 -27468
rect 33792 -27548 39164 -27532
rect 33792 -27612 39080 -27548
rect 39144 -27612 39164 -27548
rect 33792 -27628 39164 -27612
rect 33792 -27692 39080 -27628
rect 39144 -27692 39164 -27628
rect 33792 -27708 39164 -27692
rect 33792 -27772 39080 -27708
rect 39144 -27772 39164 -27708
rect 33792 -27788 39164 -27772
rect 33792 -27852 39080 -27788
rect 39144 -27852 39164 -27788
rect 33792 -27868 39164 -27852
rect 33792 -27932 39080 -27868
rect 39144 -27932 39164 -27868
rect 33792 -27948 39164 -27932
rect 33792 -28012 39080 -27948
rect 39144 -28012 39164 -27948
rect 33792 -28028 39164 -28012
rect 33792 -28092 39080 -28028
rect 39144 -28092 39164 -28028
rect 33792 -28108 39164 -28092
rect 33792 -28172 39080 -28108
rect 39144 -28172 39164 -28108
rect 33792 -28188 39164 -28172
rect 33792 -28252 39080 -28188
rect 39144 -28252 39164 -28188
rect 33792 -28268 39164 -28252
rect 33792 -28332 39080 -28268
rect 39144 -28332 39164 -28268
rect 33792 -28348 39164 -28332
rect 33792 -28412 39080 -28348
rect 39144 -28412 39164 -28348
rect 33792 -28428 39164 -28412
rect 33792 -28492 39080 -28428
rect 39144 -28492 39164 -28428
rect 33792 -28508 39164 -28492
rect 33792 -28572 39080 -28508
rect 39144 -28572 39164 -28508
rect 33792 -28588 39164 -28572
rect 33792 -28652 39080 -28588
rect 39144 -28652 39164 -28588
rect 33792 -28668 39164 -28652
rect 33792 -28732 39080 -28668
rect 39144 -28732 39164 -28668
rect 33792 -28748 39164 -28732
rect 33792 -28812 39080 -28748
rect 39144 -28812 39164 -28748
rect 33792 -28828 39164 -28812
rect 33792 -28892 39080 -28828
rect 39144 -28892 39164 -28828
rect 33792 -28908 39164 -28892
rect 33792 -28972 39080 -28908
rect 39144 -28972 39164 -28908
rect 33792 -28988 39164 -28972
rect 33792 -29052 39080 -28988
rect 39144 -29052 39164 -28988
rect 33792 -29068 39164 -29052
rect 33792 -29132 39080 -29068
rect 39144 -29132 39164 -29068
rect 33792 -29148 39164 -29132
rect 33792 -29212 39080 -29148
rect 39144 -29212 39164 -29148
rect 33792 -29228 39164 -29212
rect 33792 -29292 39080 -29228
rect 39144 -29292 39164 -29228
rect 33792 -29308 39164 -29292
rect 33792 -29372 39080 -29308
rect 39144 -29372 39164 -29308
rect 33792 -29388 39164 -29372
rect 33792 -29452 39080 -29388
rect 39144 -29452 39164 -29388
rect 33792 -29468 39164 -29452
rect 33792 -29532 39080 -29468
rect 39144 -29532 39164 -29468
rect 33792 -29548 39164 -29532
rect 33792 -29612 39080 -29548
rect 39144 -29612 39164 -29548
rect 33792 -29628 39164 -29612
rect 33792 -29692 39080 -29628
rect 39144 -29692 39164 -29628
rect 33792 -29708 39164 -29692
rect 33792 -29772 39080 -29708
rect 39144 -29772 39164 -29708
rect 33792 -29788 39164 -29772
rect 33792 -29852 39080 -29788
rect 39144 -29852 39164 -29788
rect 33792 -29868 39164 -29852
rect 33792 -29932 39080 -29868
rect 39144 -29932 39164 -29868
rect 33792 -29948 39164 -29932
rect 33792 -30012 39080 -29948
rect 39144 -30012 39164 -29948
rect 33792 -30028 39164 -30012
rect 33792 -30092 39080 -30028
rect 39144 -30092 39164 -30028
rect 33792 -30108 39164 -30092
rect 33792 -30172 39080 -30108
rect 39144 -30172 39164 -30108
rect 33792 -30188 39164 -30172
rect 33792 -30252 39080 -30188
rect 39144 -30252 39164 -30188
rect 33792 -30268 39164 -30252
rect 33792 -30332 39080 -30268
rect 39144 -30332 39164 -30268
rect 33792 -30348 39164 -30332
rect 33792 -30412 39080 -30348
rect 39144 -30412 39164 -30348
rect 33792 -30428 39164 -30412
rect 33792 -30492 39080 -30428
rect 39144 -30492 39164 -30428
rect 33792 -30508 39164 -30492
rect 33792 -30572 39080 -30508
rect 39144 -30572 39164 -30508
rect 33792 -30588 39164 -30572
rect 33792 -30652 39080 -30588
rect 39144 -30652 39164 -30588
rect 33792 -30668 39164 -30652
rect 33792 -30732 39080 -30668
rect 39144 -30732 39164 -30668
rect 33792 -30748 39164 -30732
rect 33792 -30812 39080 -30748
rect 39144 -30812 39164 -30748
rect 33792 -30828 39164 -30812
rect 33792 -30892 39080 -30828
rect 39144 -30892 39164 -30828
rect 33792 -30908 39164 -30892
rect 33792 -30972 39080 -30908
rect 39144 -30972 39164 -30908
rect 33792 -30988 39164 -30972
rect 33792 -31052 39080 -30988
rect 39144 -31052 39164 -30988
rect 33792 -31068 39164 -31052
rect 33792 -31132 39080 -31068
rect 39144 -31132 39164 -31068
rect 33792 -31148 39164 -31132
rect 33792 -31212 39080 -31148
rect 39144 -31212 39164 -31148
rect 33792 -31228 39164 -31212
rect 33792 -31292 39080 -31228
rect 39144 -31292 39164 -31228
rect 33792 -31308 39164 -31292
rect 33792 -31372 39080 -31308
rect 39144 -31372 39164 -31308
rect 33792 -31388 39164 -31372
rect 33792 -31452 39080 -31388
rect 39144 -31452 39164 -31388
rect 33792 -31468 39164 -31452
rect 33792 -31532 39080 -31468
rect 39144 -31532 39164 -31468
rect 33792 -31548 39164 -31532
rect 33792 -31612 39080 -31548
rect 39144 -31612 39164 -31548
rect 33792 -31628 39164 -31612
rect 33792 -31692 39080 -31628
rect 39144 -31692 39164 -31628
rect 33792 -31708 39164 -31692
rect 33792 -31772 39080 -31708
rect 39144 -31772 39164 -31708
rect 33792 -31800 39164 -31772
rect -39164 -32068 -33792 -32040
rect -39164 -32132 -33876 -32068
rect -33812 -32132 -33792 -32068
rect -39164 -32148 -33792 -32132
rect -39164 -32212 -33876 -32148
rect -33812 -32212 -33792 -32148
rect -39164 -32228 -33792 -32212
rect -39164 -32292 -33876 -32228
rect -33812 -32292 -33792 -32228
rect -39164 -32308 -33792 -32292
rect -39164 -32372 -33876 -32308
rect -33812 -32372 -33792 -32308
rect -39164 -32388 -33792 -32372
rect -39164 -32452 -33876 -32388
rect -33812 -32452 -33792 -32388
rect -39164 -32468 -33792 -32452
rect -39164 -32532 -33876 -32468
rect -33812 -32532 -33792 -32468
rect -39164 -32548 -33792 -32532
rect -39164 -32612 -33876 -32548
rect -33812 -32612 -33792 -32548
rect -39164 -32628 -33792 -32612
rect -39164 -32692 -33876 -32628
rect -33812 -32692 -33792 -32628
rect -39164 -32708 -33792 -32692
rect -39164 -32772 -33876 -32708
rect -33812 -32772 -33792 -32708
rect -39164 -32788 -33792 -32772
rect -39164 -32852 -33876 -32788
rect -33812 -32852 -33792 -32788
rect -39164 -32868 -33792 -32852
rect -39164 -32932 -33876 -32868
rect -33812 -32932 -33792 -32868
rect -39164 -32948 -33792 -32932
rect -39164 -33012 -33876 -32948
rect -33812 -33012 -33792 -32948
rect -39164 -33028 -33792 -33012
rect -39164 -33092 -33876 -33028
rect -33812 -33092 -33792 -33028
rect -39164 -33108 -33792 -33092
rect -39164 -33172 -33876 -33108
rect -33812 -33172 -33792 -33108
rect -39164 -33188 -33792 -33172
rect -39164 -33252 -33876 -33188
rect -33812 -33252 -33792 -33188
rect -39164 -33268 -33792 -33252
rect -39164 -33332 -33876 -33268
rect -33812 -33332 -33792 -33268
rect -39164 -33348 -33792 -33332
rect -39164 -33412 -33876 -33348
rect -33812 -33412 -33792 -33348
rect -39164 -33428 -33792 -33412
rect -39164 -33492 -33876 -33428
rect -33812 -33492 -33792 -33428
rect -39164 -33508 -33792 -33492
rect -39164 -33572 -33876 -33508
rect -33812 -33572 -33792 -33508
rect -39164 -33588 -33792 -33572
rect -39164 -33652 -33876 -33588
rect -33812 -33652 -33792 -33588
rect -39164 -33668 -33792 -33652
rect -39164 -33732 -33876 -33668
rect -33812 -33732 -33792 -33668
rect -39164 -33748 -33792 -33732
rect -39164 -33812 -33876 -33748
rect -33812 -33812 -33792 -33748
rect -39164 -33828 -33792 -33812
rect -39164 -33892 -33876 -33828
rect -33812 -33892 -33792 -33828
rect -39164 -33908 -33792 -33892
rect -39164 -33972 -33876 -33908
rect -33812 -33972 -33792 -33908
rect -39164 -33988 -33792 -33972
rect -39164 -34052 -33876 -33988
rect -33812 -34052 -33792 -33988
rect -39164 -34068 -33792 -34052
rect -39164 -34132 -33876 -34068
rect -33812 -34132 -33792 -34068
rect -39164 -34148 -33792 -34132
rect -39164 -34212 -33876 -34148
rect -33812 -34212 -33792 -34148
rect -39164 -34228 -33792 -34212
rect -39164 -34292 -33876 -34228
rect -33812 -34292 -33792 -34228
rect -39164 -34308 -33792 -34292
rect -39164 -34372 -33876 -34308
rect -33812 -34372 -33792 -34308
rect -39164 -34388 -33792 -34372
rect -39164 -34452 -33876 -34388
rect -33812 -34452 -33792 -34388
rect -39164 -34468 -33792 -34452
rect -39164 -34532 -33876 -34468
rect -33812 -34532 -33792 -34468
rect -39164 -34548 -33792 -34532
rect -39164 -34612 -33876 -34548
rect -33812 -34612 -33792 -34548
rect -39164 -34628 -33792 -34612
rect -39164 -34692 -33876 -34628
rect -33812 -34692 -33792 -34628
rect -39164 -34708 -33792 -34692
rect -39164 -34772 -33876 -34708
rect -33812 -34772 -33792 -34708
rect -39164 -34788 -33792 -34772
rect -39164 -34852 -33876 -34788
rect -33812 -34852 -33792 -34788
rect -39164 -34868 -33792 -34852
rect -39164 -34932 -33876 -34868
rect -33812 -34932 -33792 -34868
rect -39164 -34948 -33792 -34932
rect -39164 -35012 -33876 -34948
rect -33812 -35012 -33792 -34948
rect -39164 -35028 -33792 -35012
rect -39164 -35092 -33876 -35028
rect -33812 -35092 -33792 -35028
rect -39164 -35108 -33792 -35092
rect -39164 -35172 -33876 -35108
rect -33812 -35172 -33792 -35108
rect -39164 -35188 -33792 -35172
rect -39164 -35252 -33876 -35188
rect -33812 -35252 -33792 -35188
rect -39164 -35268 -33792 -35252
rect -39164 -35332 -33876 -35268
rect -33812 -35332 -33792 -35268
rect -39164 -35348 -33792 -35332
rect -39164 -35412 -33876 -35348
rect -33812 -35412 -33792 -35348
rect -39164 -35428 -33792 -35412
rect -39164 -35492 -33876 -35428
rect -33812 -35492 -33792 -35428
rect -39164 -35508 -33792 -35492
rect -39164 -35572 -33876 -35508
rect -33812 -35572 -33792 -35508
rect -39164 -35588 -33792 -35572
rect -39164 -35652 -33876 -35588
rect -33812 -35652 -33792 -35588
rect -39164 -35668 -33792 -35652
rect -39164 -35732 -33876 -35668
rect -33812 -35732 -33792 -35668
rect -39164 -35748 -33792 -35732
rect -39164 -35812 -33876 -35748
rect -33812 -35812 -33792 -35748
rect -39164 -35828 -33792 -35812
rect -39164 -35892 -33876 -35828
rect -33812 -35892 -33792 -35828
rect -39164 -35908 -33792 -35892
rect -39164 -35972 -33876 -35908
rect -33812 -35972 -33792 -35908
rect -39164 -35988 -33792 -35972
rect -39164 -36052 -33876 -35988
rect -33812 -36052 -33792 -35988
rect -39164 -36068 -33792 -36052
rect -39164 -36132 -33876 -36068
rect -33812 -36132 -33792 -36068
rect -39164 -36148 -33792 -36132
rect -39164 -36212 -33876 -36148
rect -33812 -36212 -33792 -36148
rect -39164 -36228 -33792 -36212
rect -39164 -36292 -33876 -36228
rect -33812 -36292 -33792 -36228
rect -39164 -36308 -33792 -36292
rect -39164 -36372 -33876 -36308
rect -33812 -36372 -33792 -36308
rect -39164 -36388 -33792 -36372
rect -39164 -36452 -33876 -36388
rect -33812 -36452 -33792 -36388
rect -39164 -36468 -33792 -36452
rect -39164 -36532 -33876 -36468
rect -33812 -36532 -33792 -36468
rect -39164 -36548 -33792 -36532
rect -39164 -36612 -33876 -36548
rect -33812 -36612 -33792 -36548
rect -39164 -36628 -33792 -36612
rect -39164 -36692 -33876 -36628
rect -33812 -36692 -33792 -36628
rect -39164 -36708 -33792 -36692
rect -39164 -36772 -33876 -36708
rect -33812 -36772 -33792 -36708
rect -39164 -36788 -33792 -36772
rect -39164 -36852 -33876 -36788
rect -33812 -36852 -33792 -36788
rect -39164 -36868 -33792 -36852
rect -39164 -36932 -33876 -36868
rect -33812 -36932 -33792 -36868
rect -39164 -36948 -33792 -36932
rect -39164 -37012 -33876 -36948
rect -33812 -37012 -33792 -36948
rect -39164 -37028 -33792 -37012
rect -39164 -37092 -33876 -37028
rect -33812 -37092 -33792 -37028
rect -39164 -37120 -33792 -37092
rect -33552 -32068 -28180 -32040
rect -33552 -32132 -28264 -32068
rect -28200 -32132 -28180 -32068
rect -33552 -32148 -28180 -32132
rect -33552 -32212 -28264 -32148
rect -28200 -32212 -28180 -32148
rect -33552 -32228 -28180 -32212
rect -33552 -32292 -28264 -32228
rect -28200 -32292 -28180 -32228
rect -33552 -32308 -28180 -32292
rect -33552 -32372 -28264 -32308
rect -28200 -32372 -28180 -32308
rect -33552 -32388 -28180 -32372
rect -33552 -32452 -28264 -32388
rect -28200 -32452 -28180 -32388
rect -33552 -32468 -28180 -32452
rect -33552 -32532 -28264 -32468
rect -28200 -32532 -28180 -32468
rect -33552 -32548 -28180 -32532
rect -33552 -32612 -28264 -32548
rect -28200 -32612 -28180 -32548
rect -33552 -32628 -28180 -32612
rect -33552 -32692 -28264 -32628
rect -28200 -32692 -28180 -32628
rect -33552 -32708 -28180 -32692
rect -33552 -32772 -28264 -32708
rect -28200 -32772 -28180 -32708
rect -33552 -32788 -28180 -32772
rect -33552 -32852 -28264 -32788
rect -28200 -32852 -28180 -32788
rect -33552 -32868 -28180 -32852
rect -33552 -32932 -28264 -32868
rect -28200 -32932 -28180 -32868
rect -33552 -32948 -28180 -32932
rect -33552 -33012 -28264 -32948
rect -28200 -33012 -28180 -32948
rect -33552 -33028 -28180 -33012
rect -33552 -33092 -28264 -33028
rect -28200 -33092 -28180 -33028
rect -33552 -33108 -28180 -33092
rect -33552 -33172 -28264 -33108
rect -28200 -33172 -28180 -33108
rect -33552 -33188 -28180 -33172
rect -33552 -33252 -28264 -33188
rect -28200 -33252 -28180 -33188
rect -33552 -33268 -28180 -33252
rect -33552 -33332 -28264 -33268
rect -28200 -33332 -28180 -33268
rect -33552 -33348 -28180 -33332
rect -33552 -33412 -28264 -33348
rect -28200 -33412 -28180 -33348
rect -33552 -33428 -28180 -33412
rect -33552 -33492 -28264 -33428
rect -28200 -33492 -28180 -33428
rect -33552 -33508 -28180 -33492
rect -33552 -33572 -28264 -33508
rect -28200 -33572 -28180 -33508
rect -33552 -33588 -28180 -33572
rect -33552 -33652 -28264 -33588
rect -28200 -33652 -28180 -33588
rect -33552 -33668 -28180 -33652
rect -33552 -33732 -28264 -33668
rect -28200 -33732 -28180 -33668
rect -33552 -33748 -28180 -33732
rect -33552 -33812 -28264 -33748
rect -28200 -33812 -28180 -33748
rect -33552 -33828 -28180 -33812
rect -33552 -33892 -28264 -33828
rect -28200 -33892 -28180 -33828
rect -33552 -33908 -28180 -33892
rect -33552 -33972 -28264 -33908
rect -28200 -33972 -28180 -33908
rect -33552 -33988 -28180 -33972
rect -33552 -34052 -28264 -33988
rect -28200 -34052 -28180 -33988
rect -33552 -34068 -28180 -34052
rect -33552 -34132 -28264 -34068
rect -28200 -34132 -28180 -34068
rect -33552 -34148 -28180 -34132
rect -33552 -34212 -28264 -34148
rect -28200 -34212 -28180 -34148
rect -33552 -34228 -28180 -34212
rect -33552 -34292 -28264 -34228
rect -28200 -34292 -28180 -34228
rect -33552 -34308 -28180 -34292
rect -33552 -34372 -28264 -34308
rect -28200 -34372 -28180 -34308
rect -33552 -34388 -28180 -34372
rect -33552 -34452 -28264 -34388
rect -28200 -34452 -28180 -34388
rect -33552 -34468 -28180 -34452
rect -33552 -34532 -28264 -34468
rect -28200 -34532 -28180 -34468
rect -33552 -34548 -28180 -34532
rect -33552 -34612 -28264 -34548
rect -28200 -34612 -28180 -34548
rect -33552 -34628 -28180 -34612
rect -33552 -34692 -28264 -34628
rect -28200 -34692 -28180 -34628
rect -33552 -34708 -28180 -34692
rect -33552 -34772 -28264 -34708
rect -28200 -34772 -28180 -34708
rect -33552 -34788 -28180 -34772
rect -33552 -34852 -28264 -34788
rect -28200 -34852 -28180 -34788
rect -33552 -34868 -28180 -34852
rect -33552 -34932 -28264 -34868
rect -28200 -34932 -28180 -34868
rect -33552 -34948 -28180 -34932
rect -33552 -35012 -28264 -34948
rect -28200 -35012 -28180 -34948
rect -33552 -35028 -28180 -35012
rect -33552 -35092 -28264 -35028
rect -28200 -35092 -28180 -35028
rect -33552 -35108 -28180 -35092
rect -33552 -35172 -28264 -35108
rect -28200 -35172 -28180 -35108
rect -33552 -35188 -28180 -35172
rect -33552 -35252 -28264 -35188
rect -28200 -35252 -28180 -35188
rect -33552 -35268 -28180 -35252
rect -33552 -35332 -28264 -35268
rect -28200 -35332 -28180 -35268
rect -33552 -35348 -28180 -35332
rect -33552 -35412 -28264 -35348
rect -28200 -35412 -28180 -35348
rect -33552 -35428 -28180 -35412
rect -33552 -35492 -28264 -35428
rect -28200 -35492 -28180 -35428
rect -33552 -35508 -28180 -35492
rect -33552 -35572 -28264 -35508
rect -28200 -35572 -28180 -35508
rect -33552 -35588 -28180 -35572
rect -33552 -35652 -28264 -35588
rect -28200 -35652 -28180 -35588
rect -33552 -35668 -28180 -35652
rect -33552 -35732 -28264 -35668
rect -28200 -35732 -28180 -35668
rect -33552 -35748 -28180 -35732
rect -33552 -35812 -28264 -35748
rect -28200 -35812 -28180 -35748
rect -33552 -35828 -28180 -35812
rect -33552 -35892 -28264 -35828
rect -28200 -35892 -28180 -35828
rect -33552 -35908 -28180 -35892
rect -33552 -35972 -28264 -35908
rect -28200 -35972 -28180 -35908
rect -33552 -35988 -28180 -35972
rect -33552 -36052 -28264 -35988
rect -28200 -36052 -28180 -35988
rect -33552 -36068 -28180 -36052
rect -33552 -36132 -28264 -36068
rect -28200 -36132 -28180 -36068
rect -33552 -36148 -28180 -36132
rect -33552 -36212 -28264 -36148
rect -28200 -36212 -28180 -36148
rect -33552 -36228 -28180 -36212
rect -33552 -36292 -28264 -36228
rect -28200 -36292 -28180 -36228
rect -33552 -36308 -28180 -36292
rect -33552 -36372 -28264 -36308
rect -28200 -36372 -28180 -36308
rect -33552 -36388 -28180 -36372
rect -33552 -36452 -28264 -36388
rect -28200 -36452 -28180 -36388
rect -33552 -36468 -28180 -36452
rect -33552 -36532 -28264 -36468
rect -28200 -36532 -28180 -36468
rect -33552 -36548 -28180 -36532
rect -33552 -36612 -28264 -36548
rect -28200 -36612 -28180 -36548
rect -33552 -36628 -28180 -36612
rect -33552 -36692 -28264 -36628
rect -28200 -36692 -28180 -36628
rect -33552 -36708 -28180 -36692
rect -33552 -36772 -28264 -36708
rect -28200 -36772 -28180 -36708
rect -33552 -36788 -28180 -36772
rect -33552 -36852 -28264 -36788
rect -28200 -36852 -28180 -36788
rect -33552 -36868 -28180 -36852
rect -33552 -36932 -28264 -36868
rect -28200 -36932 -28180 -36868
rect -33552 -36948 -28180 -36932
rect -33552 -37012 -28264 -36948
rect -28200 -37012 -28180 -36948
rect -33552 -37028 -28180 -37012
rect -33552 -37092 -28264 -37028
rect -28200 -37092 -28180 -37028
rect -33552 -37120 -28180 -37092
rect -27940 -32068 -22568 -32040
rect -27940 -32132 -22652 -32068
rect -22588 -32132 -22568 -32068
rect -27940 -32148 -22568 -32132
rect -27940 -32212 -22652 -32148
rect -22588 -32212 -22568 -32148
rect -27940 -32228 -22568 -32212
rect -27940 -32292 -22652 -32228
rect -22588 -32292 -22568 -32228
rect -27940 -32308 -22568 -32292
rect -27940 -32372 -22652 -32308
rect -22588 -32372 -22568 -32308
rect -27940 -32388 -22568 -32372
rect -27940 -32452 -22652 -32388
rect -22588 -32452 -22568 -32388
rect -27940 -32468 -22568 -32452
rect -27940 -32532 -22652 -32468
rect -22588 -32532 -22568 -32468
rect -27940 -32548 -22568 -32532
rect -27940 -32612 -22652 -32548
rect -22588 -32612 -22568 -32548
rect -27940 -32628 -22568 -32612
rect -27940 -32692 -22652 -32628
rect -22588 -32692 -22568 -32628
rect -27940 -32708 -22568 -32692
rect -27940 -32772 -22652 -32708
rect -22588 -32772 -22568 -32708
rect -27940 -32788 -22568 -32772
rect -27940 -32852 -22652 -32788
rect -22588 -32852 -22568 -32788
rect -27940 -32868 -22568 -32852
rect -27940 -32932 -22652 -32868
rect -22588 -32932 -22568 -32868
rect -27940 -32948 -22568 -32932
rect -27940 -33012 -22652 -32948
rect -22588 -33012 -22568 -32948
rect -27940 -33028 -22568 -33012
rect -27940 -33092 -22652 -33028
rect -22588 -33092 -22568 -33028
rect -27940 -33108 -22568 -33092
rect -27940 -33172 -22652 -33108
rect -22588 -33172 -22568 -33108
rect -27940 -33188 -22568 -33172
rect -27940 -33252 -22652 -33188
rect -22588 -33252 -22568 -33188
rect -27940 -33268 -22568 -33252
rect -27940 -33332 -22652 -33268
rect -22588 -33332 -22568 -33268
rect -27940 -33348 -22568 -33332
rect -27940 -33412 -22652 -33348
rect -22588 -33412 -22568 -33348
rect -27940 -33428 -22568 -33412
rect -27940 -33492 -22652 -33428
rect -22588 -33492 -22568 -33428
rect -27940 -33508 -22568 -33492
rect -27940 -33572 -22652 -33508
rect -22588 -33572 -22568 -33508
rect -27940 -33588 -22568 -33572
rect -27940 -33652 -22652 -33588
rect -22588 -33652 -22568 -33588
rect -27940 -33668 -22568 -33652
rect -27940 -33732 -22652 -33668
rect -22588 -33732 -22568 -33668
rect -27940 -33748 -22568 -33732
rect -27940 -33812 -22652 -33748
rect -22588 -33812 -22568 -33748
rect -27940 -33828 -22568 -33812
rect -27940 -33892 -22652 -33828
rect -22588 -33892 -22568 -33828
rect -27940 -33908 -22568 -33892
rect -27940 -33972 -22652 -33908
rect -22588 -33972 -22568 -33908
rect -27940 -33988 -22568 -33972
rect -27940 -34052 -22652 -33988
rect -22588 -34052 -22568 -33988
rect -27940 -34068 -22568 -34052
rect -27940 -34132 -22652 -34068
rect -22588 -34132 -22568 -34068
rect -27940 -34148 -22568 -34132
rect -27940 -34212 -22652 -34148
rect -22588 -34212 -22568 -34148
rect -27940 -34228 -22568 -34212
rect -27940 -34292 -22652 -34228
rect -22588 -34292 -22568 -34228
rect -27940 -34308 -22568 -34292
rect -27940 -34372 -22652 -34308
rect -22588 -34372 -22568 -34308
rect -27940 -34388 -22568 -34372
rect -27940 -34452 -22652 -34388
rect -22588 -34452 -22568 -34388
rect -27940 -34468 -22568 -34452
rect -27940 -34532 -22652 -34468
rect -22588 -34532 -22568 -34468
rect -27940 -34548 -22568 -34532
rect -27940 -34612 -22652 -34548
rect -22588 -34612 -22568 -34548
rect -27940 -34628 -22568 -34612
rect -27940 -34692 -22652 -34628
rect -22588 -34692 -22568 -34628
rect -27940 -34708 -22568 -34692
rect -27940 -34772 -22652 -34708
rect -22588 -34772 -22568 -34708
rect -27940 -34788 -22568 -34772
rect -27940 -34852 -22652 -34788
rect -22588 -34852 -22568 -34788
rect -27940 -34868 -22568 -34852
rect -27940 -34932 -22652 -34868
rect -22588 -34932 -22568 -34868
rect -27940 -34948 -22568 -34932
rect -27940 -35012 -22652 -34948
rect -22588 -35012 -22568 -34948
rect -27940 -35028 -22568 -35012
rect -27940 -35092 -22652 -35028
rect -22588 -35092 -22568 -35028
rect -27940 -35108 -22568 -35092
rect -27940 -35172 -22652 -35108
rect -22588 -35172 -22568 -35108
rect -27940 -35188 -22568 -35172
rect -27940 -35252 -22652 -35188
rect -22588 -35252 -22568 -35188
rect -27940 -35268 -22568 -35252
rect -27940 -35332 -22652 -35268
rect -22588 -35332 -22568 -35268
rect -27940 -35348 -22568 -35332
rect -27940 -35412 -22652 -35348
rect -22588 -35412 -22568 -35348
rect -27940 -35428 -22568 -35412
rect -27940 -35492 -22652 -35428
rect -22588 -35492 -22568 -35428
rect -27940 -35508 -22568 -35492
rect -27940 -35572 -22652 -35508
rect -22588 -35572 -22568 -35508
rect -27940 -35588 -22568 -35572
rect -27940 -35652 -22652 -35588
rect -22588 -35652 -22568 -35588
rect -27940 -35668 -22568 -35652
rect -27940 -35732 -22652 -35668
rect -22588 -35732 -22568 -35668
rect -27940 -35748 -22568 -35732
rect -27940 -35812 -22652 -35748
rect -22588 -35812 -22568 -35748
rect -27940 -35828 -22568 -35812
rect -27940 -35892 -22652 -35828
rect -22588 -35892 -22568 -35828
rect -27940 -35908 -22568 -35892
rect -27940 -35972 -22652 -35908
rect -22588 -35972 -22568 -35908
rect -27940 -35988 -22568 -35972
rect -27940 -36052 -22652 -35988
rect -22588 -36052 -22568 -35988
rect -27940 -36068 -22568 -36052
rect -27940 -36132 -22652 -36068
rect -22588 -36132 -22568 -36068
rect -27940 -36148 -22568 -36132
rect -27940 -36212 -22652 -36148
rect -22588 -36212 -22568 -36148
rect -27940 -36228 -22568 -36212
rect -27940 -36292 -22652 -36228
rect -22588 -36292 -22568 -36228
rect -27940 -36308 -22568 -36292
rect -27940 -36372 -22652 -36308
rect -22588 -36372 -22568 -36308
rect -27940 -36388 -22568 -36372
rect -27940 -36452 -22652 -36388
rect -22588 -36452 -22568 -36388
rect -27940 -36468 -22568 -36452
rect -27940 -36532 -22652 -36468
rect -22588 -36532 -22568 -36468
rect -27940 -36548 -22568 -36532
rect -27940 -36612 -22652 -36548
rect -22588 -36612 -22568 -36548
rect -27940 -36628 -22568 -36612
rect -27940 -36692 -22652 -36628
rect -22588 -36692 -22568 -36628
rect -27940 -36708 -22568 -36692
rect -27940 -36772 -22652 -36708
rect -22588 -36772 -22568 -36708
rect -27940 -36788 -22568 -36772
rect -27940 -36852 -22652 -36788
rect -22588 -36852 -22568 -36788
rect -27940 -36868 -22568 -36852
rect -27940 -36932 -22652 -36868
rect -22588 -36932 -22568 -36868
rect -27940 -36948 -22568 -36932
rect -27940 -37012 -22652 -36948
rect -22588 -37012 -22568 -36948
rect -27940 -37028 -22568 -37012
rect -27940 -37092 -22652 -37028
rect -22588 -37092 -22568 -37028
rect -27940 -37120 -22568 -37092
rect -22328 -32068 -16956 -32040
rect -22328 -32132 -17040 -32068
rect -16976 -32132 -16956 -32068
rect -22328 -32148 -16956 -32132
rect -22328 -32212 -17040 -32148
rect -16976 -32212 -16956 -32148
rect -22328 -32228 -16956 -32212
rect -22328 -32292 -17040 -32228
rect -16976 -32292 -16956 -32228
rect -22328 -32308 -16956 -32292
rect -22328 -32372 -17040 -32308
rect -16976 -32372 -16956 -32308
rect -22328 -32388 -16956 -32372
rect -22328 -32452 -17040 -32388
rect -16976 -32452 -16956 -32388
rect -22328 -32468 -16956 -32452
rect -22328 -32532 -17040 -32468
rect -16976 -32532 -16956 -32468
rect -22328 -32548 -16956 -32532
rect -22328 -32612 -17040 -32548
rect -16976 -32612 -16956 -32548
rect -22328 -32628 -16956 -32612
rect -22328 -32692 -17040 -32628
rect -16976 -32692 -16956 -32628
rect -22328 -32708 -16956 -32692
rect -22328 -32772 -17040 -32708
rect -16976 -32772 -16956 -32708
rect -22328 -32788 -16956 -32772
rect -22328 -32852 -17040 -32788
rect -16976 -32852 -16956 -32788
rect -22328 -32868 -16956 -32852
rect -22328 -32932 -17040 -32868
rect -16976 -32932 -16956 -32868
rect -22328 -32948 -16956 -32932
rect -22328 -33012 -17040 -32948
rect -16976 -33012 -16956 -32948
rect -22328 -33028 -16956 -33012
rect -22328 -33092 -17040 -33028
rect -16976 -33092 -16956 -33028
rect -22328 -33108 -16956 -33092
rect -22328 -33172 -17040 -33108
rect -16976 -33172 -16956 -33108
rect -22328 -33188 -16956 -33172
rect -22328 -33252 -17040 -33188
rect -16976 -33252 -16956 -33188
rect -22328 -33268 -16956 -33252
rect -22328 -33332 -17040 -33268
rect -16976 -33332 -16956 -33268
rect -22328 -33348 -16956 -33332
rect -22328 -33412 -17040 -33348
rect -16976 -33412 -16956 -33348
rect -22328 -33428 -16956 -33412
rect -22328 -33492 -17040 -33428
rect -16976 -33492 -16956 -33428
rect -22328 -33508 -16956 -33492
rect -22328 -33572 -17040 -33508
rect -16976 -33572 -16956 -33508
rect -22328 -33588 -16956 -33572
rect -22328 -33652 -17040 -33588
rect -16976 -33652 -16956 -33588
rect -22328 -33668 -16956 -33652
rect -22328 -33732 -17040 -33668
rect -16976 -33732 -16956 -33668
rect -22328 -33748 -16956 -33732
rect -22328 -33812 -17040 -33748
rect -16976 -33812 -16956 -33748
rect -22328 -33828 -16956 -33812
rect -22328 -33892 -17040 -33828
rect -16976 -33892 -16956 -33828
rect -22328 -33908 -16956 -33892
rect -22328 -33972 -17040 -33908
rect -16976 -33972 -16956 -33908
rect -22328 -33988 -16956 -33972
rect -22328 -34052 -17040 -33988
rect -16976 -34052 -16956 -33988
rect -22328 -34068 -16956 -34052
rect -22328 -34132 -17040 -34068
rect -16976 -34132 -16956 -34068
rect -22328 -34148 -16956 -34132
rect -22328 -34212 -17040 -34148
rect -16976 -34212 -16956 -34148
rect -22328 -34228 -16956 -34212
rect -22328 -34292 -17040 -34228
rect -16976 -34292 -16956 -34228
rect -22328 -34308 -16956 -34292
rect -22328 -34372 -17040 -34308
rect -16976 -34372 -16956 -34308
rect -22328 -34388 -16956 -34372
rect -22328 -34452 -17040 -34388
rect -16976 -34452 -16956 -34388
rect -22328 -34468 -16956 -34452
rect -22328 -34532 -17040 -34468
rect -16976 -34532 -16956 -34468
rect -22328 -34548 -16956 -34532
rect -22328 -34612 -17040 -34548
rect -16976 -34612 -16956 -34548
rect -22328 -34628 -16956 -34612
rect -22328 -34692 -17040 -34628
rect -16976 -34692 -16956 -34628
rect -22328 -34708 -16956 -34692
rect -22328 -34772 -17040 -34708
rect -16976 -34772 -16956 -34708
rect -22328 -34788 -16956 -34772
rect -22328 -34852 -17040 -34788
rect -16976 -34852 -16956 -34788
rect -22328 -34868 -16956 -34852
rect -22328 -34932 -17040 -34868
rect -16976 -34932 -16956 -34868
rect -22328 -34948 -16956 -34932
rect -22328 -35012 -17040 -34948
rect -16976 -35012 -16956 -34948
rect -22328 -35028 -16956 -35012
rect -22328 -35092 -17040 -35028
rect -16976 -35092 -16956 -35028
rect -22328 -35108 -16956 -35092
rect -22328 -35172 -17040 -35108
rect -16976 -35172 -16956 -35108
rect -22328 -35188 -16956 -35172
rect -22328 -35252 -17040 -35188
rect -16976 -35252 -16956 -35188
rect -22328 -35268 -16956 -35252
rect -22328 -35332 -17040 -35268
rect -16976 -35332 -16956 -35268
rect -22328 -35348 -16956 -35332
rect -22328 -35412 -17040 -35348
rect -16976 -35412 -16956 -35348
rect -22328 -35428 -16956 -35412
rect -22328 -35492 -17040 -35428
rect -16976 -35492 -16956 -35428
rect -22328 -35508 -16956 -35492
rect -22328 -35572 -17040 -35508
rect -16976 -35572 -16956 -35508
rect -22328 -35588 -16956 -35572
rect -22328 -35652 -17040 -35588
rect -16976 -35652 -16956 -35588
rect -22328 -35668 -16956 -35652
rect -22328 -35732 -17040 -35668
rect -16976 -35732 -16956 -35668
rect -22328 -35748 -16956 -35732
rect -22328 -35812 -17040 -35748
rect -16976 -35812 -16956 -35748
rect -22328 -35828 -16956 -35812
rect -22328 -35892 -17040 -35828
rect -16976 -35892 -16956 -35828
rect -22328 -35908 -16956 -35892
rect -22328 -35972 -17040 -35908
rect -16976 -35972 -16956 -35908
rect -22328 -35988 -16956 -35972
rect -22328 -36052 -17040 -35988
rect -16976 -36052 -16956 -35988
rect -22328 -36068 -16956 -36052
rect -22328 -36132 -17040 -36068
rect -16976 -36132 -16956 -36068
rect -22328 -36148 -16956 -36132
rect -22328 -36212 -17040 -36148
rect -16976 -36212 -16956 -36148
rect -22328 -36228 -16956 -36212
rect -22328 -36292 -17040 -36228
rect -16976 -36292 -16956 -36228
rect -22328 -36308 -16956 -36292
rect -22328 -36372 -17040 -36308
rect -16976 -36372 -16956 -36308
rect -22328 -36388 -16956 -36372
rect -22328 -36452 -17040 -36388
rect -16976 -36452 -16956 -36388
rect -22328 -36468 -16956 -36452
rect -22328 -36532 -17040 -36468
rect -16976 -36532 -16956 -36468
rect -22328 -36548 -16956 -36532
rect -22328 -36612 -17040 -36548
rect -16976 -36612 -16956 -36548
rect -22328 -36628 -16956 -36612
rect -22328 -36692 -17040 -36628
rect -16976 -36692 -16956 -36628
rect -22328 -36708 -16956 -36692
rect -22328 -36772 -17040 -36708
rect -16976 -36772 -16956 -36708
rect -22328 -36788 -16956 -36772
rect -22328 -36852 -17040 -36788
rect -16976 -36852 -16956 -36788
rect -22328 -36868 -16956 -36852
rect -22328 -36932 -17040 -36868
rect -16976 -36932 -16956 -36868
rect -22328 -36948 -16956 -36932
rect -22328 -37012 -17040 -36948
rect -16976 -37012 -16956 -36948
rect -22328 -37028 -16956 -37012
rect -22328 -37092 -17040 -37028
rect -16976 -37092 -16956 -37028
rect -22328 -37120 -16956 -37092
rect -16716 -32068 -11344 -32040
rect -16716 -32132 -11428 -32068
rect -11364 -32132 -11344 -32068
rect -16716 -32148 -11344 -32132
rect -16716 -32212 -11428 -32148
rect -11364 -32212 -11344 -32148
rect -16716 -32228 -11344 -32212
rect -16716 -32292 -11428 -32228
rect -11364 -32292 -11344 -32228
rect -16716 -32308 -11344 -32292
rect -16716 -32372 -11428 -32308
rect -11364 -32372 -11344 -32308
rect -16716 -32388 -11344 -32372
rect -16716 -32452 -11428 -32388
rect -11364 -32452 -11344 -32388
rect -16716 -32468 -11344 -32452
rect -16716 -32532 -11428 -32468
rect -11364 -32532 -11344 -32468
rect -16716 -32548 -11344 -32532
rect -16716 -32612 -11428 -32548
rect -11364 -32612 -11344 -32548
rect -16716 -32628 -11344 -32612
rect -16716 -32692 -11428 -32628
rect -11364 -32692 -11344 -32628
rect -16716 -32708 -11344 -32692
rect -16716 -32772 -11428 -32708
rect -11364 -32772 -11344 -32708
rect -16716 -32788 -11344 -32772
rect -16716 -32852 -11428 -32788
rect -11364 -32852 -11344 -32788
rect -16716 -32868 -11344 -32852
rect -16716 -32932 -11428 -32868
rect -11364 -32932 -11344 -32868
rect -16716 -32948 -11344 -32932
rect -16716 -33012 -11428 -32948
rect -11364 -33012 -11344 -32948
rect -16716 -33028 -11344 -33012
rect -16716 -33092 -11428 -33028
rect -11364 -33092 -11344 -33028
rect -16716 -33108 -11344 -33092
rect -16716 -33172 -11428 -33108
rect -11364 -33172 -11344 -33108
rect -16716 -33188 -11344 -33172
rect -16716 -33252 -11428 -33188
rect -11364 -33252 -11344 -33188
rect -16716 -33268 -11344 -33252
rect -16716 -33332 -11428 -33268
rect -11364 -33332 -11344 -33268
rect -16716 -33348 -11344 -33332
rect -16716 -33412 -11428 -33348
rect -11364 -33412 -11344 -33348
rect -16716 -33428 -11344 -33412
rect -16716 -33492 -11428 -33428
rect -11364 -33492 -11344 -33428
rect -16716 -33508 -11344 -33492
rect -16716 -33572 -11428 -33508
rect -11364 -33572 -11344 -33508
rect -16716 -33588 -11344 -33572
rect -16716 -33652 -11428 -33588
rect -11364 -33652 -11344 -33588
rect -16716 -33668 -11344 -33652
rect -16716 -33732 -11428 -33668
rect -11364 -33732 -11344 -33668
rect -16716 -33748 -11344 -33732
rect -16716 -33812 -11428 -33748
rect -11364 -33812 -11344 -33748
rect -16716 -33828 -11344 -33812
rect -16716 -33892 -11428 -33828
rect -11364 -33892 -11344 -33828
rect -16716 -33908 -11344 -33892
rect -16716 -33972 -11428 -33908
rect -11364 -33972 -11344 -33908
rect -16716 -33988 -11344 -33972
rect -16716 -34052 -11428 -33988
rect -11364 -34052 -11344 -33988
rect -16716 -34068 -11344 -34052
rect -16716 -34132 -11428 -34068
rect -11364 -34132 -11344 -34068
rect -16716 -34148 -11344 -34132
rect -16716 -34212 -11428 -34148
rect -11364 -34212 -11344 -34148
rect -16716 -34228 -11344 -34212
rect -16716 -34292 -11428 -34228
rect -11364 -34292 -11344 -34228
rect -16716 -34308 -11344 -34292
rect -16716 -34372 -11428 -34308
rect -11364 -34372 -11344 -34308
rect -16716 -34388 -11344 -34372
rect -16716 -34452 -11428 -34388
rect -11364 -34452 -11344 -34388
rect -16716 -34468 -11344 -34452
rect -16716 -34532 -11428 -34468
rect -11364 -34532 -11344 -34468
rect -16716 -34548 -11344 -34532
rect -16716 -34612 -11428 -34548
rect -11364 -34612 -11344 -34548
rect -16716 -34628 -11344 -34612
rect -16716 -34692 -11428 -34628
rect -11364 -34692 -11344 -34628
rect -16716 -34708 -11344 -34692
rect -16716 -34772 -11428 -34708
rect -11364 -34772 -11344 -34708
rect -16716 -34788 -11344 -34772
rect -16716 -34852 -11428 -34788
rect -11364 -34852 -11344 -34788
rect -16716 -34868 -11344 -34852
rect -16716 -34932 -11428 -34868
rect -11364 -34932 -11344 -34868
rect -16716 -34948 -11344 -34932
rect -16716 -35012 -11428 -34948
rect -11364 -35012 -11344 -34948
rect -16716 -35028 -11344 -35012
rect -16716 -35092 -11428 -35028
rect -11364 -35092 -11344 -35028
rect -16716 -35108 -11344 -35092
rect -16716 -35172 -11428 -35108
rect -11364 -35172 -11344 -35108
rect -16716 -35188 -11344 -35172
rect -16716 -35252 -11428 -35188
rect -11364 -35252 -11344 -35188
rect -16716 -35268 -11344 -35252
rect -16716 -35332 -11428 -35268
rect -11364 -35332 -11344 -35268
rect -16716 -35348 -11344 -35332
rect -16716 -35412 -11428 -35348
rect -11364 -35412 -11344 -35348
rect -16716 -35428 -11344 -35412
rect -16716 -35492 -11428 -35428
rect -11364 -35492 -11344 -35428
rect -16716 -35508 -11344 -35492
rect -16716 -35572 -11428 -35508
rect -11364 -35572 -11344 -35508
rect -16716 -35588 -11344 -35572
rect -16716 -35652 -11428 -35588
rect -11364 -35652 -11344 -35588
rect -16716 -35668 -11344 -35652
rect -16716 -35732 -11428 -35668
rect -11364 -35732 -11344 -35668
rect -16716 -35748 -11344 -35732
rect -16716 -35812 -11428 -35748
rect -11364 -35812 -11344 -35748
rect -16716 -35828 -11344 -35812
rect -16716 -35892 -11428 -35828
rect -11364 -35892 -11344 -35828
rect -16716 -35908 -11344 -35892
rect -16716 -35972 -11428 -35908
rect -11364 -35972 -11344 -35908
rect -16716 -35988 -11344 -35972
rect -16716 -36052 -11428 -35988
rect -11364 -36052 -11344 -35988
rect -16716 -36068 -11344 -36052
rect -16716 -36132 -11428 -36068
rect -11364 -36132 -11344 -36068
rect -16716 -36148 -11344 -36132
rect -16716 -36212 -11428 -36148
rect -11364 -36212 -11344 -36148
rect -16716 -36228 -11344 -36212
rect -16716 -36292 -11428 -36228
rect -11364 -36292 -11344 -36228
rect -16716 -36308 -11344 -36292
rect -16716 -36372 -11428 -36308
rect -11364 -36372 -11344 -36308
rect -16716 -36388 -11344 -36372
rect -16716 -36452 -11428 -36388
rect -11364 -36452 -11344 -36388
rect -16716 -36468 -11344 -36452
rect -16716 -36532 -11428 -36468
rect -11364 -36532 -11344 -36468
rect -16716 -36548 -11344 -36532
rect -16716 -36612 -11428 -36548
rect -11364 -36612 -11344 -36548
rect -16716 -36628 -11344 -36612
rect -16716 -36692 -11428 -36628
rect -11364 -36692 -11344 -36628
rect -16716 -36708 -11344 -36692
rect -16716 -36772 -11428 -36708
rect -11364 -36772 -11344 -36708
rect -16716 -36788 -11344 -36772
rect -16716 -36852 -11428 -36788
rect -11364 -36852 -11344 -36788
rect -16716 -36868 -11344 -36852
rect -16716 -36932 -11428 -36868
rect -11364 -36932 -11344 -36868
rect -16716 -36948 -11344 -36932
rect -16716 -37012 -11428 -36948
rect -11364 -37012 -11344 -36948
rect -16716 -37028 -11344 -37012
rect -16716 -37092 -11428 -37028
rect -11364 -37092 -11344 -37028
rect -16716 -37120 -11344 -37092
rect -11104 -32068 -5732 -32040
rect -11104 -32132 -5816 -32068
rect -5752 -32132 -5732 -32068
rect -11104 -32148 -5732 -32132
rect -11104 -32212 -5816 -32148
rect -5752 -32212 -5732 -32148
rect -11104 -32228 -5732 -32212
rect -11104 -32292 -5816 -32228
rect -5752 -32292 -5732 -32228
rect -11104 -32308 -5732 -32292
rect -11104 -32372 -5816 -32308
rect -5752 -32372 -5732 -32308
rect -11104 -32388 -5732 -32372
rect -11104 -32452 -5816 -32388
rect -5752 -32452 -5732 -32388
rect -11104 -32468 -5732 -32452
rect -11104 -32532 -5816 -32468
rect -5752 -32532 -5732 -32468
rect -11104 -32548 -5732 -32532
rect -11104 -32612 -5816 -32548
rect -5752 -32612 -5732 -32548
rect -11104 -32628 -5732 -32612
rect -11104 -32692 -5816 -32628
rect -5752 -32692 -5732 -32628
rect -11104 -32708 -5732 -32692
rect -11104 -32772 -5816 -32708
rect -5752 -32772 -5732 -32708
rect -11104 -32788 -5732 -32772
rect -11104 -32852 -5816 -32788
rect -5752 -32852 -5732 -32788
rect -11104 -32868 -5732 -32852
rect -11104 -32932 -5816 -32868
rect -5752 -32932 -5732 -32868
rect -11104 -32948 -5732 -32932
rect -11104 -33012 -5816 -32948
rect -5752 -33012 -5732 -32948
rect -11104 -33028 -5732 -33012
rect -11104 -33092 -5816 -33028
rect -5752 -33092 -5732 -33028
rect -11104 -33108 -5732 -33092
rect -11104 -33172 -5816 -33108
rect -5752 -33172 -5732 -33108
rect -11104 -33188 -5732 -33172
rect -11104 -33252 -5816 -33188
rect -5752 -33252 -5732 -33188
rect -11104 -33268 -5732 -33252
rect -11104 -33332 -5816 -33268
rect -5752 -33332 -5732 -33268
rect -11104 -33348 -5732 -33332
rect -11104 -33412 -5816 -33348
rect -5752 -33412 -5732 -33348
rect -11104 -33428 -5732 -33412
rect -11104 -33492 -5816 -33428
rect -5752 -33492 -5732 -33428
rect -11104 -33508 -5732 -33492
rect -11104 -33572 -5816 -33508
rect -5752 -33572 -5732 -33508
rect -11104 -33588 -5732 -33572
rect -11104 -33652 -5816 -33588
rect -5752 -33652 -5732 -33588
rect -11104 -33668 -5732 -33652
rect -11104 -33732 -5816 -33668
rect -5752 -33732 -5732 -33668
rect -11104 -33748 -5732 -33732
rect -11104 -33812 -5816 -33748
rect -5752 -33812 -5732 -33748
rect -11104 -33828 -5732 -33812
rect -11104 -33892 -5816 -33828
rect -5752 -33892 -5732 -33828
rect -11104 -33908 -5732 -33892
rect -11104 -33972 -5816 -33908
rect -5752 -33972 -5732 -33908
rect -11104 -33988 -5732 -33972
rect -11104 -34052 -5816 -33988
rect -5752 -34052 -5732 -33988
rect -11104 -34068 -5732 -34052
rect -11104 -34132 -5816 -34068
rect -5752 -34132 -5732 -34068
rect -11104 -34148 -5732 -34132
rect -11104 -34212 -5816 -34148
rect -5752 -34212 -5732 -34148
rect -11104 -34228 -5732 -34212
rect -11104 -34292 -5816 -34228
rect -5752 -34292 -5732 -34228
rect -11104 -34308 -5732 -34292
rect -11104 -34372 -5816 -34308
rect -5752 -34372 -5732 -34308
rect -11104 -34388 -5732 -34372
rect -11104 -34452 -5816 -34388
rect -5752 -34452 -5732 -34388
rect -11104 -34468 -5732 -34452
rect -11104 -34532 -5816 -34468
rect -5752 -34532 -5732 -34468
rect -11104 -34548 -5732 -34532
rect -11104 -34612 -5816 -34548
rect -5752 -34612 -5732 -34548
rect -11104 -34628 -5732 -34612
rect -11104 -34692 -5816 -34628
rect -5752 -34692 -5732 -34628
rect -11104 -34708 -5732 -34692
rect -11104 -34772 -5816 -34708
rect -5752 -34772 -5732 -34708
rect -11104 -34788 -5732 -34772
rect -11104 -34852 -5816 -34788
rect -5752 -34852 -5732 -34788
rect -11104 -34868 -5732 -34852
rect -11104 -34932 -5816 -34868
rect -5752 -34932 -5732 -34868
rect -11104 -34948 -5732 -34932
rect -11104 -35012 -5816 -34948
rect -5752 -35012 -5732 -34948
rect -11104 -35028 -5732 -35012
rect -11104 -35092 -5816 -35028
rect -5752 -35092 -5732 -35028
rect -11104 -35108 -5732 -35092
rect -11104 -35172 -5816 -35108
rect -5752 -35172 -5732 -35108
rect -11104 -35188 -5732 -35172
rect -11104 -35252 -5816 -35188
rect -5752 -35252 -5732 -35188
rect -11104 -35268 -5732 -35252
rect -11104 -35332 -5816 -35268
rect -5752 -35332 -5732 -35268
rect -11104 -35348 -5732 -35332
rect -11104 -35412 -5816 -35348
rect -5752 -35412 -5732 -35348
rect -11104 -35428 -5732 -35412
rect -11104 -35492 -5816 -35428
rect -5752 -35492 -5732 -35428
rect -11104 -35508 -5732 -35492
rect -11104 -35572 -5816 -35508
rect -5752 -35572 -5732 -35508
rect -11104 -35588 -5732 -35572
rect -11104 -35652 -5816 -35588
rect -5752 -35652 -5732 -35588
rect -11104 -35668 -5732 -35652
rect -11104 -35732 -5816 -35668
rect -5752 -35732 -5732 -35668
rect -11104 -35748 -5732 -35732
rect -11104 -35812 -5816 -35748
rect -5752 -35812 -5732 -35748
rect -11104 -35828 -5732 -35812
rect -11104 -35892 -5816 -35828
rect -5752 -35892 -5732 -35828
rect -11104 -35908 -5732 -35892
rect -11104 -35972 -5816 -35908
rect -5752 -35972 -5732 -35908
rect -11104 -35988 -5732 -35972
rect -11104 -36052 -5816 -35988
rect -5752 -36052 -5732 -35988
rect -11104 -36068 -5732 -36052
rect -11104 -36132 -5816 -36068
rect -5752 -36132 -5732 -36068
rect -11104 -36148 -5732 -36132
rect -11104 -36212 -5816 -36148
rect -5752 -36212 -5732 -36148
rect -11104 -36228 -5732 -36212
rect -11104 -36292 -5816 -36228
rect -5752 -36292 -5732 -36228
rect -11104 -36308 -5732 -36292
rect -11104 -36372 -5816 -36308
rect -5752 -36372 -5732 -36308
rect -11104 -36388 -5732 -36372
rect -11104 -36452 -5816 -36388
rect -5752 -36452 -5732 -36388
rect -11104 -36468 -5732 -36452
rect -11104 -36532 -5816 -36468
rect -5752 -36532 -5732 -36468
rect -11104 -36548 -5732 -36532
rect -11104 -36612 -5816 -36548
rect -5752 -36612 -5732 -36548
rect -11104 -36628 -5732 -36612
rect -11104 -36692 -5816 -36628
rect -5752 -36692 -5732 -36628
rect -11104 -36708 -5732 -36692
rect -11104 -36772 -5816 -36708
rect -5752 -36772 -5732 -36708
rect -11104 -36788 -5732 -36772
rect -11104 -36852 -5816 -36788
rect -5752 -36852 -5732 -36788
rect -11104 -36868 -5732 -36852
rect -11104 -36932 -5816 -36868
rect -5752 -36932 -5732 -36868
rect -11104 -36948 -5732 -36932
rect -11104 -37012 -5816 -36948
rect -5752 -37012 -5732 -36948
rect -11104 -37028 -5732 -37012
rect -11104 -37092 -5816 -37028
rect -5752 -37092 -5732 -37028
rect -11104 -37120 -5732 -37092
rect -5492 -32068 -120 -32040
rect -5492 -32132 -204 -32068
rect -140 -32132 -120 -32068
rect -5492 -32148 -120 -32132
rect -5492 -32212 -204 -32148
rect -140 -32212 -120 -32148
rect -5492 -32228 -120 -32212
rect -5492 -32292 -204 -32228
rect -140 -32292 -120 -32228
rect -5492 -32308 -120 -32292
rect -5492 -32372 -204 -32308
rect -140 -32372 -120 -32308
rect -5492 -32388 -120 -32372
rect -5492 -32452 -204 -32388
rect -140 -32452 -120 -32388
rect -5492 -32468 -120 -32452
rect -5492 -32532 -204 -32468
rect -140 -32532 -120 -32468
rect -5492 -32548 -120 -32532
rect -5492 -32612 -204 -32548
rect -140 -32612 -120 -32548
rect -5492 -32628 -120 -32612
rect -5492 -32692 -204 -32628
rect -140 -32692 -120 -32628
rect -5492 -32708 -120 -32692
rect -5492 -32772 -204 -32708
rect -140 -32772 -120 -32708
rect -5492 -32788 -120 -32772
rect -5492 -32852 -204 -32788
rect -140 -32852 -120 -32788
rect -5492 -32868 -120 -32852
rect -5492 -32932 -204 -32868
rect -140 -32932 -120 -32868
rect -5492 -32948 -120 -32932
rect -5492 -33012 -204 -32948
rect -140 -33012 -120 -32948
rect -5492 -33028 -120 -33012
rect -5492 -33092 -204 -33028
rect -140 -33092 -120 -33028
rect -5492 -33108 -120 -33092
rect -5492 -33172 -204 -33108
rect -140 -33172 -120 -33108
rect -5492 -33188 -120 -33172
rect -5492 -33252 -204 -33188
rect -140 -33252 -120 -33188
rect -5492 -33268 -120 -33252
rect -5492 -33332 -204 -33268
rect -140 -33332 -120 -33268
rect -5492 -33348 -120 -33332
rect -5492 -33412 -204 -33348
rect -140 -33412 -120 -33348
rect -5492 -33428 -120 -33412
rect -5492 -33492 -204 -33428
rect -140 -33492 -120 -33428
rect -5492 -33508 -120 -33492
rect -5492 -33572 -204 -33508
rect -140 -33572 -120 -33508
rect -5492 -33588 -120 -33572
rect -5492 -33652 -204 -33588
rect -140 -33652 -120 -33588
rect -5492 -33668 -120 -33652
rect -5492 -33732 -204 -33668
rect -140 -33732 -120 -33668
rect -5492 -33748 -120 -33732
rect -5492 -33812 -204 -33748
rect -140 -33812 -120 -33748
rect -5492 -33828 -120 -33812
rect -5492 -33892 -204 -33828
rect -140 -33892 -120 -33828
rect -5492 -33908 -120 -33892
rect -5492 -33972 -204 -33908
rect -140 -33972 -120 -33908
rect -5492 -33988 -120 -33972
rect -5492 -34052 -204 -33988
rect -140 -34052 -120 -33988
rect -5492 -34068 -120 -34052
rect -5492 -34132 -204 -34068
rect -140 -34132 -120 -34068
rect -5492 -34148 -120 -34132
rect -5492 -34212 -204 -34148
rect -140 -34212 -120 -34148
rect -5492 -34228 -120 -34212
rect -5492 -34292 -204 -34228
rect -140 -34292 -120 -34228
rect -5492 -34308 -120 -34292
rect -5492 -34372 -204 -34308
rect -140 -34372 -120 -34308
rect -5492 -34388 -120 -34372
rect -5492 -34452 -204 -34388
rect -140 -34452 -120 -34388
rect -5492 -34468 -120 -34452
rect -5492 -34532 -204 -34468
rect -140 -34532 -120 -34468
rect -5492 -34548 -120 -34532
rect -5492 -34612 -204 -34548
rect -140 -34612 -120 -34548
rect -5492 -34628 -120 -34612
rect -5492 -34692 -204 -34628
rect -140 -34692 -120 -34628
rect -5492 -34708 -120 -34692
rect -5492 -34772 -204 -34708
rect -140 -34772 -120 -34708
rect -5492 -34788 -120 -34772
rect -5492 -34852 -204 -34788
rect -140 -34852 -120 -34788
rect -5492 -34868 -120 -34852
rect -5492 -34932 -204 -34868
rect -140 -34932 -120 -34868
rect -5492 -34948 -120 -34932
rect -5492 -35012 -204 -34948
rect -140 -35012 -120 -34948
rect -5492 -35028 -120 -35012
rect -5492 -35092 -204 -35028
rect -140 -35092 -120 -35028
rect -5492 -35108 -120 -35092
rect -5492 -35172 -204 -35108
rect -140 -35172 -120 -35108
rect -5492 -35188 -120 -35172
rect -5492 -35252 -204 -35188
rect -140 -35252 -120 -35188
rect -5492 -35268 -120 -35252
rect -5492 -35332 -204 -35268
rect -140 -35332 -120 -35268
rect -5492 -35348 -120 -35332
rect -5492 -35412 -204 -35348
rect -140 -35412 -120 -35348
rect -5492 -35428 -120 -35412
rect -5492 -35492 -204 -35428
rect -140 -35492 -120 -35428
rect -5492 -35508 -120 -35492
rect -5492 -35572 -204 -35508
rect -140 -35572 -120 -35508
rect -5492 -35588 -120 -35572
rect -5492 -35652 -204 -35588
rect -140 -35652 -120 -35588
rect -5492 -35668 -120 -35652
rect -5492 -35732 -204 -35668
rect -140 -35732 -120 -35668
rect -5492 -35748 -120 -35732
rect -5492 -35812 -204 -35748
rect -140 -35812 -120 -35748
rect -5492 -35828 -120 -35812
rect -5492 -35892 -204 -35828
rect -140 -35892 -120 -35828
rect -5492 -35908 -120 -35892
rect -5492 -35972 -204 -35908
rect -140 -35972 -120 -35908
rect -5492 -35988 -120 -35972
rect -5492 -36052 -204 -35988
rect -140 -36052 -120 -35988
rect -5492 -36068 -120 -36052
rect -5492 -36132 -204 -36068
rect -140 -36132 -120 -36068
rect -5492 -36148 -120 -36132
rect -5492 -36212 -204 -36148
rect -140 -36212 -120 -36148
rect -5492 -36228 -120 -36212
rect -5492 -36292 -204 -36228
rect -140 -36292 -120 -36228
rect -5492 -36308 -120 -36292
rect -5492 -36372 -204 -36308
rect -140 -36372 -120 -36308
rect -5492 -36388 -120 -36372
rect -5492 -36452 -204 -36388
rect -140 -36452 -120 -36388
rect -5492 -36468 -120 -36452
rect -5492 -36532 -204 -36468
rect -140 -36532 -120 -36468
rect -5492 -36548 -120 -36532
rect -5492 -36612 -204 -36548
rect -140 -36612 -120 -36548
rect -5492 -36628 -120 -36612
rect -5492 -36692 -204 -36628
rect -140 -36692 -120 -36628
rect -5492 -36708 -120 -36692
rect -5492 -36772 -204 -36708
rect -140 -36772 -120 -36708
rect -5492 -36788 -120 -36772
rect -5492 -36852 -204 -36788
rect -140 -36852 -120 -36788
rect -5492 -36868 -120 -36852
rect -5492 -36932 -204 -36868
rect -140 -36932 -120 -36868
rect -5492 -36948 -120 -36932
rect -5492 -37012 -204 -36948
rect -140 -37012 -120 -36948
rect -5492 -37028 -120 -37012
rect -5492 -37092 -204 -37028
rect -140 -37092 -120 -37028
rect -5492 -37120 -120 -37092
rect 120 -32068 5492 -32040
rect 120 -32132 5408 -32068
rect 5472 -32132 5492 -32068
rect 120 -32148 5492 -32132
rect 120 -32212 5408 -32148
rect 5472 -32212 5492 -32148
rect 120 -32228 5492 -32212
rect 120 -32292 5408 -32228
rect 5472 -32292 5492 -32228
rect 120 -32308 5492 -32292
rect 120 -32372 5408 -32308
rect 5472 -32372 5492 -32308
rect 120 -32388 5492 -32372
rect 120 -32452 5408 -32388
rect 5472 -32452 5492 -32388
rect 120 -32468 5492 -32452
rect 120 -32532 5408 -32468
rect 5472 -32532 5492 -32468
rect 120 -32548 5492 -32532
rect 120 -32612 5408 -32548
rect 5472 -32612 5492 -32548
rect 120 -32628 5492 -32612
rect 120 -32692 5408 -32628
rect 5472 -32692 5492 -32628
rect 120 -32708 5492 -32692
rect 120 -32772 5408 -32708
rect 5472 -32772 5492 -32708
rect 120 -32788 5492 -32772
rect 120 -32852 5408 -32788
rect 5472 -32852 5492 -32788
rect 120 -32868 5492 -32852
rect 120 -32932 5408 -32868
rect 5472 -32932 5492 -32868
rect 120 -32948 5492 -32932
rect 120 -33012 5408 -32948
rect 5472 -33012 5492 -32948
rect 120 -33028 5492 -33012
rect 120 -33092 5408 -33028
rect 5472 -33092 5492 -33028
rect 120 -33108 5492 -33092
rect 120 -33172 5408 -33108
rect 5472 -33172 5492 -33108
rect 120 -33188 5492 -33172
rect 120 -33252 5408 -33188
rect 5472 -33252 5492 -33188
rect 120 -33268 5492 -33252
rect 120 -33332 5408 -33268
rect 5472 -33332 5492 -33268
rect 120 -33348 5492 -33332
rect 120 -33412 5408 -33348
rect 5472 -33412 5492 -33348
rect 120 -33428 5492 -33412
rect 120 -33492 5408 -33428
rect 5472 -33492 5492 -33428
rect 120 -33508 5492 -33492
rect 120 -33572 5408 -33508
rect 5472 -33572 5492 -33508
rect 120 -33588 5492 -33572
rect 120 -33652 5408 -33588
rect 5472 -33652 5492 -33588
rect 120 -33668 5492 -33652
rect 120 -33732 5408 -33668
rect 5472 -33732 5492 -33668
rect 120 -33748 5492 -33732
rect 120 -33812 5408 -33748
rect 5472 -33812 5492 -33748
rect 120 -33828 5492 -33812
rect 120 -33892 5408 -33828
rect 5472 -33892 5492 -33828
rect 120 -33908 5492 -33892
rect 120 -33972 5408 -33908
rect 5472 -33972 5492 -33908
rect 120 -33988 5492 -33972
rect 120 -34052 5408 -33988
rect 5472 -34052 5492 -33988
rect 120 -34068 5492 -34052
rect 120 -34132 5408 -34068
rect 5472 -34132 5492 -34068
rect 120 -34148 5492 -34132
rect 120 -34212 5408 -34148
rect 5472 -34212 5492 -34148
rect 120 -34228 5492 -34212
rect 120 -34292 5408 -34228
rect 5472 -34292 5492 -34228
rect 120 -34308 5492 -34292
rect 120 -34372 5408 -34308
rect 5472 -34372 5492 -34308
rect 120 -34388 5492 -34372
rect 120 -34452 5408 -34388
rect 5472 -34452 5492 -34388
rect 120 -34468 5492 -34452
rect 120 -34532 5408 -34468
rect 5472 -34532 5492 -34468
rect 120 -34548 5492 -34532
rect 120 -34612 5408 -34548
rect 5472 -34612 5492 -34548
rect 120 -34628 5492 -34612
rect 120 -34692 5408 -34628
rect 5472 -34692 5492 -34628
rect 120 -34708 5492 -34692
rect 120 -34772 5408 -34708
rect 5472 -34772 5492 -34708
rect 120 -34788 5492 -34772
rect 120 -34852 5408 -34788
rect 5472 -34852 5492 -34788
rect 120 -34868 5492 -34852
rect 120 -34932 5408 -34868
rect 5472 -34932 5492 -34868
rect 120 -34948 5492 -34932
rect 120 -35012 5408 -34948
rect 5472 -35012 5492 -34948
rect 120 -35028 5492 -35012
rect 120 -35092 5408 -35028
rect 5472 -35092 5492 -35028
rect 120 -35108 5492 -35092
rect 120 -35172 5408 -35108
rect 5472 -35172 5492 -35108
rect 120 -35188 5492 -35172
rect 120 -35252 5408 -35188
rect 5472 -35252 5492 -35188
rect 120 -35268 5492 -35252
rect 120 -35332 5408 -35268
rect 5472 -35332 5492 -35268
rect 120 -35348 5492 -35332
rect 120 -35412 5408 -35348
rect 5472 -35412 5492 -35348
rect 120 -35428 5492 -35412
rect 120 -35492 5408 -35428
rect 5472 -35492 5492 -35428
rect 120 -35508 5492 -35492
rect 120 -35572 5408 -35508
rect 5472 -35572 5492 -35508
rect 120 -35588 5492 -35572
rect 120 -35652 5408 -35588
rect 5472 -35652 5492 -35588
rect 120 -35668 5492 -35652
rect 120 -35732 5408 -35668
rect 5472 -35732 5492 -35668
rect 120 -35748 5492 -35732
rect 120 -35812 5408 -35748
rect 5472 -35812 5492 -35748
rect 120 -35828 5492 -35812
rect 120 -35892 5408 -35828
rect 5472 -35892 5492 -35828
rect 120 -35908 5492 -35892
rect 120 -35972 5408 -35908
rect 5472 -35972 5492 -35908
rect 120 -35988 5492 -35972
rect 120 -36052 5408 -35988
rect 5472 -36052 5492 -35988
rect 120 -36068 5492 -36052
rect 120 -36132 5408 -36068
rect 5472 -36132 5492 -36068
rect 120 -36148 5492 -36132
rect 120 -36212 5408 -36148
rect 5472 -36212 5492 -36148
rect 120 -36228 5492 -36212
rect 120 -36292 5408 -36228
rect 5472 -36292 5492 -36228
rect 120 -36308 5492 -36292
rect 120 -36372 5408 -36308
rect 5472 -36372 5492 -36308
rect 120 -36388 5492 -36372
rect 120 -36452 5408 -36388
rect 5472 -36452 5492 -36388
rect 120 -36468 5492 -36452
rect 120 -36532 5408 -36468
rect 5472 -36532 5492 -36468
rect 120 -36548 5492 -36532
rect 120 -36612 5408 -36548
rect 5472 -36612 5492 -36548
rect 120 -36628 5492 -36612
rect 120 -36692 5408 -36628
rect 5472 -36692 5492 -36628
rect 120 -36708 5492 -36692
rect 120 -36772 5408 -36708
rect 5472 -36772 5492 -36708
rect 120 -36788 5492 -36772
rect 120 -36852 5408 -36788
rect 5472 -36852 5492 -36788
rect 120 -36868 5492 -36852
rect 120 -36932 5408 -36868
rect 5472 -36932 5492 -36868
rect 120 -36948 5492 -36932
rect 120 -37012 5408 -36948
rect 5472 -37012 5492 -36948
rect 120 -37028 5492 -37012
rect 120 -37092 5408 -37028
rect 5472 -37092 5492 -37028
rect 120 -37120 5492 -37092
rect 5732 -32068 11104 -32040
rect 5732 -32132 11020 -32068
rect 11084 -32132 11104 -32068
rect 5732 -32148 11104 -32132
rect 5732 -32212 11020 -32148
rect 11084 -32212 11104 -32148
rect 5732 -32228 11104 -32212
rect 5732 -32292 11020 -32228
rect 11084 -32292 11104 -32228
rect 5732 -32308 11104 -32292
rect 5732 -32372 11020 -32308
rect 11084 -32372 11104 -32308
rect 5732 -32388 11104 -32372
rect 5732 -32452 11020 -32388
rect 11084 -32452 11104 -32388
rect 5732 -32468 11104 -32452
rect 5732 -32532 11020 -32468
rect 11084 -32532 11104 -32468
rect 5732 -32548 11104 -32532
rect 5732 -32612 11020 -32548
rect 11084 -32612 11104 -32548
rect 5732 -32628 11104 -32612
rect 5732 -32692 11020 -32628
rect 11084 -32692 11104 -32628
rect 5732 -32708 11104 -32692
rect 5732 -32772 11020 -32708
rect 11084 -32772 11104 -32708
rect 5732 -32788 11104 -32772
rect 5732 -32852 11020 -32788
rect 11084 -32852 11104 -32788
rect 5732 -32868 11104 -32852
rect 5732 -32932 11020 -32868
rect 11084 -32932 11104 -32868
rect 5732 -32948 11104 -32932
rect 5732 -33012 11020 -32948
rect 11084 -33012 11104 -32948
rect 5732 -33028 11104 -33012
rect 5732 -33092 11020 -33028
rect 11084 -33092 11104 -33028
rect 5732 -33108 11104 -33092
rect 5732 -33172 11020 -33108
rect 11084 -33172 11104 -33108
rect 5732 -33188 11104 -33172
rect 5732 -33252 11020 -33188
rect 11084 -33252 11104 -33188
rect 5732 -33268 11104 -33252
rect 5732 -33332 11020 -33268
rect 11084 -33332 11104 -33268
rect 5732 -33348 11104 -33332
rect 5732 -33412 11020 -33348
rect 11084 -33412 11104 -33348
rect 5732 -33428 11104 -33412
rect 5732 -33492 11020 -33428
rect 11084 -33492 11104 -33428
rect 5732 -33508 11104 -33492
rect 5732 -33572 11020 -33508
rect 11084 -33572 11104 -33508
rect 5732 -33588 11104 -33572
rect 5732 -33652 11020 -33588
rect 11084 -33652 11104 -33588
rect 5732 -33668 11104 -33652
rect 5732 -33732 11020 -33668
rect 11084 -33732 11104 -33668
rect 5732 -33748 11104 -33732
rect 5732 -33812 11020 -33748
rect 11084 -33812 11104 -33748
rect 5732 -33828 11104 -33812
rect 5732 -33892 11020 -33828
rect 11084 -33892 11104 -33828
rect 5732 -33908 11104 -33892
rect 5732 -33972 11020 -33908
rect 11084 -33972 11104 -33908
rect 5732 -33988 11104 -33972
rect 5732 -34052 11020 -33988
rect 11084 -34052 11104 -33988
rect 5732 -34068 11104 -34052
rect 5732 -34132 11020 -34068
rect 11084 -34132 11104 -34068
rect 5732 -34148 11104 -34132
rect 5732 -34212 11020 -34148
rect 11084 -34212 11104 -34148
rect 5732 -34228 11104 -34212
rect 5732 -34292 11020 -34228
rect 11084 -34292 11104 -34228
rect 5732 -34308 11104 -34292
rect 5732 -34372 11020 -34308
rect 11084 -34372 11104 -34308
rect 5732 -34388 11104 -34372
rect 5732 -34452 11020 -34388
rect 11084 -34452 11104 -34388
rect 5732 -34468 11104 -34452
rect 5732 -34532 11020 -34468
rect 11084 -34532 11104 -34468
rect 5732 -34548 11104 -34532
rect 5732 -34612 11020 -34548
rect 11084 -34612 11104 -34548
rect 5732 -34628 11104 -34612
rect 5732 -34692 11020 -34628
rect 11084 -34692 11104 -34628
rect 5732 -34708 11104 -34692
rect 5732 -34772 11020 -34708
rect 11084 -34772 11104 -34708
rect 5732 -34788 11104 -34772
rect 5732 -34852 11020 -34788
rect 11084 -34852 11104 -34788
rect 5732 -34868 11104 -34852
rect 5732 -34932 11020 -34868
rect 11084 -34932 11104 -34868
rect 5732 -34948 11104 -34932
rect 5732 -35012 11020 -34948
rect 11084 -35012 11104 -34948
rect 5732 -35028 11104 -35012
rect 5732 -35092 11020 -35028
rect 11084 -35092 11104 -35028
rect 5732 -35108 11104 -35092
rect 5732 -35172 11020 -35108
rect 11084 -35172 11104 -35108
rect 5732 -35188 11104 -35172
rect 5732 -35252 11020 -35188
rect 11084 -35252 11104 -35188
rect 5732 -35268 11104 -35252
rect 5732 -35332 11020 -35268
rect 11084 -35332 11104 -35268
rect 5732 -35348 11104 -35332
rect 5732 -35412 11020 -35348
rect 11084 -35412 11104 -35348
rect 5732 -35428 11104 -35412
rect 5732 -35492 11020 -35428
rect 11084 -35492 11104 -35428
rect 5732 -35508 11104 -35492
rect 5732 -35572 11020 -35508
rect 11084 -35572 11104 -35508
rect 5732 -35588 11104 -35572
rect 5732 -35652 11020 -35588
rect 11084 -35652 11104 -35588
rect 5732 -35668 11104 -35652
rect 5732 -35732 11020 -35668
rect 11084 -35732 11104 -35668
rect 5732 -35748 11104 -35732
rect 5732 -35812 11020 -35748
rect 11084 -35812 11104 -35748
rect 5732 -35828 11104 -35812
rect 5732 -35892 11020 -35828
rect 11084 -35892 11104 -35828
rect 5732 -35908 11104 -35892
rect 5732 -35972 11020 -35908
rect 11084 -35972 11104 -35908
rect 5732 -35988 11104 -35972
rect 5732 -36052 11020 -35988
rect 11084 -36052 11104 -35988
rect 5732 -36068 11104 -36052
rect 5732 -36132 11020 -36068
rect 11084 -36132 11104 -36068
rect 5732 -36148 11104 -36132
rect 5732 -36212 11020 -36148
rect 11084 -36212 11104 -36148
rect 5732 -36228 11104 -36212
rect 5732 -36292 11020 -36228
rect 11084 -36292 11104 -36228
rect 5732 -36308 11104 -36292
rect 5732 -36372 11020 -36308
rect 11084 -36372 11104 -36308
rect 5732 -36388 11104 -36372
rect 5732 -36452 11020 -36388
rect 11084 -36452 11104 -36388
rect 5732 -36468 11104 -36452
rect 5732 -36532 11020 -36468
rect 11084 -36532 11104 -36468
rect 5732 -36548 11104 -36532
rect 5732 -36612 11020 -36548
rect 11084 -36612 11104 -36548
rect 5732 -36628 11104 -36612
rect 5732 -36692 11020 -36628
rect 11084 -36692 11104 -36628
rect 5732 -36708 11104 -36692
rect 5732 -36772 11020 -36708
rect 11084 -36772 11104 -36708
rect 5732 -36788 11104 -36772
rect 5732 -36852 11020 -36788
rect 11084 -36852 11104 -36788
rect 5732 -36868 11104 -36852
rect 5732 -36932 11020 -36868
rect 11084 -36932 11104 -36868
rect 5732 -36948 11104 -36932
rect 5732 -37012 11020 -36948
rect 11084 -37012 11104 -36948
rect 5732 -37028 11104 -37012
rect 5732 -37092 11020 -37028
rect 11084 -37092 11104 -37028
rect 5732 -37120 11104 -37092
rect 11344 -32068 16716 -32040
rect 11344 -32132 16632 -32068
rect 16696 -32132 16716 -32068
rect 11344 -32148 16716 -32132
rect 11344 -32212 16632 -32148
rect 16696 -32212 16716 -32148
rect 11344 -32228 16716 -32212
rect 11344 -32292 16632 -32228
rect 16696 -32292 16716 -32228
rect 11344 -32308 16716 -32292
rect 11344 -32372 16632 -32308
rect 16696 -32372 16716 -32308
rect 11344 -32388 16716 -32372
rect 11344 -32452 16632 -32388
rect 16696 -32452 16716 -32388
rect 11344 -32468 16716 -32452
rect 11344 -32532 16632 -32468
rect 16696 -32532 16716 -32468
rect 11344 -32548 16716 -32532
rect 11344 -32612 16632 -32548
rect 16696 -32612 16716 -32548
rect 11344 -32628 16716 -32612
rect 11344 -32692 16632 -32628
rect 16696 -32692 16716 -32628
rect 11344 -32708 16716 -32692
rect 11344 -32772 16632 -32708
rect 16696 -32772 16716 -32708
rect 11344 -32788 16716 -32772
rect 11344 -32852 16632 -32788
rect 16696 -32852 16716 -32788
rect 11344 -32868 16716 -32852
rect 11344 -32932 16632 -32868
rect 16696 -32932 16716 -32868
rect 11344 -32948 16716 -32932
rect 11344 -33012 16632 -32948
rect 16696 -33012 16716 -32948
rect 11344 -33028 16716 -33012
rect 11344 -33092 16632 -33028
rect 16696 -33092 16716 -33028
rect 11344 -33108 16716 -33092
rect 11344 -33172 16632 -33108
rect 16696 -33172 16716 -33108
rect 11344 -33188 16716 -33172
rect 11344 -33252 16632 -33188
rect 16696 -33252 16716 -33188
rect 11344 -33268 16716 -33252
rect 11344 -33332 16632 -33268
rect 16696 -33332 16716 -33268
rect 11344 -33348 16716 -33332
rect 11344 -33412 16632 -33348
rect 16696 -33412 16716 -33348
rect 11344 -33428 16716 -33412
rect 11344 -33492 16632 -33428
rect 16696 -33492 16716 -33428
rect 11344 -33508 16716 -33492
rect 11344 -33572 16632 -33508
rect 16696 -33572 16716 -33508
rect 11344 -33588 16716 -33572
rect 11344 -33652 16632 -33588
rect 16696 -33652 16716 -33588
rect 11344 -33668 16716 -33652
rect 11344 -33732 16632 -33668
rect 16696 -33732 16716 -33668
rect 11344 -33748 16716 -33732
rect 11344 -33812 16632 -33748
rect 16696 -33812 16716 -33748
rect 11344 -33828 16716 -33812
rect 11344 -33892 16632 -33828
rect 16696 -33892 16716 -33828
rect 11344 -33908 16716 -33892
rect 11344 -33972 16632 -33908
rect 16696 -33972 16716 -33908
rect 11344 -33988 16716 -33972
rect 11344 -34052 16632 -33988
rect 16696 -34052 16716 -33988
rect 11344 -34068 16716 -34052
rect 11344 -34132 16632 -34068
rect 16696 -34132 16716 -34068
rect 11344 -34148 16716 -34132
rect 11344 -34212 16632 -34148
rect 16696 -34212 16716 -34148
rect 11344 -34228 16716 -34212
rect 11344 -34292 16632 -34228
rect 16696 -34292 16716 -34228
rect 11344 -34308 16716 -34292
rect 11344 -34372 16632 -34308
rect 16696 -34372 16716 -34308
rect 11344 -34388 16716 -34372
rect 11344 -34452 16632 -34388
rect 16696 -34452 16716 -34388
rect 11344 -34468 16716 -34452
rect 11344 -34532 16632 -34468
rect 16696 -34532 16716 -34468
rect 11344 -34548 16716 -34532
rect 11344 -34612 16632 -34548
rect 16696 -34612 16716 -34548
rect 11344 -34628 16716 -34612
rect 11344 -34692 16632 -34628
rect 16696 -34692 16716 -34628
rect 11344 -34708 16716 -34692
rect 11344 -34772 16632 -34708
rect 16696 -34772 16716 -34708
rect 11344 -34788 16716 -34772
rect 11344 -34852 16632 -34788
rect 16696 -34852 16716 -34788
rect 11344 -34868 16716 -34852
rect 11344 -34932 16632 -34868
rect 16696 -34932 16716 -34868
rect 11344 -34948 16716 -34932
rect 11344 -35012 16632 -34948
rect 16696 -35012 16716 -34948
rect 11344 -35028 16716 -35012
rect 11344 -35092 16632 -35028
rect 16696 -35092 16716 -35028
rect 11344 -35108 16716 -35092
rect 11344 -35172 16632 -35108
rect 16696 -35172 16716 -35108
rect 11344 -35188 16716 -35172
rect 11344 -35252 16632 -35188
rect 16696 -35252 16716 -35188
rect 11344 -35268 16716 -35252
rect 11344 -35332 16632 -35268
rect 16696 -35332 16716 -35268
rect 11344 -35348 16716 -35332
rect 11344 -35412 16632 -35348
rect 16696 -35412 16716 -35348
rect 11344 -35428 16716 -35412
rect 11344 -35492 16632 -35428
rect 16696 -35492 16716 -35428
rect 11344 -35508 16716 -35492
rect 11344 -35572 16632 -35508
rect 16696 -35572 16716 -35508
rect 11344 -35588 16716 -35572
rect 11344 -35652 16632 -35588
rect 16696 -35652 16716 -35588
rect 11344 -35668 16716 -35652
rect 11344 -35732 16632 -35668
rect 16696 -35732 16716 -35668
rect 11344 -35748 16716 -35732
rect 11344 -35812 16632 -35748
rect 16696 -35812 16716 -35748
rect 11344 -35828 16716 -35812
rect 11344 -35892 16632 -35828
rect 16696 -35892 16716 -35828
rect 11344 -35908 16716 -35892
rect 11344 -35972 16632 -35908
rect 16696 -35972 16716 -35908
rect 11344 -35988 16716 -35972
rect 11344 -36052 16632 -35988
rect 16696 -36052 16716 -35988
rect 11344 -36068 16716 -36052
rect 11344 -36132 16632 -36068
rect 16696 -36132 16716 -36068
rect 11344 -36148 16716 -36132
rect 11344 -36212 16632 -36148
rect 16696 -36212 16716 -36148
rect 11344 -36228 16716 -36212
rect 11344 -36292 16632 -36228
rect 16696 -36292 16716 -36228
rect 11344 -36308 16716 -36292
rect 11344 -36372 16632 -36308
rect 16696 -36372 16716 -36308
rect 11344 -36388 16716 -36372
rect 11344 -36452 16632 -36388
rect 16696 -36452 16716 -36388
rect 11344 -36468 16716 -36452
rect 11344 -36532 16632 -36468
rect 16696 -36532 16716 -36468
rect 11344 -36548 16716 -36532
rect 11344 -36612 16632 -36548
rect 16696 -36612 16716 -36548
rect 11344 -36628 16716 -36612
rect 11344 -36692 16632 -36628
rect 16696 -36692 16716 -36628
rect 11344 -36708 16716 -36692
rect 11344 -36772 16632 -36708
rect 16696 -36772 16716 -36708
rect 11344 -36788 16716 -36772
rect 11344 -36852 16632 -36788
rect 16696 -36852 16716 -36788
rect 11344 -36868 16716 -36852
rect 11344 -36932 16632 -36868
rect 16696 -36932 16716 -36868
rect 11344 -36948 16716 -36932
rect 11344 -37012 16632 -36948
rect 16696 -37012 16716 -36948
rect 11344 -37028 16716 -37012
rect 11344 -37092 16632 -37028
rect 16696 -37092 16716 -37028
rect 11344 -37120 16716 -37092
rect 16956 -32068 22328 -32040
rect 16956 -32132 22244 -32068
rect 22308 -32132 22328 -32068
rect 16956 -32148 22328 -32132
rect 16956 -32212 22244 -32148
rect 22308 -32212 22328 -32148
rect 16956 -32228 22328 -32212
rect 16956 -32292 22244 -32228
rect 22308 -32292 22328 -32228
rect 16956 -32308 22328 -32292
rect 16956 -32372 22244 -32308
rect 22308 -32372 22328 -32308
rect 16956 -32388 22328 -32372
rect 16956 -32452 22244 -32388
rect 22308 -32452 22328 -32388
rect 16956 -32468 22328 -32452
rect 16956 -32532 22244 -32468
rect 22308 -32532 22328 -32468
rect 16956 -32548 22328 -32532
rect 16956 -32612 22244 -32548
rect 22308 -32612 22328 -32548
rect 16956 -32628 22328 -32612
rect 16956 -32692 22244 -32628
rect 22308 -32692 22328 -32628
rect 16956 -32708 22328 -32692
rect 16956 -32772 22244 -32708
rect 22308 -32772 22328 -32708
rect 16956 -32788 22328 -32772
rect 16956 -32852 22244 -32788
rect 22308 -32852 22328 -32788
rect 16956 -32868 22328 -32852
rect 16956 -32932 22244 -32868
rect 22308 -32932 22328 -32868
rect 16956 -32948 22328 -32932
rect 16956 -33012 22244 -32948
rect 22308 -33012 22328 -32948
rect 16956 -33028 22328 -33012
rect 16956 -33092 22244 -33028
rect 22308 -33092 22328 -33028
rect 16956 -33108 22328 -33092
rect 16956 -33172 22244 -33108
rect 22308 -33172 22328 -33108
rect 16956 -33188 22328 -33172
rect 16956 -33252 22244 -33188
rect 22308 -33252 22328 -33188
rect 16956 -33268 22328 -33252
rect 16956 -33332 22244 -33268
rect 22308 -33332 22328 -33268
rect 16956 -33348 22328 -33332
rect 16956 -33412 22244 -33348
rect 22308 -33412 22328 -33348
rect 16956 -33428 22328 -33412
rect 16956 -33492 22244 -33428
rect 22308 -33492 22328 -33428
rect 16956 -33508 22328 -33492
rect 16956 -33572 22244 -33508
rect 22308 -33572 22328 -33508
rect 16956 -33588 22328 -33572
rect 16956 -33652 22244 -33588
rect 22308 -33652 22328 -33588
rect 16956 -33668 22328 -33652
rect 16956 -33732 22244 -33668
rect 22308 -33732 22328 -33668
rect 16956 -33748 22328 -33732
rect 16956 -33812 22244 -33748
rect 22308 -33812 22328 -33748
rect 16956 -33828 22328 -33812
rect 16956 -33892 22244 -33828
rect 22308 -33892 22328 -33828
rect 16956 -33908 22328 -33892
rect 16956 -33972 22244 -33908
rect 22308 -33972 22328 -33908
rect 16956 -33988 22328 -33972
rect 16956 -34052 22244 -33988
rect 22308 -34052 22328 -33988
rect 16956 -34068 22328 -34052
rect 16956 -34132 22244 -34068
rect 22308 -34132 22328 -34068
rect 16956 -34148 22328 -34132
rect 16956 -34212 22244 -34148
rect 22308 -34212 22328 -34148
rect 16956 -34228 22328 -34212
rect 16956 -34292 22244 -34228
rect 22308 -34292 22328 -34228
rect 16956 -34308 22328 -34292
rect 16956 -34372 22244 -34308
rect 22308 -34372 22328 -34308
rect 16956 -34388 22328 -34372
rect 16956 -34452 22244 -34388
rect 22308 -34452 22328 -34388
rect 16956 -34468 22328 -34452
rect 16956 -34532 22244 -34468
rect 22308 -34532 22328 -34468
rect 16956 -34548 22328 -34532
rect 16956 -34612 22244 -34548
rect 22308 -34612 22328 -34548
rect 16956 -34628 22328 -34612
rect 16956 -34692 22244 -34628
rect 22308 -34692 22328 -34628
rect 16956 -34708 22328 -34692
rect 16956 -34772 22244 -34708
rect 22308 -34772 22328 -34708
rect 16956 -34788 22328 -34772
rect 16956 -34852 22244 -34788
rect 22308 -34852 22328 -34788
rect 16956 -34868 22328 -34852
rect 16956 -34932 22244 -34868
rect 22308 -34932 22328 -34868
rect 16956 -34948 22328 -34932
rect 16956 -35012 22244 -34948
rect 22308 -35012 22328 -34948
rect 16956 -35028 22328 -35012
rect 16956 -35092 22244 -35028
rect 22308 -35092 22328 -35028
rect 16956 -35108 22328 -35092
rect 16956 -35172 22244 -35108
rect 22308 -35172 22328 -35108
rect 16956 -35188 22328 -35172
rect 16956 -35252 22244 -35188
rect 22308 -35252 22328 -35188
rect 16956 -35268 22328 -35252
rect 16956 -35332 22244 -35268
rect 22308 -35332 22328 -35268
rect 16956 -35348 22328 -35332
rect 16956 -35412 22244 -35348
rect 22308 -35412 22328 -35348
rect 16956 -35428 22328 -35412
rect 16956 -35492 22244 -35428
rect 22308 -35492 22328 -35428
rect 16956 -35508 22328 -35492
rect 16956 -35572 22244 -35508
rect 22308 -35572 22328 -35508
rect 16956 -35588 22328 -35572
rect 16956 -35652 22244 -35588
rect 22308 -35652 22328 -35588
rect 16956 -35668 22328 -35652
rect 16956 -35732 22244 -35668
rect 22308 -35732 22328 -35668
rect 16956 -35748 22328 -35732
rect 16956 -35812 22244 -35748
rect 22308 -35812 22328 -35748
rect 16956 -35828 22328 -35812
rect 16956 -35892 22244 -35828
rect 22308 -35892 22328 -35828
rect 16956 -35908 22328 -35892
rect 16956 -35972 22244 -35908
rect 22308 -35972 22328 -35908
rect 16956 -35988 22328 -35972
rect 16956 -36052 22244 -35988
rect 22308 -36052 22328 -35988
rect 16956 -36068 22328 -36052
rect 16956 -36132 22244 -36068
rect 22308 -36132 22328 -36068
rect 16956 -36148 22328 -36132
rect 16956 -36212 22244 -36148
rect 22308 -36212 22328 -36148
rect 16956 -36228 22328 -36212
rect 16956 -36292 22244 -36228
rect 22308 -36292 22328 -36228
rect 16956 -36308 22328 -36292
rect 16956 -36372 22244 -36308
rect 22308 -36372 22328 -36308
rect 16956 -36388 22328 -36372
rect 16956 -36452 22244 -36388
rect 22308 -36452 22328 -36388
rect 16956 -36468 22328 -36452
rect 16956 -36532 22244 -36468
rect 22308 -36532 22328 -36468
rect 16956 -36548 22328 -36532
rect 16956 -36612 22244 -36548
rect 22308 -36612 22328 -36548
rect 16956 -36628 22328 -36612
rect 16956 -36692 22244 -36628
rect 22308 -36692 22328 -36628
rect 16956 -36708 22328 -36692
rect 16956 -36772 22244 -36708
rect 22308 -36772 22328 -36708
rect 16956 -36788 22328 -36772
rect 16956 -36852 22244 -36788
rect 22308 -36852 22328 -36788
rect 16956 -36868 22328 -36852
rect 16956 -36932 22244 -36868
rect 22308 -36932 22328 -36868
rect 16956 -36948 22328 -36932
rect 16956 -37012 22244 -36948
rect 22308 -37012 22328 -36948
rect 16956 -37028 22328 -37012
rect 16956 -37092 22244 -37028
rect 22308 -37092 22328 -37028
rect 16956 -37120 22328 -37092
rect 22568 -32068 27940 -32040
rect 22568 -32132 27856 -32068
rect 27920 -32132 27940 -32068
rect 22568 -32148 27940 -32132
rect 22568 -32212 27856 -32148
rect 27920 -32212 27940 -32148
rect 22568 -32228 27940 -32212
rect 22568 -32292 27856 -32228
rect 27920 -32292 27940 -32228
rect 22568 -32308 27940 -32292
rect 22568 -32372 27856 -32308
rect 27920 -32372 27940 -32308
rect 22568 -32388 27940 -32372
rect 22568 -32452 27856 -32388
rect 27920 -32452 27940 -32388
rect 22568 -32468 27940 -32452
rect 22568 -32532 27856 -32468
rect 27920 -32532 27940 -32468
rect 22568 -32548 27940 -32532
rect 22568 -32612 27856 -32548
rect 27920 -32612 27940 -32548
rect 22568 -32628 27940 -32612
rect 22568 -32692 27856 -32628
rect 27920 -32692 27940 -32628
rect 22568 -32708 27940 -32692
rect 22568 -32772 27856 -32708
rect 27920 -32772 27940 -32708
rect 22568 -32788 27940 -32772
rect 22568 -32852 27856 -32788
rect 27920 -32852 27940 -32788
rect 22568 -32868 27940 -32852
rect 22568 -32932 27856 -32868
rect 27920 -32932 27940 -32868
rect 22568 -32948 27940 -32932
rect 22568 -33012 27856 -32948
rect 27920 -33012 27940 -32948
rect 22568 -33028 27940 -33012
rect 22568 -33092 27856 -33028
rect 27920 -33092 27940 -33028
rect 22568 -33108 27940 -33092
rect 22568 -33172 27856 -33108
rect 27920 -33172 27940 -33108
rect 22568 -33188 27940 -33172
rect 22568 -33252 27856 -33188
rect 27920 -33252 27940 -33188
rect 22568 -33268 27940 -33252
rect 22568 -33332 27856 -33268
rect 27920 -33332 27940 -33268
rect 22568 -33348 27940 -33332
rect 22568 -33412 27856 -33348
rect 27920 -33412 27940 -33348
rect 22568 -33428 27940 -33412
rect 22568 -33492 27856 -33428
rect 27920 -33492 27940 -33428
rect 22568 -33508 27940 -33492
rect 22568 -33572 27856 -33508
rect 27920 -33572 27940 -33508
rect 22568 -33588 27940 -33572
rect 22568 -33652 27856 -33588
rect 27920 -33652 27940 -33588
rect 22568 -33668 27940 -33652
rect 22568 -33732 27856 -33668
rect 27920 -33732 27940 -33668
rect 22568 -33748 27940 -33732
rect 22568 -33812 27856 -33748
rect 27920 -33812 27940 -33748
rect 22568 -33828 27940 -33812
rect 22568 -33892 27856 -33828
rect 27920 -33892 27940 -33828
rect 22568 -33908 27940 -33892
rect 22568 -33972 27856 -33908
rect 27920 -33972 27940 -33908
rect 22568 -33988 27940 -33972
rect 22568 -34052 27856 -33988
rect 27920 -34052 27940 -33988
rect 22568 -34068 27940 -34052
rect 22568 -34132 27856 -34068
rect 27920 -34132 27940 -34068
rect 22568 -34148 27940 -34132
rect 22568 -34212 27856 -34148
rect 27920 -34212 27940 -34148
rect 22568 -34228 27940 -34212
rect 22568 -34292 27856 -34228
rect 27920 -34292 27940 -34228
rect 22568 -34308 27940 -34292
rect 22568 -34372 27856 -34308
rect 27920 -34372 27940 -34308
rect 22568 -34388 27940 -34372
rect 22568 -34452 27856 -34388
rect 27920 -34452 27940 -34388
rect 22568 -34468 27940 -34452
rect 22568 -34532 27856 -34468
rect 27920 -34532 27940 -34468
rect 22568 -34548 27940 -34532
rect 22568 -34612 27856 -34548
rect 27920 -34612 27940 -34548
rect 22568 -34628 27940 -34612
rect 22568 -34692 27856 -34628
rect 27920 -34692 27940 -34628
rect 22568 -34708 27940 -34692
rect 22568 -34772 27856 -34708
rect 27920 -34772 27940 -34708
rect 22568 -34788 27940 -34772
rect 22568 -34852 27856 -34788
rect 27920 -34852 27940 -34788
rect 22568 -34868 27940 -34852
rect 22568 -34932 27856 -34868
rect 27920 -34932 27940 -34868
rect 22568 -34948 27940 -34932
rect 22568 -35012 27856 -34948
rect 27920 -35012 27940 -34948
rect 22568 -35028 27940 -35012
rect 22568 -35092 27856 -35028
rect 27920 -35092 27940 -35028
rect 22568 -35108 27940 -35092
rect 22568 -35172 27856 -35108
rect 27920 -35172 27940 -35108
rect 22568 -35188 27940 -35172
rect 22568 -35252 27856 -35188
rect 27920 -35252 27940 -35188
rect 22568 -35268 27940 -35252
rect 22568 -35332 27856 -35268
rect 27920 -35332 27940 -35268
rect 22568 -35348 27940 -35332
rect 22568 -35412 27856 -35348
rect 27920 -35412 27940 -35348
rect 22568 -35428 27940 -35412
rect 22568 -35492 27856 -35428
rect 27920 -35492 27940 -35428
rect 22568 -35508 27940 -35492
rect 22568 -35572 27856 -35508
rect 27920 -35572 27940 -35508
rect 22568 -35588 27940 -35572
rect 22568 -35652 27856 -35588
rect 27920 -35652 27940 -35588
rect 22568 -35668 27940 -35652
rect 22568 -35732 27856 -35668
rect 27920 -35732 27940 -35668
rect 22568 -35748 27940 -35732
rect 22568 -35812 27856 -35748
rect 27920 -35812 27940 -35748
rect 22568 -35828 27940 -35812
rect 22568 -35892 27856 -35828
rect 27920 -35892 27940 -35828
rect 22568 -35908 27940 -35892
rect 22568 -35972 27856 -35908
rect 27920 -35972 27940 -35908
rect 22568 -35988 27940 -35972
rect 22568 -36052 27856 -35988
rect 27920 -36052 27940 -35988
rect 22568 -36068 27940 -36052
rect 22568 -36132 27856 -36068
rect 27920 -36132 27940 -36068
rect 22568 -36148 27940 -36132
rect 22568 -36212 27856 -36148
rect 27920 -36212 27940 -36148
rect 22568 -36228 27940 -36212
rect 22568 -36292 27856 -36228
rect 27920 -36292 27940 -36228
rect 22568 -36308 27940 -36292
rect 22568 -36372 27856 -36308
rect 27920 -36372 27940 -36308
rect 22568 -36388 27940 -36372
rect 22568 -36452 27856 -36388
rect 27920 -36452 27940 -36388
rect 22568 -36468 27940 -36452
rect 22568 -36532 27856 -36468
rect 27920 -36532 27940 -36468
rect 22568 -36548 27940 -36532
rect 22568 -36612 27856 -36548
rect 27920 -36612 27940 -36548
rect 22568 -36628 27940 -36612
rect 22568 -36692 27856 -36628
rect 27920 -36692 27940 -36628
rect 22568 -36708 27940 -36692
rect 22568 -36772 27856 -36708
rect 27920 -36772 27940 -36708
rect 22568 -36788 27940 -36772
rect 22568 -36852 27856 -36788
rect 27920 -36852 27940 -36788
rect 22568 -36868 27940 -36852
rect 22568 -36932 27856 -36868
rect 27920 -36932 27940 -36868
rect 22568 -36948 27940 -36932
rect 22568 -37012 27856 -36948
rect 27920 -37012 27940 -36948
rect 22568 -37028 27940 -37012
rect 22568 -37092 27856 -37028
rect 27920 -37092 27940 -37028
rect 22568 -37120 27940 -37092
rect 28180 -32068 33552 -32040
rect 28180 -32132 33468 -32068
rect 33532 -32132 33552 -32068
rect 28180 -32148 33552 -32132
rect 28180 -32212 33468 -32148
rect 33532 -32212 33552 -32148
rect 28180 -32228 33552 -32212
rect 28180 -32292 33468 -32228
rect 33532 -32292 33552 -32228
rect 28180 -32308 33552 -32292
rect 28180 -32372 33468 -32308
rect 33532 -32372 33552 -32308
rect 28180 -32388 33552 -32372
rect 28180 -32452 33468 -32388
rect 33532 -32452 33552 -32388
rect 28180 -32468 33552 -32452
rect 28180 -32532 33468 -32468
rect 33532 -32532 33552 -32468
rect 28180 -32548 33552 -32532
rect 28180 -32612 33468 -32548
rect 33532 -32612 33552 -32548
rect 28180 -32628 33552 -32612
rect 28180 -32692 33468 -32628
rect 33532 -32692 33552 -32628
rect 28180 -32708 33552 -32692
rect 28180 -32772 33468 -32708
rect 33532 -32772 33552 -32708
rect 28180 -32788 33552 -32772
rect 28180 -32852 33468 -32788
rect 33532 -32852 33552 -32788
rect 28180 -32868 33552 -32852
rect 28180 -32932 33468 -32868
rect 33532 -32932 33552 -32868
rect 28180 -32948 33552 -32932
rect 28180 -33012 33468 -32948
rect 33532 -33012 33552 -32948
rect 28180 -33028 33552 -33012
rect 28180 -33092 33468 -33028
rect 33532 -33092 33552 -33028
rect 28180 -33108 33552 -33092
rect 28180 -33172 33468 -33108
rect 33532 -33172 33552 -33108
rect 28180 -33188 33552 -33172
rect 28180 -33252 33468 -33188
rect 33532 -33252 33552 -33188
rect 28180 -33268 33552 -33252
rect 28180 -33332 33468 -33268
rect 33532 -33332 33552 -33268
rect 28180 -33348 33552 -33332
rect 28180 -33412 33468 -33348
rect 33532 -33412 33552 -33348
rect 28180 -33428 33552 -33412
rect 28180 -33492 33468 -33428
rect 33532 -33492 33552 -33428
rect 28180 -33508 33552 -33492
rect 28180 -33572 33468 -33508
rect 33532 -33572 33552 -33508
rect 28180 -33588 33552 -33572
rect 28180 -33652 33468 -33588
rect 33532 -33652 33552 -33588
rect 28180 -33668 33552 -33652
rect 28180 -33732 33468 -33668
rect 33532 -33732 33552 -33668
rect 28180 -33748 33552 -33732
rect 28180 -33812 33468 -33748
rect 33532 -33812 33552 -33748
rect 28180 -33828 33552 -33812
rect 28180 -33892 33468 -33828
rect 33532 -33892 33552 -33828
rect 28180 -33908 33552 -33892
rect 28180 -33972 33468 -33908
rect 33532 -33972 33552 -33908
rect 28180 -33988 33552 -33972
rect 28180 -34052 33468 -33988
rect 33532 -34052 33552 -33988
rect 28180 -34068 33552 -34052
rect 28180 -34132 33468 -34068
rect 33532 -34132 33552 -34068
rect 28180 -34148 33552 -34132
rect 28180 -34212 33468 -34148
rect 33532 -34212 33552 -34148
rect 28180 -34228 33552 -34212
rect 28180 -34292 33468 -34228
rect 33532 -34292 33552 -34228
rect 28180 -34308 33552 -34292
rect 28180 -34372 33468 -34308
rect 33532 -34372 33552 -34308
rect 28180 -34388 33552 -34372
rect 28180 -34452 33468 -34388
rect 33532 -34452 33552 -34388
rect 28180 -34468 33552 -34452
rect 28180 -34532 33468 -34468
rect 33532 -34532 33552 -34468
rect 28180 -34548 33552 -34532
rect 28180 -34612 33468 -34548
rect 33532 -34612 33552 -34548
rect 28180 -34628 33552 -34612
rect 28180 -34692 33468 -34628
rect 33532 -34692 33552 -34628
rect 28180 -34708 33552 -34692
rect 28180 -34772 33468 -34708
rect 33532 -34772 33552 -34708
rect 28180 -34788 33552 -34772
rect 28180 -34852 33468 -34788
rect 33532 -34852 33552 -34788
rect 28180 -34868 33552 -34852
rect 28180 -34932 33468 -34868
rect 33532 -34932 33552 -34868
rect 28180 -34948 33552 -34932
rect 28180 -35012 33468 -34948
rect 33532 -35012 33552 -34948
rect 28180 -35028 33552 -35012
rect 28180 -35092 33468 -35028
rect 33532 -35092 33552 -35028
rect 28180 -35108 33552 -35092
rect 28180 -35172 33468 -35108
rect 33532 -35172 33552 -35108
rect 28180 -35188 33552 -35172
rect 28180 -35252 33468 -35188
rect 33532 -35252 33552 -35188
rect 28180 -35268 33552 -35252
rect 28180 -35332 33468 -35268
rect 33532 -35332 33552 -35268
rect 28180 -35348 33552 -35332
rect 28180 -35412 33468 -35348
rect 33532 -35412 33552 -35348
rect 28180 -35428 33552 -35412
rect 28180 -35492 33468 -35428
rect 33532 -35492 33552 -35428
rect 28180 -35508 33552 -35492
rect 28180 -35572 33468 -35508
rect 33532 -35572 33552 -35508
rect 28180 -35588 33552 -35572
rect 28180 -35652 33468 -35588
rect 33532 -35652 33552 -35588
rect 28180 -35668 33552 -35652
rect 28180 -35732 33468 -35668
rect 33532 -35732 33552 -35668
rect 28180 -35748 33552 -35732
rect 28180 -35812 33468 -35748
rect 33532 -35812 33552 -35748
rect 28180 -35828 33552 -35812
rect 28180 -35892 33468 -35828
rect 33532 -35892 33552 -35828
rect 28180 -35908 33552 -35892
rect 28180 -35972 33468 -35908
rect 33532 -35972 33552 -35908
rect 28180 -35988 33552 -35972
rect 28180 -36052 33468 -35988
rect 33532 -36052 33552 -35988
rect 28180 -36068 33552 -36052
rect 28180 -36132 33468 -36068
rect 33532 -36132 33552 -36068
rect 28180 -36148 33552 -36132
rect 28180 -36212 33468 -36148
rect 33532 -36212 33552 -36148
rect 28180 -36228 33552 -36212
rect 28180 -36292 33468 -36228
rect 33532 -36292 33552 -36228
rect 28180 -36308 33552 -36292
rect 28180 -36372 33468 -36308
rect 33532 -36372 33552 -36308
rect 28180 -36388 33552 -36372
rect 28180 -36452 33468 -36388
rect 33532 -36452 33552 -36388
rect 28180 -36468 33552 -36452
rect 28180 -36532 33468 -36468
rect 33532 -36532 33552 -36468
rect 28180 -36548 33552 -36532
rect 28180 -36612 33468 -36548
rect 33532 -36612 33552 -36548
rect 28180 -36628 33552 -36612
rect 28180 -36692 33468 -36628
rect 33532 -36692 33552 -36628
rect 28180 -36708 33552 -36692
rect 28180 -36772 33468 -36708
rect 33532 -36772 33552 -36708
rect 28180 -36788 33552 -36772
rect 28180 -36852 33468 -36788
rect 33532 -36852 33552 -36788
rect 28180 -36868 33552 -36852
rect 28180 -36932 33468 -36868
rect 33532 -36932 33552 -36868
rect 28180 -36948 33552 -36932
rect 28180 -37012 33468 -36948
rect 33532 -37012 33552 -36948
rect 28180 -37028 33552 -37012
rect 28180 -37092 33468 -37028
rect 33532 -37092 33552 -37028
rect 28180 -37120 33552 -37092
rect 33792 -32068 39164 -32040
rect 33792 -32132 39080 -32068
rect 39144 -32132 39164 -32068
rect 33792 -32148 39164 -32132
rect 33792 -32212 39080 -32148
rect 39144 -32212 39164 -32148
rect 33792 -32228 39164 -32212
rect 33792 -32292 39080 -32228
rect 39144 -32292 39164 -32228
rect 33792 -32308 39164 -32292
rect 33792 -32372 39080 -32308
rect 39144 -32372 39164 -32308
rect 33792 -32388 39164 -32372
rect 33792 -32452 39080 -32388
rect 39144 -32452 39164 -32388
rect 33792 -32468 39164 -32452
rect 33792 -32532 39080 -32468
rect 39144 -32532 39164 -32468
rect 33792 -32548 39164 -32532
rect 33792 -32612 39080 -32548
rect 39144 -32612 39164 -32548
rect 33792 -32628 39164 -32612
rect 33792 -32692 39080 -32628
rect 39144 -32692 39164 -32628
rect 33792 -32708 39164 -32692
rect 33792 -32772 39080 -32708
rect 39144 -32772 39164 -32708
rect 33792 -32788 39164 -32772
rect 33792 -32852 39080 -32788
rect 39144 -32852 39164 -32788
rect 33792 -32868 39164 -32852
rect 33792 -32932 39080 -32868
rect 39144 -32932 39164 -32868
rect 33792 -32948 39164 -32932
rect 33792 -33012 39080 -32948
rect 39144 -33012 39164 -32948
rect 33792 -33028 39164 -33012
rect 33792 -33092 39080 -33028
rect 39144 -33092 39164 -33028
rect 33792 -33108 39164 -33092
rect 33792 -33172 39080 -33108
rect 39144 -33172 39164 -33108
rect 33792 -33188 39164 -33172
rect 33792 -33252 39080 -33188
rect 39144 -33252 39164 -33188
rect 33792 -33268 39164 -33252
rect 33792 -33332 39080 -33268
rect 39144 -33332 39164 -33268
rect 33792 -33348 39164 -33332
rect 33792 -33412 39080 -33348
rect 39144 -33412 39164 -33348
rect 33792 -33428 39164 -33412
rect 33792 -33492 39080 -33428
rect 39144 -33492 39164 -33428
rect 33792 -33508 39164 -33492
rect 33792 -33572 39080 -33508
rect 39144 -33572 39164 -33508
rect 33792 -33588 39164 -33572
rect 33792 -33652 39080 -33588
rect 39144 -33652 39164 -33588
rect 33792 -33668 39164 -33652
rect 33792 -33732 39080 -33668
rect 39144 -33732 39164 -33668
rect 33792 -33748 39164 -33732
rect 33792 -33812 39080 -33748
rect 39144 -33812 39164 -33748
rect 33792 -33828 39164 -33812
rect 33792 -33892 39080 -33828
rect 39144 -33892 39164 -33828
rect 33792 -33908 39164 -33892
rect 33792 -33972 39080 -33908
rect 39144 -33972 39164 -33908
rect 33792 -33988 39164 -33972
rect 33792 -34052 39080 -33988
rect 39144 -34052 39164 -33988
rect 33792 -34068 39164 -34052
rect 33792 -34132 39080 -34068
rect 39144 -34132 39164 -34068
rect 33792 -34148 39164 -34132
rect 33792 -34212 39080 -34148
rect 39144 -34212 39164 -34148
rect 33792 -34228 39164 -34212
rect 33792 -34292 39080 -34228
rect 39144 -34292 39164 -34228
rect 33792 -34308 39164 -34292
rect 33792 -34372 39080 -34308
rect 39144 -34372 39164 -34308
rect 33792 -34388 39164 -34372
rect 33792 -34452 39080 -34388
rect 39144 -34452 39164 -34388
rect 33792 -34468 39164 -34452
rect 33792 -34532 39080 -34468
rect 39144 -34532 39164 -34468
rect 33792 -34548 39164 -34532
rect 33792 -34612 39080 -34548
rect 39144 -34612 39164 -34548
rect 33792 -34628 39164 -34612
rect 33792 -34692 39080 -34628
rect 39144 -34692 39164 -34628
rect 33792 -34708 39164 -34692
rect 33792 -34772 39080 -34708
rect 39144 -34772 39164 -34708
rect 33792 -34788 39164 -34772
rect 33792 -34852 39080 -34788
rect 39144 -34852 39164 -34788
rect 33792 -34868 39164 -34852
rect 33792 -34932 39080 -34868
rect 39144 -34932 39164 -34868
rect 33792 -34948 39164 -34932
rect 33792 -35012 39080 -34948
rect 39144 -35012 39164 -34948
rect 33792 -35028 39164 -35012
rect 33792 -35092 39080 -35028
rect 39144 -35092 39164 -35028
rect 33792 -35108 39164 -35092
rect 33792 -35172 39080 -35108
rect 39144 -35172 39164 -35108
rect 33792 -35188 39164 -35172
rect 33792 -35252 39080 -35188
rect 39144 -35252 39164 -35188
rect 33792 -35268 39164 -35252
rect 33792 -35332 39080 -35268
rect 39144 -35332 39164 -35268
rect 33792 -35348 39164 -35332
rect 33792 -35412 39080 -35348
rect 39144 -35412 39164 -35348
rect 33792 -35428 39164 -35412
rect 33792 -35492 39080 -35428
rect 39144 -35492 39164 -35428
rect 33792 -35508 39164 -35492
rect 33792 -35572 39080 -35508
rect 39144 -35572 39164 -35508
rect 33792 -35588 39164 -35572
rect 33792 -35652 39080 -35588
rect 39144 -35652 39164 -35588
rect 33792 -35668 39164 -35652
rect 33792 -35732 39080 -35668
rect 39144 -35732 39164 -35668
rect 33792 -35748 39164 -35732
rect 33792 -35812 39080 -35748
rect 39144 -35812 39164 -35748
rect 33792 -35828 39164 -35812
rect 33792 -35892 39080 -35828
rect 39144 -35892 39164 -35828
rect 33792 -35908 39164 -35892
rect 33792 -35972 39080 -35908
rect 39144 -35972 39164 -35908
rect 33792 -35988 39164 -35972
rect 33792 -36052 39080 -35988
rect 39144 -36052 39164 -35988
rect 33792 -36068 39164 -36052
rect 33792 -36132 39080 -36068
rect 39144 -36132 39164 -36068
rect 33792 -36148 39164 -36132
rect 33792 -36212 39080 -36148
rect 39144 -36212 39164 -36148
rect 33792 -36228 39164 -36212
rect 33792 -36292 39080 -36228
rect 39144 -36292 39164 -36228
rect 33792 -36308 39164 -36292
rect 33792 -36372 39080 -36308
rect 39144 -36372 39164 -36308
rect 33792 -36388 39164 -36372
rect 33792 -36452 39080 -36388
rect 39144 -36452 39164 -36388
rect 33792 -36468 39164 -36452
rect 33792 -36532 39080 -36468
rect 39144 -36532 39164 -36468
rect 33792 -36548 39164 -36532
rect 33792 -36612 39080 -36548
rect 39144 -36612 39164 -36548
rect 33792 -36628 39164 -36612
rect 33792 -36692 39080 -36628
rect 39144 -36692 39164 -36628
rect 33792 -36708 39164 -36692
rect 33792 -36772 39080 -36708
rect 39144 -36772 39164 -36708
rect 33792 -36788 39164 -36772
rect 33792 -36852 39080 -36788
rect 39144 -36852 39164 -36788
rect 33792 -36868 39164 -36852
rect 33792 -36932 39080 -36868
rect 39144 -36932 39164 -36868
rect 33792 -36948 39164 -36932
rect 33792 -37012 39080 -36948
rect 39144 -37012 39164 -36948
rect 33792 -37028 39164 -37012
rect 33792 -37092 39080 -37028
rect 39144 -37092 39164 -37028
rect 33792 -37120 39164 -37092
<< via3 >>
rect -33876 37028 -33812 37092
rect -33876 36948 -33812 37012
rect -33876 36868 -33812 36932
rect -33876 36788 -33812 36852
rect -33876 36708 -33812 36772
rect -33876 36628 -33812 36692
rect -33876 36548 -33812 36612
rect -33876 36468 -33812 36532
rect -33876 36388 -33812 36452
rect -33876 36308 -33812 36372
rect -33876 36228 -33812 36292
rect -33876 36148 -33812 36212
rect -33876 36068 -33812 36132
rect -33876 35988 -33812 36052
rect -33876 35908 -33812 35972
rect -33876 35828 -33812 35892
rect -33876 35748 -33812 35812
rect -33876 35668 -33812 35732
rect -33876 35588 -33812 35652
rect -33876 35508 -33812 35572
rect -33876 35428 -33812 35492
rect -33876 35348 -33812 35412
rect -33876 35268 -33812 35332
rect -33876 35188 -33812 35252
rect -33876 35108 -33812 35172
rect -33876 35028 -33812 35092
rect -33876 34948 -33812 35012
rect -33876 34868 -33812 34932
rect -33876 34788 -33812 34852
rect -33876 34708 -33812 34772
rect -33876 34628 -33812 34692
rect -33876 34548 -33812 34612
rect -33876 34468 -33812 34532
rect -33876 34388 -33812 34452
rect -33876 34308 -33812 34372
rect -33876 34228 -33812 34292
rect -33876 34148 -33812 34212
rect -33876 34068 -33812 34132
rect -33876 33988 -33812 34052
rect -33876 33908 -33812 33972
rect -33876 33828 -33812 33892
rect -33876 33748 -33812 33812
rect -33876 33668 -33812 33732
rect -33876 33588 -33812 33652
rect -33876 33508 -33812 33572
rect -33876 33428 -33812 33492
rect -33876 33348 -33812 33412
rect -33876 33268 -33812 33332
rect -33876 33188 -33812 33252
rect -33876 33108 -33812 33172
rect -33876 33028 -33812 33092
rect -33876 32948 -33812 33012
rect -33876 32868 -33812 32932
rect -33876 32788 -33812 32852
rect -33876 32708 -33812 32772
rect -33876 32628 -33812 32692
rect -33876 32548 -33812 32612
rect -33876 32468 -33812 32532
rect -33876 32388 -33812 32452
rect -33876 32308 -33812 32372
rect -33876 32228 -33812 32292
rect -33876 32148 -33812 32212
rect -33876 32068 -33812 32132
rect -28264 37028 -28200 37092
rect -28264 36948 -28200 37012
rect -28264 36868 -28200 36932
rect -28264 36788 -28200 36852
rect -28264 36708 -28200 36772
rect -28264 36628 -28200 36692
rect -28264 36548 -28200 36612
rect -28264 36468 -28200 36532
rect -28264 36388 -28200 36452
rect -28264 36308 -28200 36372
rect -28264 36228 -28200 36292
rect -28264 36148 -28200 36212
rect -28264 36068 -28200 36132
rect -28264 35988 -28200 36052
rect -28264 35908 -28200 35972
rect -28264 35828 -28200 35892
rect -28264 35748 -28200 35812
rect -28264 35668 -28200 35732
rect -28264 35588 -28200 35652
rect -28264 35508 -28200 35572
rect -28264 35428 -28200 35492
rect -28264 35348 -28200 35412
rect -28264 35268 -28200 35332
rect -28264 35188 -28200 35252
rect -28264 35108 -28200 35172
rect -28264 35028 -28200 35092
rect -28264 34948 -28200 35012
rect -28264 34868 -28200 34932
rect -28264 34788 -28200 34852
rect -28264 34708 -28200 34772
rect -28264 34628 -28200 34692
rect -28264 34548 -28200 34612
rect -28264 34468 -28200 34532
rect -28264 34388 -28200 34452
rect -28264 34308 -28200 34372
rect -28264 34228 -28200 34292
rect -28264 34148 -28200 34212
rect -28264 34068 -28200 34132
rect -28264 33988 -28200 34052
rect -28264 33908 -28200 33972
rect -28264 33828 -28200 33892
rect -28264 33748 -28200 33812
rect -28264 33668 -28200 33732
rect -28264 33588 -28200 33652
rect -28264 33508 -28200 33572
rect -28264 33428 -28200 33492
rect -28264 33348 -28200 33412
rect -28264 33268 -28200 33332
rect -28264 33188 -28200 33252
rect -28264 33108 -28200 33172
rect -28264 33028 -28200 33092
rect -28264 32948 -28200 33012
rect -28264 32868 -28200 32932
rect -28264 32788 -28200 32852
rect -28264 32708 -28200 32772
rect -28264 32628 -28200 32692
rect -28264 32548 -28200 32612
rect -28264 32468 -28200 32532
rect -28264 32388 -28200 32452
rect -28264 32308 -28200 32372
rect -28264 32228 -28200 32292
rect -28264 32148 -28200 32212
rect -28264 32068 -28200 32132
rect -22652 37028 -22588 37092
rect -22652 36948 -22588 37012
rect -22652 36868 -22588 36932
rect -22652 36788 -22588 36852
rect -22652 36708 -22588 36772
rect -22652 36628 -22588 36692
rect -22652 36548 -22588 36612
rect -22652 36468 -22588 36532
rect -22652 36388 -22588 36452
rect -22652 36308 -22588 36372
rect -22652 36228 -22588 36292
rect -22652 36148 -22588 36212
rect -22652 36068 -22588 36132
rect -22652 35988 -22588 36052
rect -22652 35908 -22588 35972
rect -22652 35828 -22588 35892
rect -22652 35748 -22588 35812
rect -22652 35668 -22588 35732
rect -22652 35588 -22588 35652
rect -22652 35508 -22588 35572
rect -22652 35428 -22588 35492
rect -22652 35348 -22588 35412
rect -22652 35268 -22588 35332
rect -22652 35188 -22588 35252
rect -22652 35108 -22588 35172
rect -22652 35028 -22588 35092
rect -22652 34948 -22588 35012
rect -22652 34868 -22588 34932
rect -22652 34788 -22588 34852
rect -22652 34708 -22588 34772
rect -22652 34628 -22588 34692
rect -22652 34548 -22588 34612
rect -22652 34468 -22588 34532
rect -22652 34388 -22588 34452
rect -22652 34308 -22588 34372
rect -22652 34228 -22588 34292
rect -22652 34148 -22588 34212
rect -22652 34068 -22588 34132
rect -22652 33988 -22588 34052
rect -22652 33908 -22588 33972
rect -22652 33828 -22588 33892
rect -22652 33748 -22588 33812
rect -22652 33668 -22588 33732
rect -22652 33588 -22588 33652
rect -22652 33508 -22588 33572
rect -22652 33428 -22588 33492
rect -22652 33348 -22588 33412
rect -22652 33268 -22588 33332
rect -22652 33188 -22588 33252
rect -22652 33108 -22588 33172
rect -22652 33028 -22588 33092
rect -22652 32948 -22588 33012
rect -22652 32868 -22588 32932
rect -22652 32788 -22588 32852
rect -22652 32708 -22588 32772
rect -22652 32628 -22588 32692
rect -22652 32548 -22588 32612
rect -22652 32468 -22588 32532
rect -22652 32388 -22588 32452
rect -22652 32308 -22588 32372
rect -22652 32228 -22588 32292
rect -22652 32148 -22588 32212
rect -22652 32068 -22588 32132
rect -17040 37028 -16976 37092
rect -17040 36948 -16976 37012
rect -17040 36868 -16976 36932
rect -17040 36788 -16976 36852
rect -17040 36708 -16976 36772
rect -17040 36628 -16976 36692
rect -17040 36548 -16976 36612
rect -17040 36468 -16976 36532
rect -17040 36388 -16976 36452
rect -17040 36308 -16976 36372
rect -17040 36228 -16976 36292
rect -17040 36148 -16976 36212
rect -17040 36068 -16976 36132
rect -17040 35988 -16976 36052
rect -17040 35908 -16976 35972
rect -17040 35828 -16976 35892
rect -17040 35748 -16976 35812
rect -17040 35668 -16976 35732
rect -17040 35588 -16976 35652
rect -17040 35508 -16976 35572
rect -17040 35428 -16976 35492
rect -17040 35348 -16976 35412
rect -17040 35268 -16976 35332
rect -17040 35188 -16976 35252
rect -17040 35108 -16976 35172
rect -17040 35028 -16976 35092
rect -17040 34948 -16976 35012
rect -17040 34868 -16976 34932
rect -17040 34788 -16976 34852
rect -17040 34708 -16976 34772
rect -17040 34628 -16976 34692
rect -17040 34548 -16976 34612
rect -17040 34468 -16976 34532
rect -17040 34388 -16976 34452
rect -17040 34308 -16976 34372
rect -17040 34228 -16976 34292
rect -17040 34148 -16976 34212
rect -17040 34068 -16976 34132
rect -17040 33988 -16976 34052
rect -17040 33908 -16976 33972
rect -17040 33828 -16976 33892
rect -17040 33748 -16976 33812
rect -17040 33668 -16976 33732
rect -17040 33588 -16976 33652
rect -17040 33508 -16976 33572
rect -17040 33428 -16976 33492
rect -17040 33348 -16976 33412
rect -17040 33268 -16976 33332
rect -17040 33188 -16976 33252
rect -17040 33108 -16976 33172
rect -17040 33028 -16976 33092
rect -17040 32948 -16976 33012
rect -17040 32868 -16976 32932
rect -17040 32788 -16976 32852
rect -17040 32708 -16976 32772
rect -17040 32628 -16976 32692
rect -17040 32548 -16976 32612
rect -17040 32468 -16976 32532
rect -17040 32388 -16976 32452
rect -17040 32308 -16976 32372
rect -17040 32228 -16976 32292
rect -17040 32148 -16976 32212
rect -17040 32068 -16976 32132
rect -11428 37028 -11364 37092
rect -11428 36948 -11364 37012
rect -11428 36868 -11364 36932
rect -11428 36788 -11364 36852
rect -11428 36708 -11364 36772
rect -11428 36628 -11364 36692
rect -11428 36548 -11364 36612
rect -11428 36468 -11364 36532
rect -11428 36388 -11364 36452
rect -11428 36308 -11364 36372
rect -11428 36228 -11364 36292
rect -11428 36148 -11364 36212
rect -11428 36068 -11364 36132
rect -11428 35988 -11364 36052
rect -11428 35908 -11364 35972
rect -11428 35828 -11364 35892
rect -11428 35748 -11364 35812
rect -11428 35668 -11364 35732
rect -11428 35588 -11364 35652
rect -11428 35508 -11364 35572
rect -11428 35428 -11364 35492
rect -11428 35348 -11364 35412
rect -11428 35268 -11364 35332
rect -11428 35188 -11364 35252
rect -11428 35108 -11364 35172
rect -11428 35028 -11364 35092
rect -11428 34948 -11364 35012
rect -11428 34868 -11364 34932
rect -11428 34788 -11364 34852
rect -11428 34708 -11364 34772
rect -11428 34628 -11364 34692
rect -11428 34548 -11364 34612
rect -11428 34468 -11364 34532
rect -11428 34388 -11364 34452
rect -11428 34308 -11364 34372
rect -11428 34228 -11364 34292
rect -11428 34148 -11364 34212
rect -11428 34068 -11364 34132
rect -11428 33988 -11364 34052
rect -11428 33908 -11364 33972
rect -11428 33828 -11364 33892
rect -11428 33748 -11364 33812
rect -11428 33668 -11364 33732
rect -11428 33588 -11364 33652
rect -11428 33508 -11364 33572
rect -11428 33428 -11364 33492
rect -11428 33348 -11364 33412
rect -11428 33268 -11364 33332
rect -11428 33188 -11364 33252
rect -11428 33108 -11364 33172
rect -11428 33028 -11364 33092
rect -11428 32948 -11364 33012
rect -11428 32868 -11364 32932
rect -11428 32788 -11364 32852
rect -11428 32708 -11364 32772
rect -11428 32628 -11364 32692
rect -11428 32548 -11364 32612
rect -11428 32468 -11364 32532
rect -11428 32388 -11364 32452
rect -11428 32308 -11364 32372
rect -11428 32228 -11364 32292
rect -11428 32148 -11364 32212
rect -11428 32068 -11364 32132
rect -5816 37028 -5752 37092
rect -5816 36948 -5752 37012
rect -5816 36868 -5752 36932
rect -5816 36788 -5752 36852
rect -5816 36708 -5752 36772
rect -5816 36628 -5752 36692
rect -5816 36548 -5752 36612
rect -5816 36468 -5752 36532
rect -5816 36388 -5752 36452
rect -5816 36308 -5752 36372
rect -5816 36228 -5752 36292
rect -5816 36148 -5752 36212
rect -5816 36068 -5752 36132
rect -5816 35988 -5752 36052
rect -5816 35908 -5752 35972
rect -5816 35828 -5752 35892
rect -5816 35748 -5752 35812
rect -5816 35668 -5752 35732
rect -5816 35588 -5752 35652
rect -5816 35508 -5752 35572
rect -5816 35428 -5752 35492
rect -5816 35348 -5752 35412
rect -5816 35268 -5752 35332
rect -5816 35188 -5752 35252
rect -5816 35108 -5752 35172
rect -5816 35028 -5752 35092
rect -5816 34948 -5752 35012
rect -5816 34868 -5752 34932
rect -5816 34788 -5752 34852
rect -5816 34708 -5752 34772
rect -5816 34628 -5752 34692
rect -5816 34548 -5752 34612
rect -5816 34468 -5752 34532
rect -5816 34388 -5752 34452
rect -5816 34308 -5752 34372
rect -5816 34228 -5752 34292
rect -5816 34148 -5752 34212
rect -5816 34068 -5752 34132
rect -5816 33988 -5752 34052
rect -5816 33908 -5752 33972
rect -5816 33828 -5752 33892
rect -5816 33748 -5752 33812
rect -5816 33668 -5752 33732
rect -5816 33588 -5752 33652
rect -5816 33508 -5752 33572
rect -5816 33428 -5752 33492
rect -5816 33348 -5752 33412
rect -5816 33268 -5752 33332
rect -5816 33188 -5752 33252
rect -5816 33108 -5752 33172
rect -5816 33028 -5752 33092
rect -5816 32948 -5752 33012
rect -5816 32868 -5752 32932
rect -5816 32788 -5752 32852
rect -5816 32708 -5752 32772
rect -5816 32628 -5752 32692
rect -5816 32548 -5752 32612
rect -5816 32468 -5752 32532
rect -5816 32388 -5752 32452
rect -5816 32308 -5752 32372
rect -5816 32228 -5752 32292
rect -5816 32148 -5752 32212
rect -5816 32068 -5752 32132
rect -204 37028 -140 37092
rect -204 36948 -140 37012
rect -204 36868 -140 36932
rect -204 36788 -140 36852
rect -204 36708 -140 36772
rect -204 36628 -140 36692
rect -204 36548 -140 36612
rect -204 36468 -140 36532
rect -204 36388 -140 36452
rect -204 36308 -140 36372
rect -204 36228 -140 36292
rect -204 36148 -140 36212
rect -204 36068 -140 36132
rect -204 35988 -140 36052
rect -204 35908 -140 35972
rect -204 35828 -140 35892
rect -204 35748 -140 35812
rect -204 35668 -140 35732
rect -204 35588 -140 35652
rect -204 35508 -140 35572
rect -204 35428 -140 35492
rect -204 35348 -140 35412
rect -204 35268 -140 35332
rect -204 35188 -140 35252
rect -204 35108 -140 35172
rect -204 35028 -140 35092
rect -204 34948 -140 35012
rect -204 34868 -140 34932
rect -204 34788 -140 34852
rect -204 34708 -140 34772
rect -204 34628 -140 34692
rect -204 34548 -140 34612
rect -204 34468 -140 34532
rect -204 34388 -140 34452
rect -204 34308 -140 34372
rect -204 34228 -140 34292
rect -204 34148 -140 34212
rect -204 34068 -140 34132
rect -204 33988 -140 34052
rect -204 33908 -140 33972
rect -204 33828 -140 33892
rect -204 33748 -140 33812
rect -204 33668 -140 33732
rect -204 33588 -140 33652
rect -204 33508 -140 33572
rect -204 33428 -140 33492
rect -204 33348 -140 33412
rect -204 33268 -140 33332
rect -204 33188 -140 33252
rect -204 33108 -140 33172
rect -204 33028 -140 33092
rect -204 32948 -140 33012
rect -204 32868 -140 32932
rect -204 32788 -140 32852
rect -204 32708 -140 32772
rect -204 32628 -140 32692
rect -204 32548 -140 32612
rect -204 32468 -140 32532
rect -204 32388 -140 32452
rect -204 32308 -140 32372
rect -204 32228 -140 32292
rect -204 32148 -140 32212
rect -204 32068 -140 32132
rect 5408 37028 5472 37092
rect 5408 36948 5472 37012
rect 5408 36868 5472 36932
rect 5408 36788 5472 36852
rect 5408 36708 5472 36772
rect 5408 36628 5472 36692
rect 5408 36548 5472 36612
rect 5408 36468 5472 36532
rect 5408 36388 5472 36452
rect 5408 36308 5472 36372
rect 5408 36228 5472 36292
rect 5408 36148 5472 36212
rect 5408 36068 5472 36132
rect 5408 35988 5472 36052
rect 5408 35908 5472 35972
rect 5408 35828 5472 35892
rect 5408 35748 5472 35812
rect 5408 35668 5472 35732
rect 5408 35588 5472 35652
rect 5408 35508 5472 35572
rect 5408 35428 5472 35492
rect 5408 35348 5472 35412
rect 5408 35268 5472 35332
rect 5408 35188 5472 35252
rect 5408 35108 5472 35172
rect 5408 35028 5472 35092
rect 5408 34948 5472 35012
rect 5408 34868 5472 34932
rect 5408 34788 5472 34852
rect 5408 34708 5472 34772
rect 5408 34628 5472 34692
rect 5408 34548 5472 34612
rect 5408 34468 5472 34532
rect 5408 34388 5472 34452
rect 5408 34308 5472 34372
rect 5408 34228 5472 34292
rect 5408 34148 5472 34212
rect 5408 34068 5472 34132
rect 5408 33988 5472 34052
rect 5408 33908 5472 33972
rect 5408 33828 5472 33892
rect 5408 33748 5472 33812
rect 5408 33668 5472 33732
rect 5408 33588 5472 33652
rect 5408 33508 5472 33572
rect 5408 33428 5472 33492
rect 5408 33348 5472 33412
rect 5408 33268 5472 33332
rect 5408 33188 5472 33252
rect 5408 33108 5472 33172
rect 5408 33028 5472 33092
rect 5408 32948 5472 33012
rect 5408 32868 5472 32932
rect 5408 32788 5472 32852
rect 5408 32708 5472 32772
rect 5408 32628 5472 32692
rect 5408 32548 5472 32612
rect 5408 32468 5472 32532
rect 5408 32388 5472 32452
rect 5408 32308 5472 32372
rect 5408 32228 5472 32292
rect 5408 32148 5472 32212
rect 5408 32068 5472 32132
rect 11020 37028 11084 37092
rect 11020 36948 11084 37012
rect 11020 36868 11084 36932
rect 11020 36788 11084 36852
rect 11020 36708 11084 36772
rect 11020 36628 11084 36692
rect 11020 36548 11084 36612
rect 11020 36468 11084 36532
rect 11020 36388 11084 36452
rect 11020 36308 11084 36372
rect 11020 36228 11084 36292
rect 11020 36148 11084 36212
rect 11020 36068 11084 36132
rect 11020 35988 11084 36052
rect 11020 35908 11084 35972
rect 11020 35828 11084 35892
rect 11020 35748 11084 35812
rect 11020 35668 11084 35732
rect 11020 35588 11084 35652
rect 11020 35508 11084 35572
rect 11020 35428 11084 35492
rect 11020 35348 11084 35412
rect 11020 35268 11084 35332
rect 11020 35188 11084 35252
rect 11020 35108 11084 35172
rect 11020 35028 11084 35092
rect 11020 34948 11084 35012
rect 11020 34868 11084 34932
rect 11020 34788 11084 34852
rect 11020 34708 11084 34772
rect 11020 34628 11084 34692
rect 11020 34548 11084 34612
rect 11020 34468 11084 34532
rect 11020 34388 11084 34452
rect 11020 34308 11084 34372
rect 11020 34228 11084 34292
rect 11020 34148 11084 34212
rect 11020 34068 11084 34132
rect 11020 33988 11084 34052
rect 11020 33908 11084 33972
rect 11020 33828 11084 33892
rect 11020 33748 11084 33812
rect 11020 33668 11084 33732
rect 11020 33588 11084 33652
rect 11020 33508 11084 33572
rect 11020 33428 11084 33492
rect 11020 33348 11084 33412
rect 11020 33268 11084 33332
rect 11020 33188 11084 33252
rect 11020 33108 11084 33172
rect 11020 33028 11084 33092
rect 11020 32948 11084 33012
rect 11020 32868 11084 32932
rect 11020 32788 11084 32852
rect 11020 32708 11084 32772
rect 11020 32628 11084 32692
rect 11020 32548 11084 32612
rect 11020 32468 11084 32532
rect 11020 32388 11084 32452
rect 11020 32308 11084 32372
rect 11020 32228 11084 32292
rect 11020 32148 11084 32212
rect 11020 32068 11084 32132
rect 16632 37028 16696 37092
rect 16632 36948 16696 37012
rect 16632 36868 16696 36932
rect 16632 36788 16696 36852
rect 16632 36708 16696 36772
rect 16632 36628 16696 36692
rect 16632 36548 16696 36612
rect 16632 36468 16696 36532
rect 16632 36388 16696 36452
rect 16632 36308 16696 36372
rect 16632 36228 16696 36292
rect 16632 36148 16696 36212
rect 16632 36068 16696 36132
rect 16632 35988 16696 36052
rect 16632 35908 16696 35972
rect 16632 35828 16696 35892
rect 16632 35748 16696 35812
rect 16632 35668 16696 35732
rect 16632 35588 16696 35652
rect 16632 35508 16696 35572
rect 16632 35428 16696 35492
rect 16632 35348 16696 35412
rect 16632 35268 16696 35332
rect 16632 35188 16696 35252
rect 16632 35108 16696 35172
rect 16632 35028 16696 35092
rect 16632 34948 16696 35012
rect 16632 34868 16696 34932
rect 16632 34788 16696 34852
rect 16632 34708 16696 34772
rect 16632 34628 16696 34692
rect 16632 34548 16696 34612
rect 16632 34468 16696 34532
rect 16632 34388 16696 34452
rect 16632 34308 16696 34372
rect 16632 34228 16696 34292
rect 16632 34148 16696 34212
rect 16632 34068 16696 34132
rect 16632 33988 16696 34052
rect 16632 33908 16696 33972
rect 16632 33828 16696 33892
rect 16632 33748 16696 33812
rect 16632 33668 16696 33732
rect 16632 33588 16696 33652
rect 16632 33508 16696 33572
rect 16632 33428 16696 33492
rect 16632 33348 16696 33412
rect 16632 33268 16696 33332
rect 16632 33188 16696 33252
rect 16632 33108 16696 33172
rect 16632 33028 16696 33092
rect 16632 32948 16696 33012
rect 16632 32868 16696 32932
rect 16632 32788 16696 32852
rect 16632 32708 16696 32772
rect 16632 32628 16696 32692
rect 16632 32548 16696 32612
rect 16632 32468 16696 32532
rect 16632 32388 16696 32452
rect 16632 32308 16696 32372
rect 16632 32228 16696 32292
rect 16632 32148 16696 32212
rect 16632 32068 16696 32132
rect 22244 37028 22308 37092
rect 22244 36948 22308 37012
rect 22244 36868 22308 36932
rect 22244 36788 22308 36852
rect 22244 36708 22308 36772
rect 22244 36628 22308 36692
rect 22244 36548 22308 36612
rect 22244 36468 22308 36532
rect 22244 36388 22308 36452
rect 22244 36308 22308 36372
rect 22244 36228 22308 36292
rect 22244 36148 22308 36212
rect 22244 36068 22308 36132
rect 22244 35988 22308 36052
rect 22244 35908 22308 35972
rect 22244 35828 22308 35892
rect 22244 35748 22308 35812
rect 22244 35668 22308 35732
rect 22244 35588 22308 35652
rect 22244 35508 22308 35572
rect 22244 35428 22308 35492
rect 22244 35348 22308 35412
rect 22244 35268 22308 35332
rect 22244 35188 22308 35252
rect 22244 35108 22308 35172
rect 22244 35028 22308 35092
rect 22244 34948 22308 35012
rect 22244 34868 22308 34932
rect 22244 34788 22308 34852
rect 22244 34708 22308 34772
rect 22244 34628 22308 34692
rect 22244 34548 22308 34612
rect 22244 34468 22308 34532
rect 22244 34388 22308 34452
rect 22244 34308 22308 34372
rect 22244 34228 22308 34292
rect 22244 34148 22308 34212
rect 22244 34068 22308 34132
rect 22244 33988 22308 34052
rect 22244 33908 22308 33972
rect 22244 33828 22308 33892
rect 22244 33748 22308 33812
rect 22244 33668 22308 33732
rect 22244 33588 22308 33652
rect 22244 33508 22308 33572
rect 22244 33428 22308 33492
rect 22244 33348 22308 33412
rect 22244 33268 22308 33332
rect 22244 33188 22308 33252
rect 22244 33108 22308 33172
rect 22244 33028 22308 33092
rect 22244 32948 22308 33012
rect 22244 32868 22308 32932
rect 22244 32788 22308 32852
rect 22244 32708 22308 32772
rect 22244 32628 22308 32692
rect 22244 32548 22308 32612
rect 22244 32468 22308 32532
rect 22244 32388 22308 32452
rect 22244 32308 22308 32372
rect 22244 32228 22308 32292
rect 22244 32148 22308 32212
rect 22244 32068 22308 32132
rect 27856 37028 27920 37092
rect 27856 36948 27920 37012
rect 27856 36868 27920 36932
rect 27856 36788 27920 36852
rect 27856 36708 27920 36772
rect 27856 36628 27920 36692
rect 27856 36548 27920 36612
rect 27856 36468 27920 36532
rect 27856 36388 27920 36452
rect 27856 36308 27920 36372
rect 27856 36228 27920 36292
rect 27856 36148 27920 36212
rect 27856 36068 27920 36132
rect 27856 35988 27920 36052
rect 27856 35908 27920 35972
rect 27856 35828 27920 35892
rect 27856 35748 27920 35812
rect 27856 35668 27920 35732
rect 27856 35588 27920 35652
rect 27856 35508 27920 35572
rect 27856 35428 27920 35492
rect 27856 35348 27920 35412
rect 27856 35268 27920 35332
rect 27856 35188 27920 35252
rect 27856 35108 27920 35172
rect 27856 35028 27920 35092
rect 27856 34948 27920 35012
rect 27856 34868 27920 34932
rect 27856 34788 27920 34852
rect 27856 34708 27920 34772
rect 27856 34628 27920 34692
rect 27856 34548 27920 34612
rect 27856 34468 27920 34532
rect 27856 34388 27920 34452
rect 27856 34308 27920 34372
rect 27856 34228 27920 34292
rect 27856 34148 27920 34212
rect 27856 34068 27920 34132
rect 27856 33988 27920 34052
rect 27856 33908 27920 33972
rect 27856 33828 27920 33892
rect 27856 33748 27920 33812
rect 27856 33668 27920 33732
rect 27856 33588 27920 33652
rect 27856 33508 27920 33572
rect 27856 33428 27920 33492
rect 27856 33348 27920 33412
rect 27856 33268 27920 33332
rect 27856 33188 27920 33252
rect 27856 33108 27920 33172
rect 27856 33028 27920 33092
rect 27856 32948 27920 33012
rect 27856 32868 27920 32932
rect 27856 32788 27920 32852
rect 27856 32708 27920 32772
rect 27856 32628 27920 32692
rect 27856 32548 27920 32612
rect 27856 32468 27920 32532
rect 27856 32388 27920 32452
rect 27856 32308 27920 32372
rect 27856 32228 27920 32292
rect 27856 32148 27920 32212
rect 27856 32068 27920 32132
rect 33468 37028 33532 37092
rect 33468 36948 33532 37012
rect 33468 36868 33532 36932
rect 33468 36788 33532 36852
rect 33468 36708 33532 36772
rect 33468 36628 33532 36692
rect 33468 36548 33532 36612
rect 33468 36468 33532 36532
rect 33468 36388 33532 36452
rect 33468 36308 33532 36372
rect 33468 36228 33532 36292
rect 33468 36148 33532 36212
rect 33468 36068 33532 36132
rect 33468 35988 33532 36052
rect 33468 35908 33532 35972
rect 33468 35828 33532 35892
rect 33468 35748 33532 35812
rect 33468 35668 33532 35732
rect 33468 35588 33532 35652
rect 33468 35508 33532 35572
rect 33468 35428 33532 35492
rect 33468 35348 33532 35412
rect 33468 35268 33532 35332
rect 33468 35188 33532 35252
rect 33468 35108 33532 35172
rect 33468 35028 33532 35092
rect 33468 34948 33532 35012
rect 33468 34868 33532 34932
rect 33468 34788 33532 34852
rect 33468 34708 33532 34772
rect 33468 34628 33532 34692
rect 33468 34548 33532 34612
rect 33468 34468 33532 34532
rect 33468 34388 33532 34452
rect 33468 34308 33532 34372
rect 33468 34228 33532 34292
rect 33468 34148 33532 34212
rect 33468 34068 33532 34132
rect 33468 33988 33532 34052
rect 33468 33908 33532 33972
rect 33468 33828 33532 33892
rect 33468 33748 33532 33812
rect 33468 33668 33532 33732
rect 33468 33588 33532 33652
rect 33468 33508 33532 33572
rect 33468 33428 33532 33492
rect 33468 33348 33532 33412
rect 33468 33268 33532 33332
rect 33468 33188 33532 33252
rect 33468 33108 33532 33172
rect 33468 33028 33532 33092
rect 33468 32948 33532 33012
rect 33468 32868 33532 32932
rect 33468 32788 33532 32852
rect 33468 32708 33532 32772
rect 33468 32628 33532 32692
rect 33468 32548 33532 32612
rect 33468 32468 33532 32532
rect 33468 32388 33532 32452
rect 33468 32308 33532 32372
rect 33468 32228 33532 32292
rect 33468 32148 33532 32212
rect 33468 32068 33532 32132
rect 39080 37028 39144 37092
rect 39080 36948 39144 37012
rect 39080 36868 39144 36932
rect 39080 36788 39144 36852
rect 39080 36708 39144 36772
rect 39080 36628 39144 36692
rect 39080 36548 39144 36612
rect 39080 36468 39144 36532
rect 39080 36388 39144 36452
rect 39080 36308 39144 36372
rect 39080 36228 39144 36292
rect 39080 36148 39144 36212
rect 39080 36068 39144 36132
rect 39080 35988 39144 36052
rect 39080 35908 39144 35972
rect 39080 35828 39144 35892
rect 39080 35748 39144 35812
rect 39080 35668 39144 35732
rect 39080 35588 39144 35652
rect 39080 35508 39144 35572
rect 39080 35428 39144 35492
rect 39080 35348 39144 35412
rect 39080 35268 39144 35332
rect 39080 35188 39144 35252
rect 39080 35108 39144 35172
rect 39080 35028 39144 35092
rect 39080 34948 39144 35012
rect 39080 34868 39144 34932
rect 39080 34788 39144 34852
rect 39080 34708 39144 34772
rect 39080 34628 39144 34692
rect 39080 34548 39144 34612
rect 39080 34468 39144 34532
rect 39080 34388 39144 34452
rect 39080 34308 39144 34372
rect 39080 34228 39144 34292
rect 39080 34148 39144 34212
rect 39080 34068 39144 34132
rect 39080 33988 39144 34052
rect 39080 33908 39144 33972
rect 39080 33828 39144 33892
rect 39080 33748 39144 33812
rect 39080 33668 39144 33732
rect 39080 33588 39144 33652
rect 39080 33508 39144 33572
rect 39080 33428 39144 33492
rect 39080 33348 39144 33412
rect 39080 33268 39144 33332
rect 39080 33188 39144 33252
rect 39080 33108 39144 33172
rect 39080 33028 39144 33092
rect 39080 32948 39144 33012
rect 39080 32868 39144 32932
rect 39080 32788 39144 32852
rect 39080 32708 39144 32772
rect 39080 32628 39144 32692
rect 39080 32548 39144 32612
rect 39080 32468 39144 32532
rect 39080 32388 39144 32452
rect 39080 32308 39144 32372
rect 39080 32228 39144 32292
rect 39080 32148 39144 32212
rect 39080 32068 39144 32132
rect -33876 31708 -33812 31772
rect -33876 31628 -33812 31692
rect -33876 31548 -33812 31612
rect -33876 31468 -33812 31532
rect -33876 31388 -33812 31452
rect -33876 31308 -33812 31372
rect -33876 31228 -33812 31292
rect -33876 31148 -33812 31212
rect -33876 31068 -33812 31132
rect -33876 30988 -33812 31052
rect -33876 30908 -33812 30972
rect -33876 30828 -33812 30892
rect -33876 30748 -33812 30812
rect -33876 30668 -33812 30732
rect -33876 30588 -33812 30652
rect -33876 30508 -33812 30572
rect -33876 30428 -33812 30492
rect -33876 30348 -33812 30412
rect -33876 30268 -33812 30332
rect -33876 30188 -33812 30252
rect -33876 30108 -33812 30172
rect -33876 30028 -33812 30092
rect -33876 29948 -33812 30012
rect -33876 29868 -33812 29932
rect -33876 29788 -33812 29852
rect -33876 29708 -33812 29772
rect -33876 29628 -33812 29692
rect -33876 29548 -33812 29612
rect -33876 29468 -33812 29532
rect -33876 29388 -33812 29452
rect -33876 29308 -33812 29372
rect -33876 29228 -33812 29292
rect -33876 29148 -33812 29212
rect -33876 29068 -33812 29132
rect -33876 28988 -33812 29052
rect -33876 28908 -33812 28972
rect -33876 28828 -33812 28892
rect -33876 28748 -33812 28812
rect -33876 28668 -33812 28732
rect -33876 28588 -33812 28652
rect -33876 28508 -33812 28572
rect -33876 28428 -33812 28492
rect -33876 28348 -33812 28412
rect -33876 28268 -33812 28332
rect -33876 28188 -33812 28252
rect -33876 28108 -33812 28172
rect -33876 28028 -33812 28092
rect -33876 27948 -33812 28012
rect -33876 27868 -33812 27932
rect -33876 27788 -33812 27852
rect -33876 27708 -33812 27772
rect -33876 27628 -33812 27692
rect -33876 27548 -33812 27612
rect -33876 27468 -33812 27532
rect -33876 27388 -33812 27452
rect -33876 27308 -33812 27372
rect -33876 27228 -33812 27292
rect -33876 27148 -33812 27212
rect -33876 27068 -33812 27132
rect -33876 26988 -33812 27052
rect -33876 26908 -33812 26972
rect -33876 26828 -33812 26892
rect -33876 26748 -33812 26812
rect -28264 31708 -28200 31772
rect -28264 31628 -28200 31692
rect -28264 31548 -28200 31612
rect -28264 31468 -28200 31532
rect -28264 31388 -28200 31452
rect -28264 31308 -28200 31372
rect -28264 31228 -28200 31292
rect -28264 31148 -28200 31212
rect -28264 31068 -28200 31132
rect -28264 30988 -28200 31052
rect -28264 30908 -28200 30972
rect -28264 30828 -28200 30892
rect -28264 30748 -28200 30812
rect -28264 30668 -28200 30732
rect -28264 30588 -28200 30652
rect -28264 30508 -28200 30572
rect -28264 30428 -28200 30492
rect -28264 30348 -28200 30412
rect -28264 30268 -28200 30332
rect -28264 30188 -28200 30252
rect -28264 30108 -28200 30172
rect -28264 30028 -28200 30092
rect -28264 29948 -28200 30012
rect -28264 29868 -28200 29932
rect -28264 29788 -28200 29852
rect -28264 29708 -28200 29772
rect -28264 29628 -28200 29692
rect -28264 29548 -28200 29612
rect -28264 29468 -28200 29532
rect -28264 29388 -28200 29452
rect -28264 29308 -28200 29372
rect -28264 29228 -28200 29292
rect -28264 29148 -28200 29212
rect -28264 29068 -28200 29132
rect -28264 28988 -28200 29052
rect -28264 28908 -28200 28972
rect -28264 28828 -28200 28892
rect -28264 28748 -28200 28812
rect -28264 28668 -28200 28732
rect -28264 28588 -28200 28652
rect -28264 28508 -28200 28572
rect -28264 28428 -28200 28492
rect -28264 28348 -28200 28412
rect -28264 28268 -28200 28332
rect -28264 28188 -28200 28252
rect -28264 28108 -28200 28172
rect -28264 28028 -28200 28092
rect -28264 27948 -28200 28012
rect -28264 27868 -28200 27932
rect -28264 27788 -28200 27852
rect -28264 27708 -28200 27772
rect -28264 27628 -28200 27692
rect -28264 27548 -28200 27612
rect -28264 27468 -28200 27532
rect -28264 27388 -28200 27452
rect -28264 27308 -28200 27372
rect -28264 27228 -28200 27292
rect -28264 27148 -28200 27212
rect -28264 27068 -28200 27132
rect -28264 26988 -28200 27052
rect -28264 26908 -28200 26972
rect -28264 26828 -28200 26892
rect -28264 26748 -28200 26812
rect -22652 31708 -22588 31772
rect -22652 31628 -22588 31692
rect -22652 31548 -22588 31612
rect -22652 31468 -22588 31532
rect -22652 31388 -22588 31452
rect -22652 31308 -22588 31372
rect -22652 31228 -22588 31292
rect -22652 31148 -22588 31212
rect -22652 31068 -22588 31132
rect -22652 30988 -22588 31052
rect -22652 30908 -22588 30972
rect -22652 30828 -22588 30892
rect -22652 30748 -22588 30812
rect -22652 30668 -22588 30732
rect -22652 30588 -22588 30652
rect -22652 30508 -22588 30572
rect -22652 30428 -22588 30492
rect -22652 30348 -22588 30412
rect -22652 30268 -22588 30332
rect -22652 30188 -22588 30252
rect -22652 30108 -22588 30172
rect -22652 30028 -22588 30092
rect -22652 29948 -22588 30012
rect -22652 29868 -22588 29932
rect -22652 29788 -22588 29852
rect -22652 29708 -22588 29772
rect -22652 29628 -22588 29692
rect -22652 29548 -22588 29612
rect -22652 29468 -22588 29532
rect -22652 29388 -22588 29452
rect -22652 29308 -22588 29372
rect -22652 29228 -22588 29292
rect -22652 29148 -22588 29212
rect -22652 29068 -22588 29132
rect -22652 28988 -22588 29052
rect -22652 28908 -22588 28972
rect -22652 28828 -22588 28892
rect -22652 28748 -22588 28812
rect -22652 28668 -22588 28732
rect -22652 28588 -22588 28652
rect -22652 28508 -22588 28572
rect -22652 28428 -22588 28492
rect -22652 28348 -22588 28412
rect -22652 28268 -22588 28332
rect -22652 28188 -22588 28252
rect -22652 28108 -22588 28172
rect -22652 28028 -22588 28092
rect -22652 27948 -22588 28012
rect -22652 27868 -22588 27932
rect -22652 27788 -22588 27852
rect -22652 27708 -22588 27772
rect -22652 27628 -22588 27692
rect -22652 27548 -22588 27612
rect -22652 27468 -22588 27532
rect -22652 27388 -22588 27452
rect -22652 27308 -22588 27372
rect -22652 27228 -22588 27292
rect -22652 27148 -22588 27212
rect -22652 27068 -22588 27132
rect -22652 26988 -22588 27052
rect -22652 26908 -22588 26972
rect -22652 26828 -22588 26892
rect -22652 26748 -22588 26812
rect -17040 31708 -16976 31772
rect -17040 31628 -16976 31692
rect -17040 31548 -16976 31612
rect -17040 31468 -16976 31532
rect -17040 31388 -16976 31452
rect -17040 31308 -16976 31372
rect -17040 31228 -16976 31292
rect -17040 31148 -16976 31212
rect -17040 31068 -16976 31132
rect -17040 30988 -16976 31052
rect -17040 30908 -16976 30972
rect -17040 30828 -16976 30892
rect -17040 30748 -16976 30812
rect -17040 30668 -16976 30732
rect -17040 30588 -16976 30652
rect -17040 30508 -16976 30572
rect -17040 30428 -16976 30492
rect -17040 30348 -16976 30412
rect -17040 30268 -16976 30332
rect -17040 30188 -16976 30252
rect -17040 30108 -16976 30172
rect -17040 30028 -16976 30092
rect -17040 29948 -16976 30012
rect -17040 29868 -16976 29932
rect -17040 29788 -16976 29852
rect -17040 29708 -16976 29772
rect -17040 29628 -16976 29692
rect -17040 29548 -16976 29612
rect -17040 29468 -16976 29532
rect -17040 29388 -16976 29452
rect -17040 29308 -16976 29372
rect -17040 29228 -16976 29292
rect -17040 29148 -16976 29212
rect -17040 29068 -16976 29132
rect -17040 28988 -16976 29052
rect -17040 28908 -16976 28972
rect -17040 28828 -16976 28892
rect -17040 28748 -16976 28812
rect -17040 28668 -16976 28732
rect -17040 28588 -16976 28652
rect -17040 28508 -16976 28572
rect -17040 28428 -16976 28492
rect -17040 28348 -16976 28412
rect -17040 28268 -16976 28332
rect -17040 28188 -16976 28252
rect -17040 28108 -16976 28172
rect -17040 28028 -16976 28092
rect -17040 27948 -16976 28012
rect -17040 27868 -16976 27932
rect -17040 27788 -16976 27852
rect -17040 27708 -16976 27772
rect -17040 27628 -16976 27692
rect -17040 27548 -16976 27612
rect -17040 27468 -16976 27532
rect -17040 27388 -16976 27452
rect -17040 27308 -16976 27372
rect -17040 27228 -16976 27292
rect -17040 27148 -16976 27212
rect -17040 27068 -16976 27132
rect -17040 26988 -16976 27052
rect -17040 26908 -16976 26972
rect -17040 26828 -16976 26892
rect -17040 26748 -16976 26812
rect -11428 31708 -11364 31772
rect -11428 31628 -11364 31692
rect -11428 31548 -11364 31612
rect -11428 31468 -11364 31532
rect -11428 31388 -11364 31452
rect -11428 31308 -11364 31372
rect -11428 31228 -11364 31292
rect -11428 31148 -11364 31212
rect -11428 31068 -11364 31132
rect -11428 30988 -11364 31052
rect -11428 30908 -11364 30972
rect -11428 30828 -11364 30892
rect -11428 30748 -11364 30812
rect -11428 30668 -11364 30732
rect -11428 30588 -11364 30652
rect -11428 30508 -11364 30572
rect -11428 30428 -11364 30492
rect -11428 30348 -11364 30412
rect -11428 30268 -11364 30332
rect -11428 30188 -11364 30252
rect -11428 30108 -11364 30172
rect -11428 30028 -11364 30092
rect -11428 29948 -11364 30012
rect -11428 29868 -11364 29932
rect -11428 29788 -11364 29852
rect -11428 29708 -11364 29772
rect -11428 29628 -11364 29692
rect -11428 29548 -11364 29612
rect -11428 29468 -11364 29532
rect -11428 29388 -11364 29452
rect -11428 29308 -11364 29372
rect -11428 29228 -11364 29292
rect -11428 29148 -11364 29212
rect -11428 29068 -11364 29132
rect -11428 28988 -11364 29052
rect -11428 28908 -11364 28972
rect -11428 28828 -11364 28892
rect -11428 28748 -11364 28812
rect -11428 28668 -11364 28732
rect -11428 28588 -11364 28652
rect -11428 28508 -11364 28572
rect -11428 28428 -11364 28492
rect -11428 28348 -11364 28412
rect -11428 28268 -11364 28332
rect -11428 28188 -11364 28252
rect -11428 28108 -11364 28172
rect -11428 28028 -11364 28092
rect -11428 27948 -11364 28012
rect -11428 27868 -11364 27932
rect -11428 27788 -11364 27852
rect -11428 27708 -11364 27772
rect -11428 27628 -11364 27692
rect -11428 27548 -11364 27612
rect -11428 27468 -11364 27532
rect -11428 27388 -11364 27452
rect -11428 27308 -11364 27372
rect -11428 27228 -11364 27292
rect -11428 27148 -11364 27212
rect -11428 27068 -11364 27132
rect -11428 26988 -11364 27052
rect -11428 26908 -11364 26972
rect -11428 26828 -11364 26892
rect -11428 26748 -11364 26812
rect -5816 31708 -5752 31772
rect -5816 31628 -5752 31692
rect -5816 31548 -5752 31612
rect -5816 31468 -5752 31532
rect -5816 31388 -5752 31452
rect -5816 31308 -5752 31372
rect -5816 31228 -5752 31292
rect -5816 31148 -5752 31212
rect -5816 31068 -5752 31132
rect -5816 30988 -5752 31052
rect -5816 30908 -5752 30972
rect -5816 30828 -5752 30892
rect -5816 30748 -5752 30812
rect -5816 30668 -5752 30732
rect -5816 30588 -5752 30652
rect -5816 30508 -5752 30572
rect -5816 30428 -5752 30492
rect -5816 30348 -5752 30412
rect -5816 30268 -5752 30332
rect -5816 30188 -5752 30252
rect -5816 30108 -5752 30172
rect -5816 30028 -5752 30092
rect -5816 29948 -5752 30012
rect -5816 29868 -5752 29932
rect -5816 29788 -5752 29852
rect -5816 29708 -5752 29772
rect -5816 29628 -5752 29692
rect -5816 29548 -5752 29612
rect -5816 29468 -5752 29532
rect -5816 29388 -5752 29452
rect -5816 29308 -5752 29372
rect -5816 29228 -5752 29292
rect -5816 29148 -5752 29212
rect -5816 29068 -5752 29132
rect -5816 28988 -5752 29052
rect -5816 28908 -5752 28972
rect -5816 28828 -5752 28892
rect -5816 28748 -5752 28812
rect -5816 28668 -5752 28732
rect -5816 28588 -5752 28652
rect -5816 28508 -5752 28572
rect -5816 28428 -5752 28492
rect -5816 28348 -5752 28412
rect -5816 28268 -5752 28332
rect -5816 28188 -5752 28252
rect -5816 28108 -5752 28172
rect -5816 28028 -5752 28092
rect -5816 27948 -5752 28012
rect -5816 27868 -5752 27932
rect -5816 27788 -5752 27852
rect -5816 27708 -5752 27772
rect -5816 27628 -5752 27692
rect -5816 27548 -5752 27612
rect -5816 27468 -5752 27532
rect -5816 27388 -5752 27452
rect -5816 27308 -5752 27372
rect -5816 27228 -5752 27292
rect -5816 27148 -5752 27212
rect -5816 27068 -5752 27132
rect -5816 26988 -5752 27052
rect -5816 26908 -5752 26972
rect -5816 26828 -5752 26892
rect -5816 26748 -5752 26812
rect -204 31708 -140 31772
rect -204 31628 -140 31692
rect -204 31548 -140 31612
rect -204 31468 -140 31532
rect -204 31388 -140 31452
rect -204 31308 -140 31372
rect -204 31228 -140 31292
rect -204 31148 -140 31212
rect -204 31068 -140 31132
rect -204 30988 -140 31052
rect -204 30908 -140 30972
rect -204 30828 -140 30892
rect -204 30748 -140 30812
rect -204 30668 -140 30732
rect -204 30588 -140 30652
rect -204 30508 -140 30572
rect -204 30428 -140 30492
rect -204 30348 -140 30412
rect -204 30268 -140 30332
rect -204 30188 -140 30252
rect -204 30108 -140 30172
rect -204 30028 -140 30092
rect -204 29948 -140 30012
rect -204 29868 -140 29932
rect -204 29788 -140 29852
rect -204 29708 -140 29772
rect -204 29628 -140 29692
rect -204 29548 -140 29612
rect -204 29468 -140 29532
rect -204 29388 -140 29452
rect -204 29308 -140 29372
rect -204 29228 -140 29292
rect -204 29148 -140 29212
rect -204 29068 -140 29132
rect -204 28988 -140 29052
rect -204 28908 -140 28972
rect -204 28828 -140 28892
rect -204 28748 -140 28812
rect -204 28668 -140 28732
rect -204 28588 -140 28652
rect -204 28508 -140 28572
rect -204 28428 -140 28492
rect -204 28348 -140 28412
rect -204 28268 -140 28332
rect -204 28188 -140 28252
rect -204 28108 -140 28172
rect -204 28028 -140 28092
rect -204 27948 -140 28012
rect -204 27868 -140 27932
rect -204 27788 -140 27852
rect -204 27708 -140 27772
rect -204 27628 -140 27692
rect -204 27548 -140 27612
rect -204 27468 -140 27532
rect -204 27388 -140 27452
rect -204 27308 -140 27372
rect -204 27228 -140 27292
rect -204 27148 -140 27212
rect -204 27068 -140 27132
rect -204 26988 -140 27052
rect -204 26908 -140 26972
rect -204 26828 -140 26892
rect -204 26748 -140 26812
rect 5408 31708 5472 31772
rect 5408 31628 5472 31692
rect 5408 31548 5472 31612
rect 5408 31468 5472 31532
rect 5408 31388 5472 31452
rect 5408 31308 5472 31372
rect 5408 31228 5472 31292
rect 5408 31148 5472 31212
rect 5408 31068 5472 31132
rect 5408 30988 5472 31052
rect 5408 30908 5472 30972
rect 5408 30828 5472 30892
rect 5408 30748 5472 30812
rect 5408 30668 5472 30732
rect 5408 30588 5472 30652
rect 5408 30508 5472 30572
rect 5408 30428 5472 30492
rect 5408 30348 5472 30412
rect 5408 30268 5472 30332
rect 5408 30188 5472 30252
rect 5408 30108 5472 30172
rect 5408 30028 5472 30092
rect 5408 29948 5472 30012
rect 5408 29868 5472 29932
rect 5408 29788 5472 29852
rect 5408 29708 5472 29772
rect 5408 29628 5472 29692
rect 5408 29548 5472 29612
rect 5408 29468 5472 29532
rect 5408 29388 5472 29452
rect 5408 29308 5472 29372
rect 5408 29228 5472 29292
rect 5408 29148 5472 29212
rect 5408 29068 5472 29132
rect 5408 28988 5472 29052
rect 5408 28908 5472 28972
rect 5408 28828 5472 28892
rect 5408 28748 5472 28812
rect 5408 28668 5472 28732
rect 5408 28588 5472 28652
rect 5408 28508 5472 28572
rect 5408 28428 5472 28492
rect 5408 28348 5472 28412
rect 5408 28268 5472 28332
rect 5408 28188 5472 28252
rect 5408 28108 5472 28172
rect 5408 28028 5472 28092
rect 5408 27948 5472 28012
rect 5408 27868 5472 27932
rect 5408 27788 5472 27852
rect 5408 27708 5472 27772
rect 5408 27628 5472 27692
rect 5408 27548 5472 27612
rect 5408 27468 5472 27532
rect 5408 27388 5472 27452
rect 5408 27308 5472 27372
rect 5408 27228 5472 27292
rect 5408 27148 5472 27212
rect 5408 27068 5472 27132
rect 5408 26988 5472 27052
rect 5408 26908 5472 26972
rect 5408 26828 5472 26892
rect 5408 26748 5472 26812
rect 11020 31708 11084 31772
rect 11020 31628 11084 31692
rect 11020 31548 11084 31612
rect 11020 31468 11084 31532
rect 11020 31388 11084 31452
rect 11020 31308 11084 31372
rect 11020 31228 11084 31292
rect 11020 31148 11084 31212
rect 11020 31068 11084 31132
rect 11020 30988 11084 31052
rect 11020 30908 11084 30972
rect 11020 30828 11084 30892
rect 11020 30748 11084 30812
rect 11020 30668 11084 30732
rect 11020 30588 11084 30652
rect 11020 30508 11084 30572
rect 11020 30428 11084 30492
rect 11020 30348 11084 30412
rect 11020 30268 11084 30332
rect 11020 30188 11084 30252
rect 11020 30108 11084 30172
rect 11020 30028 11084 30092
rect 11020 29948 11084 30012
rect 11020 29868 11084 29932
rect 11020 29788 11084 29852
rect 11020 29708 11084 29772
rect 11020 29628 11084 29692
rect 11020 29548 11084 29612
rect 11020 29468 11084 29532
rect 11020 29388 11084 29452
rect 11020 29308 11084 29372
rect 11020 29228 11084 29292
rect 11020 29148 11084 29212
rect 11020 29068 11084 29132
rect 11020 28988 11084 29052
rect 11020 28908 11084 28972
rect 11020 28828 11084 28892
rect 11020 28748 11084 28812
rect 11020 28668 11084 28732
rect 11020 28588 11084 28652
rect 11020 28508 11084 28572
rect 11020 28428 11084 28492
rect 11020 28348 11084 28412
rect 11020 28268 11084 28332
rect 11020 28188 11084 28252
rect 11020 28108 11084 28172
rect 11020 28028 11084 28092
rect 11020 27948 11084 28012
rect 11020 27868 11084 27932
rect 11020 27788 11084 27852
rect 11020 27708 11084 27772
rect 11020 27628 11084 27692
rect 11020 27548 11084 27612
rect 11020 27468 11084 27532
rect 11020 27388 11084 27452
rect 11020 27308 11084 27372
rect 11020 27228 11084 27292
rect 11020 27148 11084 27212
rect 11020 27068 11084 27132
rect 11020 26988 11084 27052
rect 11020 26908 11084 26972
rect 11020 26828 11084 26892
rect 11020 26748 11084 26812
rect 16632 31708 16696 31772
rect 16632 31628 16696 31692
rect 16632 31548 16696 31612
rect 16632 31468 16696 31532
rect 16632 31388 16696 31452
rect 16632 31308 16696 31372
rect 16632 31228 16696 31292
rect 16632 31148 16696 31212
rect 16632 31068 16696 31132
rect 16632 30988 16696 31052
rect 16632 30908 16696 30972
rect 16632 30828 16696 30892
rect 16632 30748 16696 30812
rect 16632 30668 16696 30732
rect 16632 30588 16696 30652
rect 16632 30508 16696 30572
rect 16632 30428 16696 30492
rect 16632 30348 16696 30412
rect 16632 30268 16696 30332
rect 16632 30188 16696 30252
rect 16632 30108 16696 30172
rect 16632 30028 16696 30092
rect 16632 29948 16696 30012
rect 16632 29868 16696 29932
rect 16632 29788 16696 29852
rect 16632 29708 16696 29772
rect 16632 29628 16696 29692
rect 16632 29548 16696 29612
rect 16632 29468 16696 29532
rect 16632 29388 16696 29452
rect 16632 29308 16696 29372
rect 16632 29228 16696 29292
rect 16632 29148 16696 29212
rect 16632 29068 16696 29132
rect 16632 28988 16696 29052
rect 16632 28908 16696 28972
rect 16632 28828 16696 28892
rect 16632 28748 16696 28812
rect 16632 28668 16696 28732
rect 16632 28588 16696 28652
rect 16632 28508 16696 28572
rect 16632 28428 16696 28492
rect 16632 28348 16696 28412
rect 16632 28268 16696 28332
rect 16632 28188 16696 28252
rect 16632 28108 16696 28172
rect 16632 28028 16696 28092
rect 16632 27948 16696 28012
rect 16632 27868 16696 27932
rect 16632 27788 16696 27852
rect 16632 27708 16696 27772
rect 16632 27628 16696 27692
rect 16632 27548 16696 27612
rect 16632 27468 16696 27532
rect 16632 27388 16696 27452
rect 16632 27308 16696 27372
rect 16632 27228 16696 27292
rect 16632 27148 16696 27212
rect 16632 27068 16696 27132
rect 16632 26988 16696 27052
rect 16632 26908 16696 26972
rect 16632 26828 16696 26892
rect 16632 26748 16696 26812
rect 22244 31708 22308 31772
rect 22244 31628 22308 31692
rect 22244 31548 22308 31612
rect 22244 31468 22308 31532
rect 22244 31388 22308 31452
rect 22244 31308 22308 31372
rect 22244 31228 22308 31292
rect 22244 31148 22308 31212
rect 22244 31068 22308 31132
rect 22244 30988 22308 31052
rect 22244 30908 22308 30972
rect 22244 30828 22308 30892
rect 22244 30748 22308 30812
rect 22244 30668 22308 30732
rect 22244 30588 22308 30652
rect 22244 30508 22308 30572
rect 22244 30428 22308 30492
rect 22244 30348 22308 30412
rect 22244 30268 22308 30332
rect 22244 30188 22308 30252
rect 22244 30108 22308 30172
rect 22244 30028 22308 30092
rect 22244 29948 22308 30012
rect 22244 29868 22308 29932
rect 22244 29788 22308 29852
rect 22244 29708 22308 29772
rect 22244 29628 22308 29692
rect 22244 29548 22308 29612
rect 22244 29468 22308 29532
rect 22244 29388 22308 29452
rect 22244 29308 22308 29372
rect 22244 29228 22308 29292
rect 22244 29148 22308 29212
rect 22244 29068 22308 29132
rect 22244 28988 22308 29052
rect 22244 28908 22308 28972
rect 22244 28828 22308 28892
rect 22244 28748 22308 28812
rect 22244 28668 22308 28732
rect 22244 28588 22308 28652
rect 22244 28508 22308 28572
rect 22244 28428 22308 28492
rect 22244 28348 22308 28412
rect 22244 28268 22308 28332
rect 22244 28188 22308 28252
rect 22244 28108 22308 28172
rect 22244 28028 22308 28092
rect 22244 27948 22308 28012
rect 22244 27868 22308 27932
rect 22244 27788 22308 27852
rect 22244 27708 22308 27772
rect 22244 27628 22308 27692
rect 22244 27548 22308 27612
rect 22244 27468 22308 27532
rect 22244 27388 22308 27452
rect 22244 27308 22308 27372
rect 22244 27228 22308 27292
rect 22244 27148 22308 27212
rect 22244 27068 22308 27132
rect 22244 26988 22308 27052
rect 22244 26908 22308 26972
rect 22244 26828 22308 26892
rect 22244 26748 22308 26812
rect 27856 31708 27920 31772
rect 27856 31628 27920 31692
rect 27856 31548 27920 31612
rect 27856 31468 27920 31532
rect 27856 31388 27920 31452
rect 27856 31308 27920 31372
rect 27856 31228 27920 31292
rect 27856 31148 27920 31212
rect 27856 31068 27920 31132
rect 27856 30988 27920 31052
rect 27856 30908 27920 30972
rect 27856 30828 27920 30892
rect 27856 30748 27920 30812
rect 27856 30668 27920 30732
rect 27856 30588 27920 30652
rect 27856 30508 27920 30572
rect 27856 30428 27920 30492
rect 27856 30348 27920 30412
rect 27856 30268 27920 30332
rect 27856 30188 27920 30252
rect 27856 30108 27920 30172
rect 27856 30028 27920 30092
rect 27856 29948 27920 30012
rect 27856 29868 27920 29932
rect 27856 29788 27920 29852
rect 27856 29708 27920 29772
rect 27856 29628 27920 29692
rect 27856 29548 27920 29612
rect 27856 29468 27920 29532
rect 27856 29388 27920 29452
rect 27856 29308 27920 29372
rect 27856 29228 27920 29292
rect 27856 29148 27920 29212
rect 27856 29068 27920 29132
rect 27856 28988 27920 29052
rect 27856 28908 27920 28972
rect 27856 28828 27920 28892
rect 27856 28748 27920 28812
rect 27856 28668 27920 28732
rect 27856 28588 27920 28652
rect 27856 28508 27920 28572
rect 27856 28428 27920 28492
rect 27856 28348 27920 28412
rect 27856 28268 27920 28332
rect 27856 28188 27920 28252
rect 27856 28108 27920 28172
rect 27856 28028 27920 28092
rect 27856 27948 27920 28012
rect 27856 27868 27920 27932
rect 27856 27788 27920 27852
rect 27856 27708 27920 27772
rect 27856 27628 27920 27692
rect 27856 27548 27920 27612
rect 27856 27468 27920 27532
rect 27856 27388 27920 27452
rect 27856 27308 27920 27372
rect 27856 27228 27920 27292
rect 27856 27148 27920 27212
rect 27856 27068 27920 27132
rect 27856 26988 27920 27052
rect 27856 26908 27920 26972
rect 27856 26828 27920 26892
rect 27856 26748 27920 26812
rect 33468 31708 33532 31772
rect 33468 31628 33532 31692
rect 33468 31548 33532 31612
rect 33468 31468 33532 31532
rect 33468 31388 33532 31452
rect 33468 31308 33532 31372
rect 33468 31228 33532 31292
rect 33468 31148 33532 31212
rect 33468 31068 33532 31132
rect 33468 30988 33532 31052
rect 33468 30908 33532 30972
rect 33468 30828 33532 30892
rect 33468 30748 33532 30812
rect 33468 30668 33532 30732
rect 33468 30588 33532 30652
rect 33468 30508 33532 30572
rect 33468 30428 33532 30492
rect 33468 30348 33532 30412
rect 33468 30268 33532 30332
rect 33468 30188 33532 30252
rect 33468 30108 33532 30172
rect 33468 30028 33532 30092
rect 33468 29948 33532 30012
rect 33468 29868 33532 29932
rect 33468 29788 33532 29852
rect 33468 29708 33532 29772
rect 33468 29628 33532 29692
rect 33468 29548 33532 29612
rect 33468 29468 33532 29532
rect 33468 29388 33532 29452
rect 33468 29308 33532 29372
rect 33468 29228 33532 29292
rect 33468 29148 33532 29212
rect 33468 29068 33532 29132
rect 33468 28988 33532 29052
rect 33468 28908 33532 28972
rect 33468 28828 33532 28892
rect 33468 28748 33532 28812
rect 33468 28668 33532 28732
rect 33468 28588 33532 28652
rect 33468 28508 33532 28572
rect 33468 28428 33532 28492
rect 33468 28348 33532 28412
rect 33468 28268 33532 28332
rect 33468 28188 33532 28252
rect 33468 28108 33532 28172
rect 33468 28028 33532 28092
rect 33468 27948 33532 28012
rect 33468 27868 33532 27932
rect 33468 27788 33532 27852
rect 33468 27708 33532 27772
rect 33468 27628 33532 27692
rect 33468 27548 33532 27612
rect 33468 27468 33532 27532
rect 33468 27388 33532 27452
rect 33468 27308 33532 27372
rect 33468 27228 33532 27292
rect 33468 27148 33532 27212
rect 33468 27068 33532 27132
rect 33468 26988 33532 27052
rect 33468 26908 33532 26972
rect 33468 26828 33532 26892
rect 33468 26748 33532 26812
rect 39080 31708 39144 31772
rect 39080 31628 39144 31692
rect 39080 31548 39144 31612
rect 39080 31468 39144 31532
rect 39080 31388 39144 31452
rect 39080 31308 39144 31372
rect 39080 31228 39144 31292
rect 39080 31148 39144 31212
rect 39080 31068 39144 31132
rect 39080 30988 39144 31052
rect 39080 30908 39144 30972
rect 39080 30828 39144 30892
rect 39080 30748 39144 30812
rect 39080 30668 39144 30732
rect 39080 30588 39144 30652
rect 39080 30508 39144 30572
rect 39080 30428 39144 30492
rect 39080 30348 39144 30412
rect 39080 30268 39144 30332
rect 39080 30188 39144 30252
rect 39080 30108 39144 30172
rect 39080 30028 39144 30092
rect 39080 29948 39144 30012
rect 39080 29868 39144 29932
rect 39080 29788 39144 29852
rect 39080 29708 39144 29772
rect 39080 29628 39144 29692
rect 39080 29548 39144 29612
rect 39080 29468 39144 29532
rect 39080 29388 39144 29452
rect 39080 29308 39144 29372
rect 39080 29228 39144 29292
rect 39080 29148 39144 29212
rect 39080 29068 39144 29132
rect 39080 28988 39144 29052
rect 39080 28908 39144 28972
rect 39080 28828 39144 28892
rect 39080 28748 39144 28812
rect 39080 28668 39144 28732
rect 39080 28588 39144 28652
rect 39080 28508 39144 28572
rect 39080 28428 39144 28492
rect 39080 28348 39144 28412
rect 39080 28268 39144 28332
rect 39080 28188 39144 28252
rect 39080 28108 39144 28172
rect 39080 28028 39144 28092
rect 39080 27948 39144 28012
rect 39080 27868 39144 27932
rect 39080 27788 39144 27852
rect 39080 27708 39144 27772
rect 39080 27628 39144 27692
rect 39080 27548 39144 27612
rect 39080 27468 39144 27532
rect 39080 27388 39144 27452
rect 39080 27308 39144 27372
rect 39080 27228 39144 27292
rect 39080 27148 39144 27212
rect 39080 27068 39144 27132
rect 39080 26988 39144 27052
rect 39080 26908 39144 26972
rect 39080 26828 39144 26892
rect 39080 26748 39144 26812
rect -33876 26388 -33812 26452
rect -33876 26308 -33812 26372
rect -33876 26228 -33812 26292
rect -33876 26148 -33812 26212
rect -33876 26068 -33812 26132
rect -33876 25988 -33812 26052
rect -33876 25908 -33812 25972
rect -33876 25828 -33812 25892
rect -33876 25748 -33812 25812
rect -33876 25668 -33812 25732
rect -33876 25588 -33812 25652
rect -33876 25508 -33812 25572
rect -33876 25428 -33812 25492
rect -33876 25348 -33812 25412
rect -33876 25268 -33812 25332
rect -33876 25188 -33812 25252
rect -33876 25108 -33812 25172
rect -33876 25028 -33812 25092
rect -33876 24948 -33812 25012
rect -33876 24868 -33812 24932
rect -33876 24788 -33812 24852
rect -33876 24708 -33812 24772
rect -33876 24628 -33812 24692
rect -33876 24548 -33812 24612
rect -33876 24468 -33812 24532
rect -33876 24388 -33812 24452
rect -33876 24308 -33812 24372
rect -33876 24228 -33812 24292
rect -33876 24148 -33812 24212
rect -33876 24068 -33812 24132
rect -33876 23988 -33812 24052
rect -33876 23908 -33812 23972
rect -33876 23828 -33812 23892
rect -33876 23748 -33812 23812
rect -33876 23668 -33812 23732
rect -33876 23588 -33812 23652
rect -33876 23508 -33812 23572
rect -33876 23428 -33812 23492
rect -33876 23348 -33812 23412
rect -33876 23268 -33812 23332
rect -33876 23188 -33812 23252
rect -33876 23108 -33812 23172
rect -33876 23028 -33812 23092
rect -33876 22948 -33812 23012
rect -33876 22868 -33812 22932
rect -33876 22788 -33812 22852
rect -33876 22708 -33812 22772
rect -33876 22628 -33812 22692
rect -33876 22548 -33812 22612
rect -33876 22468 -33812 22532
rect -33876 22388 -33812 22452
rect -33876 22308 -33812 22372
rect -33876 22228 -33812 22292
rect -33876 22148 -33812 22212
rect -33876 22068 -33812 22132
rect -33876 21988 -33812 22052
rect -33876 21908 -33812 21972
rect -33876 21828 -33812 21892
rect -33876 21748 -33812 21812
rect -33876 21668 -33812 21732
rect -33876 21588 -33812 21652
rect -33876 21508 -33812 21572
rect -33876 21428 -33812 21492
rect -28264 26388 -28200 26452
rect -28264 26308 -28200 26372
rect -28264 26228 -28200 26292
rect -28264 26148 -28200 26212
rect -28264 26068 -28200 26132
rect -28264 25988 -28200 26052
rect -28264 25908 -28200 25972
rect -28264 25828 -28200 25892
rect -28264 25748 -28200 25812
rect -28264 25668 -28200 25732
rect -28264 25588 -28200 25652
rect -28264 25508 -28200 25572
rect -28264 25428 -28200 25492
rect -28264 25348 -28200 25412
rect -28264 25268 -28200 25332
rect -28264 25188 -28200 25252
rect -28264 25108 -28200 25172
rect -28264 25028 -28200 25092
rect -28264 24948 -28200 25012
rect -28264 24868 -28200 24932
rect -28264 24788 -28200 24852
rect -28264 24708 -28200 24772
rect -28264 24628 -28200 24692
rect -28264 24548 -28200 24612
rect -28264 24468 -28200 24532
rect -28264 24388 -28200 24452
rect -28264 24308 -28200 24372
rect -28264 24228 -28200 24292
rect -28264 24148 -28200 24212
rect -28264 24068 -28200 24132
rect -28264 23988 -28200 24052
rect -28264 23908 -28200 23972
rect -28264 23828 -28200 23892
rect -28264 23748 -28200 23812
rect -28264 23668 -28200 23732
rect -28264 23588 -28200 23652
rect -28264 23508 -28200 23572
rect -28264 23428 -28200 23492
rect -28264 23348 -28200 23412
rect -28264 23268 -28200 23332
rect -28264 23188 -28200 23252
rect -28264 23108 -28200 23172
rect -28264 23028 -28200 23092
rect -28264 22948 -28200 23012
rect -28264 22868 -28200 22932
rect -28264 22788 -28200 22852
rect -28264 22708 -28200 22772
rect -28264 22628 -28200 22692
rect -28264 22548 -28200 22612
rect -28264 22468 -28200 22532
rect -28264 22388 -28200 22452
rect -28264 22308 -28200 22372
rect -28264 22228 -28200 22292
rect -28264 22148 -28200 22212
rect -28264 22068 -28200 22132
rect -28264 21988 -28200 22052
rect -28264 21908 -28200 21972
rect -28264 21828 -28200 21892
rect -28264 21748 -28200 21812
rect -28264 21668 -28200 21732
rect -28264 21588 -28200 21652
rect -28264 21508 -28200 21572
rect -28264 21428 -28200 21492
rect -22652 26388 -22588 26452
rect -22652 26308 -22588 26372
rect -22652 26228 -22588 26292
rect -22652 26148 -22588 26212
rect -22652 26068 -22588 26132
rect -22652 25988 -22588 26052
rect -22652 25908 -22588 25972
rect -22652 25828 -22588 25892
rect -22652 25748 -22588 25812
rect -22652 25668 -22588 25732
rect -22652 25588 -22588 25652
rect -22652 25508 -22588 25572
rect -22652 25428 -22588 25492
rect -22652 25348 -22588 25412
rect -22652 25268 -22588 25332
rect -22652 25188 -22588 25252
rect -22652 25108 -22588 25172
rect -22652 25028 -22588 25092
rect -22652 24948 -22588 25012
rect -22652 24868 -22588 24932
rect -22652 24788 -22588 24852
rect -22652 24708 -22588 24772
rect -22652 24628 -22588 24692
rect -22652 24548 -22588 24612
rect -22652 24468 -22588 24532
rect -22652 24388 -22588 24452
rect -22652 24308 -22588 24372
rect -22652 24228 -22588 24292
rect -22652 24148 -22588 24212
rect -22652 24068 -22588 24132
rect -22652 23988 -22588 24052
rect -22652 23908 -22588 23972
rect -22652 23828 -22588 23892
rect -22652 23748 -22588 23812
rect -22652 23668 -22588 23732
rect -22652 23588 -22588 23652
rect -22652 23508 -22588 23572
rect -22652 23428 -22588 23492
rect -22652 23348 -22588 23412
rect -22652 23268 -22588 23332
rect -22652 23188 -22588 23252
rect -22652 23108 -22588 23172
rect -22652 23028 -22588 23092
rect -22652 22948 -22588 23012
rect -22652 22868 -22588 22932
rect -22652 22788 -22588 22852
rect -22652 22708 -22588 22772
rect -22652 22628 -22588 22692
rect -22652 22548 -22588 22612
rect -22652 22468 -22588 22532
rect -22652 22388 -22588 22452
rect -22652 22308 -22588 22372
rect -22652 22228 -22588 22292
rect -22652 22148 -22588 22212
rect -22652 22068 -22588 22132
rect -22652 21988 -22588 22052
rect -22652 21908 -22588 21972
rect -22652 21828 -22588 21892
rect -22652 21748 -22588 21812
rect -22652 21668 -22588 21732
rect -22652 21588 -22588 21652
rect -22652 21508 -22588 21572
rect -22652 21428 -22588 21492
rect -17040 26388 -16976 26452
rect -17040 26308 -16976 26372
rect -17040 26228 -16976 26292
rect -17040 26148 -16976 26212
rect -17040 26068 -16976 26132
rect -17040 25988 -16976 26052
rect -17040 25908 -16976 25972
rect -17040 25828 -16976 25892
rect -17040 25748 -16976 25812
rect -17040 25668 -16976 25732
rect -17040 25588 -16976 25652
rect -17040 25508 -16976 25572
rect -17040 25428 -16976 25492
rect -17040 25348 -16976 25412
rect -17040 25268 -16976 25332
rect -17040 25188 -16976 25252
rect -17040 25108 -16976 25172
rect -17040 25028 -16976 25092
rect -17040 24948 -16976 25012
rect -17040 24868 -16976 24932
rect -17040 24788 -16976 24852
rect -17040 24708 -16976 24772
rect -17040 24628 -16976 24692
rect -17040 24548 -16976 24612
rect -17040 24468 -16976 24532
rect -17040 24388 -16976 24452
rect -17040 24308 -16976 24372
rect -17040 24228 -16976 24292
rect -17040 24148 -16976 24212
rect -17040 24068 -16976 24132
rect -17040 23988 -16976 24052
rect -17040 23908 -16976 23972
rect -17040 23828 -16976 23892
rect -17040 23748 -16976 23812
rect -17040 23668 -16976 23732
rect -17040 23588 -16976 23652
rect -17040 23508 -16976 23572
rect -17040 23428 -16976 23492
rect -17040 23348 -16976 23412
rect -17040 23268 -16976 23332
rect -17040 23188 -16976 23252
rect -17040 23108 -16976 23172
rect -17040 23028 -16976 23092
rect -17040 22948 -16976 23012
rect -17040 22868 -16976 22932
rect -17040 22788 -16976 22852
rect -17040 22708 -16976 22772
rect -17040 22628 -16976 22692
rect -17040 22548 -16976 22612
rect -17040 22468 -16976 22532
rect -17040 22388 -16976 22452
rect -17040 22308 -16976 22372
rect -17040 22228 -16976 22292
rect -17040 22148 -16976 22212
rect -17040 22068 -16976 22132
rect -17040 21988 -16976 22052
rect -17040 21908 -16976 21972
rect -17040 21828 -16976 21892
rect -17040 21748 -16976 21812
rect -17040 21668 -16976 21732
rect -17040 21588 -16976 21652
rect -17040 21508 -16976 21572
rect -17040 21428 -16976 21492
rect -11428 26388 -11364 26452
rect -11428 26308 -11364 26372
rect -11428 26228 -11364 26292
rect -11428 26148 -11364 26212
rect -11428 26068 -11364 26132
rect -11428 25988 -11364 26052
rect -11428 25908 -11364 25972
rect -11428 25828 -11364 25892
rect -11428 25748 -11364 25812
rect -11428 25668 -11364 25732
rect -11428 25588 -11364 25652
rect -11428 25508 -11364 25572
rect -11428 25428 -11364 25492
rect -11428 25348 -11364 25412
rect -11428 25268 -11364 25332
rect -11428 25188 -11364 25252
rect -11428 25108 -11364 25172
rect -11428 25028 -11364 25092
rect -11428 24948 -11364 25012
rect -11428 24868 -11364 24932
rect -11428 24788 -11364 24852
rect -11428 24708 -11364 24772
rect -11428 24628 -11364 24692
rect -11428 24548 -11364 24612
rect -11428 24468 -11364 24532
rect -11428 24388 -11364 24452
rect -11428 24308 -11364 24372
rect -11428 24228 -11364 24292
rect -11428 24148 -11364 24212
rect -11428 24068 -11364 24132
rect -11428 23988 -11364 24052
rect -11428 23908 -11364 23972
rect -11428 23828 -11364 23892
rect -11428 23748 -11364 23812
rect -11428 23668 -11364 23732
rect -11428 23588 -11364 23652
rect -11428 23508 -11364 23572
rect -11428 23428 -11364 23492
rect -11428 23348 -11364 23412
rect -11428 23268 -11364 23332
rect -11428 23188 -11364 23252
rect -11428 23108 -11364 23172
rect -11428 23028 -11364 23092
rect -11428 22948 -11364 23012
rect -11428 22868 -11364 22932
rect -11428 22788 -11364 22852
rect -11428 22708 -11364 22772
rect -11428 22628 -11364 22692
rect -11428 22548 -11364 22612
rect -11428 22468 -11364 22532
rect -11428 22388 -11364 22452
rect -11428 22308 -11364 22372
rect -11428 22228 -11364 22292
rect -11428 22148 -11364 22212
rect -11428 22068 -11364 22132
rect -11428 21988 -11364 22052
rect -11428 21908 -11364 21972
rect -11428 21828 -11364 21892
rect -11428 21748 -11364 21812
rect -11428 21668 -11364 21732
rect -11428 21588 -11364 21652
rect -11428 21508 -11364 21572
rect -11428 21428 -11364 21492
rect -5816 26388 -5752 26452
rect -5816 26308 -5752 26372
rect -5816 26228 -5752 26292
rect -5816 26148 -5752 26212
rect -5816 26068 -5752 26132
rect -5816 25988 -5752 26052
rect -5816 25908 -5752 25972
rect -5816 25828 -5752 25892
rect -5816 25748 -5752 25812
rect -5816 25668 -5752 25732
rect -5816 25588 -5752 25652
rect -5816 25508 -5752 25572
rect -5816 25428 -5752 25492
rect -5816 25348 -5752 25412
rect -5816 25268 -5752 25332
rect -5816 25188 -5752 25252
rect -5816 25108 -5752 25172
rect -5816 25028 -5752 25092
rect -5816 24948 -5752 25012
rect -5816 24868 -5752 24932
rect -5816 24788 -5752 24852
rect -5816 24708 -5752 24772
rect -5816 24628 -5752 24692
rect -5816 24548 -5752 24612
rect -5816 24468 -5752 24532
rect -5816 24388 -5752 24452
rect -5816 24308 -5752 24372
rect -5816 24228 -5752 24292
rect -5816 24148 -5752 24212
rect -5816 24068 -5752 24132
rect -5816 23988 -5752 24052
rect -5816 23908 -5752 23972
rect -5816 23828 -5752 23892
rect -5816 23748 -5752 23812
rect -5816 23668 -5752 23732
rect -5816 23588 -5752 23652
rect -5816 23508 -5752 23572
rect -5816 23428 -5752 23492
rect -5816 23348 -5752 23412
rect -5816 23268 -5752 23332
rect -5816 23188 -5752 23252
rect -5816 23108 -5752 23172
rect -5816 23028 -5752 23092
rect -5816 22948 -5752 23012
rect -5816 22868 -5752 22932
rect -5816 22788 -5752 22852
rect -5816 22708 -5752 22772
rect -5816 22628 -5752 22692
rect -5816 22548 -5752 22612
rect -5816 22468 -5752 22532
rect -5816 22388 -5752 22452
rect -5816 22308 -5752 22372
rect -5816 22228 -5752 22292
rect -5816 22148 -5752 22212
rect -5816 22068 -5752 22132
rect -5816 21988 -5752 22052
rect -5816 21908 -5752 21972
rect -5816 21828 -5752 21892
rect -5816 21748 -5752 21812
rect -5816 21668 -5752 21732
rect -5816 21588 -5752 21652
rect -5816 21508 -5752 21572
rect -5816 21428 -5752 21492
rect -204 26388 -140 26452
rect -204 26308 -140 26372
rect -204 26228 -140 26292
rect -204 26148 -140 26212
rect -204 26068 -140 26132
rect -204 25988 -140 26052
rect -204 25908 -140 25972
rect -204 25828 -140 25892
rect -204 25748 -140 25812
rect -204 25668 -140 25732
rect -204 25588 -140 25652
rect -204 25508 -140 25572
rect -204 25428 -140 25492
rect -204 25348 -140 25412
rect -204 25268 -140 25332
rect -204 25188 -140 25252
rect -204 25108 -140 25172
rect -204 25028 -140 25092
rect -204 24948 -140 25012
rect -204 24868 -140 24932
rect -204 24788 -140 24852
rect -204 24708 -140 24772
rect -204 24628 -140 24692
rect -204 24548 -140 24612
rect -204 24468 -140 24532
rect -204 24388 -140 24452
rect -204 24308 -140 24372
rect -204 24228 -140 24292
rect -204 24148 -140 24212
rect -204 24068 -140 24132
rect -204 23988 -140 24052
rect -204 23908 -140 23972
rect -204 23828 -140 23892
rect -204 23748 -140 23812
rect -204 23668 -140 23732
rect -204 23588 -140 23652
rect -204 23508 -140 23572
rect -204 23428 -140 23492
rect -204 23348 -140 23412
rect -204 23268 -140 23332
rect -204 23188 -140 23252
rect -204 23108 -140 23172
rect -204 23028 -140 23092
rect -204 22948 -140 23012
rect -204 22868 -140 22932
rect -204 22788 -140 22852
rect -204 22708 -140 22772
rect -204 22628 -140 22692
rect -204 22548 -140 22612
rect -204 22468 -140 22532
rect -204 22388 -140 22452
rect -204 22308 -140 22372
rect -204 22228 -140 22292
rect -204 22148 -140 22212
rect -204 22068 -140 22132
rect -204 21988 -140 22052
rect -204 21908 -140 21972
rect -204 21828 -140 21892
rect -204 21748 -140 21812
rect -204 21668 -140 21732
rect -204 21588 -140 21652
rect -204 21508 -140 21572
rect -204 21428 -140 21492
rect 5408 26388 5472 26452
rect 5408 26308 5472 26372
rect 5408 26228 5472 26292
rect 5408 26148 5472 26212
rect 5408 26068 5472 26132
rect 5408 25988 5472 26052
rect 5408 25908 5472 25972
rect 5408 25828 5472 25892
rect 5408 25748 5472 25812
rect 5408 25668 5472 25732
rect 5408 25588 5472 25652
rect 5408 25508 5472 25572
rect 5408 25428 5472 25492
rect 5408 25348 5472 25412
rect 5408 25268 5472 25332
rect 5408 25188 5472 25252
rect 5408 25108 5472 25172
rect 5408 25028 5472 25092
rect 5408 24948 5472 25012
rect 5408 24868 5472 24932
rect 5408 24788 5472 24852
rect 5408 24708 5472 24772
rect 5408 24628 5472 24692
rect 5408 24548 5472 24612
rect 5408 24468 5472 24532
rect 5408 24388 5472 24452
rect 5408 24308 5472 24372
rect 5408 24228 5472 24292
rect 5408 24148 5472 24212
rect 5408 24068 5472 24132
rect 5408 23988 5472 24052
rect 5408 23908 5472 23972
rect 5408 23828 5472 23892
rect 5408 23748 5472 23812
rect 5408 23668 5472 23732
rect 5408 23588 5472 23652
rect 5408 23508 5472 23572
rect 5408 23428 5472 23492
rect 5408 23348 5472 23412
rect 5408 23268 5472 23332
rect 5408 23188 5472 23252
rect 5408 23108 5472 23172
rect 5408 23028 5472 23092
rect 5408 22948 5472 23012
rect 5408 22868 5472 22932
rect 5408 22788 5472 22852
rect 5408 22708 5472 22772
rect 5408 22628 5472 22692
rect 5408 22548 5472 22612
rect 5408 22468 5472 22532
rect 5408 22388 5472 22452
rect 5408 22308 5472 22372
rect 5408 22228 5472 22292
rect 5408 22148 5472 22212
rect 5408 22068 5472 22132
rect 5408 21988 5472 22052
rect 5408 21908 5472 21972
rect 5408 21828 5472 21892
rect 5408 21748 5472 21812
rect 5408 21668 5472 21732
rect 5408 21588 5472 21652
rect 5408 21508 5472 21572
rect 5408 21428 5472 21492
rect 11020 26388 11084 26452
rect 11020 26308 11084 26372
rect 11020 26228 11084 26292
rect 11020 26148 11084 26212
rect 11020 26068 11084 26132
rect 11020 25988 11084 26052
rect 11020 25908 11084 25972
rect 11020 25828 11084 25892
rect 11020 25748 11084 25812
rect 11020 25668 11084 25732
rect 11020 25588 11084 25652
rect 11020 25508 11084 25572
rect 11020 25428 11084 25492
rect 11020 25348 11084 25412
rect 11020 25268 11084 25332
rect 11020 25188 11084 25252
rect 11020 25108 11084 25172
rect 11020 25028 11084 25092
rect 11020 24948 11084 25012
rect 11020 24868 11084 24932
rect 11020 24788 11084 24852
rect 11020 24708 11084 24772
rect 11020 24628 11084 24692
rect 11020 24548 11084 24612
rect 11020 24468 11084 24532
rect 11020 24388 11084 24452
rect 11020 24308 11084 24372
rect 11020 24228 11084 24292
rect 11020 24148 11084 24212
rect 11020 24068 11084 24132
rect 11020 23988 11084 24052
rect 11020 23908 11084 23972
rect 11020 23828 11084 23892
rect 11020 23748 11084 23812
rect 11020 23668 11084 23732
rect 11020 23588 11084 23652
rect 11020 23508 11084 23572
rect 11020 23428 11084 23492
rect 11020 23348 11084 23412
rect 11020 23268 11084 23332
rect 11020 23188 11084 23252
rect 11020 23108 11084 23172
rect 11020 23028 11084 23092
rect 11020 22948 11084 23012
rect 11020 22868 11084 22932
rect 11020 22788 11084 22852
rect 11020 22708 11084 22772
rect 11020 22628 11084 22692
rect 11020 22548 11084 22612
rect 11020 22468 11084 22532
rect 11020 22388 11084 22452
rect 11020 22308 11084 22372
rect 11020 22228 11084 22292
rect 11020 22148 11084 22212
rect 11020 22068 11084 22132
rect 11020 21988 11084 22052
rect 11020 21908 11084 21972
rect 11020 21828 11084 21892
rect 11020 21748 11084 21812
rect 11020 21668 11084 21732
rect 11020 21588 11084 21652
rect 11020 21508 11084 21572
rect 11020 21428 11084 21492
rect 16632 26388 16696 26452
rect 16632 26308 16696 26372
rect 16632 26228 16696 26292
rect 16632 26148 16696 26212
rect 16632 26068 16696 26132
rect 16632 25988 16696 26052
rect 16632 25908 16696 25972
rect 16632 25828 16696 25892
rect 16632 25748 16696 25812
rect 16632 25668 16696 25732
rect 16632 25588 16696 25652
rect 16632 25508 16696 25572
rect 16632 25428 16696 25492
rect 16632 25348 16696 25412
rect 16632 25268 16696 25332
rect 16632 25188 16696 25252
rect 16632 25108 16696 25172
rect 16632 25028 16696 25092
rect 16632 24948 16696 25012
rect 16632 24868 16696 24932
rect 16632 24788 16696 24852
rect 16632 24708 16696 24772
rect 16632 24628 16696 24692
rect 16632 24548 16696 24612
rect 16632 24468 16696 24532
rect 16632 24388 16696 24452
rect 16632 24308 16696 24372
rect 16632 24228 16696 24292
rect 16632 24148 16696 24212
rect 16632 24068 16696 24132
rect 16632 23988 16696 24052
rect 16632 23908 16696 23972
rect 16632 23828 16696 23892
rect 16632 23748 16696 23812
rect 16632 23668 16696 23732
rect 16632 23588 16696 23652
rect 16632 23508 16696 23572
rect 16632 23428 16696 23492
rect 16632 23348 16696 23412
rect 16632 23268 16696 23332
rect 16632 23188 16696 23252
rect 16632 23108 16696 23172
rect 16632 23028 16696 23092
rect 16632 22948 16696 23012
rect 16632 22868 16696 22932
rect 16632 22788 16696 22852
rect 16632 22708 16696 22772
rect 16632 22628 16696 22692
rect 16632 22548 16696 22612
rect 16632 22468 16696 22532
rect 16632 22388 16696 22452
rect 16632 22308 16696 22372
rect 16632 22228 16696 22292
rect 16632 22148 16696 22212
rect 16632 22068 16696 22132
rect 16632 21988 16696 22052
rect 16632 21908 16696 21972
rect 16632 21828 16696 21892
rect 16632 21748 16696 21812
rect 16632 21668 16696 21732
rect 16632 21588 16696 21652
rect 16632 21508 16696 21572
rect 16632 21428 16696 21492
rect 22244 26388 22308 26452
rect 22244 26308 22308 26372
rect 22244 26228 22308 26292
rect 22244 26148 22308 26212
rect 22244 26068 22308 26132
rect 22244 25988 22308 26052
rect 22244 25908 22308 25972
rect 22244 25828 22308 25892
rect 22244 25748 22308 25812
rect 22244 25668 22308 25732
rect 22244 25588 22308 25652
rect 22244 25508 22308 25572
rect 22244 25428 22308 25492
rect 22244 25348 22308 25412
rect 22244 25268 22308 25332
rect 22244 25188 22308 25252
rect 22244 25108 22308 25172
rect 22244 25028 22308 25092
rect 22244 24948 22308 25012
rect 22244 24868 22308 24932
rect 22244 24788 22308 24852
rect 22244 24708 22308 24772
rect 22244 24628 22308 24692
rect 22244 24548 22308 24612
rect 22244 24468 22308 24532
rect 22244 24388 22308 24452
rect 22244 24308 22308 24372
rect 22244 24228 22308 24292
rect 22244 24148 22308 24212
rect 22244 24068 22308 24132
rect 22244 23988 22308 24052
rect 22244 23908 22308 23972
rect 22244 23828 22308 23892
rect 22244 23748 22308 23812
rect 22244 23668 22308 23732
rect 22244 23588 22308 23652
rect 22244 23508 22308 23572
rect 22244 23428 22308 23492
rect 22244 23348 22308 23412
rect 22244 23268 22308 23332
rect 22244 23188 22308 23252
rect 22244 23108 22308 23172
rect 22244 23028 22308 23092
rect 22244 22948 22308 23012
rect 22244 22868 22308 22932
rect 22244 22788 22308 22852
rect 22244 22708 22308 22772
rect 22244 22628 22308 22692
rect 22244 22548 22308 22612
rect 22244 22468 22308 22532
rect 22244 22388 22308 22452
rect 22244 22308 22308 22372
rect 22244 22228 22308 22292
rect 22244 22148 22308 22212
rect 22244 22068 22308 22132
rect 22244 21988 22308 22052
rect 22244 21908 22308 21972
rect 22244 21828 22308 21892
rect 22244 21748 22308 21812
rect 22244 21668 22308 21732
rect 22244 21588 22308 21652
rect 22244 21508 22308 21572
rect 22244 21428 22308 21492
rect 27856 26388 27920 26452
rect 27856 26308 27920 26372
rect 27856 26228 27920 26292
rect 27856 26148 27920 26212
rect 27856 26068 27920 26132
rect 27856 25988 27920 26052
rect 27856 25908 27920 25972
rect 27856 25828 27920 25892
rect 27856 25748 27920 25812
rect 27856 25668 27920 25732
rect 27856 25588 27920 25652
rect 27856 25508 27920 25572
rect 27856 25428 27920 25492
rect 27856 25348 27920 25412
rect 27856 25268 27920 25332
rect 27856 25188 27920 25252
rect 27856 25108 27920 25172
rect 27856 25028 27920 25092
rect 27856 24948 27920 25012
rect 27856 24868 27920 24932
rect 27856 24788 27920 24852
rect 27856 24708 27920 24772
rect 27856 24628 27920 24692
rect 27856 24548 27920 24612
rect 27856 24468 27920 24532
rect 27856 24388 27920 24452
rect 27856 24308 27920 24372
rect 27856 24228 27920 24292
rect 27856 24148 27920 24212
rect 27856 24068 27920 24132
rect 27856 23988 27920 24052
rect 27856 23908 27920 23972
rect 27856 23828 27920 23892
rect 27856 23748 27920 23812
rect 27856 23668 27920 23732
rect 27856 23588 27920 23652
rect 27856 23508 27920 23572
rect 27856 23428 27920 23492
rect 27856 23348 27920 23412
rect 27856 23268 27920 23332
rect 27856 23188 27920 23252
rect 27856 23108 27920 23172
rect 27856 23028 27920 23092
rect 27856 22948 27920 23012
rect 27856 22868 27920 22932
rect 27856 22788 27920 22852
rect 27856 22708 27920 22772
rect 27856 22628 27920 22692
rect 27856 22548 27920 22612
rect 27856 22468 27920 22532
rect 27856 22388 27920 22452
rect 27856 22308 27920 22372
rect 27856 22228 27920 22292
rect 27856 22148 27920 22212
rect 27856 22068 27920 22132
rect 27856 21988 27920 22052
rect 27856 21908 27920 21972
rect 27856 21828 27920 21892
rect 27856 21748 27920 21812
rect 27856 21668 27920 21732
rect 27856 21588 27920 21652
rect 27856 21508 27920 21572
rect 27856 21428 27920 21492
rect 33468 26388 33532 26452
rect 33468 26308 33532 26372
rect 33468 26228 33532 26292
rect 33468 26148 33532 26212
rect 33468 26068 33532 26132
rect 33468 25988 33532 26052
rect 33468 25908 33532 25972
rect 33468 25828 33532 25892
rect 33468 25748 33532 25812
rect 33468 25668 33532 25732
rect 33468 25588 33532 25652
rect 33468 25508 33532 25572
rect 33468 25428 33532 25492
rect 33468 25348 33532 25412
rect 33468 25268 33532 25332
rect 33468 25188 33532 25252
rect 33468 25108 33532 25172
rect 33468 25028 33532 25092
rect 33468 24948 33532 25012
rect 33468 24868 33532 24932
rect 33468 24788 33532 24852
rect 33468 24708 33532 24772
rect 33468 24628 33532 24692
rect 33468 24548 33532 24612
rect 33468 24468 33532 24532
rect 33468 24388 33532 24452
rect 33468 24308 33532 24372
rect 33468 24228 33532 24292
rect 33468 24148 33532 24212
rect 33468 24068 33532 24132
rect 33468 23988 33532 24052
rect 33468 23908 33532 23972
rect 33468 23828 33532 23892
rect 33468 23748 33532 23812
rect 33468 23668 33532 23732
rect 33468 23588 33532 23652
rect 33468 23508 33532 23572
rect 33468 23428 33532 23492
rect 33468 23348 33532 23412
rect 33468 23268 33532 23332
rect 33468 23188 33532 23252
rect 33468 23108 33532 23172
rect 33468 23028 33532 23092
rect 33468 22948 33532 23012
rect 33468 22868 33532 22932
rect 33468 22788 33532 22852
rect 33468 22708 33532 22772
rect 33468 22628 33532 22692
rect 33468 22548 33532 22612
rect 33468 22468 33532 22532
rect 33468 22388 33532 22452
rect 33468 22308 33532 22372
rect 33468 22228 33532 22292
rect 33468 22148 33532 22212
rect 33468 22068 33532 22132
rect 33468 21988 33532 22052
rect 33468 21908 33532 21972
rect 33468 21828 33532 21892
rect 33468 21748 33532 21812
rect 33468 21668 33532 21732
rect 33468 21588 33532 21652
rect 33468 21508 33532 21572
rect 33468 21428 33532 21492
rect 39080 26388 39144 26452
rect 39080 26308 39144 26372
rect 39080 26228 39144 26292
rect 39080 26148 39144 26212
rect 39080 26068 39144 26132
rect 39080 25988 39144 26052
rect 39080 25908 39144 25972
rect 39080 25828 39144 25892
rect 39080 25748 39144 25812
rect 39080 25668 39144 25732
rect 39080 25588 39144 25652
rect 39080 25508 39144 25572
rect 39080 25428 39144 25492
rect 39080 25348 39144 25412
rect 39080 25268 39144 25332
rect 39080 25188 39144 25252
rect 39080 25108 39144 25172
rect 39080 25028 39144 25092
rect 39080 24948 39144 25012
rect 39080 24868 39144 24932
rect 39080 24788 39144 24852
rect 39080 24708 39144 24772
rect 39080 24628 39144 24692
rect 39080 24548 39144 24612
rect 39080 24468 39144 24532
rect 39080 24388 39144 24452
rect 39080 24308 39144 24372
rect 39080 24228 39144 24292
rect 39080 24148 39144 24212
rect 39080 24068 39144 24132
rect 39080 23988 39144 24052
rect 39080 23908 39144 23972
rect 39080 23828 39144 23892
rect 39080 23748 39144 23812
rect 39080 23668 39144 23732
rect 39080 23588 39144 23652
rect 39080 23508 39144 23572
rect 39080 23428 39144 23492
rect 39080 23348 39144 23412
rect 39080 23268 39144 23332
rect 39080 23188 39144 23252
rect 39080 23108 39144 23172
rect 39080 23028 39144 23092
rect 39080 22948 39144 23012
rect 39080 22868 39144 22932
rect 39080 22788 39144 22852
rect 39080 22708 39144 22772
rect 39080 22628 39144 22692
rect 39080 22548 39144 22612
rect 39080 22468 39144 22532
rect 39080 22388 39144 22452
rect 39080 22308 39144 22372
rect 39080 22228 39144 22292
rect 39080 22148 39144 22212
rect 39080 22068 39144 22132
rect 39080 21988 39144 22052
rect 39080 21908 39144 21972
rect 39080 21828 39144 21892
rect 39080 21748 39144 21812
rect 39080 21668 39144 21732
rect 39080 21588 39144 21652
rect 39080 21508 39144 21572
rect 39080 21428 39144 21492
rect -33876 21068 -33812 21132
rect -33876 20988 -33812 21052
rect -33876 20908 -33812 20972
rect -33876 20828 -33812 20892
rect -33876 20748 -33812 20812
rect -33876 20668 -33812 20732
rect -33876 20588 -33812 20652
rect -33876 20508 -33812 20572
rect -33876 20428 -33812 20492
rect -33876 20348 -33812 20412
rect -33876 20268 -33812 20332
rect -33876 20188 -33812 20252
rect -33876 20108 -33812 20172
rect -33876 20028 -33812 20092
rect -33876 19948 -33812 20012
rect -33876 19868 -33812 19932
rect -33876 19788 -33812 19852
rect -33876 19708 -33812 19772
rect -33876 19628 -33812 19692
rect -33876 19548 -33812 19612
rect -33876 19468 -33812 19532
rect -33876 19388 -33812 19452
rect -33876 19308 -33812 19372
rect -33876 19228 -33812 19292
rect -33876 19148 -33812 19212
rect -33876 19068 -33812 19132
rect -33876 18988 -33812 19052
rect -33876 18908 -33812 18972
rect -33876 18828 -33812 18892
rect -33876 18748 -33812 18812
rect -33876 18668 -33812 18732
rect -33876 18588 -33812 18652
rect -33876 18508 -33812 18572
rect -33876 18428 -33812 18492
rect -33876 18348 -33812 18412
rect -33876 18268 -33812 18332
rect -33876 18188 -33812 18252
rect -33876 18108 -33812 18172
rect -33876 18028 -33812 18092
rect -33876 17948 -33812 18012
rect -33876 17868 -33812 17932
rect -33876 17788 -33812 17852
rect -33876 17708 -33812 17772
rect -33876 17628 -33812 17692
rect -33876 17548 -33812 17612
rect -33876 17468 -33812 17532
rect -33876 17388 -33812 17452
rect -33876 17308 -33812 17372
rect -33876 17228 -33812 17292
rect -33876 17148 -33812 17212
rect -33876 17068 -33812 17132
rect -33876 16988 -33812 17052
rect -33876 16908 -33812 16972
rect -33876 16828 -33812 16892
rect -33876 16748 -33812 16812
rect -33876 16668 -33812 16732
rect -33876 16588 -33812 16652
rect -33876 16508 -33812 16572
rect -33876 16428 -33812 16492
rect -33876 16348 -33812 16412
rect -33876 16268 -33812 16332
rect -33876 16188 -33812 16252
rect -33876 16108 -33812 16172
rect -28264 21068 -28200 21132
rect -28264 20988 -28200 21052
rect -28264 20908 -28200 20972
rect -28264 20828 -28200 20892
rect -28264 20748 -28200 20812
rect -28264 20668 -28200 20732
rect -28264 20588 -28200 20652
rect -28264 20508 -28200 20572
rect -28264 20428 -28200 20492
rect -28264 20348 -28200 20412
rect -28264 20268 -28200 20332
rect -28264 20188 -28200 20252
rect -28264 20108 -28200 20172
rect -28264 20028 -28200 20092
rect -28264 19948 -28200 20012
rect -28264 19868 -28200 19932
rect -28264 19788 -28200 19852
rect -28264 19708 -28200 19772
rect -28264 19628 -28200 19692
rect -28264 19548 -28200 19612
rect -28264 19468 -28200 19532
rect -28264 19388 -28200 19452
rect -28264 19308 -28200 19372
rect -28264 19228 -28200 19292
rect -28264 19148 -28200 19212
rect -28264 19068 -28200 19132
rect -28264 18988 -28200 19052
rect -28264 18908 -28200 18972
rect -28264 18828 -28200 18892
rect -28264 18748 -28200 18812
rect -28264 18668 -28200 18732
rect -28264 18588 -28200 18652
rect -28264 18508 -28200 18572
rect -28264 18428 -28200 18492
rect -28264 18348 -28200 18412
rect -28264 18268 -28200 18332
rect -28264 18188 -28200 18252
rect -28264 18108 -28200 18172
rect -28264 18028 -28200 18092
rect -28264 17948 -28200 18012
rect -28264 17868 -28200 17932
rect -28264 17788 -28200 17852
rect -28264 17708 -28200 17772
rect -28264 17628 -28200 17692
rect -28264 17548 -28200 17612
rect -28264 17468 -28200 17532
rect -28264 17388 -28200 17452
rect -28264 17308 -28200 17372
rect -28264 17228 -28200 17292
rect -28264 17148 -28200 17212
rect -28264 17068 -28200 17132
rect -28264 16988 -28200 17052
rect -28264 16908 -28200 16972
rect -28264 16828 -28200 16892
rect -28264 16748 -28200 16812
rect -28264 16668 -28200 16732
rect -28264 16588 -28200 16652
rect -28264 16508 -28200 16572
rect -28264 16428 -28200 16492
rect -28264 16348 -28200 16412
rect -28264 16268 -28200 16332
rect -28264 16188 -28200 16252
rect -28264 16108 -28200 16172
rect -22652 21068 -22588 21132
rect -22652 20988 -22588 21052
rect -22652 20908 -22588 20972
rect -22652 20828 -22588 20892
rect -22652 20748 -22588 20812
rect -22652 20668 -22588 20732
rect -22652 20588 -22588 20652
rect -22652 20508 -22588 20572
rect -22652 20428 -22588 20492
rect -22652 20348 -22588 20412
rect -22652 20268 -22588 20332
rect -22652 20188 -22588 20252
rect -22652 20108 -22588 20172
rect -22652 20028 -22588 20092
rect -22652 19948 -22588 20012
rect -22652 19868 -22588 19932
rect -22652 19788 -22588 19852
rect -22652 19708 -22588 19772
rect -22652 19628 -22588 19692
rect -22652 19548 -22588 19612
rect -22652 19468 -22588 19532
rect -22652 19388 -22588 19452
rect -22652 19308 -22588 19372
rect -22652 19228 -22588 19292
rect -22652 19148 -22588 19212
rect -22652 19068 -22588 19132
rect -22652 18988 -22588 19052
rect -22652 18908 -22588 18972
rect -22652 18828 -22588 18892
rect -22652 18748 -22588 18812
rect -22652 18668 -22588 18732
rect -22652 18588 -22588 18652
rect -22652 18508 -22588 18572
rect -22652 18428 -22588 18492
rect -22652 18348 -22588 18412
rect -22652 18268 -22588 18332
rect -22652 18188 -22588 18252
rect -22652 18108 -22588 18172
rect -22652 18028 -22588 18092
rect -22652 17948 -22588 18012
rect -22652 17868 -22588 17932
rect -22652 17788 -22588 17852
rect -22652 17708 -22588 17772
rect -22652 17628 -22588 17692
rect -22652 17548 -22588 17612
rect -22652 17468 -22588 17532
rect -22652 17388 -22588 17452
rect -22652 17308 -22588 17372
rect -22652 17228 -22588 17292
rect -22652 17148 -22588 17212
rect -22652 17068 -22588 17132
rect -22652 16988 -22588 17052
rect -22652 16908 -22588 16972
rect -22652 16828 -22588 16892
rect -22652 16748 -22588 16812
rect -22652 16668 -22588 16732
rect -22652 16588 -22588 16652
rect -22652 16508 -22588 16572
rect -22652 16428 -22588 16492
rect -22652 16348 -22588 16412
rect -22652 16268 -22588 16332
rect -22652 16188 -22588 16252
rect -22652 16108 -22588 16172
rect -17040 21068 -16976 21132
rect -17040 20988 -16976 21052
rect -17040 20908 -16976 20972
rect -17040 20828 -16976 20892
rect -17040 20748 -16976 20812
rect -17040 20668 -16976 20732
rect -17040 20588 -16976 20652
rect -17040 20508 -16976 20572
rect -17040 20428 -16976 20492
rect -17040 20348 -16976 20412
rect -17040 20268 -16976 20332
rect -17040 20188 -16976 20252
rect -17040 20108 -16976 20172
rect -17040 20028 -16976 20092
rect -17040 19948 -16976 20012
rect -17040 19868 -16976 19932
rect -17040 19788 -16976 19852
rect -17040 19708 -16976 19772
rect -17040 19628 -16976 19692
rect -17040 19548 -16976 19612
rect -17040 19468 -16976 19532
rect -17040 19388 -16976 19452
rect -17040 19308 -16976 19372
rect -17040 19228 -16976 19292
rect -17040 19148 -16976 19212
rect -17040 19068 -16976 19132
rect -17040 18988 -16976 19052
rect -17040 18908 -16976 18972
rect -17040 18828 -16976 18892
rect -17040 18748 -16976 18812
rect -17040 18668 -16976 18732
rect -17040 18588 -16976 18652
rect -17040 18508 -16976 18572
rect -17040 18428 -16976 18492
rect -17040 18348 -16976 18412
rect -17040 18268 -16976 18332
rect -17040 18188 -16976 18252
rect -17040 18108 -16976 18172
rect -17040 18028 -16976 18092
rect -17040 17948 -16976 18012
rect -17040 17868 -16976 17932
rect -17040 17788 -16976 17852
rect -17040 17708 -16976 17772
rect -17040 17628 -16976 17692
rect -17040 17548 -16976 17612
rect -17040 17468 -16976 17532
rect -17040 17388 -16976 17452
rect -17040 17308 -16976 17372
rect -17040 17228 -16976 17292
rect -17040 17148 -16976 17212
rect -17040 17068 -16976 17132
rect -17040 16988 -16976 17052
rect -17040 16908 -16976 16972
rect -17040 16828 -16976 16892
rect -17040 16748 -16976 16812
rect -17040 16668 -16976 16732
rect -17040 16588 -16976 16652
rect -17040 16508 -16976 16572
rect -17040 16428 -16976 16492
rect -17040 16348 -16976 16412
rect -17040 16268 -16976 16332
rect -17040 16188 -16976 16252
rect -17040 16108 -16976 16172
rect -11428 21068 -11364 21132
rect -11428 20988 -11364 21052
rect -11428 20908 -11364 20972
rect -11428 20828 -11364 20892
rect -11428 20748 -11364 20812
rect -11428 20668 -11364 20732
rect -11428 20588 -11364 20652
rect -11428 20508 -11364 20572
rect -11428 20428 -11364 20492
rect -11428 20348 -11364 20412
rect -11428 20268 -11364 20332
rect -11428 20188 -11364 20252
rect -11428 20108 -11364 20172
rect -11428 20028 -11364 20092
rect -11428 19948 -11364 20012
rect -11428 19868 -11364 19932
rect -11428 19788 -11364 19852
rect -11428 19708 -11364 19772
rect -11428 19628 -11364 19692
rect -11428 19548 -11364 19612
rect -11428 19468 -11364 19532
rect -11428 19388 -11364 19452
rect -11428 19308 -11364 19372
rect -11428 19228 -11364 19292
rect -11428 19148 -11364 19212
rect -11428 19068 -11364 19132
rect -11428 18988 -11364 19052
rect -11428 18908 -11364 18972
rect -11428 18828 -11364 18892
rect -11428 18748 -11364 18812
rect -11428 18668 -11364 18732
rect -11428 18588 -11364 18652
rect -11428 18508 -11364 18572
rect -11428 18428 -11364 18492
rect -11428 18348 -11364 18412
rect -11428 18268 -11364 18332
rect -11428 18188 -11364 18252
rect -11428 18108 -11364 18172
rect -11428 18028 -11364 18092
rect -11428 17948 -11364 18012
rect -11428 17868 -11364 17932
rect -11428 17788 -11364 17852
rect -11428 17708 -11364 17772
rect -11428 17628 -11364 17692
rect -11428 17548 -11364 17612
rect -11428 17468 -11364 17532
rect -11428 17388 -11364 17452
rect -11428 17308 -11364 17372
rect -11428 17228 -11364 17292
rect -11428 17148 -11364 17212
rect -11428 17068 -11364 17132
rect -11428 16988 -11364 17052
rect -11428 16908 -11364 16972
rect -11428 16828 -11364 16892
rect -11428 16748 -11364 16812
rect -11428 16668 -11364 16732
rect -11428 16588 -11364 16652
rect -11428 16508 -11364 16572
rect -11428 16428 -11364 16492
rect -11428 16348 -11364 16412
rect -11428 16268 -11364 16332
rect -11428 16188 -11364 16252
rect -11428 16108 -11364 16172
rect -5816 21068 -5752 21132
rect -5816 20988 -5752 21052
rect -5816 20908 -5752 20972
rect -5816 20828 -5752 20892
rect -5816 20748 -5752 20812
rect -5816 20668 -5752 20732
rect -5816 20588 -5752 20652
rect -5816 20508 -5752 20572
rect -5816 20428 -5752 20492
rect -5816 20348 -5752 20412
rect -5816 20268 -5752 20332
rect -5816 20188 -5752 20252
rect -5816 20108 -5752 20172
rect -5816 20028 -5752 20092
rect -5816 19948 -5752 20012
rect -5816 19868 -5752 19932
rect -5816 19788 -5752 19852
rect -5816 19708 -5752 19772
rect -5816 19628 -5752 19692
rect -5816 19548 -5752 19612
rect -5816 19468 -5752 19532
rect -5816 19388 -5752 19452
rect -5816 19308 -5752 19372
rect -5816 19228 -5752 19292
rect -5816 19148 -5752 19212
rect -5816 19068 -5752 19132
rect -5816 18988 -5752 19052
rect -5816 18908 -5752 18972
rect -5816 18828 -5752 18892
rect -5816 18748 -5752 18812
rect -5816 18668 -5752 18732
rect -5816 18588 -5752 18652
rect -5816 18508 -5752 18572
rect -5816 18428 -5752 18492
rect -5816 18348 -5752 18412
rect -5816 18268 -5752 18332
rect -5816 18188 -5752 18252
rect -5816 18108 -5752 18172
rect -5816 18028 -5752 18092
rect -5816 17948 -5752 18012
rect -5816 17868 -5752 17932
rect -5816 17788 -5752 17852
rect -5816 17708 -5752 17772
rect -5816 17628 -5752 17692
rect -5816 17548 -5752 17612
rect -5816 17468 -5752 17532
rect -5816 17388 -5752 17452
rect -5816 17308 -5752 17372
rect -5816 17228 -5752 17292
rect -5816 17148 -5752 17212
rect -5816 17068 -5752 17132
rect -5816 16988 -5752 17052
rect -5816 16908 -5752 16972
rect -5816 16828 -5752 16892
rect -5816 16748 -5752 16812
rect -5816 16668 -5752 16732
rect -5816 16588 -5752 16652
rect -5816 16508 -5752 16572
rect -5816 16428 -5752 16492
rect -5816 16348 -5752 16412
rect -5816 16268 -5752 16332
rect -5816 16188 -5752 16252
rect -5816 16108 -5752 16172
rect -204 21068 -140 21132
rect -204 20988 -140 21052
rect -204 20908 -140 20972
rect -204 20828 -140 20892
rect -204 20748 -140 20812
rect -204 20668 -140 20732
rect -204 20588 -140 20652
rect -204 20508 -140 20572
rect -204 20428 -140 20492
rect -204 20348 -140 20412
rect -204 20268 -140 20332
rect -204 20188 -140 20252
rect -204 20108 -140 20172
rect -204 20028 -140 20092
rect -204 19948 -140 20012
rect -204 19868 -140 19932
rect -204 19788 -140 19852
rect -204 19708 -140 19772
rect -204 19628 -140 19692
rect -204 19548 -140 19612
rect -204 19468 -140 19532
rect -204 19388 -140 19452
rect -204 19308 -140 19372
rect -204 19228 -140 19292
rect -204 19148 -140 19212
rect -204 19068 -140 19132
rect -204 18988 -140 19052
rect -204 18908 -140 18972
rect -204 18828 -140 18892
rect -204 18748 -140 18812
rect -204 18668 -140 18732
rect -204 18588 -140 18652
rect -204 18508 -140 18572
rect -204 18428 -140 18492
rect -204 18348 -140 18412
rect -204 18268 -140 18332
rect -204 18188 -140 18252
rect -204 18108 -140 18172
rect -204 18028 -140 18092
rect -204 17948 -140 18012
rect -204 17868 -140 17932
rect -204 17788 -140 17852
rect -204 17708 -140 17772
rect -204 17628 -140 17692
rect -204 17548 -140 17612
rect -204 17468 -140 17532
rect -204 17388 -140 17452
rect -204 17308 -140 17372
rect -204 17228 -140 17292
rect -204 17148 -140 17212
rect -204 17068 -140 17132
rect -204 16988 -140 17052
rect -204 16908 -140 16972
rect -204 16828 -140 16892
rect -204 16748 -140 16812
rect -204 16668 -140 16732
rect -204 16588 -140 16652
rect -204 16508 -140 16572
rect -204 16428 -140 16492
rect -204 16348 -140 16412
rect -204 16268 -140 16332
rect -204 16188 -140 16252
rect -204 16108 -140 16172
rect 5408 21068 5472 21132
rect 5408 20988 5472 21052
rect 5408 20908 5472 20972
rect 5408 20828 5472 20892
rect 5408 20748 5472 20812
rect 5408 20668 5472 20732
rect 5408 20588 5472 20652
rect 5408 20508 5472 20572
rect 5408 20428 5472 20492
rect 5408 20348 5472 20412
rect 5408 20268 5472 20332
rect 5408 20188 5472 20252
rect 5408 20108 5472 20172
rect 5408 20028 5472 20092
rect 5408 19948 5472 20012
rect 5408 19868 5472 19932
rect 5408 19788 5472 19852
rect 5408 19708 5472 19772
rect 5408 19628 5472 19692
rect 5408 19548 5472 19612
rect 5408 19468 5472 19532
rect 5408 19388 5472 19452
rect 5408 19308 5472 19372
rect 5408 19228 5472 19292
rect 5408 19148 5472 19212
rect 5408 19068 5472 19132
rect 5408 18988 5472 19052
rect 5408 18908 5472 18972
rect 5408 18828 5472 18892
rect 5408 18748 5472 18812
rect 5408 18668 5472 18732
rect 5408 18588 5472 18652
rect 5408 18508 5472 18572
rect 5408 18428 5472 18492
rect 5408 18348 5472 18412
rect 5408 18268 5472 18332
rect 5408 18188 5472 18252
rect 5408 18108 5472 18172
rect 5408 18028 5472 18092
rect 5408 17948 5472 18012
rect 5408 17868 5472 17932
rect 5408 17788 5472 17852
rect 5408 17708 5472 17772
rect 5408 17628 5472 17692
rect 5408 17548 5472 17612
rect 5408 17468 5472 17532
rect 5408 17388 5472 17452
rect 5408 17308 5472 17372
rect 5408 17228 5472 17292
rect 5408 17148 5472 17212
rect 5408 17068 5472 17132
rect 5408 16988 5472 17052
rect 5408 16908 5472 16972
rect 5408 16828 5472 16892
rect 5408 16748 5472 16812
rect 5408 16668 5472 16732
rect 5408 16588 5472 16652
rect 5408 16508 5472 16572
rect 5408 16428 5472 16492
rect 5408 16348 5472 16412
rect 5408 16268 5472 16332
rect 5408 16188 5472 16252
rect 5408 16108 5472 16172
rect 11020 21068 11084 21132
rect 11020 20988 11084 21052
rect 11020 20908 11084 20972
rect 11020 20828 11084 20892
rect 11020 20748 11084 20812
rect 11020 20668 11084 20732
rect 11020 20588 11084 20652
rect 11020 20508 11084 20572
rect 11020 20428 11084 20492
rect 11020 20348 11084 20412
rect 11020 20268 11084 20332
rect 11020 20188 11084 20252
rect 11020 20108 11084 20172
rect 11020 20028 11084 20092
rect 11020 19948 11084 20012
rect 11020 19868 11084 19932
rect 11020 19788 11084 19852
rect 11020 19708 11084 19772
rect 11020 19628 11084 19692
rect 11020 19548 11084 19612
rect 11020 19468 11084 19532
rect 11020 19388 11084 19452
rect 11020 19308 11084 19372
rect 11020 19228 11084 19292
rect 11020 19148 11084 19212
rect 11020 19068 11084 19132
rect 11020 18988 11084 19052
rect 11020 18908 11084 18972
rect 11020 18828 11084 18892
rect 11020 18748 11084 18812
rect 11020 18668 11084 18732
rect 11020 18588 11084 18652
rect 11020 18508 11084 18572
rect 11020 18428 11084 18492
rect 11020 18348 11084 18412
rect 11020 18268 11084 18332
rect 11020 18188 11084 18252
rect 11020 18108 11084 18172
rect 11020 18028 11084 18092
rect 11020 17948 11084 18012
rect 11020 17868 11084 17932
rect 11020 17788 11084 17852
rect 11020 17708 11084 17772
rect 11020 17628 11084 17692
rect 11020 17548 11084 17612
rect 11020 17468 11084 17532
rect 11020 17388 11084 17452
rect 11020 17308 11084 17372
rect 11020 17228 11084 17292
rect 11020 17148 11084 17212
rect 11020 17068 11084 17132
rect 11020 16988 11084 17052
rect 11020 16908 11084 16972
rect 11020 16828 11084 16892
rect 11020 16748 11084 16812
rect 11020 16668 11084 16732
rect 11020 16588 11084 16652
rect 11020 16508 11084 16572
rect 11020 16428 11084 16492
rect 11020 16348 11084 16412
rect 11020 16268 11084 16332
rect 11020 16188 11084 16252
rect 11020 16108 11084 16172
rect 16632 21068 16696 21132
rect 16632 20988 16696 21052
rect 16632 20908 16696 20972
rect 16632 20828 16696 20892
rect 16632 20748 16696 20812
rect 16632 20668 16696 20732
rect 16632 20588 16696 20652
rect 16632 20508 16696 20572
rect 16632 20428 16696 20492
rect 16632 20348 16696 20412
rect 16632 20268 16696 20332
rect 16632 20188 16696 20252
rect 16632 20108 16696 20172
rect 16632 20028 16696 20092
rect 16632 19948 16696 20012
rect 16632 19868 16696 19932
rect 16632 19788 16696 19852
rect 16632 19708 16696 19772
rect 16632 19628 16696 19692
rect 16632 19548 16696 19612
rect 16632 19468 16696 19532
rect 16632 19388 16696 19452
rect 16632 19308 16696 19372
rect 16632 19228 16696 19292
rect 16632 19148 16696 19212
rect 16632 19068 16696 19132
rect 16632 18988 16696 19052
rect 16632 18908 16696 18972
rect 16632 18828 16696 18892
rect 16632 18748 16696 18812
rect 16632 18668 16696 18732
rect 16632 18588 16696 18652
rect 16632 18508 16696 18572
rect 16632 18428 16696 18492
rect 16632 18348 16696 18412
rect 16632 18268 16696 18332
rect 16632 18188 16696 18252
rect 16632 18108 16696 18172
rect 16632 18028 16696 18092
rect 16632 17948 16696 18012
rect 16632 17868 16696 17932
rect 16632 17788 16696 17852
rect 16632 17708 16696 17772
rect 16632 17628 16696 17692
rect 16632 17548 16696 17612
rect 16632 17468 16696 17532
rect 16632 17388 16696 17452
rect 16632 17308 16696 17372
rect 16632 17228 16696 17292
rect 16632 17148 16696 17212
rect 16632 17068 16696 17132
rect 16632 16988 16696 17052
rect 16632 16908 16696 16972
rect 16632 16828 16696 16892
rect 16632 16748 16696 16812
rect 16632 16668 16696 16732
rect 16632 16588 16696 16652
rect 16632 16508 16696 16572
rect 16632 16428 16696 16492
rect 16632 16348 16696 16412
rect 16632 16268 16696 16332
rect 16632 16188 16696 16252
rect 16632 16108 16696 16172
rect 22244 21068 22308 21132
rect 22244 20988 22308 21052
rect 22244 20908 22308 20972
rect 22244 20828 22308 20892
rect 22244 20748 22308 20812
rect 22244 20668 22308 20732
rect 22244 20588 22308 20652
rect 22244 20508 22308 20572
rect 22244 20428 22308 20492
rect 22244 20348 22308 20412
rect 22244 20268 22308 20332
rect 22244 20188 22308 20252
rect 22244 20108 22308 20172
rect 22244 20028 22308 20092
rect 22244 19948 22308 20012
rect 22244 19868 22308 19932
rect 22244 19788 22308 19852
rect 22244 19708 22308 19772
rect 22244 19628 22308 19692
rect 22244 19548 22308 19612
rect 22244 19468 22308 19532
rect 22244 19388 22308 19452
rect 22244 19308 22308 19372
rect 22244 19228 22308 19292
rect 22244 19148 22308 19212
rect 22244 19068 22308 19132
rect 22244 18988 22308 19052
rect 22244 18908 22308 18972
rect 22244 18828 22308 18892
rect 22244 18748 22308 18812
rect 22244 18668 22308 18732
rect 22244 18588 22308 18652
rect 22244 18508 22308 18572
rect 22244 18428 22308 18492
rect 22244 18348 22308 18412
rect 22244 18268 22308 18332
rect 22244 18188 22308 18252
rect 22244 18108 22308 18172
rect 22244 18028 22308 18092
rect 22244 17948 22308 18012
rect 22244 17868 22308 17932
rect 22244 17788 22308 17852
rect 22244 17708 22308 17772
rect 22244 17628 22308 17692
rect 22244 17548 22308 17612
rect 22244 17468 22308 17532
rect 22244 17388 22308 17452
rect 22244 17308 22308 17372
rect 22244 17228 22308 17292
rect 22244 17148 22308 17212
rect 22244 17068 22308 17132
rect 22244 16988 22308 17052
rect 22244 16908 22308 16972
rect 22244 16828 22308 16892
rect 22244 16748 22308 16812
rect 22244 16668 22308 16732
rect 22244 16588 22308 16652
rect 22244 16508 22308 16572
rect 22244 16428 22308 16492
rect 22244 16348 22308 16412
rect 22244 16268 22308 16332
rect 22244 16188 22308 16252
rect 22244 16108 22308 16172
rect 27856 21068 27920 21132
rect 27856 20988 27920 21052
rect 27856 20908 27920 20972
rect 27856 20828 27920 20892
rect 27856 20748 27920 20812
rect 27856 20668 27920 20732
rect 27856 20588 27920 20652
rect 27856 20508 27920 20572
rect 27856 20428 27920 20492
rect 27856 20348 27920 20412
rect 27856 20268 27920 20332
rect 27856 20188 27920 20252
rect 27856 20108 27920 20172
rect 27856 20028 27920 20092
rect 27856 19948 27920 20012
rect 27856 19868 27920 19932
rect 27856 19788 27920 19852
rect 27856 19708 27920 19772
rect 27856 19628 27920 19692
rect 27856 19548 27920 19612
rect 27856 19468 27920 19532
rect 27856 19388 27920 19452
rect 27856 19308 27920 19372
rect 27856 19228 27920 19292
rect 27856 19148 27920 19212
rect 27856 19068 27920 19132
rect 27856 18988 27920 19052
rect 27856 18908 27920 18972
rect 27856 18828 27920 18892
rect 27856 18748 27920 18812
rect 27856 18668 27920 18732
rect 27856 18588 27920 18652
rect 27856 18508 27920 18572
rect 27856 18428 27920 18492
rect 27856 18348 27920 18412
rect 27856 18268 27920 18332
rect 27856 18188 27920 18252
rect 27856 18108 27920 18172
rect 27856 18028 27920 18092
rect 27856 17948 27920 18012
rect 27856 17868 27920 17932
rect 27856 17788 27920 17852
rect 27856 17708 27920 17772
rect 27856 17628 27920 17692
rect 27856 17548 27920 17612
rect 27856 17468 27920 17532
rect 27856 17388 27920 17452
rect 27856 17308 27920 17372
rect 27856 17228 27920 17292
rect 27856 17148 27920 17212
rect 27856 17068 27920 17132
rect 27856 16988 27920 17052
rect 27856 16908 27920 16972
rect 27856 16828 27920 16892
rect 27856 16748 27920 16812
rect 27856 16668 27920 16732
rect 27856 16588 27920 16652
rect 27856 16508 27920 16572
rect 27856 16428 27920 16492
rect 27856 16348 27920 16412
rect 27856 16268 27920 16332
rect 27856 16188 27920 16252
rect 27856 16108 27920 16172
rect 33468 21068 33532 21132
rect 33468 20988 33532 21052
rect 33468 20908 33532 20972
rect 33468 20828 33532 20892
rect 33468 20748 33532 20812
rect 33468 20668 33532 20732
rect 33468 20588 33532 20652
rect 33468 20508 33532 20572
rect 33468 20428 33532 20492
rect 33468 20348 33532 20412
rect 33468 20268 33532 20332
rect 33468 20188 33532 20252
rect 33468 20108 33532 20172
rect 33468 20028 33532 20092
rect 33468 19948 33532 20012
rect 33468 19868 33532 19932
rect 33468 19788 33532 19852
rect 33468 19708 33532 19772
rect 33468 19628 33532 19692
rect 33468 19548 33532 19612
rect 33468 19468 33532 19532
rect 33468 19388 33532 19452
rect 33468 19308 33532 19372
rect 33468 19228 33532 19292
rect 33468 19148 33532 19212
rect 33468 19068 33532 19132
rect 33468 18988 33532 19052
rect 33468 18908 33532 18972
rect 33468 18828 33532 18892
rect 33468 18748 33532 18812
rect 33468 18668 33532 18732
rect 33468 18588 33532 18652
rect 33468 18508 33532 18572
rect 33468 18428 33532 18492
rect 33468 18348 33532 18412
rect 33468 18268 33532 18332
rect 33468 18188 33532 18252
rect 33468 18108 33532 18172
rect 33468 18028 33532 18092
rect 33468 17948 33532 18012
rect 33468 17868 33532 17932
rect 33468 17788 33532 17852
rect 33468 17708 33532 17772
rect 33468 17628 33532 17692
rect 33468 17548 33532 17612
rect 33468 17468 33532 17532
rect 33468 17388 33532 17452
rect 33468 17308 33532 17372
rect 33468 17228 33532 17292
rect 33468 17148 33532 17212
rect 33468 17068 33532 17132
rect 33468 16988 33532 17052
rect 33468 16908 33532 16972
rect 33468 16828 33532 16892
rect 33468 16748 33532 16812
rect 33468 16668 33532 16732
rect 33468 16588 33532 16652
rect 33468 16508 33532 16572
rect 33468 16428 33532 16492
rect 33468 16348 33532 16412
rect 33468 16268 33532 16332
rect 33468 16188 33532 16252
rect 33468 16108 33532 16172
rect 39080 21068 39144 21132
rect 39080 20988 39144 21052
rect 39080 20908 39144 20972
rect 39080 20828 39144 20892
rect 39080 20748 39144 20812
rect 39080 20668 39144 20732
rect 39080 20588 39144 20652
rect 39080 20508 39144 20572
rect 39080 20428 39144 20492
rect 39080 20348 39144 20412
rect 39080 20268 39144 20332
rect 39080 20188 39144 20252
rect 39080 20108 39144 20172
rect 39080 20028 39144 20092
rect 39080 19948 39144 20012
rect 39080 19868 39144 19932
rect 39080 19788 39144 19852
rect 39080 19708 39144 19772
rect 39080 19628 39144 19692
rect 39080 19548 39144 19612
rect 39080 19468 39144 19532
rect 39080 19388 39144 19452
rect 39080 19308 39144 19372
rect 39080 19228 39144 19292
rect 39080 19148 39144 19212
rect 39080 19068 39144 19132
rect 39080 18988 39144 19052
rect 39080 18908 39144 18972
rect 39080 18828 39144 18892
rect 39080 18748 39144 18812
rect 39080 18668 39144 18732
rect 39080 18588 39144 18652
rect 39080 18508 39144 18572
rect 39080 18428 39144 18492
rect 39080 18348 39144 18412
rect 39080 18268 39144 18332
rect 39080 18188 39144 18252
rect 39080 18108 39144 18172
rect 39080 18028 39144 18092
rect 39080 17948 39144 18012
rect 39080 17868 39144 17932
rect 39080 17788 39144 17852
rect 39080 17708 39144 17772
rect 39080 17628 39144 17692
rect 39080 17548 39144 17612
rect 39080 17468 39144 17532
rect 39080 17388 39144 17452
rect 39080 17308 39144 17372
rect 39080 17228 39144 17292
rect 39080 17148 39144 17212
rect 39080 17068 39144 17132
rect 39080 16988 39144 17052
rect 39080 16908 39144 16972
rect 39080 16828 39144 16892
rect 39080 16748 39144 16812
rect 39080 16668 39144 16732
rect 39080 16588 39144 16652
rect 39080 16508 39144 16572
rect 39080 16428 39144 16492
rect 39080 16348 39144 16412
rect 39080 16268 39144 16332
rect 39080 16188 39144 16252
rect 39080 16108 39144 16172
rect -33876 15748 -33812 15812
rect -33876 15668 -33812 15732
rect -33876 15588 -33812 15652
rect -33876 15508 -33812 15572
rect -33876 15428 -33812 15492
rect -33876 15348 -33812 15412
rect -33876 15268 -33812 15332
rect -33876 15188 -33812 15252
rect -33876 15108 -33812 15172
rect -33876 15028 -33812 15092
rect -33876 14948 -33812 15012
rect -33876 14868 -33812 14932
rect -33876 14788 -33812 14852
rect -33876 14708 -33812 14772
rect -33876 14628 -33812 14692
rect -33876 14548 -33812 14612
rect -33876 14468 -33812 14532
rect -33876 14388 -33812 14452
rect -33876 14308 -33812 14372
rect -33876 14228 -33812 14292
rect -33876 14148 -33812 14212
rect -33876 14068 -33812 14132
rect -33876 13988 -33812 14052
rect -33876 13908 -33812 13972
rect -33876 13828 -33812 13892
rect -33876 13748 -33812 13812
rect -33876 13668 -33812 13732
rect -33876 13588 -33812 13652
rect -33876 13508 -33812 13572
rect -33876 13428 -33812 13492
rect -33876 13348 -33812 13412
rect -33876 13268 -33812 13332
rect -33876 13188 -33812 13252
rect -33876 13108 -33812 13172
rect -33876 13028 -33812 13092
rect -33876 12948 -33812 13012
rect -33876 12868 -33812 12932
rect -33876 12788 -33812 12852
rect -33876 12708 -33812 12772
rect -33876 12628 -33812 12692
rect -33876 12548 -33812 12612
rect -33876 12468 -33812 12532
rect -33876 12388 -33812 12452
rect -33876 12308 -33812 12372
rect -33876 12228 -33812 12292
rect -33876 12148 -33812 12212
rect -33876 12068 -33812 12132
rect -33876 11988 -33812 12052
rect -33876 11908 -33812 11972
rect -33876 11828 -33812 11892
rect -33876 11748 -33812 11812
rect -33876 11668 -33812 11732
rect -33876 11588 -33812 11652
rect -33876 11508 -33812 11572
rect -33876 11428 -33812 11492
rect -33876 11348 -33812 11412
rect -33876 11268 -33812 11332
rect -33876 11188 -33812 11252
rect -33876 11108 -33812 11172
rect -33876 11028 -33812 11092
rect -33876 10948 -33812 11012
rect -33876 10868 -33812 10932
rect -33876 10788 -33812 10852
rect -28264 15748 -28200 15812
rect -28264 15668 -28200 15732
rect -28264 15588 -28200 15652
rect -28264 15508 -28200 15572
rect -28264 15428 -28200 15492
rect -28264 15348 -28200 15412
rect -28264 15268 -28200 15332
rect -28264 15188 -28200 15252
rect -28264 15108 -28200 15172
rect -28264 15028 -28200 15092
rect -28264 14948 -28200 15012
rect -28264 14868 -28200 14932
rect -28264 14788 -28200 14852
rect -28264 14708 -28200 14772
rect -28264 14628 -28200 14692
rect -28264 14548 -28200 14612
rect -28264 14468 -28200 14532
rect -28264 14388 -28200 14452
rect -28264 14308 -28200 14372
rect -28264 14228 -28200 14292
rect -28264 14148 -28200 14212
rect -28264 14068 -28200 14132
rect -28264 13988 -28200 14052
rect -28264 13908 -28200 13972
rect -28264 13828 -28200 13892
rect -28264 13748 -28200 13812
rect -28264 13668 -28200 13732
rect -28264 13588 -28200 13652
rect -28264 13508 -28200 13572
rect -28264 13428 -28200 13492
rect -28264 13348 -28200 13412
rect -28264 13268 -28200 13332
rect -28264 13188 -28200 13252
rect -28264 13108 -28200 13172
rect -28264 13028 -28200 13092
rect -28264 12948 -28200 13012
rect -28264 12868 -28200 12932
rect -28264 12788 -28200 12852
rect -28264 12708 -28200 12772
rect -28264 12628 -28200 12692
rect -28264 12548 -28200 12612
rect -28264 12468 -28200 12532
rect -28264 12388 -28200 12452
rect -28264 12308 -28200 12372
rect -28264 12228 -28200 12292
rect -28264 12148 -28200 12212
rect -28264 12068 -28200 12132
rect -28264 11988 -28200 12052
rect -28264 11908 -28200 11972
rect -28264 11828 -28200 11892
rect -28264 11748 -28200 11812
rect -28264 11668 -28200 11732
rect -28264 11588 -28200 11652
rect -28264 11508 -28200 11572
rect -28264 11428 -28200 11492
rect -28264 11348 -28200 11412
rect -28264 11268 -28200 11332
rect -28264 11188 -28200 11252
rect -28264 11108 -28200 11172
rect -28264 11028 -28200 11092
rect -28264 10948 -28200 11012
rect -28264 10868 -28200 10932
rect -28264 10788 -28200 10852
rect -22652 15748 -22588 15812
rect -22652 15668 -22588 15732
rect -22652 15588 -22588 15652
rect -22652 15508 -22588 15572
rect -22652 15428 -22588 15492
rect -22652 15348 -22588 15412
rect -22652 15268 -22588 15332
rect -22652 15188 -22588 15252
rect -22652 15108 -22588 15172
rect -22652 15028 -22588 15092
rect -22652 14948 -22588 15012
rect -22652 14868 -22588 14932
rect -22652 14788 -22588 14852
rect -22652 14708 -22588 14772
rect -22652 14628 -22588 14692
rect -22652 14548 -22588 14612
rect -22652 14468 -22588 14532
rect -22652 14388 -22588 14452
rect -22652 14308 -22588 14372
rect -22652 14228 -22588 14292
rect -22652 14148 -22588 14212
rect -22652 14068 -22588 14132
rect -22652 13988 -22588 14052
rect -22652 13908 -22588 13972
rect -22652 13828 -22588 13892
rect -22652 13748 -22588 13812
rect -22652 13668 -22588 13732
rect -22652 13588 -22588 13652
rect -22652 13508 -22588 13572
rect -22652 13428 -22588 13492
rect -22652 13348 -22588 13412
rect -22652 13268 -22588 13332
rect -22652 13188 -22588 13252
rect -22652 13108 -22588 13172
rect -22652 13028 -22588 13092
rect -22652 12948 -22588 13012
rect -22652 12868 -22588 12932
rect -22652 12788 -22588 12852
rect -22652 12708 -22588 12772
rect -22652 12628 -22588 12692
rect -22652 12548 -22588 12612
rect -22652 12468 -22588 12532
rect -22652 12388 -22588 12452
rect -22652 12308 -22588 12372
rect -22652 12228 -22588 12292
rect -22652 12148 -22588 12212
rect -22652 12068 -22588 12132
rect -22652 11988 -22588 12052
rect -22652 11908 -22588 11972
rect -22652 11828 -22588 11892
rect -22652 11748 -22588 11812
rect -22652 11668 -22588 11732
rect -22652 11588 -22588 11652
rect -22652 11508 -22588 11572
rect -22652 11428 -22588 11492
rect -22652 11348 -22588 11412
rect -22652 11268 -22588 11332
rect -22652 11188 -22588 11252
rect -22652 11108 -22588 11172
rect -22652 11028 -22588 11092
rect -22652 10948 -22588 11012
rect -22652 10868 -22588 10932
rect -22652 10788 -22588 10852
rect -17040 15748 -16976 15812
rect -17040 15668 -16976 15732
rect -17040 15588 -16976 15652
rect -17040 15508 -16976 15572
rect -17040 15428 -16976 15492
rect -17040 15348 -16976 15412
rect -17040 15268 -16976 15332
rect -17040 15188 -16976 15252
rect -17040 15108 -16976 15172
rect -17040 15028 -16976 15092
rect -17040 14948 -16976 15012
rect -17040 14868 -16976 14932
rect -17040 14788 -16976 14852
rect -17040 14708 -16976 14772
rect -17040 14628 -16976 14692
rect -17040 14548 -16976 14612
rect -17040 14468 -16976 14532
rect -17040 14388 -16976 14452
rect -17040 14308 -16976 14372
rect -17040 14228 -16976 14292
rect -17040 14148 -16976 14212
rect -17040 14068 -16976 14132
rect -17040 13988 -16976 14052
rect -17040 13908 -16976 13972
rect -17040 13828 -16976 13892
rect -17040 13748 -16976 13812
rect -17040 13668 -16976 13732
rect -17040 13588 -16976 13652
rect -17040 13508 -16976 13572
rect -17040 13428 -16976 13492
rect -17040 13348 -16976 13412
rect -17040 13268 -16976 13332
rect -17040 13188 -16976 13252
rect -17040 13108 -16976 13172
rect -17040 13028 -16976 13092
rect -17040 12948 -16976 13012
rect -17040 12868 -16976 12932
rect -17040 12788 -16976 12852
rect -17040 12708 -16976 12772
rect -17040 12628 -16976 12692
rect -17040 12548 -16976 12612
rect -17040 12468 -16976 12532
rect -17040 12388 -16976 12452
rect -17040 12308 -16976 12372
rect -17040 12228 -16976 12292
rect -17040 12148 -16976 12212
rect -17040 12068 -16976 12132
rect -17040 11988 -16976 12052
rect -17040 11908 -16976 11972
rect -17040 11828 -16976 11892
rect -17040 11748 -16976 11812
rect -17040 11668 -16976 11732
rect -17040 11588 -16976 11652
rect -17040 11508 -16976 11572
rect -17040 11428 -16976 11492
rect -17040 11348 -16976 11412
rect -17040 11268 -16976 11332
rect -17040 11188 -16976 11252
rect -17040 11108 -16976 11172
rect -17040 11028 -16976 11092
rect -17040 10948 -16976 11012
rect -17040 10868 -16976 10932
rect -17040 10788 -16976 10852
rect -11428 15748 -11364 15812
rect -11428 15668 -11364 15732
rect -11428 15588 -11364 15652
rect -11428 15508 -11364 15572
rect -11428 15428 -11364 15492
rect -11428 15348 -11364 15412
rect -11428 15268 -11364 15332
rect -11428 15188 -11364 15252
rect -11428 15108 -11364 15172
rect -11428 15028 -11364 15092
rect -11428 14948 -11364 15012
rect -11428 14868 -11364 14932
rect -11428 14788 -11364 14852
rect -11428 14708 -11364 14772
rect -11428 14628 -11364 14692
rect -11428 14548 -11364 14612
rect -11428 14468 -11364 14532
rect -11428 14388 -11364 14452
rect -11428 14308 -11364 14372
rect -11428 14228 -11364 14292
rect -11428 14148 -11364 14212
rect -11428 14068 -11364 14132
rect -11428 13988 -11364 14052
rect -11428 13908 -11364 13972
rect -11428 13828 -11364 13892
rect -11428 13748 -11364 13812
rect -11428 13668 -11364 13732
rect -11428 13588 -11364 13652
rect -11428 13508 -11364 13572
rect -11428 13428 -11364 13492
rect -11428 13348 -11364 13412
rect -11428 13268 -11364 13332
rect -11428 13188 -11364 13252
rect -11428 13108 -11364 13172
rect -11428 13028 -11364 13092
rect -11428 12948 -11364 13012
rect -11428 12868 -11364 12932
rect -11428 12788 -11364 12852
rect -11428 12708 -11364 12772
rect -11428 12628 -11364 12692
rect -11428 12548 -11364 12612
rect -11428 12468 -11364 12532
rect -11428 12388 -11364 12452
rect -11428 12308 -11364 12372
rect -11428 12228 -11364 12292
rect -11428 12148 -11364 12212
rect -11428 12068 -11364 12132
rect -11428 11988 -11364 12052
rect -11428 11908 -11364 11972
rect -11428 11828 -11364 11892
rect -11428 11748 -11364 11812
rect -11428 11668 -11364 11732
rect -11428 11588 -11364 11652
rect -11428 11508 -11364 11572
rect -11428 11428 -11364 11492
rect -11428 11348 -11364 11412
rect -11428 11268 -11364 11332
rect -11428 11188 -11364 11252
rect -11428 11108 -11364 11172
rect -11428 11028 -11364 11092
rect -11428 10948 -11364 11012
rect -11428 10868 -11364 10932
rect -11428 10788 -11364 10852
rect -5816 15748 -5752 15812
rect -5816 15668 -5752 15732
rect -5816 15588 -5752 15652
rect -5816 15508 -5752 15572
rect -5816 15428 -5752 15492
rect -5816 15348 -5752 15412
rect -5816 15268 -5752 15332
rect -5816 15188 -5752 15252
rect -5816 15108 -5752 15172
rect -5816 15028 -5752 15092
rect -5816 14948 -5752 15012
rect -5816 14868 -5752 14932
rect -5816 14788 -5752 14852
rect -5816 14708 -5752 14772
rect -5816 14628 -5752 14692
rect -5816 14548 -5752 14612
rect -5816 14468 -5752 14532
rect -5816 14388 -5752 14452
rect -5816 14308 -5752 14372
rect -5816 14228 -5752 14292
rect -5816 14148 -5752 14212
rect -5816 14068 -5752 14132
rect -5816 13988 -5752 14052
rect -5816 13908 -5752 13972
rect -5816 13828 -5752 13892
rect -5816 13748 -5752 13812
rect -5816 13668 -5752 13732
rect -5816 13588 -5752 13652
rect -5816 13508 -5752 13572
rect -5816 13428 -5752 13492
rect -5816 13348 -5752 13412
rect -5816 13268 -5752 13332
rect -5816 13188 -5752 13252
rect -5816 13108 -5752 13172
rect -5816 13028 -5752 13092
rect -5816 12948 -5752 13012
rect -5816 12868 -5752 12932
rect -5816 12788 -5752 12852
rect -5816 12708 -5752 12772
rect -5816 12628 -5752 12692
rect -5816 12548 -5752 12612
rect -5816 12468 -5752 12532
rect -5816 12388 -5752 12452
rect -5816 12308 -5752 12372
rect -5816 12228 -5752 12292
rect -5816 12148 -5752 12212
rect -5816 12068 -5752 12132
rect -5816 11988 -5752 12052
rect -5816 11908 -5752 11972
rect -5816 11828 -5752 11892
rect -5816 11748 -5752 11812
rect -5816 11668 -5752 11732
rect -5816 11588 -5752 11652
rect -5816 11508 -5752 11572
rect -5816 11428 -5752 11492
rect -5816 11348 -5752 11412
rect -5816 11268 -5752 11332
rect -5816 11188 -5752 11252
rect -5816 11108 -5752 11172
rect -5816 11028 -5752 11092
rect -5816 10948 -5752 11012
rect -5816 10868 -5752 10932
rect -5816 10788 -5752 10852
rect -204 15748 -140 15812
rect -204 15668 -140 15732
rect -204 15588 -140 15652
rect -204 15508 -140 15572
rect -204 15428 -140 15492
rect -204 15348 -140 15412
rect -204 15268 -140 15332
rect -204 15188 -140 15252
rect -204 15108 -140 15172
rect -204 15028 -140 15092
rect -204 14948 -140 15012
rect -204 14868 -140 14932
rect -204 14788 -140 14852
rect -204 14708 -140 14772
rect -204 14628 -140 14692
rect -204 14548 -140 14612
rect -204 14468 -140 14532
rect -204 14388 -140 14452
rect -204 14308 -140 14372
rect -204 14228 -140 14292
rect -204 14148 -140 14212
rect -204 14068 -140 14132
rect -204 13988 -140 14052
rect -204 13908 -140 13972
rect -204 13828 -140 13892
rect -204 13748 -140 13812
rect -204 13668 -140 13732
rect -204 13588 -140 13652
rect -204 13508 -140 13572
rect -204 13428 -140 13492
rect -204 13348 -140 13412
rect -204 13268 -140 13332
rect -204 13188 -140 13252
rect -204 13108 -140 13172
rect -204 13028 -140 13092
rect -204 12948 -140 13012
rect -204 12868 -140 12932
rect -204 12788 -140 12852
rect -204 12708 -140 12772
rect -204 12628 -140 12692
rect -204 12548 -140 12612
rect -204 12468 -140 12532
rect -204 12388 -140 12452
rect -204 12308 -140 12372
rect -204 12228 -140 12292
rect -204 12148 -140 12212
rect -204 12068 -140 12132
rect -204 11988 -140 12052
rect -204 11908 -140 11972
rect -204 11828 -140 11892
rect -204 11748 -140 11812
rect -204 11668 -140 11732
rect -204 11588 -140 11652
rect -204 11508 -140 11572
rect -204 11428 -140 11492
rect -204 11348 -140 11412
rect -204 11268 -140 11332
rect -204 11188 -140 11252
rect -204 11108 -140 11172
rect -204 11028 -140 11092
rect -204 10948 -140 11012
rect -204 10868 -140 10932
rect -204 10788 -140 10852
rect 5408 15748 5472 15812
rect 5408 15668 5472 15732
rect 5408 15588 5472 15652
rect 5408 15508 5472 15572
rect 5408 15428 5472 15492
rect 5408 15348 5472 15412
rect 5408 15268 5472 15332
rect 5408 15188 5472 15252
rect 5408 15108 5472 15172
rect 5408 15028 5472 15092
rect 5408 14948 5472 15012
rect 5408 14868 5472 14932
rect 5408 14788 5472 14852
rect 5408 14708 5472 14772
rect 5408 14628 5472 14692
rect 5408 14548 5472 14612
rect 5408 14468 5472 14532
rect 5408 14388 5472 14452
rect 5408 14308 5472 14372
rect 5408 14228 5472 14292
rect 5408 14148 5472 14212
rect 5408 14068 5472 14132
rect 5408 13988 5472 14052
rect 5408 13908 5472 13972
rect 5408 13828 5472 13892
rect 5408 13748 5472 13812
rect 5408 13668 5472 13732
rect 5408 13588 5472 13652
rect 5408 13508 5472 13572
rect 5408 13428 5472 13492
rect 5408 13348 5472 13412
rect 5408 13268 5472 13332
rect 5408 13188 5472 13252
rect 5408 13108 5472 13172
rect 5408 13028 5472 13092
rect 5408 12948 5472 13012
rect 5408 12868 5472 12932
rect 5408 12788 5472 12852
rect 5408 12708 5472 12772
rect 5408 12628 5472 12692
rect 5408 12548 5472 12612
rect 5408 12468 5472 12532
rect 5408 12388 5472 12452
rect 5408 12308 5472 12372
rect 5408 12228 5472 12292
rect 5408 12148 5472 12212
rect 5408 12068 5472 12132
rect 5408 11988 5472 12052
rect 5408 11908 5472 11972
rect 5408 11828 5472 11892
rect 5408 11748 5472 11812
rect 5408 11668 5472 11732
rect 5408 11588 5472 11652
rect 5408 11508 5472 11572
rect 5408 11428 5472 11492
rect 5408 11348 5472 11412
rect 5408 11268 5472 11332
rect 5408 11188 5472 11252
rect 5408 11108 5472 11172
rect 5408 11028 5472 11092
rect 5408 10948 5472 11012
rect 5408 10868 5472 10932
rect 5408 10788 5472 10852
rect 11020 15748 11084 15812
rect 11020 15668 11084 15732
rect 11020 15588 11084 15652
rect 11020 15508 11084 15572
rect 11020 15428 11084 15492
rect 11020 15348 11084 15412
rect 11020 15268 11084 15332
rect 11020 15188 11084 15252
rect 11020 15108 11084 15172
rect 11020 15028 11084 15092
rect 11020 14948 11084 15012
rect 11020 14868 11084 14932
rect 11020 14788 11084 14852
rect 11020 14708 11084 14772
rect 11020 14628 11084 14692
rect 11020 14548 11084 14612
rect 11020 14468 11084 14532
rect 11020 14388 11084 14452
rect 11020 14308 11084 14372
rect 11020 14228 11084 14292
rect 11020 14148 11084 14212
rect 11020 14068 11084 14132
rect 11020 13988 11084 14052
rect 11020 13908 11084 13972
rect 11020 13828 11084 13892
rect 11020 13748 11084 13812
rect 11020 13668 11084 13732
rect 11020 13588 11084 13652
rect 11020 13508 11084 13572
rect 11020 13428 11084 13492
rect 11020 13348 11084 13412
rect 11020 13268 11084 13332
rect 11020 13188 11084 13252
rect 11020 13108 11084 13172
rect 11020 13028 11084 13092
rect 11020 12948 11084 13012
rect 11020 12868 11084 12932
rect 11020 12788 11084 12852
rect 11020 12708 11084 12772
rect 11020 12628 11084 12692
rect 11020 12548 11084 12612
rect 11020 12468 11084 12532
rect 11020 12388 11084 12452
rect 11020 12308 11084 12372
rect 11020 12228 11084 12292
rect 11020 12148 11084 12212
rect 11020 12068 11084 12132
rect 11020 11988 11084 12052
rect 11020 11908 11084 11972
rect 11020 11828 11084 11892
rect 11020 11748 11084 11812
rect 11020 11668 11084 11732
rect 11020 11588 11084 11652
rect 11020 11508 11084 11572
rect 11020 11428 11084 11492
rect 11020 11348 11084 11412
rect 11020 11268 11084 11332
rect 11020 11188 11084 11252
rect 11020 11108 11084 11172
rect 11020 11028 11084 11092
rect 11020 10948 11084 11012
rect 11020 10868 11084 10932
rect 11020 10788 11084 10852
rect 16632 15748 16696 15812
rect 16632 15668 16696 15732
rect 16632 15588 16696 15652
rect 16632 15508 16696 15572
rect 16632 15428 16696 15492
rect 16632 15348 16696 15412
rect 16632 15268 16696 15332
rect 16632 15188 16696 15252
rect 16632 15108 16696 15172
rect 16632 15028 16696 15092
rect 16632 14948 16696 15012
rect 16632 14868 16696 14932
rect 16632 14788 16696 14852
rect 16632 14708 16696 14772
rect 16632 14628 16696 14692
rect 16632 14548 16696 14612
rect 16632 14468 16696 14532
rect 16632 14388 16696 14452
rect 16632 14308 16696 14372
rect 16632 14228 16696 14292
rect 16632 14148 16696 14212
rect 16632 14068 16696 14132
rect 16632 13988 16696 14052
rect 16632 13908 16696 13972
rect 16632 13828 16696 13892
rect 16632 13748 16696 13812
rect 16632 13668 16696 13732
rect 16632 13588 16696 13652
rect 16632 13508 16696 13572
rect 16632 13428 16696 13492
rect 16632 13348 16696 13412
rect 16632 13268 16696 13332
rect 16632 13188 16696 13252
rect 16632 13108 16696 13172
rect 16632 13028 16696 13092
rect 16632 12948 16696 13012
rect 16632 12868 16696 12932
rect 16632 12788 16696 12852
rect 16632 12708 16696 12772
rect 16632 12628 16696 12692
rect 16632 12548 16696 12612
rect 16632 12468 16696 12532
rect 16632 12388 16696 12452
rect 16632 12308 16696 12372
rect 16632 12228 16696 12292
rect 16632 12148 16696 12212
rect 16632 12068 16696 12132
rect 16632 11988 16696 12052
rect 16632 11908 16696 11972
rect 16632 11828 16696 11892
rect 16632 11748 16696 11812
rect 16632 11668 16696 11732
rect 16632 11588 16696 11652
rect 16632 11508 16696 11572
rect 16632 11428 16696 11492
rect 16632 11348 16696 11412
rect 16632 11268 16696 11332
rect 16632 11188 16696 11252
rect 16632 11108 16696 11172
rect 16632 11028 16696 11092
rect 16632 10948 16696 11012
rect 16632 10868 16696 10932
rect 16632 10788 16696 10852
rect 22244 15748 22308 15812
rect 22244 15668 22308 15732
rect 22244 15588 22308 15652
rect 22244 15508 22308 15572
rect 22244 15428 22308 15492
rect 22244 15348 22308 15412
rect 22244 15268 22308 15332
rect 22244 15188 22308 15252
rect 22244 15108 22308 15172
rect 22244 15028 22308 15092
rect 22244 14948 22308 15012
rect 22244 14868 22308 14932
rect 22244 14788 22308 14852
rect 22244 14708 22308 14772
rect 22244 14628 22308 14692
rect 22244 14548 22308 14612
rect 22244 14468 22308 14532
rect 22244 14388 22308 14452
rect 22244 14308 22308 14372
rect 22244 14228 22308 14292
rect 22244 14148 22308 14212
rect 22244 14068 22308 14132
rect 22244 13988 22308 14052
rect 22244 13908 22308 13972
rect 22244 13828 22308 13892
rect 22244 13748 22308 13812
rect 22244 13668 22308 13732
rect 22244 13588 22308 13652
rect 22244 13508 22308 13572
rect 22244 13428 22308 13492
rect 22244 13348 22308 13412
rect 22244 13268 22308 13332
rect 22244 13188 22308 13252
rect 22244 13108 22308 13172
rect 22244 13028 22308 13092
rect 22244 12948 22308 13012
rect 22244 12868 22308 12932
rect 22244 12788 22308 12852
rect 22244 12708 22308 12772
rect 22244 12628 22308 12692
rect 22244 12548 22308 12612
rect 22244 12468 22308 12532
rect 22244 12388 22308 12452
rect 22244 12308 22308 12372
rect 22244 12228 22308 12292
rect 22244 12148 22308 12212
rect 22244 12068 22308 12132
rect 22244 11988 22308 12052
rect 22244 11908 22308 11972
rect 22244 11828 22308 11892
rect 22244 11748 22308 11812
rect 22244 11668 22308 11732
rect 22244 11588 22308 11652
rect 22244 11508 22308 11572
rect 22244 11428 22308 11492
rect 22244 11348 22308 11412
rect 22244 11268 22308 11332
rect 22244 11188 22308 11252
rect 22244 11108 22308 11172
rect 22244 11028 22308 11092
rect 22244 10948 22308 11012
rect 22244 10868 22308 10932
rect 22244 10788 22308 10852
rect 27856 15748 27920 15812
rect 27856 15668 27920 15732
rect 27856 15588 27920 15652
rect 27856 15508 27920 15572
rect 27856 15428 27920 15492
rect 27856 15348 27920 15412
rect 27856 15268 27920 15332
rect 27856 15188 27920 15252
rect 27856 15108 27920 15172
rect 27856 15028 27920 15092
rect 27856 14948 27920 15012
rect 27856 14868 27920 14932
rect 27856 14788 27920 14852
rect 27856 14708 27920 14772
rect 27856 14628 27920 14692
rect 27856 14548 27920 14612
rect 27856 14468 27920 14532
rect 27856 14388 27920 14452
rect 27856 14308 27920 14372
rect 27856 14228 27920 14292
rect 27856 14148 27920 14212
rect 27856 14068 27920 14132
rect 27856 13988 27920 14052
rect 27856 13908 27920 13972
rect 27856 13828 27920 13892
rect 27856 13748 27920 13812
rect 27856 13668 27920 13732
rect 27856 13588 27920 13652
rect 27856 13508 27920 13572
rect 27856 13428 27920 13492
rect 27856 13348 27920 13412
rect 27856 13268 27920 13332
rect 27856 13188 27920 13252
rect 27856 13108 27920 13172
rect 27856 13028 27920 13092
rect 27856 12948 27920 13012
rect 27856 12868 27920 12932
rect 27856 12788 27920 12852
rect 27856 12708 27920 12772
rect 27856 12628 27920 12692
rect 27856 12548 27920 12612
rect 27856 12468 27920 12532
rect 27856 12388 27920 12452
rect 27856 12308 27920 12372
rect 27856 12228 27920 12292
rect 27856 12148 27920 12212
rect 27856 12068 27920 12132
rect 27856 11988 27920 12052
rect 27856 11908 27920 11972
rect 27856 11828 27920 11892
rect 27856 11748 27920 11812
rect 27856 11668 27920 11732
rect 27856 11588 27920 11652
rect 27856 11508 27920 11572
rect 27856 11428 27920 11492
rect 27856 11348 27920 11412
rect 27856 11268 27920 11332
rect 27856 11188 27920 11252
rect 27856 11108 27920 11172
rect 27856 11028 27920 11092
rect 27856 10948 27920 11012
rect 27856 10868 27920 10932
rect 27856 10788 27920 10852
rect 33468 15748 33532 15812
rect 33468 15668 33532 15732
rect 33468 15588 33532 15652
rect 33468 15508 33532 15572
rect 33468 15428 33532 15492
rect 33468 15348 33532 15412
rect 33468 15268 33532 15332
rect 33468 15188 33532 15252
rect 33468 15108 33532 15172
rect 33468 15028 33532 15092
rect 33468 14948 33532 15012
rect 33468 14868 33532 14932
rect 33468 14788 33532 14852
rect 33468 14708 33532 14772
rect 33468 14628 33532 14692
rect 33468 14548 33532 14612
rect 33468 14468 33532 14532
rect 33468 14388 33532 14452
rect 33468 14308 33532 14372
rect 33468 14228 33532 14292
rect 33468 14148 33532 14212
rect 33468 14068 33532 14132
rect 33468 13988 33532 14052
rect 33468 13908 33532 13972
rect 33468 13828 33532 13892
rect 33468 13748 33532 13812
rect 33468 13668 33532 13732
rect 33468 13588 33532 13652
rect 33468 13508 33532 13572
rect 33468 13428 33532 13492
rect 33468 13348 33532 13412
rect 33468 13268 33532 13332
rect 33468 13188 33532 13252
rect 33468 13108 33532 13172
rect 33468 13028 33532 13092
rect 33468 12948 33532 13012
rect 33468 12868 33532 12932
rect 33468 12788 33532 12852
rect 33468 12708 33532 12772
rect 33468 12628 33532 12692
rect 33468 12548 33532 12612
rect 33468 12468 33532 12532
rect 33468 12388 33532 12452
rect 33468 12308 33532 12372
rect 33468 12228 33532 12292
rect 33468 12148 33532 12212
rect 33468 12068 33532 12132
rect 33468 11988 33532 12052
rect 33468 11908 33532 11972
rect 33468 11828 33532 11892
rect 33468 11748 33532 11812
rect 33468 11668 33532 11732
rect 33468 11588 33532 11652
rect 33468 11508 33532 11572
rect 33468 11428 33532 11492
rect 33468 11348 33532 11412
rect 33468 11268 33532 11332
rect 33468 11188 33532 11252
rect 33468 11108 33532 11172
rect 33468 11028 33532 11092
rect 33468 10948 33532 11012
rect 33468 10868 33532 10932
rect 33468 10788 33532 10852
rect 39080 15748 39144 15812
rect 39080 15668 39144 15732
rect 39080 15588 39144 15652
rect 39080 15508 39144 15572
rect 39080 15428 39144 15492
rect 39080 15348 39144 15412
rect 39080 15268 39144 15332
rect 39080 15188 39144 15252
rect 39080 15108 39144 15172
rect 39080 15028 39144 15092
rect 39080 14948 39144 15012
rect 39080 14868 39144 14932
rect 39080 14788 39144 14852
rect 39080 14708 39144 14772
rect 39080 14628 39144 14692
rect 39080 14548 39144 14612
rect 39080 14468 39144 14532
rect 39080 14388 39144 14452
rect 39080 14308 39144 14372
rect 39080 14228 39144 14292
rect 39080 14148 39144 14212
rect 39080 14068 39144 14132
rect 39080 13988 39144 14052
rect 39080 13908 39144 13972
rect 39080 13828 39144 13892
rect 39080 13748 39144 13812
rect 39080 13668 39144 13732
rect 39080 13588 39144 13652
rect 39080 13508 39144 13572
rect 39080 13428 39144 13492
rect 39080 13348 39144 13412
rect 39080 13268 39144 13332
rect 39080 13188 39144 13252
rect 39080 13108 39144 13172
rect 39080 13028 39144 13092
rect 39080 12948 39144 13012
rect 39080 12868 39144 12932
rect 39080 12788 39144 12852
rect 39080 12708 39144 12772
rect 39080 12628 39144 12692
rect 39080 12548 39144 12612
rect 39080 12468 39144 12532
rect 39080 12388 39144 12452
rect 39080 12308 39144 12372
rect 39080 12228 39144 12292
rect 39080 12148 39144 12212
rect 39080 12068 39144 12132
rect 39080 11988 39144 12052
rect 39080 11908 39144 11972
rect 39080 11828 39144 11892
rect 39080 11748 39144 11812
rect 39080 11668 39144 11732
rect 39080 11588 39144 11652
rect 39080 11508 39144 11572
rect 39080 11428 39144 11492
rect 39080 11348 39144 11412
rect 39080 11268 39144 11332
rect 39080 11188 39144 11252
rect 39080 11108 39144 11172
rect 39080 11028 39144 11092
rect 39080 10948 39144 11012
rect 39080 10868 39144 10932
rect 39080 10788 39144 10852
rect -33876 10428 -33812 10492
rect -33876 10348 -33812 10412
rect -33876 10268 -33812 10332
rect -33876 10188 -33812 10252
rect -33876 10108 -33812 10172
rect -33876 10028 -33812 10092
rect -33876 9948 -33812 10012
rect -33876 9868 -33812 9932
rect -33876 9788 -33812 9852
rect -33876 9708 -33812 9772
rect -33876 9628 -33812 9692
rect -33876 9548 -33812 9612
rect -33876 9468 -33812 9532
rect -33876 9388 -33812 9452
rect -33876 9308 -33812 9372
rect -33876 9228 -33812 9292
rect -33876 9148 -33812 9212
rect -33876 9068 -33812 9132
rect -33876 8988 -33812 9052
rect -33876 8908 -33812 8972
rect -33876 8828 -33812 8892
rect -33876 8748 -33812 8812
rect -33876 8668 -33812 8732
rect -33876 8588 -33812 8652
rect -33876 8508 -33812 8572
rect -33876 8428 -33812 8492
rect -33876 8348 -33812 8412
rect -33876 8268 -33812 8332
rect -33876 8188 -33812 8252
rect -33876 8108 -33812 8172
rect -33876 8028 -33812 8092
rect -33876 7948 -33812 8012
rect -33876 7868 -33812 7932
rect -33876 7788 -33812 7852
rect -33876 7708 -33812 7772
rect -33876 7628 -33812 7692
rect -33876 7548 -33812 7612
rect -33876 7468 -33812 7532
rect -33876 7388 -33812 7452
rect -33876 7308 -33812 7372
rect -33876 7228 -33812 7292
rect -33876 7148 -33812 7212
rect -33876 7068 -33812 7132
rect -33876 6988 -33812 7052
rect -33876 6908 -33812 6972
rect -33876 6828 -33812 6892
rect -33876 6748 -33812 6812
rect -33876 6668 -33812 6732
rect -33876 6588 -33812 6652
rect -33876 6508 -33812 6572
rect -33876 6428 -33812 6492
rect -33876 6348 -33812 6412
rect -33876 6268 -33812 6332
rect -33876 6188 -33812 6252
rect -33876 6108 -33812 6172
rect -33876 6028 -33812 6092
rect -33876 5948 -33812 6012
rect -33876 5868 -33812 5932
rect -33876 5788 -33812 5852
rect -33876 5708 -33812 5772
rect -33876 5628 -33812 5692
rect -33876 5548 -33812 5612
rect -33876 5468 -33812 5532
rect -28264 10428 -28200 10492
rect -28264 10348 -28200 10412
rect -28264 10268 -28200 10332
rect -28264 10188 -28200 10252
rect -28264 10108 -28200 10172
rect -28264 10028 -28200 10092
rect -28264 9948 -28200 10012
rect -28264 9868 -28200 9932
rect -28264 9788 -28200 9852
rect -28264 9708 -28200 9772
rect -28264 9628 -28200 9692
rect -28264 9548 -28200 9612
rect -28264 9468 -28200 9532
rect -28264 9388 -28200 9452
rect -28264 9308 -28200 9372
rect -28264 9228 -28200 9292
rect -28264 9148 -28200 9212
rect -28264 9068 -28200 9132
rect -28264 8988 -28200 9052
rect -28264 8908 -28200 8972
rect -28264 8828 -28200 8892
rect -28264 8748 -28200 8812
rect -28264 8668 -28200 8732
rect -28264 8588 -28200 8652
rect -28264 8508 -28200 8572
rect -28264 8428 -28200 8492
rect -28264 8348 -28200 8412
rect -28264 8268 -28200 8332
rect -28264 8188 -28200 8252
rect -28264 8108 -28200 8172
rect -28264 8028 -28200 8092
rect -28264 7948 -28200 8012
rect -28264 7868 -28200 7932
rect -28264 7788 -28200 7852
rect -28264 7708 -28200 7772
rect -28264 7628 -28200 7692
rect -28264 7548 -28200 7612
rect -28264 7468 -28200 7532
rect -28264 7388 -28200 7452
rect -28264 7308 -28200 7372
rect -28264 7228 -28200 7292
rect -28264 7148 -28200 7212
rect -28264 7068 -28200 7132
rect -28264 6988 -28200 7052
rect -28264 6908 -28200 6972
rect -28264 6828 -28200 6892
rect -28264 6748 -28200 6812
rect -28264 6668 -28200 6732
rect -28264 6588 -28200 6652
rect -28264 6508 -28200 6572
rect -28264 6428 -28200 6492
rect -28264 6348 -28200 6412
rect -28264 6268 -28200 6332
rect -28264 6188 -28200 6252
rect -28264 6108 -28200 6172
rect -28264 6028 -28200 6092
rect -28264 5948 -28200 6012
rect -28264 5868 -28200 5932
rect -28264 5788 -28200 5852
rect -28264 5708 -28200 5772
rect -28264 5628 -28200 5692
rect -28264 5548 -28200 5612
rect -28264 5468 -28200 5532
rect -22652 10428 -22588 10492
rect -22652 10348 -22588 10412
rect -22652 10268 -22588 10332
rect -22652 10188 -22588 10252
rect -22652 10108 -22588 10172
rect -22652 10028 -22588 10092
rect -22652 9948 -22588 10012
rect -22652 9868 -22588 9932
rect -22652 9788 -22588 9852
rect -22652 9708 -22588 9772
rect -22652 9628 -22588 9692
rect -22652 9548 -22588 9612
rect -22652 9468 -22588 9532
rect -22652 9388 -22588 9452
rect -22652 9308 -22588 9372
rect -22652 9228 -22588 9292
rect -22652 9148 -22588 9212
rect -22652 9068 -22588 9132
rect -22652 8988 -22588 9052
rect -22652 8908 -22588 8972
rect -22652 8828 -22588 8892
rect -22652 8748 -22588 8812
rect -22652 8668 -22588 8732
rect -22652 8588 -22588 8652
rect -22652 8508 -22588 8572
rect -22652 8428 -22588 8492
rect -22652 8348 -22588 8412
rect -22652 8268 -22588 8332
rect -22652 8188 -22588 8252
rect -22652 8108 -22588 8172
rect -22652 8028 -22588 8092
rect -22652 7948 -22588 8012
rect -22652 7868 -22588 7932
rect -22652 7788 -22588 7852
rect -22652 7708 -22588 7772
rect -22652 7628 -22588 7692
rect -22652 7548 -22588 7612
rect -22652 7468 -22588 7532
rect -22652 7388 -22588 7452
rect -22652 7308 -22588 7372
rect -22652 7228 -22588 7292
rect -22652 7148 -22588 7212
rect -22652 7068 -22588 7132
rect -22652 6988 -22588 7052
rect -22652 6908 -22588 6972
rect -22652 6828 -22588 6892
rect -22652 6748 -22588 6812
rect -22652 6668 -22588 6732
rect -22652 6588 -22588 6652
rect -22652 6508 -22588 6572
rect -22652 6428 -22588 6492
rect -22652 6348 -22588 6412
rect -22652 6268 -22588 6332
rect -22652 6188 -22588 6252
rect -22652 6108 -22588 6172
rect -22652 6028 -22588 6092
rect -22652 5948 -22588 6012
rect -22652 5868 -22588 5932
rect -22652 5788 -22588 5852
rect -22652 5708 -22588 5772
rect -22652 5628 -22588 5692
rect -22652 5548 -22588 5612
rect -22652 5468 -22588 5532
rect -17040 10428 -16976 10492
rect -17040 10348 -16976 10412
rect -17040 10268 -16976 10332
rect -17040 10188 -16976 10252
rect -17040 10108 -16976 10172
rect -17040 10028 -16976 10092
rect -17040 9948 -16976 10012
rect -17040 9868 -16976 9932
rect -17040 9788 -16976 9852
rect -17040 9708 -16976 9772
rect -17040 9628 -16976 9692
rect -17040 9548 -16976 9612
rect -17040 9468 -16976 9532
rect -17040 9388 -16976 9452
rect -17040 9308 -16976 9372
rect -17040 9228 -16976 9292
rect -17040 9148 -16976 9212
rect -17040 9068 -16976 9132
rect -17040 8988 -16976 9052
rect -17040 8908 -16976 8972
rect -17040 8828 -16976 8892
rect -17040 8748 -16976 8812
rect -17040 8668 -16976 8732
rect -17040 8588 -16976 8652
rect -17040 8508 -16976 8572
rect -17040 8428 -16976 8492
rect -17040 8348 -16976 8412
rect -17040 8268 -16976 8332
rect -17040 8188 -16976 8252
rect -17040 8108 -16976 8172
rect -17040 8028 -16976 8092
rect -17040 7948 -16976 8012
rect -17040 7868 -16976 7932
rect -17040 7788 -16976 7852
rect -17040 7708 -16976 7772
rect -17040 7628 -16976 7692
rect -17040 7548 -16976 7612
rect -17040 7468 -16976 7532
rect -17040 7388 -16976 7452
rect -17040 7308 -16976 7372
rect -17040 7228 -16976 7292
rect -17040 7148 -16976 7212
rect -17040 7068 -16976 7132
rect -17040 6988 -16976 7052
rect -17040 6908 -16976 6972
rect -17040 6828 -16976 6892
rect -17040 6748 -16976 6812
rect -17040 6668 -16976 6732
rect -17040 6588 -16976 6652
rect -17040 6508 -16976 6572
rect -17040 6428 -16976 6492
rect -17040 6348 -16976 6412
rect -17040 6268 -16976 6332
rect -17040 6188 -16976 6252
rect -17040 6108 -16976 6172
rect -17040 6028 -16976 6092
rect -17040 5948 -16976 6012
rect -17040 5868 -16976 5932
rect -17040 5788 -16976 5852
rect -17040 5708 -16976 5772
rect -17040 5628 -16976 5692
rect -17040 5548 -16976 5612
rect -17040 5468 -16976 5532
rect -11428 10428 -11364 10492
rect -11428 10348 -11364 10412
rect -11428 10268 -11364 10332
rect -11428 10188 -11364 10252
rect -11428 10108 -11364 10172
rect -11428 10028 -11364 10092
rect -11428 9948 -11364 10012
rect -11428 9868 -11364 9932
rect -11428 9788 -11364 9852
rect -11428 9708 -11364 9772
rect -11428 9628 -11364 9692
rect -11428 9548 -11364 9612
rect -11428 9468 -11364 9532
rect -11428 9388 -11364 9452
rect -11428 9308 -11364 9372
rect -11428 9228 -11364 9292
rect -11428 9148 -11364 9212
rect -11428 9068 -11364 9132
rect -11428 8988 -11364 9052
rect -11428 8908 -11364 8972
rect -11428 8828 -11364 8892
rect -11428 8748 -11364 8812
rect -11428 8668 -11364 8732
rect -11428 8588 -11364 8652
rect -11428 8508 -11364 8572
rect -11428 8428 -11364 8492
rect -11428 8348 -11364 8412
rect -11428 8268 -11364 8332
rect -11428 8188 -11364 8252
rect -11428 8108 -11364 8172
rect -11428 8028 -11364 8092
rect -11428 7948 -11364 8012
rect -11428 7868 -11364 7932
rect -11428 7788 -11364 7852
rect -11428 7708 -11364 7772
rect -11428 7628 -11364 7692
rect -11428 7548 -11364 7612
rect -11428 7468 -11364 7532
rect -11428 7388 -11364 7452
rect -11428 7308 -11364 7372
rect -11428 7228 -11364 7292
rect -11428 7148 -11364 7212
rect -11428 7068 -11364 7132
rect -11428 6988 -11364 7052
rect -11428 6908 -11364 6972
rect -11428 6828 -11364 6892
rect -11428 6748 -11364 6812
rect -11428 6668 -11364 6732
rect -11428 6588 -11364 6652
rect -11428 6508 -11364 6572
rect -11428 6428 -11364 6492
rect -11428 6348 -11364 6412
rect -11428 6268 -11364 6332
rect -11428 6188 -11364 6252
rect -11428 6108 -11364 6172
rect -11428 6028 -11364 6092
rect -11428 5948 -11364 6012
rect -11428 5868 -11364 5932
rect -11428 5788 -11364 5852
rect -11428 5708 -11364 5772
rect -11428 5628 -11364 5692
rect -11428 5548 -11364 5612
rect -11428 5468 -11364 5532
rect -5816 10428 -5752 10492
rect -5816 10348 -5752 10412
rect -5816 10268 -5752 10332
rect -5816 10188 -5752 10252
rect -5816 10108 -5752 10172
rect -5816 10028 -5752 10092
rect -5816 9948 -5752 10012
rect -5816 9868 -5752 9932
rect -5816 9788 -5752 9852
rect -5816 9708 -5752 9772
rect -5816 9628 -5752 9692
rect -5816 9548 -5752 9612
rect -5816 9468 -5752 9532
rect -5816 9388 -5752 9452
rect -5816 9308 -5752 9372
rect -5816 9228 -5752 9292
rect -5816 9148 -5752 9212
rect -5816 9068 -5752 9132
rect -5816 8988 -5752 9052
rect -5816 8908 -5752 8972
rect -5816 8828 -5752 8892
rect -5816 8748 -5752 8812
rect -5816 8668 -5752 8732
rect -5816 8588 -5752 8652
rect -5816 8508 -5752 8572
rect -5816 8428 -5752 8492
rect -5816 8348 -5752 8412
rect -5816 8268 -5752 8332
rect -5816 8188 -5752 8252
rect -5816 8108 -5752 8172
rect -5816 8028 -5752 8092
rect -5816 7948 -5752 8012
rect -5816 7868 -5752 7932
rect -5816 7788 -5752 7852
rect -5816 7708 -5752 7772
rect -5816 7628 -5752 7692
rect -5816 7548 -5752 7612
rect -5816 7468 -5752 7532
rect -5816 7388 -5752 7452
rect -5816 7308 -5752 7372
rect -5816 7228 -5752 7292
rect -5816 7148 -5752 7212
rect -5816 7068 -5752 7132
rect -5816 6988 -5752 7052
rect -5816 6908 -5752 6972
rect -5816 6828 -5752 6892
rect -5816 6748 -5752 6812
rect -5816 6668 -5752 6732
rect -5816 6588 -5752 6652
rect -5816 6508 -5752 6572
rect -5816 6428 -5752 6492
rect -5816 6348 -5752 6412
rect -5816 6268 -5752 6332
rect -5816 6188 -5752 6252
rect -5816 6108 -5752 6172
rect -5816 6028 -5752 6092
rect -5816 5948 -5752 6012
rect -5816 5868 -5752 5932
rect -5816 5788 -5752 5852
rect -5816 5708 -5752 5772
rect -5816 5628 -5752 5692
rect -5816 5548 -5752 5612
rect -5816 5468 -5752 5532
rect -204 10428 -140 10492
rect -204 10348 -140 10412
rect -204 10268 -140 10332
rect -204 10188 -140 10252
rect -204 10108 -140 10172
rect -204 10028 -140 10092
rect -204 9948 -140 10012
rect -204 9868 -140 9932
rect -204 9788 -140 9852
rect -204 9708 -140 9772
rect -204 9628 -140 9692
rect -204 9548 -140 9612
rect -204 9468 -140 9532
rect -204 9388 -140 9452
rect -204 9308 -140 9372
rect -204 9228 -140 9292
rect -204 9148 -140 9212
rect -204 9068 -140 9132
rect -204 8988 -140 9052
rect -204 8908 -140 8972
rect -204 8828 -140 8892
rect -204 8748 -140 8812
rect -204 8668 -140 8732
rect -204 8588 -140 8652
rect -204 8508 -140 8572
rect -204 8428 -140 8492
rect -204 8348 -140 8412
rect -204 8268 -140 8332
rect -204 8188 -140 8252
rect -204 8108 -140 8172
rect -204 8028 -140 8092
rect -204 7948 -140 8012
rect -204 7868 -140 7932
rect -204 7788 -140 7852
rect -204 7708 -140 7772
rect -204 7628 -140 7692
rect -204 7548 -140 7612
rect -204 7468 -140 7532
rect -204 7388 -140 7452
rect -204 7308 -140 7372
rect -204 7228 -140 7292
rect -204 7148 -140 7212
rect -204 7068 -140 7132
rect -204 6988 -140 7052
rect -204 6908 -140 6972
rect -204 6828 -140 6892
rect -204 6748 -140 6812
rect -204 6668 -140 6732
rect -204 6588 -140 6652
rect -204 6508 -140 6572
rect -204 6428 -140 6492
rect -204 6348 -140 6412
rect -204 6268 -140 6332
rect -204 6188 -140 6252
rect -204 6108 -140 6172
rect -204 6028 -140 6092
rect -204 5948 -140 6012
rect -204 5868 -140 5932
rect -204 5788 -140 5852
rect -204 5708 -140 5772
rect -204 5628 -140 5692
rect -204 5548 -140 5612
rect -204 5468 -140 5532
rect 5408 10428 5472 10492
rect 5408 10348 5472 10412
rect 5408 10268 5472 10332
rect 5408 10188 5472 10252
rect 5408 10108 5472 10172
rect 5408 10028 5472 10092
rect 5408 9948 5472 10012
rect 5408 9868 5472 9932
rect 5408 9788 5472 9852
rect 5408 9708 5472 9772
rect 5408 9628 5472 9692
rect 5408 9548 5472 9612
rect 5408 9468 5472 9532
rect 5408 9388 5472 9452
rect 5408 9308 5472 9372
rect 5408 9228 5472 9292
rect 5408 9148 5472 9212
rect 5408 9068 5472 9132
rect 5408 8988 5472 9052
rect 5408 8908 5472 8972
rect 5408 8828 5472 8892
rect 5408 8748 5472 8812
rect 5408 8668 5472 8732
rect 5408 8588 5472 8652
rect 5408 8508 5472 8572
rect 5408 8428 5472 8492
rect 5408 8348 5472 8412
rect 5408 8268 5472 8332
rect 5408 8188 5472 8252
rect 5408 8108 5472 8172
rect 5408 8028 5472 8092
rect 5408 7948 5472 8012
rect 5408 7868 5472 7932
rect 5408 7788 5472 7852
rect 5408 7708 5472 7772
rect 5408 7628 5472 7692
rect 5408 7548 5472 7612
rect 5408 7468 5472 7532
rect 5408 7388 5472 7452
rect 5408 7308 5472 7372
rect 5408 7228 5472 7292
rect 5408 7148 5472 7212
rect 5408 7068 5472 7132
rect 5408 6988 5472 7052
rect 5408 6908 5472 6972
rect 5408 6828 5472 6892
rect 5408 6748 5472 6812
rect 5408 6668 5472 6732
rect 5408 6588 5472 6652
rect 5408 6508 5472 6572
rect 5408 6428 5472 6492
rect 5408 6348 5472 6412
rect 5408 6268 5472 6332
rect 5408 6188 5472 6252
rect 5408 6108 5472 6172
rect 5408 6028 5472 6092
rect 5408 5948 5472 6012
rect 5408 5868 5472 5932
rect 5408 5788 5472 5852
rect 5408 5708 5472 5772
rect 5408 5628 5472 5692
rect 5408 5548 5472 5612
rect 5408 5468 5472 5532
rect 11020 10428 11084 10492
rect 11020 10348 11084 10412
rect 11020 10268 11084 10332
rect 11020 10188 11084 10252
rect 11020 10108 11084 10172
rect 11020 10028 11084 10092
rect 11020 9948 11084 10012
rect 11020 9868 11084 9932
rect 11020 9788 11084 9852
rect 11020 9708 11084 9772
rect 11020 9628 11084 9692
rect 11020 9548 11084 9612
rect 11020 9468 11084 9532
rect 11020 9388 11084 9452
rect 11020 9308 11084 9372
rect 11020 9228 11084 9292
rect 11020 9148 11084 9212
rect 11020 9068 11084 9132
rect 11020 8988 11084 9052
rect 11020 8908 11084 8972
rect 11020 8828 11084 8892
rect 11020 8748 11084 8812
rect 11020 8668 11084 8732
rect 11020 8588 11084 8652
rect 11020 8508 11084 8572
rect 11020 8428 11084 8492
rect 11020 8348 11084 8412
rect 11020 8268 11084 8332
rect 11020 8188 11084 8252
rect 11020 8108 11084 8172
rect 11020 8028 11084 8092
rect 11020 7948 11084 8012
rect 11020 7868 11084 7932
rect 11020 7788 11084 7852
rect 11020 7708 11084 7772
rect 11020 7628 11084 7692
rect 11020 7548 11084 7612
rect 11020 7468 11084 7532
rect 11020 7388 11084 7452
rect 11020 7308 11084 7372
rect 11020 7228 11084 7292
rect 11020 7148 11084 7212
rect 11020 7068 11084 7132
rect 11020 6988 11084 7052
rect 11020 6908 11084 6972
rect 11020 6828 11084 6892
rect 11020 6748 11084 6812
rect 11020 6668 11084 6732
rect 11020 6588 11084 6652
rect 11020 6508 11084 6572
rect 11020 6428 11084 6492
rect 11020 6348 11084 6412
rect 11020 6268 11084 6332
rect 11020 6188 11084 6252
rect 11020 6108 11084 6172
rect 11020 6028 11084 6092
rect 11020 5948 11084 6012
rect 11020 5868 11084 5932
rect 11020 5788 11084 5852
rect 11020 5708 11084 5772
rect 11020 5628 11084 5692
rect 11020 5548 11084 5612
rect 11020 5468 11084 5532
rect 16632 10428 16696 10492
rect 16632 10348 16696 10412
rect 16632 10268 16696 10332
rect 16632 10188 16696 10252
rect 16632 10108 16696 10172
rect 16632 10028 16696 10092
rect 16632 9948 16696 10012
rect 16632 9868 16696 9932
rect 16632 9788 16696 9852
rect 16632 9708 16696 9772
rect 16632 9628 16696 9692
rect 16632 9548 16696 9612
rect 16632 9468 16696 9532
rect 16632 9388 16696 9452
rect 16632 9308 16696 9372
rect 16632 9228 16696 9292
rect 16632 9148 16696 9212
rect 16632 9068 16696 9132
rect 16632 8988 16696 9052
rect 16632 8908 16696 8972
rect 16632 8828 16696 8892
rect 16632 8748 16696 8812
rect 16632 8668 16696 8732
rect 16632 8588 16696 8652
rect 16632 8508 16696 8572
rect 16632 8428 16696 8492
rect 16632 8348 16696 8412
rect 16632 8268 16696 8332
rect 16632 8188 16696 8252
rect 16632 8108 16696 8172
rect 16632 8028 16696 8092
rect 16632 7948 16696 8012
rect 16632 7868 16696 7932
rect 16632 7788 16696 7852
rect 16632 7708 16696 7772
rect 16632 7628 16696 7692
rect 16632 7548 16696 7612
rect 16632 7468 16696 7532
rect 16632 7388 16696 7452
rect 16632 7308 16696 7372
rect 16632 7228 16696 7292
rect 16632 7148 16696 7212
rect 16632 7068 16696 7132
rect 16632 6988 16696 7052
rect 16632 6908 16696 6972
rect 16632 6828 16696 6892
rect 16632 6748 16696 6812
rect 16632 6668 16696 6732
rect 16632 6588 16696 6652
rect 16632 6508 16696 6572
rect 16632 6428 16696 6492
rect 16632 6348 16696 6412
rect 16632 6268 16696 6332
rect 16632 6188 16696 6252
rect 16632 6108 16696 6172
rect 16632 6028 16696 6092
rect 16632 5948 16696 6012
rect 16632 5868 16696 5932
rect 16632 5788 16696 5852
rect 16632 5708 16696 5772
rect 16632 5628 16696 5692
rect 16632 5548 16696 5612
rect 16632 5468 16696 5532
rect 22244 10428 22308 10492
rect 22244 10348 22308 10412
rect 22244 10268 22308 10332
rect 22244 10188 22308 10252
rect 22244 10108 22308 10172
rect 22244 10028 22308 10092
rect 22244 9948 22308 10012
rect 22244 9868 22308 9932
rect 22244 9788 22308 9852
rect 22244 9708 22308 9772
rect 22244 9628 22308 9692
rect 22244 9548 22308 9612
rect 22244 9468 22308 9532
rect 22244 9388 22308 9452
rect 22244 9308 22308 9372
rect 22244 9228 22308 9292
rect 22244 9148 22308 9212
rect 22244 9068 22308 9132
rect 22244 8988 22308 9052
rect 22244 8908 22308 8972
rect 22244 8828 22308 8892
rect 22244 8748 22308 8812
rect 22244 8668 22308 8732
rect 22244 8588 22308 8652
rect 22244 8508 22308 8572
rect 22244 8428 22308 8492
rect 22244 8348 22308 8412
rect 22244 8268 22308 8332
rect 22244 8188 22308 8252
rect 22244 8108 22308 8172
rect 22244 8028 22308 8092
rect 22244 7948 22308 8012
rect 22244 7868 22308 7932
rect 22244 7788 22308 7852
rect 22244 7708 22308 7772
rect 22244 7628 22308 7692
rect 22244 7548 22308 7612
rect 22244 7468 22308 7532
rect 22244 7388 22308 7452
rect 22244 7308 22308 7372
rect 22244 7228 22308 7292
rect 22244 7148 22308 7212
rect 22244 7068 22308 7132
rect 22244 6988 22308 7052
rect 22244 6908 22308 6972
rect 22244 6828 22308 6892
rect 22244 6748 22308 6812
rect 22244 6668 22308 6732
rect 22244 6588 22308 6652
rect 22244 6508 22308 6572
rect 22244 6428 22308 6492
rect 22244 6348 22308 6412
rect 22244 6268 22308 6332
rect 22244 6188 22308 6252
rect 22244 6108 22308 6172
rect 22244 6028 22308 6092
rect 22244 5948 22308 6012
rect 22244 5868 22308 5932
rect 22244 5788 22308 5852
rect 22244 5708 22308 5772
rect 22244 5628 22308 5692
rect 22244 5548 22308 5612
rect 22244 5468 22308 5532
rect 27856 10428 27920 10492
rect 27856 10348 27920 10412
rect 27856 10268 27920 10332
rect 27856 10188 27920 10252
rect 27856 10108 27920 10172
rect 27856 10028 27920 10092
rect 27856 9948 27920 10012
rect 27856 9868 27920 9932
rect 27856 9788 27920 9852
rect 27856 9708 27920 9772
rect 27856 9628 27920 9692
rect 27856 9548 27920 9612
rect 27856 9468 27920 9532
rect 27856 9388 27920 9452
rect 27856 9308 27920 9372
rect 27856 9228 27920 9292
rect 27856 9148 27920 9212
rect 27856 9068 27920 9132
rect 27856 8988 27920 9052
rect 27856 8908 27920 8972
rect 27856 8828 27920 8892
rect 27856 8748 27920 8812
rect 27856 8668 27920 8732
rect 27856 8588 27920 8652
rect 27856 8508 27920 8572
rect 27856 8428 27920 8492
rect 27856 8348 27920 8412
rect 27856 8268 27920 8332
rect 27856 8188 27920 8252
rect 27856 8108 27920 8172
rect 27856 8028 27920 8092
rect 27856 7948 27920 8012
rect 27856 7868 27920 7932
rect 27856 7788 27920 7852
rect 27856 7708 27920 7772
rect 27856 7628 27920 7692
rect 27856 7548 27920 7612
rect 27856 7468 27920 7532
rect 27856 7388 27920 7452
rect 27856 7308 27920 7372
rect 27856 7228 27920 7292
rect 27856 7148 27920 7212
rect 27856 7068 27920 7132
rect 27856 6988 27920 7052
rect 27856 6908 27920 6972
rect 27856 6828 27920 6892
rect 27856 6748 27920 6812
rect 27856 6668 27920 6732
rect 27856 6588 27920 6652
rect 27856 6508 27920 6572
rect 27856 6428 27920 6492
rect 27856 6348 27920 6412
rect 27856 6268 27920 6332
rect 27856 6188 27920 6252
rect 27856 6108 27920 6172
rect 27856 6028 27920 6092
rect 27856 5948 27920 6012
rect 27856 5868 27920 5932
rect 27856 5788 27920 5852
rect 27856 5708 27920 5772
rect 27856 5628 27920 5692
rect 27856 5548 27920 5612
rect 27856 5468 27920 5532
rect 33468 10428 33532 10492
rect 33468 10348 33532 10412
rect 33468 10268 33532 10332
rect 33468 10188 33532 10252
rect 33468 10108 33532 10172
rect 33468 10028 33532 10092
rect 33468 9948 33532 10012
rect 33468 9868 33532 9932
rect 33468 9788 33532 9852
rect 33468 9708 33532 9772
rect 33468 9628 33532 9692
rect 33468 9548 33532 9612
rect 33468 9468 33532 9532
rect 33468 9388 33532 9452
rect 33468 9308 33532 9372
rect 33468 9228 33532 9292
rect 33468 9148 33532 9212
rect 33468 9068 33532 9132
rect 33468 8988 33532 9052
rect 33468 8908 33532 8972
rect 33468 8828 33532 8892
rect 33468 8748 33532 8812
rect 33468 8668 33532 8732
rect 33468 8588 33532 8652
rect 33468 8508 33532 8572
rect 33468 8428 33532 8492
rect 33468 8348 33532 8412
rect 33468 8268 33532 8332
rect 33468 8188 33532 8252
rect 33468 8108 33532 8172
rect 33468 8028 33532 8092
rect 33468 7948 33532 8012
rect 33468 7868 33532 7932
rect 33468 7788 33532 7852
rect 33468 7708 33532 7772
rect 33468 7628 33532 7692
rect 33468 7548 33532 7612
rect 33468 7468 33532 7532
rect 33468 7388 33532 7452
rect 33468 7308 33532 7372
rect 33468 7228 33532 7292
rect 33468 7148 33532 7212
rect 33468 7068 33532 7132
rect 33468 6988 33532 7052
rect 33468 6908 33532 6972
rect 33468 6828 33532 6892
rect 33468 6748 33532 6812
rect 33468 6668 33532 6732
rect 33468 6588 33532 6652
rect 33468 6508 33532 6572
rect 33468 6428 33532 6492
rect 33468 6348 33532 6412
rect 33468 6268 33532 6332
rect 33468 6188 33532 6252
rect 33468 6108 33532 6172
rect 33468 6028 33532 6092
rect 33468 5948 33532 6012
rect 33468 5868 33532 5932
rect 33468 5788 33532 5852
rect 33468 5708 33532 5772
rect 33468 5628 33532 5692
rect 33468 5548 33532 5612
rect 33468 5468 33532 5532
rect 39080 10428 39144 10492
rect 39080 10348 39144 10412
rect 39080 10268 39144 10332
rect 39080 10188 39144 10252
rect 39080 10108 39144 10172
rect 39080 10028 39144 10092
rect 39080 9948 39144 10012
rect 39080 9868 39144 9932
rect 39080 9788 39144 9852
rect 39080 9708 39144 9772
rect 39080 9628 39144 9692
rect 39080 9548 39144 9612
rect 39080 9468 39144 9532
rect 39080 9388 39144 9452
rect 39080 9308 39144 9372
rect 39080 9228 39144 9292
rect 39080 9148 39144 9212
rect 39080 9068 39144 9132
rect 39080 8988 39144 9052
rect 39080 8908 39144 8972
rect 39080 8828 39144 8892
rect 39080 8748 39144 8812
rect 39080 8668 39144 8732
rect 39080 8588 39144 8652
rect 39080 8508 39144 8572
rect 39080 8428 39144 8492
rect 39080 8348 39144 8412
rect 39080 8268 39144 8332
rect 39080 8188 39144 8252
rect 39080 8108 39144 8172
rect 39080 8028 39144 8092
rect 39080 7948 39144 8012
rect 39080 7868 39144 7932
rect 39080 7788 39144 7852
rect 39080 7708 39144 7772
rect 39080 7628 39144 7692
rect 39080 7548 39144 7612
rect 39080 7468 39144 7532
rect 39080 7388 39144 7452
rect 39080 7308 39144 7372
rect 39080 7228 39144 7292
rect 39080 7148 39144 7212
rect 39080 7068 39144 7132
rect 39080 6988 39144 7052
rect 39080 6908 39144 6972
rect 39080 6828 39144 6892
rect 39080 6748 39144 6812
rect 39080 6668 39144 6732
rect 39080 6588 39144 6652
rect 39080 6508 39144 6572
rect 39080 6428 39144 6492
rect 39080 6348 39144 6412
rect 39080 6268 39144 6332
rect 39080 6188 39144 6252
rect 39080 6108 39144 6172
rect 39080 6028 39144 6092
rect 39080 5948 39144 6012
rect 39080 5868 39144 5932
rect 39080 5788 39144 5852
rect 39080 5708 39144 5772
rect 39080 5628 39144 5692
rect 39080 5548 39144 5612
rect 39080 5468 39144 5532
rect -33876 5108 -33812 5172
rect -33876 5028 -33812 5092
rect -33876 4948 -33812 5012
rect -33876 4868 -33812 4932
rect -33876 4788 -33812 4852
rect -33876 4708 -33812 4772
rect -33876 4628 -33812 4692
rect -33876 4548 -33812 4612
rect -33876 4468 -33812 4532
rect -33876 4388 -33812 4452
rect -33876 4308 -33812 4372
rect -33876 4228 -33812 4292
rect -33876 4148 -33812 4212
rect -33876 4068 -33812 4132
rect -33876 3988 -33812 4052
rect -33876 3908 -33812 3972
rect -33876 3828 -33812 3892
rect -33876 3748 -33812 3812
rect -33876 3668 -33812 3732
rect -33876 3588 -33812 3652
rect -33876 3508 -33812 3572
rect -33876 3428 -33812 3492
rect -33876 3348 -33812 3412
rect -33876 3268 -33812 3332
rect -33876 3188 -33812 3252
rect -33876 3108 -33812 3172
rect -33876 3028 -33812 3092
rect -33876 2948 -33812 3012
rect -33876 2868 -33812 2932
rect -33876 2788 -33812 2852
rect -33876 2708 -33812 2772
rect -33876 2628 -33812 2692
rect -33876 2548 -33812 2612
rect -33876 2468 -33812 2532
rect -33876 2388 -33812 2452
rect -33876 2308 -33812 2372
rect -33876 2228 -33812 2292
rect -33876 2148 -33812 2212
rect -33876 2068 -33812 2132
rect -33876 1988 -33812 2052
rect -33876 1908 -33812 1972
rect -33876 1828 -33812 1892
rect -33876 1748 -33812 1812
rect -33876 1668 -33812 1732
rect -33876 1588 -33812 1652
rect -33876 1508 -33812 1572
rect -33876 1428 -33812 1492
rect -33876 1348 -33812 1412
rect -33876 1268 -33812 1332
rect -33876 1188 -33812 1252
rect -33876 1108 -33812 1172
rect -33876 1028 -33812 1092
rect -33876 948 -33812 1012
rect -33876 868 -33812 932
rect -33876 788 -33812 852
rect -33876 708 -33812 772
rect -33876 628 -33812 692
rect -33876 548 -33812 612
rect -33876 468 -33812 532
rect -33876 388 -33812 452
rect -33876 308 -33812 372
rect -33876 228 -33812 292
rect -33876 148 -33812 212
rect -28264 5108 -28200 5172
rect -28264 5028 -28200 5092
rect -28264 4948 -28200 5012
rect -28264 4868 -28200 4932
rect -28264 4788 -28200 4852
rect -28264 4708 -28200 4772
rect -28264 4628 -28200 4692
rect -28264 4548 -28200 4612
rect -28264 4468 -28200 4532
rect -28264 4388 -28200 4452
rect -28264 4308 -28200 4372
rect -28264 4228 -28200 4292
rect -28264 4148 -28200 4212
rect -28264 4068 -28200 4132
rect -28264 3988 -28200 4052
rect -28264 3908 -28200 3972
rect -28264 3828 -28200 3892
rect -28264 3748 -28200 3812
rect -28264 3668 -28200 3732
rect -28264 3588 -28200 3652
rect -28264 3508 -28200 3572
rect -28264 3428 -28200 3492
rect -28264 3348 -28200 3412
rect -28264 3268 -28200 3332
rect -28264 3188 -28200 3252
rect -28264 3108 -28200 3172
rect -28264 3028 -28200 3092
rect -28264 2948 -28200 3012
rect -28264 2868 -28200 2932
rect -28264 2788 -28200 2852
rect -28264 2708 -28200 2772
rect -28264 2628 -28200 2692
rect -28264 2548 -28200 2612
rect -28264 2468 -28200 2532
rect -28264 2388 -28200 2452
rect -28264 2308 -28200 2372
rect -28264 2228 -28200 2292
rect -28264 2148 -28200 2212
rect -28264 2068 -28200 2132
rect -28264 1988 -28200 2052
rect -28264 1908 -28200 1972
rect -28264 1828 -28200 1892
rect -28264 1748 -28200 1812
rect -28264 1668 -28200 1732
rect -28264 1588 -28200 1652
rect -28264 1508 -28200 1572
rect -28264 1428 -28200 1492
rect -28264 1348 -28200 1412
rect -28264 1268 -28200 1332
rect -28264 1188 -28200 1252
rect -28264 1108 -28200 1172
rect -28264 1028 -28200 1092
rect -28264 948 -28200 1012
rect -28264 868 -28200 932
rect -28264 788 -28200 852
rect -28264 708 -28200 772
rect -28264 628 -28200 692
rect -28264 548 -28200 612
rect -28264 468 -28200 532
rect -28264 388 -28200 452
rect -28264 308 -28200 372
rect -28264 228 -28200 292
rect -28264 148 -28200 212
rect -22652 5108 -22588 5172
rect -22652 5028 -22588 5092
rect -22652 4948 -22588 5012
rect -22652 4868 -22588 4932
rect -22652 4788 -22588 4852
rect -22652 4708 -22588 4772
rect -22652 4628 -22588 4692
rect -22652 4548 -22588 4612
rect -22652 4468 -22588 4532
rect -22652 4388 -22588 4452
rect -22652 4308 -22588 4372
rect -22652 4228 -22588 4292
rect -22652 4148 -22588 4212
rect -22652 4068 -22588 4132
rect -22652 3988 -22588 4052
rect -22652 3908 -22588 3972
rect -22652 3828 -22588 3892
rect -22652 3748 -22588 3812
rect -22652 3668 -22588 3732
rect -22652 3588 -22588 3652
rect -22652 3508 -22588 3572
rect -22652 3428 -22588 3492
rect -22652 3348 -22588 3412
rect -22652 3268 -22588 3332
rect -22652 3188 -22588 3252
rect -22652 3108 -22588 3172
rect -22652 3028 -22588 3092
rect -22652 2948 -22588 3012
rect -22652 2868 -22588 2932
rect -22652 2788 -22588 2852
rect -22652 2708 -22588 2772
rect -22652 2628 -22588 2692
rect -22652 2548 -22588 2612
rect -22652 2468 -22588 2532
rect -22652 2388 -22588 2452
rect -22652 2308 -22588 2372
rect -22652 2228 -22588 2292
rect -22652 2148 -22588 2212
rect -22652 2068 -22588 2132
rect -22652 1988 -22588 2052
rect -22652 1908 -22588 1972
rect -22652 1828 -22588 1892
rect -22652 1748 -22588 1812
rect -22652 1668 -22588 1732
rect -22652 1588 -22588 1652
rect -22652 1508 -22588 1572
rect -22652 1428 -22588 1492
rect -22652 1348 -22588 1412
rect -22652 1268 -22588 1332
rect -22652 1188 -22588 1252
rect -22652 1108 -22588 1172
rect -22652 1028 -22588 1092
rect -22652 948 -22588 1012
rect -22652 868 -22588 932
rect -22652 788 -22588 852
rect -22652 708 -22588 772
rect -22652 628 -22588 692
rect -22652 548 -22588 612
rect -22652 468 -22588 532
rect -22652 388 -22588 452
rect -22652 308 -22588 372
rect -22652 228 -22588 292
rect -22652 148 -22588 212
rect -17040 5108 -16976 5172
rect -17040 5028 -16976 5092
rect -17040 4948 -16976 5012
rect -17040 4868 -16976 4932
rect -17040 4788 -16976 4852
rect -17040 4708 -16976 4772
rect -17040 4628 -16976 4692
rect -17040 4548 -16976 4612
rect -17040 4468 -16976 4532
rect -17040 4388 -16976 4452
rect -17040 4308 -16976 4372
rect -17040 4228 -16976 4292
rect -17040 4148 -16976 4212
rect -17040 4068 -16976 4132
rect -17040 3988 -16976 4052
rect -17040 3908 -16976 3972
rect -17040 3828 -16976 3892
rect -17040 3748 -16976 3812
rect -17040 3668 -16976 3732
rect -17040 3588 -16976 3652
rect -17040 3508 -16976 3572
rect -17040 3428 -16976 3492
rect -17040 3348 -16976 3412
rect -17040 3268 -16976 3332
rect -17040 3188 -16976 3252
rect -17040 3108 -16976 3172
rect -17040 3028 -16976 3092
rect -17040 2948 -16976 3012
rect -17040 2868 -16976 2932
rect -17040 2788 -16976 2852
rect -17040 2708 -16976 2772
rect -17040 2628 -16976 2692
rect -17040 2548 -16976 2612
rect -17040 2468 -16976 2532
rect -17040 2388 -16976 2452
rect -17040 2308 -16976 2372
rect -17040 2228 -16976 2292
rect -17040 2148 -16976 2212
rect -17040 2068 -16976 2132
rect -17040 1988 -16976 2052
rect -17040 1908 -16976 1972
rect -17040 1828 -16976 1892
rect -17040 1748 -16976 1812
rect -17040 1668 -16976 1732
rect -17040 1588 -16976 1652
rect -17040 1508 -16976 1572
rect -17040 1428 -16976 1492
rect -17040 1348 -16976 1412
rect -17040 1268 -16976 1332
rect -17040 1188 -16976 1252
rect -17040 1108 -16976 1172
rect -17040 1028 -16976 1092
rect -17040 948 -16976 1012
rect -17040 868 -16976 932
rect -17040 788 -16976 852
rect -17040 708 -16976 772
rect -17040 628 -16976 692
rect -17040 548 -16976 612
rect -17040 468 -16976 532
rect -17040 388 -16976 452
rect -17040 308 -16976 372
rect -17040 228 -16976 292
rect -17040 148 -16976 212
rect -11428 5108 -11364 5172
rect -11428 5028 -11364 5092
rect -11428 4948 -11364 5012
rect -11428 4868 -11364 4932
rect -11428 4788 -11364 4852
rect -11428 4708 -11364 4772
rect -11428 4628 -11364 4692
rect -11428 4548 -11364 4612
rect -11428 4468 -11364 4532
rect -11428 4388 -11364 4452
rect -11428 4308 -11364 4372
rect -11428 4228 -11364 4292
rect -11428 4148 -11364 4212
rect -11428 4068 -11364 4132
rect -11428 3988 -11364 4052
rect -11428 3908 -11364 3972
rect -11428 3828 -11364 3892
rect -11428 3748 -11364 3812
rect -11428 3668 -11364 3732
rect -11428 3588 -11364 3652
rect -11428 3508 -11364 3572
rect -11428 3428 -11364 3492
rect -11428 3348 -11364 3412
rect -11428 3268 -11364 3332
rect -11428 3188 -11364 3252
rect -11428 3108 -11364 3172
rect -11428 3028 -11364 3092
rect -11428 2948 -11364 3012
rect -11428 2868 -11364 2932
rect -11428 2788 -11364 2852
rect -11428 2708 -11364 2772
rect -11428 2628 -11364 2692
rect -11428 2548 -11364 2612
rect -11428 2468 -11364 2532
rect -11428 2388 -11364 2452
rect -11428 2308 -11364 2372
rect -11428 2228 -11364 2292
rect -11428 2148 -11364 2212
rect -11428 2068 -11364 2132
rect -11428 1988 -11364 2052
rect -11428 1908 -11364 1972
rect -11428 1828 -11364 1892
rect -11428 1748 -11364 1812
rect -11428 1668 -11364 1732
rect -11428 1588 -11364 1652
rect -11428 1508 -11364 1572
rect -11428 1428 -11364 1492
rect -11428 1348 -11364 1412
rect -11428 1268 -11364 1332
rect -11428 1188 -11364 1252
rect -11428 1108 -11364 1172
rect -11428 1028 -11364 1092
rect -11428 948 -11364 1012
rect -11428 868 -11364 932
rect -11428 788 -11364 852
rect -11428 708 -11364 772
rect -11428 628 -11364 692
rect -11428 548 -11364 612
rect -11428 468 -11364 532
rect -11428 388 -11364 452
rect -11428 308 -11364 372
rect -11428 228 -11364 292
rect -11428 148 -11364 212
rect -5816 5108 -5752 5172
rect -5816 5028 -5752 5092
rect -5816 4948 -5752 5012
rect -5816 4868 -5752 4932
rect -5816 4788 -5752 4852
rect -5816 4708 -5752 4772
rect -5816 4628 -5752 4692
rect -5816 4548 -5752 4612
rect -5816 4468 -5752 4532
rect -5816 4388 -5752 4452
rect -5816 4308 -5752 4372
rect -5816 4228 -5752 4292
rect -5816 4148 -5752 4212
rect -5816 4068 -5752 4132
rect -5816 3988 -5752 4052
rect -5816 3908 -5752 3972
rect -5816 3828 -5752 3892
rect -5816 3748 -5752 3812
rect -5816 3668 -5752 3732
rect -5816 3588 -5752 3652
rect -5816 3508 -5752 3572
rect -5816 3428 -5752 3492
rect -5816 3348 -5752 3412
rect -5816 3268 -5752 3332
rect -5816 3188 -5752 3252
rect -5816 3108 -5752 3172
rect -5816 3028 -5752 3092
rect -5816 2948 -5752 3012
rect -5816 2868 -5752 2932
rect -5816 2788 -5752 2852
rect -5816 2708 -5752 2772
rect -5816 2628 -5752 2692
rect -5816 2548 -5752 2612
rect -5816 2468 -5752 2532
rect -5816 2388 -5752 2452
rect -5816 2308 -5752 2372
rect -5816 2228 -5752 2292
rect -5816 2148 -5752 2212
rect -5816 2068 -5752 2132
rect -5816 1988 -5752 2052
rect -5816 1908 -5752 1972
rect -5816 1828 -5752 1892
rect -5816 1748 -5752 1812
rect -5816 1668 -5752 1732
rect -5816 1588 -5752 1652
rect -5816 1508 -5752 1572
rect -5816 1428 -5752 1492
rect -5816 1348 -5752 1412
rect -5816 1268 -5752 1332
rect -5816 1188 -5752 1252
rect -5816 1108 -5752 1172
rect -5816 1028 -5752 1092
rect -5816 948 -5752 1012
rect -5816 868 -5752 932
rect -5816 788 -5752 852
rect -5816 708 -5752 772
rect -5816 628 -5752 692
rect -5816 548 -5752 612
rect -5816 468 -5752 532
rect -5816 388 -5752 452
rect -5816 308 -5752 372
rect -5816 228 -5752 292
rect -5816 148 -5752 212
rect -204 5108 -140 5172
rect -204 5028 -140 5092
rect -204 4948 -140 5012
rect -204 4868 -140 4932
rect -204 4788 -140 4852
rect -204 4708 -140 4772
rect -204 4628 -140 4692
rect -204 4548 -140 4612
rect -204 4468 -140 4532
rect -204 4388 -140 4452
rect -204 4308 -140 4372
rect -204 4228 -140 4292
rect -204 4148 -140 4212
rect -204 4068 -140 4132
rect -204 3988 -140 4052
rect -204 3908 -140 3972
rect -204 3828 -140 3892
rect -204 3748 -140 3812
rect -204 3668 -140 3732
rect -204 3588 -140 3652
rect -204 3508 -140 3572
rect -204 3428 -140 3492
rect -204 3348 -140 3412
rect -204 3268 -140 3332
rect -204 3188 -140 3252
rect -204 3108 -140 3172
rect -204 3028 -140 3092
rect -204 2948 -140 3012
rect -204 2868 -140 2932
rect -204 2788 -140 2852
rect -204 2708 -140 2772
rect -204 2628 -140 2692
rect -204 2548 -140 2612
rect -204 2468 -140 2532
rect -204 2388 -140 2452
rect -204 2308 -140 2372
rect -204 2228 -140 2292
rect -204 2148 -140 2212
rect -204 2068 -140 2132
rect -204 1988 -140 2052
rect -204 1908 -140 1972
rect -204 1828 -140 1892
rect -204 1748 -140 1812
rect -204 1668 -140 1732
rect -204 1588 -140 1652
rect -204 1508 -140 1572
rect -204 1428 -140 1492
rect -204 1348 -140 1412
rect -204 1268 -140 1332
rect -204 1188 -140 1252
rect -204 1108 -140 1172
rect -204 1028 -140 1092
rect -204 948 -140 1012
rect -204 868 -140 932
rect -204 788 -140 852
rect -204 708 -140 772
rect -204 628 -140 692
rect -204 548 -140 612
rect -204 468 -140 532
rect -204 388 -140 452
rect -204 308 -140 372
rect -204 228 -140 292
rect -204 148 -140 212
rect 5408 5108 5472 5172
rect 5408 5028 5472 5092
rect 5408 4948 5472 5012
rect 5408 4868 5472 4932
rect 5408 4788 5472 4852
rect 5408 4708 5472 4772
rect 5408 4628 5472 4692
rect 5408 4548 5472 4612
rect 5408 4468 5472 4532
rect 5408 4388 5472 4452
rect 5408 4308 5472 4372
rect 5408 4228 5472 4292
rect 5408 4148 5472 4212
rect 5408 4068 5472 4132
rect 5408 3988 5472 4052
rect 5408 3908 5472 3972
rect 5408 3828 5472 3892
rect 5408 3748 5472 3812
rect 5408 3668 5472 3732
rect 5408 3588 5472 3652
rect 5408 3508 5472 3572
rect 5408 3428 5472 3492
rect 5408 3348 5472 3412
rect 5408 3268 5472 3332
rect 5408 3188 5472 3252
rect 5408 3108 5472 3172
rect 5408 3028 5472 3092
rect 5408 2948 5472 3012
rect 5408 2868 5472 2932
rect 5408 2788 5472 2852
rect 5408 2708 5472 2772
rect 5408 2628 5472 2692
rect 5408 2548 5472 2612
rect 5408 2468 5472 2532
rect 5408 2388 5472 2452
rect 5408 2308 5472 2372
rect 5408 2228 5472 2292
rect 5408 2148 5472 2212
rect 5408 2068 5472 2132
rect 5408 1988 5472 2052
rect 5408 1908 5472 1972
rect 5408 1828 5472 1892
rect 5408 1748 5472 1812
rect 5408 1668 5472 1732
rect 5408 1588 5472 1652
rect 5408 1508 5472 1572
rect 5408 1428 5472 1492
rect 5408 1348 5472 1412
rect 5408 1268 5472 1332
rect 5408 1188 5472 1252
rect 5408 1108 5472 1172
rect 5408 1028 5472 1092
rect 5408 948 5472 1012
rect 5408 868 5472 932
rect 5408 788 5472 852
rect 5408 708 5472 772
rect 5408 628 5472 692
rect 5408 548 5472 612
rect 5408 468 5472 532
rect 5408 388 5472 452
rect 5408 308 5472 372
rect 5408 228 5472 292
rect 5408 148 5472 212
rect 11020 5108 11084 5172
rect 11020 5028 11084 5092
rect 11020 4948 11084 5012
rect 11020 4868 11084 4932
rect 11020 4788 11084 4852
rect 11020 4708 11084 4772
rect 11020 4628 11084 4692
rect 11020 4548 11084 4612
rect 11020 4468 11084 4532
rect 11020 4388 11084 4452
rect 11020 4308 11084 4372
rect 11020 4228 11084 4292
rect 11020 4148 11084 4212
rect 11020 4068 11084 4132
rect 11020 3988 11084 4052
rect 11020 3908 11084 3972
rect 11020 3828 11084 3892
rect 11020 3748 11084 3812
rect 11020 3668 11084 3732
rect 11020 3588 11084 3652
rect 11020 3508 11084 3572
rect 11020 3428 11084 3492
rect 11020 3348 11084 3412
rect 11020 3268 11084 3332
rect 11020 3188 11084 3252
rect 11020 3108 11084 3172
rect 11020 3028 11084 3092
rect 11020 2948 11084 3012
rect 11020 2868 11084 2932
rect 11020 2788 11084 2852
rect 11020 2708 11084 2772
rect 11020 2628 11084 2692
rect 11020 2548 11084 2612
rect 11020 2468 11084 2532
rect 11020 2388 11084 2452
rect 11020 2308 11084 2372
rect 11020 2228 11084 2292
rect 11020 2148 11084 2212
rect 11020 2068 11084 2132
rect 11020 1988 11084 2052
rect 11020 1908 11084 1972
rect 11020 1828 11084 1892
rect 11020 1748 11084 1812
rect 11020 1668 11084 1732
rect 11020 1588 11084 1652
rect 11020 1508 11084 1572
rect 11020 1428 11084 1492
rect 11020 1348 11084 1412
rect 11020 1268 11084 1332
rect 11020 1188 11084 1252
rect 11020 1108 11084 1172
rect 11020 1028 11084 1092
rect 11020 948 11084 1012
rect 11020 868 11084 932
rect 11020 788 11084 852
rect 11020 708 11084 772
rect 11020 628 11084 692
rect 11020 548 11084 612
rect 11020 468 11084 532
rect 11020 388 11084 452
rect 11020 308 11084 372
rect 11020 228 11084 292
rect 11020 148 11084 212
rect 16632 5108 16696 5172
rect 16632 5028 16696 5092
rect 16632 4948 16696 5012
rect 16632 4868 16696 4932
rect 16632 4788 16696 4852
rect 16632 4708 16696 4772
rect 16632 4628 16696 4692
rect 16632 4548 16696 4612
rect 16632 4468 16696 4532
rect 16632 4388 16696 4452
rect 16632 4308 16696 4372
rect 16632 4228 16696 4292
rect 16632 4148 16696 4212
rect 16632 4068 16696 4132
rect 16632 3988 16696 4052
rect 16632 3908 16696 3972
rect 16632 3828 16696 3892
rect 16632 3748 16696 3812
rect 16632 3668 16696 3732
rect 16632 3588 16696 3652
rect 16632 3508 16696 3572
rect 16632 3428 16696 3492
rect 16632 3348 16696 3412
rect 16632 3268 16696 3332
rect 16632 3188 16696 3252
rect 16632 3108 16696 3172
rect 16632 3028 16696 3092
rect 16632 2948 16696 3012
rect 16632 2868 16696 2932
rect 16632 2788 16696 2852
rect 16632 2708 16696 2772
rect 16632 2628 16696 2692
rect 16632 2548 16696 2612
rect 16632 2468 16696 2532
rect 16632 2388 16696 2452
rect 16632 2308 16696 2372
rect 16632 2228 16696 2292
rect 16632 2148 16696 2212
rect 16632 2068 16696 2132
rect 16632 1988 16696 2052
rect 16632 1908 16696 1972
rect 16632 1828 16696 1892
rect 16632 1748 16696 1812
rect 16632 1668 16696 1732
rect 16632 1588 16696 1652
rect 16632 1508 16696 1572
rect 16632 1428 16696 1492
rect 16632 1348 16696 1412
rect 16632 1268 16696 1332
rect 16632 1188 16696 1252
rect 16632 1108 16696 1172
rect 16632 1028 16696 1092
rect 16632 948 16696 1012
rect 16632 868 16696 932
rect 16632 788 16696 852
rect 16632 708 16696 772
rect 16632 628 16696 692
rect 16632 548 16696 612
rect 16632 468 16696 532
rect 16632 388 16696 452
rect 16632 308 16696 372
rect 16632 228 16696 292
rect 16632 148 16696 212
rect 22244 5108 22308 5172
rect 22244 5028 22308 5092
rect 22244 4948 22308 5012
rect 22244 4868 22308 4932
rect 22244 4788 22308 4852
rect 22244 4708 22308 4772
rect 22244 4628 22308 4692
rect 22244 4548 22308 4612
rect 22244 4468 22308 4532
rect 22244 4388 22308 4452
rect 22244 4308 22308 4372
rect 22244 4228 22308 4292
rect 22244 4148 22308 4212
rect 22244 4068 22308 4132
rect 22244 3988 22308 4052
rect 22244 3908 22308 3972
rect 22244 3828 22308 3892
rect 22244 3748 22308 3812
rect 22244 3668 22308 3732
rect 22244 3588 22308 3652
rect 22244 3508 22308 3572
rect 22244 3428 22308 3492
rect 22244 3348 22308 3412
rect 22244 3268 22308 3332
rect 22244 3188 22308 3252
rect 22244 3108 22308 3172
rect 22244 3028 22308 3092
rect 22244 2948 22308 3012
rect 22244 2868 22308 2932
rect 22244 2788 22308 2852
rect 22244 2708 22308 2772
rect 22244 2628 22308 2692
rect 22244 2548 22308 2612
rect 22244 2468 22308 2532
rect 22244 2388 22308 2452
rect 22244 2308 22308 2372
rect 22244 2228 22308 2292
rect 22244 2148 22308 2212
rect 22244 2068 22308 2132
rect 22244 1988 22308 2052
rect 22244 1908 22308 1972
rect 22244 1828 22308 1892
rect 22244 1748 22308 1812
rect 22244 1668 22308 1732
rect 22244 1588 22308 1652
rect 22244 1508 22308 1572
rect 22244 1428 22308 1492
rect 22244 1348 22308 1412
rect 22244 1268 22308 1332
rect 22244 1188 22308 1252
rect 22244 1108 22308 1172
rect 22244 1028 22308 1092
rect 22244 948 22308 1012
rect 22244 868 22308 932
rect 22244 788 22308 852
rect 22244 708 22308 772
rect 22244 628 22308 692
rect 22244 548 22308 612
rect 22244 468 22308 532
rect 22244 388 22308 452
rect 22244 308 22308 372
rect 22244 228 22308 292
rect 22244 148 22308 212
rect 27856 5108 27920 5172
rect 27856 5028 27920 5092
rect 27856 4948 27920 5012
rect 27856 4868 27920 4932
rect 27856 4788 27920 4852
rect 27856 4708 27920 4772
rect 27856 4628 27920 4692
rect 27856 4548 27920 4612
rect 27856 4468 27920 4532
rect 27856 4388 27920 4452
rect 27856 4308 27920 4372
rect 27856 4228 27920 4292
rect 27856 4148 27920 4212
rect 27856 4068 27920 4132
rect 27856 3988 27920 4052
rect 27856 3908 27920 3972
rect 27856 3828 27920 3892
rect 27856 3748 27920 3812
rect 27856 3668 27920 3732
rect 27856 3588 27920 3652
rect 27856 3508 27920 3572
rect 27856 3428 27920 3492
rect 27856 3348 27920 3412
rect 27856 3268 27920 3332
rect 27856 3188 27920 3252
rect 27856 3108 27920 3172
rect 27856 3028 27920 3092
rect 27856 2948 27920 3012
rect 27856 2868 27920 2932
rect 27856 2788 27920 2852
rect 27856 2708 27920 2772
rect 27856 2628 27920 2692
rect 27856 2548 27920 2612
rect 27856 2468 27920 2532
rect 27856 2388 27920 2452
rect 27856 2308 27920 2372
rect 27856 2228 27920 2292
rect 27856 2148 27920 2212
rect 27856 2068 27920 2132
rect 27856 1988 27920 2052
rect 27856 1908 27920 1972
rect 27856 1828 27920 1892
rect 27856 1748 27920 1812
rect 27856 1668 27920 1732
rect 27856 1588 27920 1652
rect 27856 1508 27920 1572
rect 27856 1428 27920 1492
rect 27856 1348 27920 1412
rect 27856 1268 27920 1332
rect 27856 1188 27920 1252
rect 27856 1108 27920 1172
rect 27856 1028 27920 1092
rect 27856 948 27920 1012
rect 27856 868 27920 932
rect 27856 788 27920 852
rect 27856 708 27920 772
rect 27856 628 27920 692
rect 27856 548 27920 612
rect 27856 468 27920 532
rect 27856 388 27920 452
rect 27856 308 27920 372
rect 27856 228 27920 292
rect 27856 148 27920 212
rect 33468 5108 33532 5172
rect 33468 5028 33532 5092
rect 33468 4948 33532 5012
rect 33468 4868 33532 4932
rect 33468 4788 33532 4852
rect 33468 4708 33532 4772
rect 33468 4628 33532 4692
rect 33468 4548 33532 4612
rect 33468 4468 33532 4532
rect 33468 4388 33532 4452
rect 33468 4308 33532 4372
rect 33468 4228 33532 4292
rect 33468 4148 33532 4212
rect 33468 4068 33532 4132
rect 33468 3988 33532 4052
rect 33468 3908 33532 3972
rect 33468 3828 33532 3892
rect 33468 3748 33532 3812
rect 33468 3668 33532 3732
rect 33468 3588 33532 3652
rect 33468 3508 33532 3572
rect 33468 3428 33532 3492
rect 33468 3348 33532 3412
rect 33468 3268 33532 3332
rect 33468 3188 33532 3252
rect 33468 3108 33532 3172
rect 33468 3028 33532 3092
rect 33468 2948 33532 3012
rect 33468 2868 33532 2932
rect 33468 2788 33532 2852
rect 33468 2708 33532 2772
rect 33468 2628 33532 2692
rect 33468 2548 33532 2612
rect 33468 2468 33532 2532
rect 33468 2388 33532 2452
rect 33468 2308 33532 2372
rect 33468 2228 33532 2292
rect 33468 2148 33532 2212
rect 33468 2068 33532 2132
rect 33468 1988 33532 2052
rect 33468 1908 33532 1972
rect 33468 1828 33532 1892
rect 33468 1748 33532 1812
rect 33468 1668 33532 1732
rect 33468 1588 33532 1652
rect 33468 1508 33532 1572
rect 33468 1428 33532 1492
rect 33468 1348 33532 1412
rect 33468 1268 33532 1332
rect 33468 1188 33532 1252
rect 33468 1108 33532 1172
rect 33468 1028 33532 1092
rect 33468 948 33532 1012
rect 33468 868 33532 932
rect 33468 788 33532 852
rect 33468 708 33532 772
rect 33468 628 33532 692
rect 33468 548 33532 612
rect 33468 468 33532 532
rect 33468 388 33532 452
rect 33468 308 33532 372
rect 33468 228 33532 292
rect 33468 148 33532 212
rect 39080 5108 39144 5172
rect 39080 5028 39144 5092
rect 39080 4948 39144 5012
rect 39080 4868 39144 4932
rect 39080 4788 39144 4852
rect 39080 4708 39144 4772
rect 39080 4628 39144 4692
rect 39080 4548 39144 4612
rect 39080 4468 39144 4532
rect 39080 4388 39144 4452
rect 39080 4308 39144 4372
rect 39080 4228 39144 4292
rect 39080 4148 39144 4212
rect 39080 4068 39144 4132
rect 39080 3988 39144 4052
rect 39080 3908 39144 3972
rect 39080 3828 39144 3892
rect 39080 3748 39144 3812
rect 39080 3668 39144 3732
rect 39080 3588 39144 3652
rect 39080 3508 39144 3572
rect 39080 3428 39144 3492
rect 39080 3348 39144 3412
rect 39080 3268 39144 3332
rect 39080 3188 39144 3252
rect 39080 3108 39144 3172
rect 39080 3028 39144 3092
rect 39080 2948 39144 3012
rect 39080 2868 39144 2932
rect 39080 2788 39144 2852
rect 39080 2708 39144 2772
rect 39080 2628 39144 2692
rect 39080 2548 39144 2612
rect 39080 2468 39144 2532
rect 39080 2388 39144 2452
rect 39080 2308 39144 2372
rect 39080 2228 39144 2292
rect 39080 2148 39144 2212
rect 39080 2068 39144 2132
rect 39080 1988 39144 2052
rect 39080 1908 39144 1972
rect 39080 1828 39144 1892
rect 39080 1748 39144 1812
rect 39080 1668 39144 1732
rect 39080 1588 39144 1652
rect 39080 1508 39144 1572
rect 39080 1428 39144 1492
rect 39080 1348 39144 1412
rect 39080 1268 39144 1332
rect 39080 1188 39144 1252
rect 39080 1108 39144 1172
rect 39080 1028 39144 1092
rect 39080 948 39144 1012
rect 39080 868 39144 932
rect 39080 788 39144 852
rect 39080 708 39144 772
rect 39080 628 39144 692
rect 39080 548 39144 612
rect 39080 468 39144 532
rect 39080 388 39144 452
rect 39080 308 39144 372
rect 39080 228 39144 292
rect 39080 148 39144 212
rect -33876 -212 -33812 -148
rect -33876 -292 -33812 -228
rect -33876 -372 -33812 -308
rect -33876 -452 -33812 -388
rect -33876 -532 -33812 -468
rect -33876 -612 -33812 -548
rect -33876 -692 -33812 -628
rect -33876 -772 -33812 -708
rect -33876 -852 -33812 -788
rect -33876 -932 -33812 -868
rect -33876 -1012 -33812 -948
rect -33876 -1092 -33812 -1028
rect -33876 -1172 -33812 -1108
rect -33876 -1252 -33812 -1188
rect -33876 -1332 -33812 -1268
rect -33876 -1412 -33812 -1348
rect -33876 -1492 -33812 -1428
rect -33876 -1572 -33812 -1508
rect -33876 -1652 -33812 -1588
rect -33876 -1732 -33812 -1668
rect -33876 -1812 -33812 -1748
rect -33876 -1892 -33812 -1828
rect -33876 -1972 -33812 -1908
rect -33876 -2052 -33812 -1988
rect -33876 -2132 -33812 -2068
rect -33876 -2212 -33812 -2148
rect -33876 -2292 -33812 -2228
rect -33876 -2372 -33812 -2308
rect -33876 -2452 -33812 -2388
rect -33876 -2532 -33812 -2468
rect -33876 -2612 -33812 -2548
rect -33876 -2692 -33812 -2628
rect -33876 -2772 -33812 -2708
rect -33876 -2852 -33812 -2788
rect -33876 -2932 -33812 -2868
rect -33876 -3012 -33812 -2948
rect -33876 -3092 -33812 -3028
rect -33876 -3172 -33812 -3108
rect -33876 -3252 -33812 -3188
rect -33876 -3332 -33812 -3268
rect -33876 -3412 -33812 -3348
rect -33876 -3492 -33812 -3428
rect -33876 -3572 -33812 -3508
rect -33876 -3652 -33812 -3588
rect -33876 -3732 -33812 -3668
rect -33876 -3812 -33812 -3748
rect -33876 -3892 -33812 -3828
rect -33876 -3972 -33812 -3908
rect -33876 -4052 -33812 -3988
rect -33876 -4132 -33812 -4068
rect -33876 -4212 -33812 -4148
rect -33876 -4292 -33812 -4228
rect -33876 -4372 -33812 -4308
rect -33876 -4452 -33812 -4388
rect -33876 -4532 -33812 -4468
rect -33876 -4612 -33812 -4548
rect -33876 -4692 -33812 -4628
rect -33876 -4772 -33812 -4708
rect -33876 -4852 -33812 -4788
rect -33876 -4932 -33812 -4868
rect -33876 -5012 -33812 -4948
rect -33876 -5092 -33812 -5028
rect -33876 -5172 -33812 -5108
rect -28264 -212 -28200 -148
rect -28264 -292 -28200 -228
rect -28264 -372 -28200 -308
rect -28264 -452 -28200 -388
rect -28264 -532 -28200 -468
rect -28264 -612 -28200 -548
rect -28264 -692 -28200 -628
rect -28264 -772 -28200 -708
rect -28264 -852 -28200 -788
rect -28264 -932 -28200 -868
rect -28264 -1012 -28200 -948
rect -28264 -1092 -28200 -1028
rect -28264 -1172 -28200 -1108
rect -28264 -1252 -28200 -1188
rect -28264 -1332 -28200 -1268
rect -28264 -1412 -28200 -1348
rect -28264 -1492 -28200 -1428
rect -28264 -1572 -28200 -1508
rect -28264 -1652 -28200 -1588
rect -28264 -1732 -28200 -1668
rect -28264 -1812 -28200 -1748
rect -28264 -1892 -28200 -1828
rect -28264 -1972 -28200 -1908
rect -28264 -2052 -28200 -1988
rect -28264 -2132 -28200 -2068
rect -28264 -2212 -28200 -2148
rect -28264 -2292 -28200 -2228
rect -28264 -2372 -28200 -2308
rect -28264 -2452 -28200 -2388
rect -28264 -2532 -28200 -2468
rect -28264 -2612 -28200 -2548
rect -28264 -2692 -28200 -2628
rect -28264 -2772 -28200 -2708
rect -28264 -2852 -28200 -2788
rect -28264 -2932 -28200 -2868
rect -28264 -3012 -28200 -2948
rect -28264 -3092 -28200 -3028
rect -28264 -3172 -28200 -3108
rect -28264 -3252 -28200 -3188
rect -28264 -3332 -28200 -3268
rect -28264 -3412 -28200 -3348
rect -28264 -3492 -28200 -3428
rect -28264 -3572 -28200 -3508
rect -28264 -3652 -28200 -3588
rect -28264 -3732 -28200 -3668
rect -28264 -3812 -28200 -3748
rect -28264 -3892 -28200 -3828
rect -28264 -3972 -28200 -3908
rect -28264 -4052 -28200 -3988
rect -28264 -4132 -28200 -4068
rect -28264 -4212 -28200 -4148
rect -28264 -4292 -28200 -4228
rect -28264 -4372 -28200 -4308
rect -28264 -4452 -28200 -4388
rect -28264 -4532 -28200 -4468
rect -28264 -4612 -28200 -4548
rect -28264 -4692 -28200 -4628
rect -28264 -4772 -28200 -4708
rect -28264 -4852 -28200 -4788
rect -28264 -4932 -28200 -4868
rect -28264 -5012 -28200 -4948
rect -28264 -5092 -28200 -5028
rect -28264 -5172 -28200 -5108
rect -22652 -212 -22588 -148
rect -22652 -292 -22588 -228
rect -22652 -372 -22588 -308
rect -22652 -452 -22588 -388
rect -22652 -532 -22588 -468
rect -22652 -612 -22588 -548
rect -22652 -692 -22588 -628
rect -22652 -772 -22588 -708
rect -22652 -852 -22588 -788
rect -22652 -932 -22588 -868
rect -22652 -1012 -22588 -948
rect -22652 -1092 -22588 -1028
rect -22652 -1172 -22588 -1108
rect -22652 -1252 -22588 -1188
rect -22652 -1332 -22588 -1268
rect -22652 -1412 -22588 -1348
rect -22652 -1492 -22588 -1428
rect -22652 -1572 -22588 -1508
rect -22652 -1652 -22588 -1588
rect -22652 -1732 -22588 -1668
rect -22652 -1812 -22588 -1748
rect -22652 -1892 -22588 -1828
rect -22652 -1972 -22588 -1908
rect -22652 -2052 -22588 -1988
rect -22652 -2132 -22588 -2068
rect -22652 -2212 -22588 -2148
rect -22652 -2292 -22588 -2228
rect -22652 -2372 -22588 -2308
rect -22652 -2452 -22588 -2388
rect -22652 -2532 -22588 -2468
rect -22652 -2612 -22588 -2548
rect -22652 -2692 -22588 -2628
rect -22652 -2772 -22588 -2708
rect -22652 -2852 -22588 -2788
rect -22652 -2932 -22588 -2868
rect -22652 -3012 -22588 -2948
rect -22652 -3092 -22588 -3028
rect -22652 -3172 -22588 -3108
rect -22652 -3252 -22588 -3188
rect -22652 -3332 -22588 -3268
rect -22652 -3412 -22588 -3348
rect -22652 -3492 -22588 -3428
rect -22652 -3572 -22588 -3508
rect -22652 -3652 -22588 -3588
rect -22652 -3732 -22588 -3668
rect -22652 -3812 -22588 -3748
rect -22652 -3892 -22588 -3828
rect -22652 -3972 -22588 -3908
rect -22652 -4052 -22588 -3988
rect -22652 -4132 -22588 -4068
rect -22652 -4212 -22588 -4148
rect -22652 -4292 -22588 -4228
rect -22652 -4372 -22588 -4308
rect -22652 -4452 -22588 -4388
rect -22652 -4532 -22588 -4468
rect -22652 -4612 -22588 -4548
rect -22652 -4692 -22588 -4628
rect -22652 -4772 -22588 -4708
rect -22652 -4852 -22588 -4788
rect -22652 -4932 -22588 -4868
rect -22652 -5012 -22588 -4948
rect -22652 -5092 -22588 -5028
rect -22652 -5172 -22588 -5108
rect -17040 -212 -16976 -148
rect -17040 -292 -16976 -228
rect -17040 -372 -16976 -308
rect -17040 -452 -16976 -388
rect -17040 -532 -16976 -468
rect -17040 -612 -16976 -548
rect -17040 -692 -16976 -628
rect -17040 -772 -16976 -708
rect -17040 -852 -16976 -788
rect -17040 -932 -16976 -868
rect -17040 -1012 -16976 -948
rect -17040 -1092 -16976 -1028
rect -17040 -1172 -16976 -1108
rect -17040 -1252 -16976 -1188
rect -17040 -1332 -16976 -1268
rect -17040 -1412 -16976 -1348
rect -17040 -1492 -16976 -1428
rect -17040 -1572 -16976 -1508
rect -17040 -1652 -16976 -1588
rect -17040 -1732 -16976 -1668
rect -17040 -1812 -16976 -1748
rect -17040 -1892 -16976 -1828
rect -17040 -1972 -16976 -1908
rect -17040 -2052 -16976 -1988
rect -17040 -2132 -16976 -2068
rect -17040 -2212 -16976 -2148
rect -17040 -2292 -16976 -2228
rect -17040 -2372 -16976 -2308
rect -17040 -2452 -16976 -2388
rect -17040 -2532 -16976 -2468
rect -17040 -2612 -16976 -2548
rect -17040 -2692 -16976 -2628
rect -17040 -2772 -16976 -2708
rect -17040 -2852 -16976 -2788
rect -17040 -2932 -16976 -2868
rect -17040 -3012 -16976 -2948
rect -17040 -3092 -16976 -3028
rect -17040 -3172 -16976 -3108
rect -17040 -3252 -16976 -3188
rect -17040 -3332 -16976 -3268
rect -17040 -3412 -16976 -3348
rect -17040 -3492 -16976 -3428
rect -17040 -3572 -16976 -3508
rect -17040 -3652 -16976 -3588
rect -17040 -3732 -16976 -3668
rect -17040 -3812 -16976 -3748
rect -17040 -3892 -16976 -3828
rect -17040 -3972 -16976 -3908
rect -17040 -4052 -16976 -3988
rect -17040 -4132 -16976 -4068
rect -17040 -4212 -16976 -4148
rect -17040 -4292 -16976 -4228
rect -17040 -4372 -16976 -4308
rect -17040 -4452 -16976 -4388
rect -17040 -4532 -16976 -4468
rect -17040 -4612 -16976 -4548
rect -17040 -4692 -16976 -4628
rect -17040 -4772 -16976 -4708
rect -17040 -4852 -16976 -4788
rect -17040 -4932 -16976 -4868
rect -17040 -5012 -16976 -4948
rect -17040 -5092 -16976 -5028
rect -17040 -5172 -16976 -5108
rect -11428 -212 -11364 -148
rect -11428 -292 -11364 -228
rect -11428 -372 -11364 -308
rect -11428 -452 -11364 -388
rect -11428 -532 -11364 -468
rect -11428 -612 -11364 -548
rect -11428 -692 -11364 -628
rect -11428 -772 -11364 -708
rect -11428 -852 -11364 -788
rect -11428 -932 -11364 -868
rect -11428 -1012 -11364 -948
rect -11428 -1092 -11364 -1028
rect -11428 -1172 -11364 -1108
rect -11428 -1252 -11364 -1188
rect -11428 -1332 -11364 -1268
rect -11428 -1412 -11364 -1348
rect -11428 -1492 -11364 -1428
rect -11428 -1572 -11364 -1508
rect -11428 -1652 -11364 -1588
rect -11428 -1732 -11364 -1668
rect -11428 -1812 -11364 -1748
rect -11428 -1892 -11364 -1828
rect -11428 -1972 -11364 -1908
rect -11428 -2052 -11364 -1988
rect -11428 -2132 -11364 -2068
rect -11428 -2212 -11364 -2148
rect -11428 -2292 -11364 -2228
rect -11428 -2372 -11364 -2308
rect -11428 -2452 -11364 -2388
rect -11428 -2532 -11364 -2468
rect -11428 -2612 -11364 -2548
rect -11428 -2692 -11364 -2628
rect -11428 -2772 -11364 -2708
rect -11428 -2852 -11364 -2788
rect -11428 -2932 -11364 -2868
rect -11428 -3012 -11364 -2948
rect -11428 -3092 -11364 -3028
rect -11428 -3172 -11364 -3108
rect -11428 -3252 -11364 -3188
rect -11428 -3332 -11364 -3268
rect -11428 -3412 -11364 -3348
rect -11428 -3492 -11364 -3428
rect -11428 -3572 -11364 -3508
rect -11428 -3652 -11364 -3588
rect -11428 -3732 -11364 -3668
rect -11428 -3812 -11364 -3748
rect -11428 -3892 -11364 -3828
rect -11428 -3972 -11364 -3908
rect -11428 -4052 -11364 -3988
rect -11428 -4132 -11364 -4068
rect -11428 -4212 -11364 -4148
rect -11428 -4292 -11364 -4228
rect -11428 -4372 -11364 -4308
rect -11428 -4452 -11364 -4388
rect -11428 -4532 -11364 -4468
rect -11428 -4612 -11364 -4548
rect -11428 -4692 -11364 -4628
rect -11428 -4772 -11364 -4708
rect -11428 -4852 -11364 -4788
rect -11428 -4932 -11364 -4868
rect -11428 -5012 -11364 -4948
rect -11428 -5092 -11364 -5028
rect -11428 -5172 -11364 -5108
rect -5816 -212 -5752 -148
rect -5816 -292 -5752 -228
rect -5816 -372 -5752 -308
rect -5816 -452 -5752 -388
rect -5816 -532 -5752 -468
rect -5816 -612 -5752 -548
rect -5816 -692 -5752 -628
rect -5816 -772 -5752 -708
rect -5816 -852 -5752 -788
rect -5816 -932 -5752 -868
rect -5816 -1012 -5752 -948
rect -5816 -1092 -5752 -1028
rect -5816 -1172 -5752 -1108
rect -5816 -1252 -5752 -1188
rect -5816 -1332 -5752 -1268
rect -5816 -1412 -5752 -1348
rect -5816 -1492 -5752 -1428
rect -5816 -1572 -5752 -1508
rect -5816 -1652 -5752 -1588
rect -5816 -1732 -5752 -1668
rect -5816 -1812 -5752 -1748
rect -5816 -1892 -5752 -1828
rect -5816 -1972 -5752 -1908
rect -5816 -2052 -5752 -1988
rect -5816 -2132 -5752 -2068
rect -5816 -2212 -5752 -2148
rect -5816 -2292 -5752 -2228
rect -5816 -2372 -5752 -2308
rect -5816 -2452 -5752 -2388
rect -5816 -2532 -5752 -2468
rect -5816 -2612 -5752 -2548
rect -5816 -2692 -5752 -2628
rect -5816 -2772 -5752 -2708
rect -5816 -2852 -5752 -2788
rect -5816 -2932 -5752 -2868
rect -5816 -3012 -5752 -2948
rect -5816 -3092 -5752 -3028
rect -5816 -3172 -5752 -3108
rect -5816 -3252 -5752 -3188
rect -5816 -3332 -5752 -3268
rect -5816 -3412 -5752 -3348
rect -5816 -3492 -5752 -3428
rect -5816 -3572 -5752 -3508
rect -5816 -3652 -5752 -3588
rect -5816 -3732 -5752 -3668
rect -5816 -3812 -5752 -3748
rect -5816 -3892 -5752 -3828
rect -5816 -3972 -5752 -3908
rect -5816 -4052 -5752 -3988
rect -5816 -4132 -5752 -4068
rect -5816 -4212 -5752 -4148
rect -5816 -4292 -5752 -4228
rect -5816 -4372 -5752 -4308
rect -5816 -4452 -5752 -4388
rect -5816 -4532 -5752 -4468
rect -5816 -4612 -5752 -4548
rect -5816 -4692 -5752 -4628
rect -5816 -4772 -5752 -4708
rect -5816 -4852 -5752 -4788
rect -5816 -4932 -5752 -4868
rect -5816 -5012 -5752 -4948
rect -5816 -5092 -5752 -5028
rect -5816 -5172 -5752 -5108
rect -204 -212 -140 -148
rect -204 -292 -140 -228
rect -204 -372 -140 -308
rect -204 -452 -140 -388
rect -204 -532 -140 -468
rect -204 -612 -140 -548
rect -204 -692 -140 -628
rect -204 -772 -140 -708
rect -204 -852 -140 -788
rect -204 -932 -140 -868
rect -204 -1012 -140 -948
rect -204 -1092 -140 -1028
rect -204 -1172 -140 -1108
rect -204 -1252 -140 -1188
rect -204 -1332 -140 -1268
rect -204 -1412 -140 -1348
rect -204 -1492 -140 -1428
rect -204 -1572 -140 -1508
rect -204 -1652 -140 -1588
rect -204 -1732 -140 -1668
rect -204 -1812 -140 -1748
rect -204 -1892 -140 -1828
rect -204 -1972 -140 -1908
rect -204 -2052 -140 -1988
rect -204 -2132 -140 -2068
rect -204 -2212 -140 -2148
rect -204 -2292 -140 -2228
rect -204 -2372 -140 -2308
rect -204 -2452 -140 -2388
rect -204 -2532 -140 -2468
rect -204 -2612 -140 -2548
rect -204 -2692 -140 -2628
rect -204 -2772 -140 -2708
rect -204 -2852 -140 -2788
rect -204 -2932 -140 -2868
rect -204 -3012 -140 -2948
rect -204 -3092 -140 -3028
rect -204 -3172 -140 -3108
rect -204 -3252 -140 -3188
rect -204 -3332 -140 -3268
rect -204 -3412 -140 -3348
rect -204 -3492 -140 -3428
rect -204 -3572 -140 -3508
rect -204 -3652 -140 -3588
rect -204 -3732 -140 -3668
rect -204 -3812 -140 -3748
rect -204 -3892 -140 -3828
rect -204 -3972 -140 -3908
rect -204 -4052 -140 -3988
rect -204 -4132 -140 -4068
rect -204 -4212 -140 -4148
rect -204 -4292 -140 -4228
rect -204 -4372 -140 -4308
rect -204 -4452 -140 -4388
rect -204 -4532 -140 -4468
rect -204 -4612 -140 -4548
rect -204 -4692 -140 -4628
rect -204 -4772 -140 -4708
rect -204 -4852 -140 -4788
rect -204 -4932 -140 -4868
rect -204 -5012 -140 -4948
rect -204 -5092 -140 -5028
rect -204 -5172 -140 -5108
rect 5408 -212 5472 -148
rect 5408 -292 5472 -228
rect 5408 -372 5472 -308
rect 5408 -452 5472 -388
rect 5408 -532 5472 -468
rect 5408 -612 5472 -548
rect 5408 -692 5472 -628
rect 5408 -772 5472 -708
rect 5408 -852 5472 -788
rect 5408 -932 5472 -868
rect 5408 -1012 5472 -948
rect 5408 -1092 5472 -1028
rect 5408 -1172 5472 -1108
rect 5408 -1252 5472 -1188
rect 5408 -1332 5472 -1268
rect 5408 -1412 5472 -1348
rect 5408 -1492 5472 -1428
rect 5408 -1572 5472 -1508
rect 5408 -1652 5472 -1588
rect 5408 -1732 5472 -1668
rect 5408 -1812 5472 -1748
rect 5408 -1892 5472 -1828
rect 5408 -1972 5472 -1908
rect 5408 -2052 5472 -1988
rect 5408 -2132 5472 -2068
rect 5408 -2212 5472 -2148
rect 5408 -2292 5472 -2228
rect 5408 -2372 5472 -2308
rect 5408 -2452 5472 -2388
rect 5408 -2532 5472 -2468
rect 5408 -2612 5472 -2548
rect 5408 -2692 5472 -2628
rect 5408 -2772 5472 -2708
rect 5408 -2852 5472 -2788
rect 5408 -2932 5472 -2868
rect 5408 -3012 5472 -2948
rect 5408 -3092 5472 -3028
rect 5408 -3172 5472 -3108
rect 5408 -3252 5472 -3188
rect 5408 -3332 5472 -3268
rect 5408 -3412 5472 -3348
rect 5408 -3492 5472 -3428
rect 5408 -3572 5472 -3508
rect 5408 -3652 5472 -3588
rect 5408 -3732 5472 -3668
rect 5408 -3812 5472 -3748
rect 5408 -3892 5472 -3828
rect 5408 -3972 5472 -3908
rect 5408 -4052 5472 -3988
rect 5408 -4132 5472 -4068
rect 5408 -4212 5472 -4148
rect 5408 -4292 5472 -4228
rect 5408 -4372 5472 -4308
rect 5408 -4452 5472 -4388
rect 5408 -4532 5472 -4468
rect 5408 -4612 5472 -4548
rect 5408 -4692 5472 -4628
rect 5408 -4772 5472 -4708
rect 5408 -4852 5472 -4788
rect 5408 -4932 5472 -4868
rect 5408 -5012 5472 -4948
rect 5408 -5092 5472 -5028
rect 5408 -5172 5472 -5108
rect 11020 -212 11084 -148
rect 11020 -292 11084 -228
rect 11020 -372 11084 -308
rect 11020 -452 11084 -388
rect 11020 -532 11084 -468
rect 11020 -612 11084 -548
rect 11020 -692 11084 -628
rect 11020 -772 11084 -708
rect 11020 -852 11084 -788
rect 11020 -932 11084 -868
rect 11020 -1012 11084 -948
rect 11020 -1092 11084 -1028
rect 11020 -1172 11084 -1108
rect 11020 -1252 11084 -1188
rect 11020 -1332 11084 -1268
rect 11020 -1412 11084 -1348
rect 11020 -1492 11084 -1428
rect 11020 -1572 11084 -1508
rect 11020 -1652 11084 -1588
rect 11020 -1732 11084 -1668
rect 11020 -1812 11084 -1748
rect 11020 -1892 11084 -1828
rect 11020 -1972 11084 -1908
rect 11020 -2052 11084 -1988
rect 11020 -2132 11084 -2068
rect 11020 -2212 11084 -2148
rect 11020 -2292 11084 -2228
rect 11020 -2372 11084 -2308
rect 11020 -2452 11084 -2388
rect 11020 -2532 11084 -2468
rect 11020 -2612 11084 -2548
rect 11020 -2692 11084 -2628
rect 11020 -2772 11084 -2708
rect 11020 -2852 11084 -2788
rect 11020 -2932 11084 -2868
rect 11020 -3012 11084 -2948
rect 11020 -3092 11084 -3028
rect 11020 -3172 11084 -3108
rect 11020 -3252 11084 -3188
rect 11020 -3332 11084 -3268
rect 11020 -3412 11084 -3348
rect 11020 -3492 11084 -3428
rect 11020 -3572 11084 -3508
rect 11020 -3652 11084 -3588
rect 11020 -3732 11084 -3668
rect 11020 -3812 11084 -3748
rect 11020 -3892 11084 -3828
rect 11020 -3972 11084 -3908
rect 11020 -4052 11084 -3988
rect 11020 -4132 11084 -4068
rect 11020 -4212 11084 -4148
rect 11020 -4292 11084 -4228
rect 11020 -4372 11084 -4308
rect 11020 -4452 11084 -4388
rect 11020 -4532 11084 -4468
rect 11020 -4612 11084 -4548
rect 11020 -4692 11084 -4628
rect 11020 -4772 11084 -4708
rect 11020 -4852 11084 -4788
rect 11020 -4932 11084 -4868
rect 11020 -5012 11084 -4948
rect 11020 -5092 11084 -5028
rect 11020 -5172 11084 -5108
rect 16632 -212 16696 -148
rect 16632 -292 16696 -228
rect 16632 -372 16696 -308
rect 16632 -452 16696 -388
rect 16632 -532 16696 -468
rect 16632 -612 16696 -548
rect 16632 -692 16696 -628
rect 16632 -772 16696 -708
rect 16632 -852 16696 -788
rect 16632 -932 16696 -868
rect 16632 -1012 16696 -948
rect 16632 -1092 16696 -1028
rect 16632 -1172 16696 -1108
rect 16632 -1252 16696 -1188
rect 16632 -1332 16696 -1268
rect 16632 -1412 16696 -1348
rect 16632 -1492 16696 -1428
rect 16632 -1572 16696 -1508
rect 16632 -1652 16696 -1588
rect 16632 -1732 16696 -1668
rect 16632 -1812 16696 -1748
rect 16632 -1892 16696 -1828
rect 16632 -1972 16696 -1908
rect 16632 -2052 16696 -1988
rect 16632 -2132 16696 -2068
rect 16632 -2212 16696 -2148
rect 16632 -2292 16696 -2228
rect 16632 -2372 16696 -2308
rect 16632 -2452 16696 -2388
rect 16632 -2532 16696 -2468
rect 16632 -2612 16696 -2548
rect 16632 -2692 16696 -2628
rect 16632 -2772 16696 -2708
rect 16632 -2852 16696 -2788
rect 16632 -2932 16696 -2868
rect 16632 -3012 16696 -2948
rect 16632 -3092 16696 -3028
rect 16632 -3172 16696 -3108
rect 16632 -3252 16696 -3188
rect 16632 -3332 16696 -3268
rect 16632 -3412 16696 -3348
rect 16632 -3492 16696 -3428
rect 16632 -3572 16696 -3508
rect 16632 -3652 16696 -3588
rect 16632 -3732 16696 -3668
rect 16632 -3812 16696 -3748
rect 16632 -3892 16696 -3828
rect 16632 -3972 16696 -3908
rect 16632 -4052 16696 -3988
rect 16632 -4132 16696 -4068
rect 16632 -4212 16696 -4148
rect 16632 -4292 16696 -4228
rect 16632 -4372 16696 -4308
rect 16632 -4452 16696 -4388
rect 16632 -4532 16696 -4468
rect 16632 -4612 16696 -4548
rect 16632 -4692 16696 -4628
rect 16632 -4772 16696 -4708
rect 16632 -4852 16696 -4788
rect 16632 -4932 16696 -4868
rect 16632 -5012 16696 -4948
rect 16632 -5092 16696 -5028
rect 16632 -5172 16696 -5108
rect 22244 -212 22308 -148
rect 22244 -292 22308 -228
rect 22244 -372 22308 -308
rect 22244 -452 22308 -388
rect 22244 -532 22308 -468
rect 22244 -612 22308 -548
rect 22244 -692 22308 -628
rect 22244 -772 22308 -708
rect 22244 -852 22308 -788
rect 22244 -932 22308 -868
rect 22244 -1012 22308 -948
rect 22244 -1092 22308 -1028
rect 22244 -1172 22308 -1108
rect 22244 -1252 22308 -1188
rect 22244 -1332 22308 -1268
rect 22244 -1412 22308 -1348
rect 22244 -1492 22308 -1428
rect 22244 -1572 22308 -1508
rect 22244 -1652 22308 -1588
rect 22244 -1732 22308 -1668
rect 22244 -1812 22308 -1748
rect 22244 -1892 22308 -1828
rect 22244 -1972 22308 -1908
rect 22244 -2052 22308 -1988
rect 22244 -2132 22308 -2068
rect 22244 -2212 22308 -2148
rect 22244 -2292 22308 -2228
rect 22244 -2372 22308 -2308
rect 22244 -2452 22308 -2388
rect 22244 -2532 22308 -2468
rect 22244 -2612 22308 -2548
rect 22244 -2692 22308 -2628
rect 22244 -2772 22308 -2708
rect 22244 -2852 22308 -2788
rect 22244 -2932 22308 -2868
rect 22244 -3012 22308 -2948
rect 22244 -3092 22308 -3028
rect 22244 -3172 22308 -3108
rect 22244 -3252 22308 -3188
rect 22244 -3332 22308 -3268
rect 22244 -3412 22308 -3348
rect 22244 -3492 22308 -3428
rect 22244 -3572 22308 -3508
rect 22244 -3652 22308 -3588
rect 22244 -3732 22308 -3668
rect 22244 -3812 22308 -3748
rect 22244 -3892 22308 -3828
rect 22244 -3972 22308 -3908
rect 22244 -4052 22308 -3988
rect 22244 -4132 22308 -4068
rect 22244 -4212 22308 -4148
rect 22244 -4292 22308 -4228
rect 22244 -4372 22308 -4308
rect 22244 -4452 22308 -4388
rect 22244 -4532 22308 -4468
rect 22244 -4612 22308 -4548
rect 22244 -4692 22308 -4628
rect 22244 -4772 22308 -4708
rect 22244 -4852 22308 -4788
rect 22244 -4932 22308 -4868
rect 22244 -5012 22308 -4948
rect 22244 -5092 22308 -5028
rect 22244 -5172 22308 -5108
rect 27856 -212 27920 -148
rect 27856 -292 27920 -228
rect 27856 -372 27920 -308
rect 27856 -452 27920 -388
rect 27856 -532 27920 -468
rect 27856 -612 27920 -548
rect 27856 -692 27920 -628
rect 27856 -772 27920 -708
rect 27856 -852 27920 -788
rect 27856 -932 27920 -868
rect 27856 -1012 27920 -948
rect 27856 -1092 27920 -1028
rect 27856 -1172 27920 -1108
rect 27856 -1252 27920 -1188
rect 27856 -1332 27920 -1268
rect 27856 -1412 27920 -1348
rect 27856 -1492 27920 -1428
rect 27856 -1572 27920 -1508
rect 27856 -1652 27920 -1588
rect 27856 -1732 27920 -1668
rect 27856 -1812 27920 -1748
rect 27856 -1892 27920 -1828
rect 27856 -1972 27920 -1908
rect 27856 -2052 27920 -1988
rect 27856 -2132 27920 -2068
rect 27856 -2212 27920 -2148
rect 27856 -2292 27920 -2228
rect 27856 -2372 27920 -2308
rect 27856 -2452 27920 -2388
rect 27856 -2532 27920 -2468
rect 27856 -2612 27920 -2548
rect 27856 -2692 27920 -2628
rect 27856 -2772 27920 -2708
rect 27856 -2852 27920 -2788
rect 27856 -2932 27920 -2868
rect 27856 -3012 27920 -2948
rect 27856 -3092 27920 -3028
rect 27856 -3172 27920 -3108
rect 27856 -3252 27920 -3188
rect 27856 -3332 27920 -3268
rect 27856 -3412 27920 -3348
rect 27856 -3492 27920 -3428
rect 27856 -3572 27920 -3508
rect 27856 -3652 27920 -3588
rect 27856 -3732 27920 -3668
rect 27856 -3812 27920 -3748
rect 27856 -3892 27920 -3828
rect 27856 -3972 27920 -3908
rect 27856 -4052 27920 -3988
rect 27856 -4132 27920 -4068
rect 27856 -4212 27920 -4148
rect 27856 -4292 27920 -4228
rect 27856 -4372 27920 -4308
rect 27856 -4452 27920 -4388
rect 27856 -4532 27920 -4468
rect 27856 -4612 27920 -4548
rect 27856 -4692 27920 -4628
rect 27856 -4772 27920 -4708
rect 27856 -4852 27920 -4788
rect 27856 -4932 27920 -4868
rect 27856 -5012 27920 -4948
rect 27856 -5092 27920 -5028
rect 27856 -5172 27920 -5108
rect 33468 -212 33532 -148
rect 33468 -292 33532 -228
rect 33468 -372 33532 -308
rect 33468 -452 33532 -388
rect 33468 -532 33532 -468
rect 33468 -612 33532 -548
rect 33468 -692 33532 -628
rect 33468 -772 33532 -708
rect 33468 -852 33532 -788
rect 33468 -932 33532 -868
rect 33468 -1012 33532 -948
rect 33468 -1092 33532 -1028
rect 33468 -1172 33532 -1108
rect 33468 -1252 33532 -1188
rect 33468 -1332 33532 -1268
rect 33468 -1412 33532 -1348
rect 33468 -1492 33532 -1428
rect 33468 -1572 33532 -1508
rect 33468 -1652 33532 -1588
rect 33468 -1732 33532 -1668
rect 33468 -1812 33532 -1748
rect 33468 -1892 33532 -1828
rect 33468 -1972 33532 -1908
rect 33468 -2052 33532 -1988
rect 33468 -2132 33532 -2068
rect 33468 -2212 33532 -2148
rect 33468 -2292 33532 -2228
rect 33468 -2372 33532 -2308
rect 33468 -2452 33532 -2388
rect 33468 -2532 33532 -2468
rect 33468 -2612 33532 -2548
rect 33468 -2692 33532 -2628
rect 33468 -2772 33532 -2708
rect 33468 -2852 33532 -2788
rect 33468 -2932 33532 -2868
rect 33468 -3012 33532 -2948
rect 33468 -3092 33532 -3028
rect 33468 -3172 33532 -3108
rect 33468 -3252 33532 -3188
rect 33468 -3332 33532 -3268
rect 33468 -3412 33532 -3348
rect 33468 -3492 33532 -3428
rect 33468 -3572 33532 -3508
rect 33468 -3652 33532 -3588
rect 33468 -3732 33532 -3668
rect 33468 -3812 33532 -3748
rect 33468 -3892 33532 -3828
rect 33468 -3972 33532 -3908
rect 33468 -4052 33532 -3988
rect 33468 -4132 33532 -4068
rect 33468 -4212 33532 -4148
rect 33468 -4292 33532 -4228
rect 33468 -4372 33532 -4308
rect 33468 -4452 33532 -4388
rect 33468 -4532 33532 -4468
rect 33468 -4612 33532 -4548
rect 33468 -4692 33532 -4628
rect 33468 -4772 33532 -4708
rect 33468 -4852 33532 -4788
rect 33468 -4932 33532 -4868
rect 33468 -5012 33532 -4948
rect 33468 -5092 33532 -5028
rect 33468 -5172 33532 -5108
rect 39080 -212 39144 -148
rect 39080 -292 39144 -228
rect 39080 -372 39144 -308
rect 39080 -452 39144 -388
rect 39080 -532 39144 -468
rect 39080 -612 39144 -548
rect 39080 -692 39144 -628
rect 39080 -772 39144 -708
rect 39080 -852 39144 -788
rect 39080 -932 39144 -868
rect 39080 -1012 39144 -948
rect 39080 -1092 39144 -1028
rect 39080 -1172 39144 -1108
rect 39080 -1252 39144 -1188
rect 39080 -1332 39144 -1268
rect 39080 -1412 39144 -1348
rect 39080 -1492 39144 -1428
rect 39080 -1572 39144 -1508
rect 39080 -1652 39144 -1588
rect 39080 -1732 39144 -1668
rect 39080 -1812 39144 -1748
rect 39080 -1892 39144 -1828
rect 39080 -1972 39144 -1908
rect 39080 -2052 39144 -1988
rect 39080 -2132 39144 -2068
rect 39080 -2212 39144 -2148
rect 39080 -2292 39144 -2228
rect 39080 -2372 39144 -2308
rect 39080 -2452 39144 -2388
rect 39080 -2532 39144 -2468
rect 39080 -2612 39144 -2548
rect 39080 -2692 39144 -2628
rect 39080 -2772 39144 -2708
rect 39080 -2852 39144 -2788
rect 39080 -2932 39144 -2868
rect 39080 -3012 39144 -2948
rect 39080 -3092 39144 -3028
rect 39080 -3172 39144 -3108
rect 39080 -3252 39144 -3188
rect 39080 -3332 39144 -3268
rect 39080 -3412 39144 -3348
rect 39080 -3492 39144 -3428
rect 39080 -3572 39144 -3508
rect 39080 -3652 39144 -3588
rect 39080 -3732 39144 -3668
rect 39080 -3812 39144 -3748
rect 39080 -3892 39144 -3828
rect 39080 -3972 39144 -3908
rect 39080 -4052 39144 -3988
rect 39080 -4132 39144 -4068
rect 39080 -4212 39144 -4148
rect 39080 -4292 39144 -4228
rect 39080 -4372 39144 -4308
rect 39080 -4452 39144 -4388
rect 39080 -4532 39144 -4468
rect 39080 -4612 39144 -4548
rect 39080 -4692 39144 -4628
rect 39080 -4772 39144 -4708
rect 39080 -4852 39144 -4788
rect 39080 -4932 39144 -4868
rect 39080 -5012 39144 -4948
rect 39080 -5092 39144 -5028
rect 39080 -5172 39144 -5108
rect -33876 -5532 -33812 -5468
rect -33876 -5612 -33812 -5548
rect -33876 -5692 -33812 -5628
rect -33876 -5772 -33812 -5708
rect -33876 -5852 -33812 -5788
rect -33876 -5932 -33812 -5868
rect -33876 -6012 -33812 -5948
rect -33876 -6092 -33812 -6028
rect -33876 -6172 -33812 -6108
rect -33876 -6252 -33812 -6188
rect -33876 -6332 -33812 -6268
rect -33876 -6412 -33812 -6348
rect -33876 -6492 -33812 -6428
rect -33876 -6572 -33812 -6508
rect -33876 -6652 -33812 -6588
rect -33876 -6732 -33812 -6668
rect -33876 -6812 -33812 -6748
rect -33876 -6892 -33812 -6828
rect -33876 -6972 -33812 -6908
rect -33876 -7052 -33812 -6988
rect -33876 -7132 -33812 -7068
rect -33876 -7212 -33812 -7148
rect -33876 -7292 -33812 -7228
rect -33876 -7372 -33812 -7308
rect -33876 -7452 -33812 -7388
rect -33876 -7532 -33812 -7468
rect -33876 -7612 -33812 -7548
rect -33876 -7692 -33812 -7628
rect -33876 -7772 -33812 -7708
rect -33876 -7852 -33812 -7788
rect -33876 -7932 -33812 -7868
rect -33876 -8012 -33812 -7948
rect -33876 -8092 -33812 -8028
rect -33876 -8172 -33812 -8108
rect -33876 -8252 -33812 -8188
rect -33876 -8332 -33812 -8268
rect -33876 -8412 -33812 -8348
rect -33876 -8492 -33812 -8428
rect -33876 -8572 -33812 -8508
rect -33876 -8652 -33812 -8588
rect -33876 -8732 -33812 -8668
rect -33876 -8812 -33812 -8748
rect -33876 -8892 -33812 -8828
rect -33876 -8972 -33812 -8908
rect -33876 -9052 -33812 -8988
rect -33876 -9132 -33812 -9068
rect -33876 -9212 -33812 -9148
rect -33876 -9292 -33812 -9228
rect -33876 -9372 -33812 -9308
rect -33876 -9452 -33812 -9388
rect -33876 -9532 -33812 -9468
rect -33876 -9612 -33812 -9548
rect -33876 -9692 -33812 -9628
rect -33876 -9772 -33812 -9708
rect -33876 -9852 -33812 -9788
rect -33876 -9932 -33812 -9868
rect -33876 -10012 -33812 -9948
rect -33876 -10092 -33812 -10028
rect -33876 -10172 -33812 -10108
rect -33876 -10252 -33812 -10188
rect -33876 -10332 -33812 -10268
rect -33876 -10412 -33812 -10348
rect -33876 -10492 -33812 -10428
rect -28264 -5532 -28200 -5468
rect -28264 -5612 -28200 -5548
rect -28264 -5692 -28200 -5628
rect -28264 -5772 -28200 -5708
rect -28264 -5852 -28200 -5788
rect -28264 -5932 -28200 -5868
rect -28264 -6012 -28200 -5948
rect -28264 -6092 -28200 -6028
rect -28264 -6172 -28200 -6108
rect -28264 -6252 -28200 -6188
rect -28264 -6332 -28200 -6268
rect -28264 -6412 -28200 -6348
rect -28264 -6492 -28200 -6428
rect -28264 -6572 -28200 -6508
rect -28264 -6652 -28200 -6588
rect -28264 -6732 -28200 -6668
rect -28264 -6812 -28200 -6748
rect -28264 -6892 -28200 -6828
rect -28264 -6972 -28200 -6908
rect -28264 -7052 -28200 -6988
rect -28264 -7132 -28200 -7068
rect -28264 -7212 -28200 -7148
rect -28264 -7292 -28200 -7228
rect -28264 -7372 -28200 -7308
rect -28264 -7452 -28200 -7388
rect -28264 -7532 -28200 -7468
rect -28264 -7612 -28200 -7548
rect -28264 -7692 -28200 -7628
rect -28264 -7772 -28200 -7708
rect -28264 -7852 -28200 -7788
rect -28264 -7932 -28200 -7868
rect -28264 -8012 -28200 -7948
rect -28264 -8092 -28200 -8028
rect -28264 -8172 -28200 -8108
rect -28264 -8252 -28200 -8188
rect -28264 -8332 -28200 -8268
rect -28264 -8412 -28200 -8348
rect -28264 -8492 -28200 -8428
rect -28264 -8572 -28200 -8508
rect -28264 -8652 -28200 -8588
rect -28264 -8732 -28200 -8668
rect -28264 -8812 -28200 -8748
rect -28264 -8892 -28200 -8828
rect -28264 -8972 -28200 -8908
rect -28264 -9052 -28200 -8988
rect -28264 -9132 -28200 -9068
rect -28264 -9212 -28200 -9148
rect -28264 -9292 -28200 -9228
rect -28264 -9372 -28200 -9308
rect -28264 -9452 -28200 -9388
rect -28264 -9532 -28200 -9468
rect -28264 -9612 -28200 -9548
rect -28264 -9692 -28200 -9628
rect -28264 -9772 -28200 -9708
rect -28264 -9852 -28200 -9788
rect -28264 -9932 -28200 -9868
rect -28264 -10012 -28200 -9948
rect -28264 -10092 -28200 -10028
rect -28264 -10172 -28200 -10108
rect -28264 -10252 -28200 -10188
rect -28264 -10332 -28200 -10268
rect -28264 -10412 -28200 -10348
rect -28264 -10492 -28200 -10428
rect -22652 -5532 -22588 -5468
rect -22652 -5612 -22588 -5548
rect -22652 -5692 -22588 -5628
rect -22652 -5772 -22588 -5708
rect -22652 -5852 -22588 -5788
rect -22652 -5932 -22588 -5868
rect -22652 -6012 -22588 -5948
rect -22652 -6092 -22588 -6028
rect -22652 -6172 -22588 -6108
rect -22652 -6252 -22588 -6188
rect -22652 -6332 -22588 -6268
rect -22652 -6412 -22588 -6348
rect -22652 -6492 -22588 -6428
rect -22652 -6572 -22588 -6508
rect -22652 -6652 -22588 -6588
rect -22652 -6732 -22588 -6668
rect -22652 -6812 -22588 -6748
rect -22652 -6892 -22588 -6828
rect -22652 -6972 -22588 -6908
rect -22652 -7052 -22588 -6988
rect -22652 -7132 -22588 -7068
rect -22652 -7212 -22588 -7148
rect -22652 -7292 -22588 -7228
rect -22652 -7372 -22588 -7308
rect -22652 -7452 -22588 -7388
rect -22652 -7532 -22588 -7468
rect -22652 -7612 -22588 -7548
rect -22652 -7692 -22588 -7628
rect -22652 -7772 -22588 -7708
rect -22652 -7852 -22588 -7788
rect -22652 -7932 -22588 -7868
rect -22652 -8012 -22588 -7948
rect -22652 -8092 -22588 -8028
rect -22652 -8172 -22588 -8108
rect -22652 -8252 -22588 -8188
rect -22652 -8332 -22588 -8268
rect -22652 -8412 -22588 -8348
rect -22652 -8492 -22588 -8428
rect -22652 -8572 -22588 -8508
rect -22652 -8652 -22588 -8588
rect -22652 -8732 -22588 -8668
rect -22652 -8812 -22588 -8748
rect -22652 -8892 -22588 -8828
rect -22652 -8972 -22588 -8908
rect -22652 -9052 -22588 -8988
rect -22652 -9132 -22588 -9068
rect -22652 -9212 -22588 -9148
rect -22652 -9292 -22588 -9228
rect -22652 -9372 -22588 -9308
rect -22652 -9452 -22588 -9388
rect -22652 -9532 -22588 -9468
rect -22652 -9612 -22588 -9548
rect -22652 -9692 -22588 -9628
rect -22652 -9772 -22588 -9708
rect -22652 -9852 -22588 -9788
rect -22652 -9932 -22588 -9868
rect -22652 -10012 -22588 -9948
rect -22652 -10092 -22588 -10028
rect -22652 -10172 -22588 -10108
rect -22652 -10252 -22588 -10188
rect -22652 -10332 -22588 -10268
rect -22652 -10412 -22588 -10348
rect -22652 -10492 -22588 -10428
rect -17040 -5532 -16976 -5468
rect -17040 -5612 -16976 -5548
rect -17040 -5692 -16976 -5628
rect -17040 -5772 -16976 -5708
rect -17040 -5852 -16976 -5788
rect -17040 -5932 -16976 -5868
rect -17040 -6012 -16976 -5948
rect -17040 -6092 -16976 -6028
rect -17040 -6172 -16976 -6108
rect -17040 -6252 -16976 -6188
rect -17040 -6332 -16976 -6268
rect -17040 -6412 -16976 -6348
rect -17040 -6492 -16976 -6428
rect -17040 -6572 -16976 -6508
rect -17040 -6652 -16976 -6588
rect -17040 -6732 -16976 -6668
rect -17040 -6812 -16976 -6748
rect -17040 -6892 -16976 -6828
rect -17040 -6972 -16976 -6908
rect -17040 -7052 -16976 -6988
rect -17040 -7132 -16976 -7068
rect -17040 -7212 -16976 -7148
rect -17040 -7292 -16976 -7228
rect -17040 -7372 -16976 -7308
rect -17040 -7452 -16976 -7388
rect -17040 -7532 -16976 -7468
rect -17040 -7612 -16976 -7548
rect -17040 -7692 -16976 -7628
rect -17040 -7772 -16976 -7708
rect -17040 -7852 -16976 -7788
rect -17040 -7932 -16976 -7868
rect -17040 -8012 -16976 -7948
rect -17040 -8092 -16976 -8028
rect -17040 -8172 -16976 -8108
rect -17040 -8252 -16976 -8188
rect -17040 -8332 -16976 -8268
rect -17040 -8412 -16976 -8348
rect -17040 -8492 -16976 -8428
rect -17040 -8572 -16976 -8508
rect -17040 -8652 -16976 -8588
rect -17040 -8732 -16976 -8668
rect -17040 -8812 -16976 -8748
rect -17040 -8892 -16976 -8828
rect -17040 -8972 -16976 -8908
rect -17040 -9052 -16976 -8988
rect -17040 -9132 -16976 -9068
rect -17040 -9212 -16976 -9148
rect -17040 -9292 -16976 -9228
rect -17040 -9372 -16976 -9308
rect -17040 -9452 -16976 -9388
rect -17040 -9532 -16976 -9468
rect -17040 -9612 -16976 -9548
rect -17040 -9692 -16976 -9628
rect -17040 -9772 -16976 -9708
rect -17040 -9852 -16976 -9788
rect -17040 -9932 -16976 -9868
rect -17040 -10012 -16976 -9948
rect -17040 -10092 -16976 -10028
rect -17040 -10172 -16976 -10108
rect -17040 -10252 -16976 -10188
rect -17040 -10332 -16976 -10268
rect -17040 -10412 -16976 -10348
rect -17040 -10492 -16976 -10428
rect -11428 -5532 -11364 -5468
rect -11428 -5612 -11364 -5548
rect -11428 -5692 -11364 -5628
rect -11428 -5772 -11364 -5708
rect -11428 -5852 -11364 -5788
rect -11428 -5932 -11364 -5868
rect -11428 -6012 -11364 -5948
rect -11428 -6092 -11364 -6028
rect -11428 -6172 -11364 -6108
rect -11428 -6252 -11364 -6188
rect -11428 -6332 -11364 -6268
rect -11428 -6412 -11364 -6348
rect -11428 -6492 -11364 -6428
rect -11428 -6572 -11364 -6508
rect -11428 -6652 -11364 -6588
rect -11428 -6732 -11364 -6668
rect -11428 -6812 -11364 -6748
rect -11428 -6892 -11364 -6828
rect -11428 -6972 -11364 -6908
rect -11428 -7052 -11364 -6988
rect -11428 -7132 -11364 -7068
rect -11428 -7212 -11364 -7148
rect -11428 -7292 -11364 -7228
rect -11428 -7372 -11364 -7308
rect -11428 -7452 -11364 -7388
rect -11428 -7532 -11364 -7468
rect -11428 -7612 -11364 -7548
rect -11428 -7692 -11364 -7628
rect -11428 -7772 -11364 -7708
rect -11428 -7852 -11364 -7788
rect -11428 -7932 -11364 -7868
rect -11428 -8012 -11364 -7948
rect -11428 -8092 -11364 -8028
rect -11428 -8172 -11364 -8108
rect -11428 -8252 -11364 -8188
rect -11428 -8332 -11364 -8268
rect -11428 -8412 -11364 -8348
rect -11428 -8492 -11364 -8428
rect -11428 -8572 -11364 -8508
rect -11428 -8652 -11364 -8588
rect -11428 -8732 -11364 -8668
rect -11428 -8812 -11364 -8748
rect -11428 -8892 -11364 -8828
rect -11428 -8972 -11364 -8908
rect -11428 -9052 -11364 -8988
rect -11428 -9132 -11364 -9068
rect -11428 -9212 -11364 -9148
rect -11428 -9292 -11364 -9228
rect -11428 -9372 -11364 -9308
rect -11428 -9452 -11364 -9388
rect -11428 -9532 -11364 -9468
rect -11428 -9612 -11364 -9548
rect -11428 -9692 -11364 -9628
rect -11428 -9772 -11364 -9708
rect -11428 -9852 -11364 -9788
rect -11428 -9932 -11364 -9868
rect -11428 -10012 -11364 -9948
rect -11428 -10092 -11364 -10028
rect -11428 -10172 -11364 -10108
rect -11428 -10252 -11364 -10188
rect -11428 -10332 -11364 -10268
rect -11428 -10412 -11364 -10348
rect -11428 -10492 -11364 -10428
rect -5816 -5532 -5752 -5468
rect -5816 -5612 -5752 -5548
rect -5816 -5692 -5752 -5628
rect -5816 -5772 -5752 -5708
rect -5816 -5852 -5752 -5788
rect -5816 -5932 -5752 -5868
rect -5816 -6012 -5752 -5948
rect -5816 -6092 -5752 -6028
rect -5816 -6172 -5752 -6108
rect -5816 -6252 -5752 -6188
rect -5816 -6332 -5752 -6268
rect -5816 -6412 -5752 -6348
rect -5816 -6492 -5752 -6428
rect -5816 -6572 -5752 -6508
rect -5816 -6652 -5752 -6588
rect -5816 -6732 -5752 -6668
rect -5816 -6812 -5752 -6748
rect -5816 -6892 -5752 -6828
rect -5816 -6972 -5752 -6908
rect -5816 -7052 -5752 -6988
rect -5816 -7132 -5752 -7068
rect -5816 -7212 -5752 -7148
rect -5816 -7292 -5752 -7228
rect -5816 -7372 -5752 -7308
rect -5816 -7452 -5752 -7388
rect -5816 -7532 -5752 -7468
rect -5816 -7612 -5752 -7548
rect -5816 -7692 -5752 -7628
rect -5816 -7772 -5752 -7708
rect -5816 -7852 -5752 -7788
rect -5816 -7932 -5752 -7868
rect -5816 -8012 -5752 -7948
rect -5816 -8092 -5752 -8028
rect -5816 -8172 -5752 -8108
rect -5816 -8252 -5752 -8188
rect -5816 -8332 -5752 -8268
rect -5816 -8412 -5752 -8348
rect -5816 -8492 -5752 -8428
rect -5816 -8572 -5752 -8508
rect -5816 -8652 -5752 -8588
rect -5816 -8732 -5752 -8668
rect -5816 -8812 -5752 -8748
rect -5816 -8892 -5752 -8828
rect -5816 -8972 -5752 -8908
rect -5816 -9052 -5752 -8988
rect -5816 -9132 -5752 -9068
rect -5816 -9212 -5752 -9148
rect -5816 -9292 -5752 -9228
rect -5816 -9372 -5752 -9308
rect -5816 -9452 -5752 -9388
rect -5816 -9532 -5752 -9468
rect -5816 -9612 -5752 -9548
rect -5816 -9692 -5752 -9628
rect -5816 -9772 -5752 -9708
rect -5816 -9852 -5752 -9788
rect -5816 -9932 -5752 -9868
rect -5816 -10012 -5752 -9948
rect -5816 -10092 -5752 -10028
rect -5816 -10172 -5752 -10108
rect -5816 -10252 -5752 -10188
rect -5816 -10332 -5752 -10268
rect -5816 -10412 -5752 -10348
rect -5816 -10492 -5752 -10428
rect -204 -5532 -140 -5468
rect -204 -5612 -140 -5548
rect -204 -5692 -140 -5628
rect -204 -5772 -140 -5708
rect -204 -5852 -140 -5788
rect -204 -5932 -140 -5868
rect -204 -6012 -140 -5948
rect -204 -6092 -140 -6028
rect -204 -6172 -140 -6108
rect -204 -6252 -140 -6188
rect -204 -6332 -140 -6268
rect -204 -6412 -140 -6348
rect -204 -6492 -140 -6428
rect -204 -6572 -140 -6508
rect -204 -6652 -140 -6588
rect -204 -6732 -140 -6668
rect -204 -6812 -140 -6748
rect -204 -6892 -140 -6828
rect -204 -6972 -140 -6908
rect -204 -7052 -140 -6988
rect -204 -7132 -140 -7068
rect -204 -7212 -140 -7148
rect -204 -7292 -140 -7228
rect -204 -7372 -140 -7308
rect -204 -7452 -140 -7388
rect -204 -7532 -140 -7468
rect -204 -7612 -140 -7548
rect -204 -7692 -140 -7628
rect -204 -7772 -140 -7708
rect -204 -7852 -140 -7788
rect -204 -7932 -140 -7868
rect -204 -8012 -140 -7948
rect -204 -8092 -140 -8028
rect -204 -8172 -140 -8108
rect -204 -8252 -140 -8188
rect -204 -8332 -140 -8268
rect -204 -8412 -140 -8348
rect -204 -8492 -140 -8428
rect -204 -8572 -140 -8508
rect -204 -8652 -140 -8588
rect -204 -8732 -140 -8668
rect -204 -8812 -140 -8748
rect -204 -8892 -140 -8828
rect -204 -8972 -140 -8908
rect -204 -9052 -140 -8988
rect -204 -9132 -140 -9068
rect -204 -9212 -140 -9148
rect -204 -9292 -140 -9228
rect -204 -9372 -140 -9308
rect -204 -9452 -140 -9388
rect -204 -9532 -140 -9468
rect -204 -9612 -140 -9548
rect -204 -9692 -140 -9628
rect -204 -9772 -140 -9708
rect -204 -9852 -140 -9788
rect -204 -9932 -140 -9868
rect -204 -10012 -140 -9948
rect -204 -10092 -140 -10028
rect -204 -10172 -140 -10108
rect -204 -10252 -140 -10188
rect -204 -10332 -140 -10268
rect -204 -10412 -140 -10348
rect -204 -10492 -140 -10428
rect 5408 -5532 5472 -5468
rect 5408 -5612 5472 -5548
rect 5408 -5692 5472 -5628
rect 5408 -5772 5472 -5708
rect 5408 -5852 5472 -5788
rect 5408 -5932 5472 -5868
rect 5408 -6012 5472 -5948
rect 5408 -6092 5472 -6028
rect 5408 -6172 5472 -6108
rect 5408 -6252 5472 -6188
rect 5408 -6332 5472 -6268
rect 5408 -6412 5472 -6348
rect 5408 -6492 5472 -6428
rect 5408 -6572 5472 -6508
rect 5408 -6652 5472 -6588
rect 5408 -6732 5472 -6668
rect 5408 -6812 5472 -6748
rect 5408 -6892 5472 -6828
rect 5408 -6972 5472 -6908
rect 5408 -7052 5472 -6988
rect 5408 -7132 5472 -7068
rect 5408 -7212 5472 -7148
rect 5408 -7292 5472 -7228
rect 5408 -7372 5472 -7308
rect 5408 -7452 5472 -7388
rect 5408 -7532 5472 -7468
rect 5408 -7612 5472 -7548
rect 5408 -7692 5472 -7628
rect 5408 -7772 5472 -7708
rect 5408 -7852 5472 -7788
rect 5408 -7932 5472 -7868
rect 5408 -8012 5472 -7948
rect 5408 -8092 5472 -8028
rect 5408 -8172 5472 -8108
rect 5408 -8252 5472 -8188
rect 5408 -8332 5472 -8268
rect 5408 -8412 5472 -8348
rect 5408 -8492 5472 -8428
rect 5408 -8572 5472 -8508
rect 5408 -8652 5472 -8588
rect 5408 -8732 5472 -8668
rect 5408 -8812 5472 -8748
rect 5408 -8892 5472 -8828
rect 5408 -8972 5472 -8908
rect 5408 -9052 5472 -8988
rect 5408 -9132 5472 -9068
rect 5408 -9212 5472 -9148
rect 5408 -9292 5472 -9228
rect 5408 -9372 5472 -9308
rect 5408 -9452 5472 -9388
rect 5408 -9532 5472 -9468
rect 5408 -9612 5472 -9548
rect 5408 -9692 5472 -9628
rect 5408 -9772 5472 -9708
rect 5408 -9852 5472 -9788
rect 5408 -9932 5472 -9868
rect 5408 -10012 5472 -9948
rect 5408 -10092 5472 -10028
rect 5408 -10172 5472 -10108
rect 5408 -10252 5472 -10188
rect 5408 -10332 5472 -10268
rect 5408 -10412 5472 -10348
rect 5408 -10492 5472 -10428
rect 11020 -5532 11084 -5468
rect 11020 -5612 11084 -5548
rect 11020 -5692 11084 -5628
rect 11020 -5772 11084 -5708
rect 11020 -5852 11084 -5788
rect 11020 -5932 11084 -5868
rect 11020 -6012 11084 -5948
rect 11020 -6092 11084 -6028
rect 11020 -6172 11084 -6108
rect 11020 -6252 11084 -6188
rect 11020 -6332 11084 -6268
rect 11020 -6412 11084 -6348
rect 11020 -6492 11084 -6428
rect 11020 -6572 11084 -6508
rect 11020 -6652 11084 -6588
rect 11020 -6732 11084 -6668
rect 11020 -6812 11084 -6748
rect 11020 -6892 11084 -6828
rect 11020 -6972 11084 -6908
rect 11020 -7052 11084 -6988
rect 11020 -7132 11084 -7068
rect 11020 -7212 11084 -7148
rect 11020 -7292 11084 -7228
rect 11020 -7372 11084 -7308
rect 11020 -7452 11084 -7388
rect 11020 -7532 11084 -7468
rect 11020 -7612 11084 -7548
rect 11020 -7692 11084 -7628
rect 11020 -7772 11084 -7708
rect 11020 -7852 11084 -7788
rect 11020 -7932 11084 -7868
rect 11020 -8012 11084 -7948
rect 11020 -8092 11084 -8028
rect 11020 -8172 11084 -8108
rect 11020 -8252 11084 -8188
rect 11020 -8332 11084 -8268
rect 11020 -8412 11084 -8348
rect 11020 -8492 11084 -8428
rect 11020 -8572 11084 -8508
rect 11020 -8652 11084 -8588
rect 11020 -8732 11084 -8668
rect 11020 -8812 11084 -8748
rect 11020 -8892 11084 -8828
rect 11020 -8972 11084 -8908
rect 11020 -9052 11084 -8988
rect 11020 -9132 11084 -9068
rect 11020 -9212 11084 -9148
rect 11020 -9292 11084 -9228
rect 11020 -9372 11084 -9308
rect 11020 -9452 11084 -9388
rect 11020 -9532 11084 -9468
rect 11020 -9612 11084 -9548
rect 11020 -9692 11084 -9628
rect 11020 -9772 11084 -9708
rect 11020 -9852 11084 -9788
rect 11020 -9932 11084 -9868
rect 11020 -10012 11084 -9948
rect 11020 -10092 11084 -10028
rect 11020 -10172 11084 -10108
rect 11020 -10252 11084 -10188
rect 11020 -10332 11084 -10268
rect 11020 -10412 11084 -10348
rect 11020 -10492 11084 -10428
rect 16632 -5532 16696 -5468
rect 16632 -5612 16696 -5548
rect 16632 -5692 16696 -5628
rect 16632 -5772 16696 -5708
rect 16632 -5852 16696 -5788
rect 16632 -5932 16696 -5868
rect 16632 -6012 16696 -5948
rect 16632 -6092 16696 -6028
rect 16632 -6172 16696 -6108
rect 16632 -6252 16696 -6188
rect 16632 -6332 16696 -6268
rect 16632 -6412 16696 -6348
rect 16632 -6492 16696 -6428
rect 16632 -6572 16696 -6508
rect 16632 -6652 16696 -6588
rect 16632 -6732 16696 -6668
rect 16632 -6812 16696 -6748
rect 16632 -6892 16696 -6828
rect 16632 -6972 16696 -6908
rect 16632 -7052 16696 -6988
rect 16632 -7132 16696 -7068
rect 16632 -7212 16696 -7148
rect 16632 -7292 16696 -7228
rect 16632 -7372 16696 -7308
rect 16632 -7452 16696 -7388
rect 16632 -7532 16696 -7468
rect 16632 -7612 16696 -7548
rect 16632 -7692 16696 -7628
rect 16632 -7772 16696 -7708
rect 16632 -7852 16696 -7788
rect 16632 -7932 16696 -7868
rect 16632 -8012 16696 -7948
rect 16632 -8092 16696 -8028
rect 16632 -8172 16696 -8108
rect 16632 -8252 16696 -8188
rect 16632 -8332 16696 -8268
rect 16632 -8412 16696 -8348
rect 16632 -8492 16696 -8428
rect 16632 -8572 16696 -8508
rect 16632 -8652 16696 -8588
rect 16632 -8732 16696 -8668
rect 16632 -8812 16696 -8748
rect 16632 -8892 16696 -8828
rect 16632 -8972 16696 -8908
rect 16632 -9052 16696 -8988
rect 16632 -9132 16696 -9068
rect 16632 -9212 16696 -9148
rect 16632 -9292 16696 -9228
rect 16632 -9372 16696 -9308
rect 16632 -9452 16696 -9388
rect 16632 -9532 16696 -9468
rect 16632 -9612 16696 -9548
rect 16632 -9692 16696 -9628
rect 16632 -9772 16696 -9708
rect 16632 -9852 16696 -9788
rect 16632 -9932 16696 -9868
rect 16632 -10012 16696 -9948
rect 16632 -10092 16696 -10028
rect 16632 -10172 16696 -10108
rect 16632 -10252 16696 -10188
rect 16632 -10332 16696 -10268
rect 16632 -10412 16696 -10348
rect 16632 -10492 16696 -10428
rect 22244 -5532 22308 -5468
rect 22244 -5612 22308 -5548
rect 22244 -5692 22308 -5628
rect 22244 -5772 22308 -5708
rect 22244 -5852 22308 -5788
rect 22244 -5932 22308 -5868
rect 22244 -6012 22308 -5948
rect 22244 -6092 22308 -6028
rect 22244 -6172 22308 -6108
rect 22244 -6252 22308 -6188
rect 22244 -6332 22308 -6268
rect 22244 -6412 22308 -6348
rect 22244 -6492 22308 -6428
rect 22244 -6572 22308 -6508
rect 22244 -6652 22308 -6588
rect 22244 -6732 22308 -6668
rect 22244 -6812 22308 -6748
rect 22244 -6892 22308 -6828
rect 22244 -6972 22308 -6908
rect 22244 -7052 22308 -6988
rect 22244 -7132 22308 -7068
rect 22244 -7212 22308 -7148
rect 22244 -7292 22308 -7228
rect 22244 -7372 22308 -7308
rect 22244 -7452 22308 -7388
rect 22244 -7532 22308 -7468
rect 22244 -7612 22308 -7548
rect 22244 -7692 22308 -7628
rect 22244 -7772 22308 -7708
rect 22244 -7852 22308 -7788
rect 22244 -7932 22308 -7868
rect 22244 -8012 22308 -7948
rect 22244 -8092 22308 -8028
rect 22244 -8172 22308 -8108
rect 22244 -8252 22308 -8188
rect 22244 -8332 22308 -8268
rect 22244 -8412 22308 -8348
rect 22244 -8492 22308 -8428
rect 22244 -8572 22308 -8508
rect 22244 -8652 22308 -8588
rect 22244 -8732 22308 -8668
rect 22244 -8812 22308 -8748
rect 22244 -8892 22308 -8828
rect 22244 -8972 22308 -8908
rect 22244 -9052 22308 -8988
rect 22244 -9132 22308 -9068
rect 22244 -9212 22308 -9148
rect 22244 -9292 22308 -9228
rect 22244 -9372 22308 -9308
rect 22244 -9452 22308 -9388
rect 22244 -9532 22308 -9468
rect 22244 -9612 22308 -9548
rect 22244 -9692 22308 -9628
rect 22244 -9772 22308 -9708
rect 22244 -9852 22308 -9788
rect 22244 -9932 22308 -9868
rect 22244 -10012 22308 -9948
rect 22244 -10092 22308 -10028
rect 22244 -10172 22308 -10108
rect 22244 -10252 22308 -10188
rect 22244 -10332 22308 -10268
rect 22244 -10412 22308 -10348
rect 22244 -10492 22308 -10428
rect 27856 -5532 27920 -5468
rect 27856 -5612 27920 -5548
rect 27856 -5692 27920 -5628
rect 27856 -5772 27920 -5708
rect 27856 -5852 27920 -5788
rect 27856 -5932 27920 -5868
rect 27856 -6012 27920 -5948
rect 27856 -6092 27920 -6028
rect 27856 -6172 27920 -6108
rect 27856 -6252 27920 -6188
rect 27856 -6332 27920 -6268
rect 27856 -6412 27920 -6348
rect 27856 -6492 27920 -6428
rect 27856 -6572 27920 -6508
rect 27856 -6652 27920 -6588
rect 27856 -6732 27920 -6668
rect 27856 -6812 27920 -6748
rect 27856 -6892 27920 -6828
rect 27856 -6972 27920 -6908
rect 27856 -7052 27920 -6988
rect 27856 -7132 27920 -7068
rect 27856 -7212 27920 -7148
rect 27856 -7292 27920 -7228
rect 27856 -7372 27920 -7308
rect 27856 -7452 27920 -7388
rect 27856 -7532 27920 -7468
rect 27856 -7612 27920 -7548
rect 27856 -7692 27920 -7628
rect 27856 -7772 27920 -7708
rect 27856 -7852 27920 -7788
rect 27856 -7932 27920 -7868
rect 27856 -8012 27920 -7948
rect 27856 -8092 27920 -8028
rect 27856 -8172 27920 -8108
rect 27856 -8252 27920 -8188
rect 27856 -8332 27920 -8268
rect 27856 -8412 27920 -8348
rect 27856 -8492 27920 -8428
rect 27856 -8572 27920 -8508
rect 27856 -8652 27920 -8588
rect 27856 -8732 27920 -8668
rect 27856 -8812 27920 -8748
rect 27856 -8892 27920 -8828
rect 27856 -8972 27920 -8908
rect 27856 -9052 27920 -8988
rect 27856 -9132 27920 -9068
rect 27856 -9212 27920 -9148
rect 27856 -9292 27920 -9228
rect 27856 -9372 27920 -9308
rect 27856 -9452 27920 -9388
rect 27856 -9532 27920 -9468
rect 27856 -9612 27920 -9548
rect 27856 -9692 27920 -9628
rect 27856 -9772 27920 -9708
rect 27856 -9852 27920 -9788
rect 27856 -9932 27920 -9868
rect 27856 -10012 27920 -9948
rect 27856 -10092 27920 -10028
rect 27856 -10172 27920 -10108
rect 27856 -10252 27920 -10188
rect 27856 -10332 27920 -10268
rect 27856 -10412 27920 -10348
rect 27856 -10492 27920 -10428
rect 33468 -5532 33532 -5468
rect 33468 -5612 33532 -5548
rect 33468 -5692 33532 -5628
rect 33468 -5772 33532 -5708
rect 33468 -5852 33532 -5788
rect 33468 -5932 33532 -5868
rect 33468 -6012 33532 -5948
rect 33468 -6092 33532 -6028
rect 33468 -6172 33532 -6108
rect 33468 -6252 33532 -6188
rect 33468 -6332 33532 -6268
rect 33468 -6412 33532 -6348
rect 33468 -6492 33532 -6428
rect 33468 -6572 33532 -6508
rect 33468 -6652 33532 -6588
rect 33468 -6732 33532 -6668
rect 33468 -6812 33532 -6748
rect 33468 -6892 33532 -6828
rect 33468 -6972 33532 -6908
rect 33468 -7052 33532 -6988
rect 33468 -7132 33532 -7068
rect 33468 -7212 33532 -7148
rect 33468 -7292 33532 -7228
rect 33468 -7372 33532 -7308
rect 33468 -7452 33532 -7388
rect 33468 -7532 33532 -7468
rect 33468 -7612 33532 -7548
rect 33468 -7692 33532 -7628
rect 33468 -7772 33532 -7708
rect 33468 -7852 33532 -7788
rect 33468 -7932 33532 -7868
rect 33468 -8012 33532 -7948
rect 33468 -8092 33532 -8028
rect 33468 -8172 33532 -8108
rect 33468 -8252 33532 -8188
rect 33468 -8332 33532 -8268
rect 33468 -8412 33532 -8348
rect 33468 -8492 33532 -8428
rect 33468 -8572 33532 -8508
rect 33468 -8652 33532 -8588
rect 33468 -8732 33532 -8668
rect 33468 -8812 33532 -8748
rect 33468 -8892 33532 -8828
rect 33468 -8972 33532 -8908
rect 33468 -9052 33532 -8988
rect 33468 -9132 33532 -9068
rect 33468 -9212 33532 -9148
rect 33468 -9292 33532 -9228
rect 33468 -9372 33532 -9308
rect 33468 -9452 33532 -9388
rect 33468 -9532 33532 -9468
rect 33468 -9612 33532 -9548
rect 33468 -9692 33532 -9628
rect 33468 -9772 33532 -9708
rect 33468 -9852 33532 -9788
rect 33468 -9932 33532 -9868
rect 33468 -10012 33532 -9948
rect 33468 -10092 33532 -10028
rect 33468 -10172 33532 -10108
rect 33468 -10252 33532 -10188
rect 33468 -10332 33532 -10268
rect 33468 -10412 33532 -10348
rect 33468 -10492 33532 -10428
rect 39080 -5532 39144 -5468
rect 39080 -5612 39144 -5548
rect 39080 -5692 39144 -5628
rect 39080 -5772 39144 -5708
rect 39080 -5852 39144 -5788
rect 39080 -5932 39144 -5868
rect 39080 -6012 39144 -5948
rect 39080 -6092 39144 -6028
rect 39080 -6172 39144 -6108
rect 39080 -6252 39144 -6188
rect 39080 -6332 39144 -6268
rect 39080 -6412 39144 -6348
rect 39080 -6492 39144 -6428
rect 39080 -6572 39144 -6508
rect 39080 -6652 39144 -6588
rect 39080 -6732 39144 -6668
rect 39080 -6812 39144 -6748
rect 39080 -6892 39144 -6828
rect 39080 -6972 39144 -6908
rect 39080 -7052 39144 -6988
rect 39080 -7132 39144 -7068
rect 39080 -7212 39144 -7148
rect 39080 -7292 39144 -7228
rect 39080 -7372 39144 -7308
rect 39080 -7452 39144 -7388
rect 39080 -7532 39144 -7468
rect 39080 -7612 39144 -7548
rect 39080 -7692 39144 -7628
rect 39080 -7772 39144 -7708
rect 39080 -7852 39144 -7788
rect 39080 -7932 39144 -7868
rect 39080 -8012 39144 -7948
rect 39080 -8092 39144 -8028
rect 39080 -8172 39144 -8108
rect 39080 -8252 39144 -8188
rect 39080 -8332 39144 -8268
rect 39080 -8412 39144 -8348
rect 39080 -8492 39144 -8428
rect 39080 -8572 39144 -8508
rect 39080 -8652 39144 -8588
rect 39080 -8732 39144 -8668
rect 39080 -8812 39144 -8748
rect 39080 -8892 39144 -8828
rect 39080 -8972 39144 -8908
rect 39080 -9052 39144 -8988
rect 39080 -9132 39144 -9068
rect 39080 -9212 39144 -9148
rect 39080 -9292 39144 -9228
rect 39080 -9372 39144 -9308
rect 39080 -9452 39144 -9388
rect 39080 -9532 39144 -9468
rect 39080 -9612 39144 -9548
rect 39080 -9692 39144 -9628
rect 39080 -9772 39144 -9708
rect 39080 -9852 39144 -9788
rect 39080 -9932 39144 -9868
rect 39080 -10012 39144 -9948
rect 39080 -10092 39144 -10028
rect 39080 -10172 39144 -10108
rect 39080 -10252 39144 -10188
rect 39080 -10332 39144 -10268
rect 39080 -10412 39144 -10348
rect 39080 -10492 39144 -10428
rect -33876 -10852 -33812 -10788
rect -33876 -10932 -33812 -10868
rect -33876 -11012 -33812 -10948
rect -33876 -11092 -33812 -11028
rect -33876 -11172 -33812 -11108
rect -33876 -11252 -33812 -11188
rect -33876 -11332 -33812 -11268
rect -33876 -11412 -33812 -11348
rect -33876 -11492 -33812 -11428
rect -33876 -11572 -33812 -11508
rect -33876 -11652 -33812 -11588
rect -33876 -11732 -33812 -11668
rect -33876 -11812 -33812 -11748
rect -33876 -11892 -33812 -11828
rect -33876 -11972 -33812 -11908
rect -33876 -12052 -33812 -11988
rect -33876 -12132 -33812 -12068
rect -33876 -12212 -33812 -12148
rect -33876 -12292 -33812 -12228
rect -33876 -12372 -33812 -12308
rect -33876 -12452 -33812 -12388
rect -33876 -12532 -33812 -12468
rect -33876 -12612 -33812 -12548
rect -33876 -12692 -33812 -12628
rect -33876 -12772 -33812 -12708
rect -33876 -12852 -33812 -12788
rect -33876 -12932 -33812 -12868
rect -33876 -13012 -33812 -12948
rect -33876 -13092 -33812 -13028
rect -33876 -13172 -33812 -13108
rect -33876 -13252 -33812 -13188
rect -33876 -13332 -33812 -13268
rect -33876 -13412 -33812 -13348
rect -33876 -13492 -33812 -13428
rect -33876 -13572 -33812 -13508
rect -33876 -13652 -33812 -13588
rect -33876 -13732 -33812 -13668
rect -33876 -13812 -33812 -13748
rect -33876 -13892 -33812 -13828
rect -33876 -13972 -33812 -13908
rect -33876 -14052 -33812 -13988
rect -33876 -14132 -33812 -14068
rect -33876 -14212 -33812 -14148
rect -33876 -14292 -33812 -14228
rect -33876 -14372 -33812 -14308
rect -33876 -14452 -33812 -14388
rect -33876 -14532 -33812 -14468
rect -33876 -14612 -33812 -14548
rect -33876 -14692 -33812 -14628
rect -33876 -14772 -33812 -14708
rect -33876 -14852 -33812 -14788
rect -33876 -14932 -33812 -14868
rect -33876 -15012 -33812 -14948
rect -33876 -15092 -33812 -15028
rect -33876 -15172 -33812 -15108
rect -33876 -15252 -33812 -15188
rect -33876 -15332 -33812 -15268
rect -33876 -15412 -33812 -15348
rect -33876 -15492 -33812 -15428
rect -33876 -15572 -33812 -15508
rect -33876 -15652 -33812 -15588
rect -33876 -15732 -33812 -15668
rect -33876 -15812 -33812 -15748
rect -28264 -10852 -28200 -10788
rect -28264 -10932 -28200 -10868
rect -28264 -11012 -28200 -10948
rect -28264 -11092 -28200 -11028
rect -28264 -11172 -28200 -11108
rect -28264 -11252 -28200 -11188
rect -28264 -11332 -28200 -11268
rect -28264 -11412 -28200 -11348
rect -28264 -11492 -28200 -11428
rect -28264 -11572 -28200 -11508
rect -28264 -11652 -28200 -11588
rect -28264 -11732 -28200 -11668
rect -28264 -11812 -28200 -11748
rect -28264 -11892 -28200 -11828
rect -28264 -11972 -28200 -11908
rect -28264 -12052 -28200 -11988
rect -28264 -12132 -28200 -12068
rect -28264 -12212 -28200 -12148
rect -28264 -12292 -28200 -12228
rect -28264 -12372 -28200 -12308
rect -28264 -12452 -28200 -12388
rect -28264 -12532 -28200 -12468
rect -28264 -12612 -28200 -12548
rect -28264 -12692 -28200 -12628
rect -28264 -12772 -28200 -12708
rect -28264 -12852 -28200 -12788
rect -28264 -12932 -28200 -12868
rect -28264 -13012 -28200 -12948
rect -28264 -13092 -28200 -13028
rect -28264 -13172 -28200 -13108
rect -28264 -13252 -28200 -13188
rect -28264 -13332 -28200 -13268
rect -28264 -13412 -28200 -13348
rect -28264 -13492 -28200 -13428
rect -28264 -13572 -28200 -13508
rect -28264 -13652 -28200 -13588
rect -28264 -13732 -28200 -13668
rect -28264 -13812 -28200 -13748
rect -28264 -13892 -28200 -13828
rect -28264 -13972 -28200 -13908
rect -28264 -14052 -28200 -13988
rect -28264 -14132 -28200 -14068
rect -28264 -14212 -28200 -14148
rect -28264 -14292 -28200 -14228
rect -28264 -14372 -28200 -14308
rect -28264 -14452 -28200 -14388
rect -28264 -14532 -28200 -14468
rect -28264 -14612 -28200 -14548
rect -28264 -14692 -28200 -14628
rect -28264 -14772 -28200 -14708
rect -28264 -14852 -28200 -14788
rect -28264 -14932 -28200 -14868
rect -28264 -15012 -28200 -14948
rect -28264 -15092 -28200 -15028
rect -28264 -15172 -28200 -15108
rect -28264 -15252 -28200 -15188
rect -28264 -15332 -28200 -15268
rect -28264 -15412 -28200 -15348
rect -28264 -15492 -28200 -15428
rect -28264 -15572 -28200 -15508
rect -28264 -15652 -28200 -15588
rect -28264 -15732 -28200 -15668
rect -28264 -15812 -28200 -15748
rect -22652 -10852 -22588 -10788
rect -22652 -10932 -22588 -10868
rect -22652 -11012 -22588 -10948
rect -22652 -11092 -22588 -11028
rect -22652 -11172 -22588 -11108
rect -22652 -11252 -22588 -11188
rect -22652 -11332 -22588 -11268
rect -22652 -11412 -22588 -11348
rect -22652 -11492 -22588 -11428
rect -22652 -11572 -22588 -11508
rect -22652 -11652 -22588 -11588
rect -22652 -11732 -22588 -11668
rect -22652 -11812 -22588 -11748
rect -22652 -11892 -22588 -11828
rect -22652 -11972 -22588 -11908
rect -22652 -12052 -22588 -11988
rect -22652 -12132 -22588 -12068
rect -22652 -12212 -22588 -12148
rect -22652 -12292 -22588 -12228
rect -22652 -12372 -22588 -12308
rect -22652 -12452 -22588 -12388
rect -22652 -12532 -22588 -12468
rect -22652 -12612 -22588 -12548
rect -22652 -12692 -22588 -12628
rect -22652 -12772 -22588 -12708
rect -22652 -12852 -22588 -12788
rect -22652 -12932 -22588 -12868
rect -22652 -13012 -22588 -12948
rect -22652 -13092 -22588 -13028
rect -22652 -13172 -22588 -13108
rect -22652 -13252 -22588 -13188
rect -22652 -13332 -22588 -13268
rect -22652 -13412 -22588 -13348
rect -22652 -13492 -22588 -13428
rect -22652 -13572 -22588 -13508
rect -22652 -13652 -22588 -13588
rect -22652 -13732 -22588 -13668
rect -22652 -13812 -22588 -13748
rect -22652 -13892 -22588 -13828
rect -22652 -13972 -22588 -13908
rect -22652 -14052 -22588 -13988
rect -22652 -14132 -22588 -14068
rect -22652 -14212 -22588 -14148
rect -22652 -14292 -22588 -14228
rect -22652 -14372 -22588 -14308
rect -22652 -14452 -22588 -14388
rect -22652 -14532 -22588 -14468
rect -22652 -14612 -22588 -14548
rect -22652 -14692 -22588 -14628
rect -22652 -14772 -22588 -14708
rect -22652 -14852 -22588 -14788
rect -22652 -14932 -22588 -14868
rect -22652 -15012 -22588 -14948
rect -22652 -15092 -22588 -15028
rect -22652 -15172 -22588 -15108
rect -22652 -15252 -22588 -15188
rect -22652 -15332 -22588 -15268
rect -22652 -15412 -22588 -15348
rect -22652 -15492 -22588 -15428
rect -22652 -15572 -22588 -15508
rect -22652 -15652 -22588 -15588
rect -22652 -15732 -22588 -15668
rect -22652 -15812 -22588 -15748
rect -17040 -10852 -16976 -10788
rect -17040 -10932 -16976 -10868
rect -17040 -11012 -16976 -10948
rect -17040 -11092 -16976 -11028
rect -17040 -11172 -16976 -11108
rect -17040 -11252 -16976 -11188
rect -17040 -11332 -16976 -11268
rect -17040 -11412 -16976 -11348
rect -17040 -11492 -16976 -11428
rect -17040 -11572 -16976 -11508
rect -17040 -11652 -16976 -11588
rect -17040 -11732 -16976 -11668
rect -17040 -11812 -16976 -11748
rect -17040 -11892 -16976 -11828
rect -17040 -11972 -16976 -11908
rect -17040 -12052 -16976 -11988
rect -17040 -12132 -16976 -12068
rect -17040 -12212 -16976 -12148
rect -17040 -12292 -16976 -12228
rect -17040 -12372 -16976 -12308
rect -17040 -12452 -16976 -12388
rect -17040 -12532 -16976 -12468
rect -17040 -12612 -16976 -12548
rect -17040 -12692 -16976 -12628
rect -17040 -12772 -16976 -12708
rect -17040 -12852 -16976 -12788
rect -17040 -12932 -16976 -12868
rect -17040 -13012 -16976 -12948
rect -17040 -13092 -16976 -13028
rect -17040 -13172 -16976 -13108
rect -17040 -13252 -16976 -13188
rect -17040 -13332 -16976 -13268
rect -17040 -13412 -16976 -13348
rect -17040 -13492 -16976 -13428
rect -17040 -13572 -16976 -13508
rect -17040 -13652 -16976 -13588
rect -17040 -13732 -16976 -13668
rect -17040 -13812 -16976 -13748
rect -17040 -13892 -16976 -13828
rect -17040 -13972 -16976 -13908
rect -17040 -14052 -16976 -13988
rect -17040 -14132 -16976 -14068
rect -17040 -14212 -16976 -14148
rect -17040 -14292 -16976 -14228
rect -17040 -14372 -16976 -14308
rect -17040 -14452 -16976 -14388
rect -17040 -14532 -16976 -14468
rect -17040 -14612 -16976 -14548
rect -17040 -14692 -16976 -14628
rect -17040 -14772 -16976 -14708
rect -17040 -14852 -16976 -14788
rect -17040 -14932 -16976 -14868
rect -17040 -15012 -16976 -14948
rect -17040 -15092 -16976 -15028
rect -17040 -15172 -16976 -15108
rect -17040 -15252 -16976 -15188
rect -17040 -15332 -16976 -15268
rect -17040 -15412 -16976 -15348
rect -17040 -15492 -16976 -15428
rect -17040 -15572 -16976 -15508
rect -17040 -15652 -16976 -15588
rect -17040 -15732 -16976 -15668
rect -17040 -15812 -16976 -15748
rect -11428 -10852 -11364 -10788
rect -11428 -10932 -11364 -10868
rect -11428 -11012 -11364 -10948
rect -11428 -11092 -11364 -11028
rect -11428 -11172 -11364 -11108
rect -11428 -11252 -11364 -11188
rect -11428 -11332 -11364 -11268
rect -11428 -11412 -11364 -11348
rect -11428 -11492 -11364 -11428
rect -11428 -11572 -11364 -11508
rect -11428 -11652 -11364 -11588
rect -11428 -11732 -11364 -11668
rect -11428 -11812 -11364 -11748
rect -11428 -11892 -11364 -11828
rect -11428 -11972 -11364 -11908
rect -11428 -12052 -11364 -11988
rect -11428 -12132 -11364 -12068
rect -11428 -12212 -11364 -12148
rect -11428 -12292 -11364 -12228
rect -11428 -12372 -11364 -12308
rect -11428 -12452 -11364 -12388
rect -11428 -12532 -11364 -12468
rect -11428 -12612 -11364 -12548
rect -11428 -12692 -11364 -12628
rect -11428 -12772 -11364 -12708
rect -11428 -12852 -11364 -12788
rect -11428 -12932 -11364 -12868
rect -11428 -13012 -11364 -12948
rect -11428 -13092 -11364 -13028
rect -11428 -13172 -11364 -13108
rect -11428 -13252 -11364 -13188
rect -11428 -13332 -11364 -13268
rect -11428 -13412 -11364 -13348
rect -11428 -13492 -11364 -13428
rect -11428 -13572 -11364 -13508
rect -11428 -13652 -11364 -13588
rect -11428 -13732 -11364 -13668
rect -11428 -13812 -11364 -13748
rect -11428 -13892 -11364 -13828
rect -11428 -13972 -11364 -13908
rect -11428 -14052 -11364 -13988
rect -11428 -14132 -11364 -14068
rect -11428 -14212 -11364 -14148
rect -11428 -14292 -11364 -14228
rect -11428 -14372 -11364 -14308
rect -11428 -14452 -11364 -14388
rect -11428 -14532 -11364 -14468
rect -11428 -14612 -11364 -14548
rect -11428 -14692 -11364 -14628
rect -11428 -14772 -11364 -14708
rect -11428 -14852 -11364 -14788
rect -11428 -14932 -11364 -14868
rect -11428 -15012 -11364 -14948
rect -11428 -15092 -11364 -15028
rect -11428 -15172 -11364 -15108
rect -11428 -15252 -11364 -15188
rect -11428 -15332 -11364 -15268
rect -11428 -15412 -11364 -15348
rect -11428 -15492 -11364 -15428
rect -11428 -15572 -11364 -15508
rect -11428 -15652 -11364 -15588
rect -11428 -15732 -11364 -15668
rect -11428 -15812 -11364 -15748
rect -5816 -10852 -5752 -10788
rect -5816 -10932 -5752 -10868
rect -5816 -11012 -5752 -10948
rect -5816 -11092 -5752 -11028
rect -5816 -11172 -5752 -11108
rect -5816 -11252 -5752 -11188
rect -5816 -11332 -5752 -11268
rect -5816 -11412 -5752 -11348
rect -5816 -11492 -5752 -11428
rect -5816 -11572 -5752 -11508
rect -5816 -11652 -5752 -11588
rect -5816 -11732 -5752 -11668
rect -5816 -11812 -5752 -11748
rect -5816 -11892 -5752 -11828
rect -5816 -11972 -5752 -11908
rect -5816 -12052 -5752 -11988
rect -5816 -12132 -5752 -12068
rect -5816 -12212 -5752 -12148
rect -5816 -12292 -5752 -12228
rect -5816 -12372 -5752 -12308
rect -5816 -12452 -5752 -12388
rect -5816 -12532 -5752 -12468
rect -5816 -12612 -5752 -12548
rect -5816 -12692 -5752 -12628
rect -5816 -12772 -5752 -12708
rect -5816 -12852 -5752 -12788
rect -5816 -12932 -5752 -12868
rect -5816 -13012 -5752 -12948
rect -5816 -13092 -5752 -13028
rect -5816 -13172 -5752 -13108
rect -5816 -13252 -5752 -13188
rect -5816 -13332 -5752 -13268
rect -5816 -13412 -5752 -13348
rect -5816 -13492 -5752 -13428
rect -5816 -13572 -5752 -13508
rect -5816 -13652 -5752 -13588
rect -5816 -13732 -5752 -13668
rect -5816 -13812 -5752 -13748
rect -5816 -13892 -5752 -13828
rect -5816 -13972 -5752 -13908
rect -5816 -14052 -5752 -13988
rect -5816 -14132 -5752 -14068
rect -5816 -14212 -5752 -14148
rect -5816 -14292 -5752 -14228
rect -5816 -14372 -5752 -14308
rect -5816 -14452 -5752 -14388
rect -5816 -14532 -5752 -14468
rect -5816 -14612 -5752 -14548
rect -5816 -14692 -5752 -14628
rect -5816 -14772 -5752 -14708
rect -5816 -14852 -5752 -14788
rect -5816 -14932 -5752 -14868
rect -5816 -15012 -5752 -14948
rect -5816 -15092 -5752 -15028
rect -5816 -15172 -5752 -15108
rect -5816 -15252 -5752 -15188
rect -5816 -15332 -5752 -15268
rect -5816 -15412 -5752 -15348
rect -5816 -15492 -5752 -15428
rect -5816 -15572 -5752 -15508
rect -5816 -15652 -5752 -15588
rect -5816 -15732 -5752 -15668
rect -5816 -15812 -5752 -15748
rect -204 -10852 -140 -10788
rect -204 -10932 -140 -10868
rect -204 -11012 -140 -10948
rect -204 -11092 -140 -11028
rect -204 -11172 -140 -11108
rect -204 -11252 -140 -11188
rect -204 -11332 -140 -11268
rect -204 -11412 -140 -11348
rect -204 -11492 -140 -11428
rect -204 -11572 -140 -11508
rect -204 -11652 -140 -11588
rect -204 -11732 -140 -11668
rect -204 -11812 -140 -11748
rect -204 -11892 -140 -11828
rect -204 -11972 -140 -11908
rect -204 -12052 -140 -11988
rect -204 -12132 -140 -12068
rect -204 -12212 -140 -12148
rect -204 -12292 -140 -12228
rect -204 -12372 -140 -12308
rect -204 -12452 -140 -12388
rect -204 -12532 -140 -12468
rect -204 -12612 -140 -12548
rect -204 -12692 -140 -12628
rect -204 -12772 -140 -12708
rect -204 -12852 -140 -12788
rect -204 -12932 -140 -12868
rect -204 -13012 -140 -12948
rect -204 -13092 -140 -13028
rect -204 -13172 -140 -13108
rect -204 -13252 -140 -13188
rect -204 -13332 -140 -13268
rect -204 -13412 -140 -13348
rect -204 -13492 -140 -13428
rect -204 -13572 -140 -13508
rect -204 -13652 -140 -13588
rect -204 -13732 -140 -13668
rect -204 -13812 -140 -13748
rect -204 -13892 -140 -13828
rect -204 -13972 -140 -13908
rect -204 -14052 -140 -13988
rect -204 -14132 -140 -14068
rect -204 -14212 -140 -14148
rect -204 -14292 -140 -14228
rect -204 -14372 -140 -14308
rect -204 -14452 -140 -14388
rect -204 -14532 -140 -14468
rect -204 -14612 -140 -14548
rect -204 -14692 -140 -14628
rect -204 -14772 -140 -14708
rect -204 -14852 -140 -14788
rect -204 -14932 -140 -14868
rect -204 -15012 -140 -14948
rect -204 -15092 -140 -15028
rect -204 -15172 -140 -15108
rect -204 -15252 -140 -15188
rect -204 -15332 -140 -15268
rect -204 -15412 -140 -15348
rect -204 -15492 -140 -15428
rect -204 -15572 -140 -15508
rect -204 -15652 -140 -15588
rect -204 -15732 -140 -15668
rect -204 -15812 -140 -15748
rect 5408 -10852 5472 -10788
rect 5408 -10932 5472 -10868
rect 5408 -11012 5472 -10948
rect 5408 -11092 5472 -11028
rect 5408 -11172 5472 -11108
rect 5408 -11252 5472 -11188
rect 5408 -11332 5472 -11268
rect 5408 -11412 5472 -11348
rect 5408 -11492 5472 -11428
rect 5408 -11572 5472 -11508
rect 5408 -11652 5472 -11588
rect 5408 -11732 5472 -11668
rect 5408 -11812 5472 -11748
rect 5408 -11892 5472 -11828
rect 5408 -11972 5472 -11908
rect 5408 -12052 5472 -11988
rect 5408 -12132 5472 -12068
rect 5408 -12212 5472 -12148
rect 5408 -12292 5472 -12228
rect 5408 -12372 5472 -12308
rect 5408 -12452 5472 -12388
rect 5408 -12532 5472 -12468
rect 5408 -12612 5472 -12548
rect 5408 -12692 5472 -12628
rect 5408 -12772 5472 -12708
rect 5408 -12852 5472 -12788
rect 5408 -12932 5472 -12868
rect 5408 -13012 5472 -12948
rect 5408 -13092 5472 -13028
rect 5408 -13172 5472 -13108
rect 5408 -13252 5472 -13188
rect 5408 -13332 5472 -13268
rect 5408 -13412 5472 -13348
rect 5408 -13492 5472 -13428
rect 5408 -13572 5472 -13508
rect 5408 -13652 5472 -13588
rect 5408 -13732 5472 -13668
rect 5408 -13812 5472 -13748
rect 5408 -13892 5472 -13828
rect 5408 -13972 5472 -13908
rect 5408 -14052 5472 -13988
rect 5408 -14132 5472 -14068
rect 5408 -14212 5472 -14148
rect 5408 -14292 5472 -14228
rect 5408 -14372 5472 -14308
rect 5408 -14452 5472 -14388
rect 5408 -14532 5472 -14468
rect 5408 -14612 5472 -14548
rect 5408 -14692 5472 -14628
rect 5408 -14772 5472 -14708
rect 5408 -14852 5472 -14788
rect 5408 -14932 5472 -14868
rect 5408 -15012 5472 -14948
rect 5408 -15092 5472 -15028
rect 5408 -15172 5472 -15108
rect 5408 -15252 5472 -15188
rect 5408 -15332 5472 -15268
rect 5408 -15412 5472 -15348
rect 5408 -15492 5472 -15428
rect 5408 -15572 5472 -15508
rect 5408 -15652 5472 -15588
rect 5408 -15732 5472 -15668
rect 5408 -15812 5472 -15748
rect 11020 -10852 11084 -10788
rect 11020 -10932 11084 -10868
rect 11020 -11012 11084 -10948
rect 11020 -11092 11084 -11028
rect 11020 -11172 11084 -11108
rect 11020 -11252 11084 -11188
rect 11020 -11332 11084 -11268
rect 11020 -11412 11084 -11348
rect 11020 -11492 11084 -11428
rect 11020 -11572 11084 -11508
rect 11020 -11652 11084 -11588
rect 11020 -11732 11084 -11668
rect 11020 -11812 11084 -11748
rect 11020 -11892 11084 -11828
rect 11020 -11972 11084 -11908
rect 11020 -12052 11084 -11988
rect 11020 -12132 11084 -12068
rect 11020 -12212 11084 -12148
rect 11020 -12292 11084 -12228
rect 11020 -12372 11084 -12308
rect 11020 -12452 11084 -12388
rect 11020 -12532 11084 -12468
rect 11020 -12612 11084 -12548
rect 11020 -12692 11084 -12628
rect 11020 -12772 11084 -12708
rect 11020 -12852 11084 -12788
rect 11020 -12932 11084 -12868
rect 11020 -13012 11084 -12948
rect 11020 -13092 11084 -13028
rect 11020 -13172 11084 -13108
rect 11020 -13252 11084 -13188
rect 11020 -13332 11084 -13268
rect 11020 -13412 11084 -13348
rect 11020 -13492 11084 -13428
rect 11020 -13572 11084 -13508
rect 11020 -13652 11084 -13588
rect 11020 -13732 11084 -13668
rect 11020 -13812 11084 -13748
rect 11020 -13892 11084 -13828
rect 11020 -13972 11084 -13908
rect 11020 -14052 11084 -13988
rect 11020 -14132 11084 -14068
rect 11020 -14212 11084 -14148
rect 11020 -14292 11084 -14228
rect 11020 -14372 11084 -14308
rect 11020 -14452 11084 -14388
rect 11020 -14532 11084 -14468
rect 11020 -14612 11084 -14548
rect 11020 -14692 11084 -14628
rect 11020 -14772 11084 -14708
rect 11020 -14852 11084 -14788
rect 11020 -14932 11084 -14868
rect 11020 -15012 11084 -14948
rect 11020 -15092 11084 -15028
rect 11020 -15172 11084 -15108
rect 11020 -15252 11084 -15188
rect 11020 -15332 11084 -15268
rect 11020 -15412 11084 -15348
rect 11020 -15492 11084 -15428
rect 11020 -15572 11084 -15508
rect 11020 -15652 11084 -15588
rect 11020 -15732 11084 -15668
rect 11020 -15812 11084 -15748
rect 16632 -10852 16696 -10788
rect 16632 -10932 16696 -10868
rect 16632 -11012 16696 -10948
rect 16632 -11092 16696 -11028
rect 16632 -11172 16696 -11108
rect 16632 -11252 16696 -11188
rect 16632 -11332 16696 -11268
rect 16632 -11412 16696 -11348
rect 16632 -11492 16696 -11428
rect 16632 -11572 16696 -11508
rect 16632 -11652 16696 -11588
rect 16632 -11732 16696 -11668
rect 16632 -11812 16696 -11748
rect 16632 -11892 16696 -11828
rect 16632 -11972 16696 -11908
rect 16632 -12052 16696 -11988
rect 16632 -12132 16696 -12068
rect 16632 -12212 16696 -12148
rect 16632 -12292 16696 -12228
rect 16632 -12372 16696 -12308
rect 16632 -12452 16696 -12388
rect 16632 -12532 16696 -12468
rect 16632 -12612 16696 -12548
rect 16632 -12692 16696 -12628
rect 16632 -12772 16696 -12708
rect 16632 -12852 16696 -12788
rect 16632 -12932 16696 -12868
rect 16632 -13012 16696 -12948
rect 16632 -13092 16696 -13028
rect 16632 -13172 16696 -13108
rect 16632 -13252 16696 -13188
rect 16632 -13332 16696 -13268
rect 16632 -13412 16696 -13348
rect 16632 -13492 16696 -13428
rect 16632 -13572 16696 -13508
rect 16632 -13652 16696 -13588
rect 16632 -13732 16696 -13668
rect 16632 -13812 16696 -13748
rect 16632 -13892 16696 -13828
rect 16632 -13972 16696 -13908
rect 16632 -14052 16696 -13988
rect 16632 -14132 16696 -14068
rect 16632 -14212 16696 -14148
rect 16632 -14292 16696 -14228
rect 16632 -14372 16696 -14308
rect 16632 -14452 16696 -14388
rect 16632 -14532 16696 -14468
rect 16632 -14612 16696 -14548
rect 16632 -14692 16696 -14628
rect 16632 -14772 16696 -14708
rect 16632 -14852 16696 -14788
rect 16632 -14932 16696 -14868
rect 16632 -15012 16696 -14948
rect 16632 -15092 16696 -15028
rect 16632 -15172 16696 -15108
rect 16632 -15252 16696 -15188
rect 16632 -15332 16696 -15268
rect 16632 -15412 16696 -15348
rect 16632 -15492 16696 -15428
rect 16632 -15572 16696 -15508
rect 16632 -15652 16696 -15588
rect 16632 -15732 16696 -15668
rect 16632 -15812 16696 -15748
rect 22244 -10852 22308 -10788
rect 22244 -10932 22308 -10868
rect 22244 -11012 22308 -10948
rect 22244 -11092 22308 -11028
rect 22244 -11172 22308 -11108
rect 22244 -11252 22308 -11188
rect 22244 -11332 22308 -11268
rect 22244 -11412 22308 -11348
rect 22244 -11492 22308 -11428
rect 22244 -11572 22308 -11508
rect 22244 -11652 22308 -11588
rect 22244 -11732 22308 -11668
rect 22244 -11812 22308 -11748
rect 22244 -11892 22308 -11828
rect 22244 -11972 22308 -11908
rect 22244 -12052 22308 -11988
rect 22244 -12132 22308 -12068
rect 22244 -12212 22308 -12148
rect 22244 -12292 22308 -12228
rect 22244 -12372 22308 -12308
rect 22244 -12452 22308 -12388
rect 22244 -12532 22308 -12468
rect 22244 -12612 22308 -12548
rect 22244 -12692 22308 -12628
rect 22244 -12772 22308 -12708
rect 22244 -12852 22308 -12788
rect 22244 -12932 22308 -12868
rect 22244 -13012 22308 -12948
rect 22244 -13092 22308 -13028
rect 22244 -13172 22308 -13108
rect 22244 -13252 22308 -13188
rect 22244 -13332 22308 -13268
rect 22244 -13412 22308 -13348
rect 22244 -13492 22308 -13428
rect 22244 -13572 22308 -13508
rect 22244 -13652 22308 -13588
rect 22244 -13732 22308 -13668
rect 22244 -13812 22308 -13748
rect 22244 -13892 22308 -13828
rect 22244 -13972 22308 -13908
rect 22244 -14052 22308 -13988
rect 22244 -14132 22308 -14068
rect 22244 -14212 22308 -14148
rect 22244 -14292 22308 -14228
rect 22244 -14372 22308 -14308
rect 22244 -14452 22308 -14388
rect 22244 -14532 22308 -14468
rect 22244 -14612 22308 -14548
rect 22244 -14692 22308 -14628
rect 22244 -14772 22308 -14708
rect 22244 -14852 22308 -14788
rect 22244 -14932 22308 -14868
rect 22244 -15012 22308 -14948
rect 22244 -15092 22308 -15028
rect 22244 -15172 22308 -15108
rect 22244 -15252 22308 -15188
rect 22244 -15332 22308 -15268
rect 22244 -15412 22308 -15348
rect 22244 -15492 22308 -15428
rect 22244 -15572 22308 -15508
rect 22244 -15652 22308 -15588
rect 22244 -15732 22308 -15668
rect 22244 -15812 22308 -15748
rect 27856 -10852 27920 -10788
rect 27856 -10932 27920 -10868
rect 27856 -11012 27920 -10948
rect 27856 -11092 27920 -11028
rect 27856 -11172 27920 -11108
rect 27856 -11252 27920 -11188
rect 27856 -11332 27920 -11268
rect 27856 -11412 27920 -11348
rect 27856 -11492 27920 -11428
rect 27856 -11572 27920 -11508
rect 27856 -11652 27920 -11588
rect 27856 -11732 27920 -11668
rect 27856 -11812 27920 -11748
rect 27856 -11892 27920 -11828
rect 27856 -11972 27920 -11908
rect 27856 -12052 27920 -11988
rect 27856 -12132 27920 -12068
rect 27856 -12212 27920 -12148
rect 27856 -12292 27920 -12228
rect 27856 -12372 27920 -12308
rect 27856 -12452 27920 -12388
rect 27856 -12532 27920 -12468
rect 27856 -12612 27920 -12548
rect 27856 -12692 27920 -12628
rect 27856 -12772 27920 -12708
rect 27856 -12852 27920 -12788
rect 27856 -12932 27920 -12868
rect 27856 -13012 27920 -12948
rect 27856 -13092 27920 -13028
rect 27856 -13172 27920 -13108
rect 27856 -13252 27920 -13188
rect 27856 -13332 27920 -13268
rect 27856 -13412 27920 -13348
rect 27856 -13492 27920 -13428
rect 27856 -13572 27920 -13508
rect 27856 -13652 27920 -13588
rect 27856 -13732 27920 -13668
rect 27856 -13812 27920 -13748
rect 27856 -13892 27920 -13828
rect 27856 -13972 27920 -13908
rect 27856 -14052 27920 -13988
rect 27856 -14132 27920 -14068
rect 27856 -14212 27920 -14148
rect 27856 -14292 27920 -14228
rect 27856 -14372 27920 -14308
rect 27856 -14452 27920 -14388
rect 27856 -14532 27920 -14468
rect 27856 -14612 27920 -14548
rect 27856 -14692 27920 -14628
rect 27856 -14772 27920 -14708
rect 27856 -14852 27920 -14788
rect 27856 -14932 27920 -14868
rect 27856 -15012 27920 -14948
rect 27856 -15092 27920 -15028
rect 27856 -15172 27920 -15108
rect 27856 -15252 27920 -15188
rect 27856 -15332 27920 -15268
rect 27856 -15412 27920 -15348
rect 27856 -15492 27920 -15428
rect 27856 -15572 27920 -15508
rect 27856 -15652 27920 -15588
rect 27856 -15732 27920 -15668
rect 27856 -15812 27920 -15748
rect 33468 -10852 33532 -10788
rect 33468 -10932 33532 -10868
rect 33468 -11012 33532 -10948
rect 33468 -11092 33532 -11028
rect 33468 -11172 33532 -11108
rect 33468 -11252 33532 -11188
rect 33468 -11332 33532 -11268
rect 33468 -11412 33532 -11348
rect 33468 -11492 33532 -11428
rect 33468 -11572 33532 -11508
rect 33468 -11652 33532 -11588
rect 33468 -11732 33532 -11668
rect 33468 -11812 33532 -11748
rect 33468 -11892 33532 -11828
rect 33468 -11972 33532 -11908
rect 33468 -12052 33532 -11988
rect 33468 -12132 33532 -12068
rect 33468 -12212 33532 -12148
rect 33468 -12292 33532 -12228
rect 33468 -12372 33532 -12308
rect 33468 -12452 33532 -12388
rect 33468 -12532 33532 -12468
rect 33468 -12612 33532 -12548
rect 33468 -12692 33532 -12628
rect 33468 -12772 33532 -12708
rect 33468 -12852 33532 -12788
rect 33468 -12932 33532 -12868
rect 33468 -13012 33532 -12948
rect 33468 -13092 33532 -13028
rect 33468 -13172 33532 -13108
rect 33468 -13252 33532 -13188
rect 33468 -13332 33532 -13268
rect 33468 -13412 33532 -13348
rect 33468 -13492 33532 -13428
rect 33468 -13572 33532 -13508
rect 33468 -13652 33532 -13588
rect 33468 -13732 33532 -13668
rect 33468 -13812 33532 -13748
rect 33468 -13892 33532 -13828
rect 33468 -13972 33532 -13908
rect 33468 -14052 33532 -13988
rect 33468 -14132 33532 -14068
rect 33468 -14212 33532 -14148
rect 33468 -14292 33532 -14228
rect 33468 -14372 33532 -14308
rect 33468 -14452 33532 -14388
rect 33468 -14532 33532 -14468
rect 33468 -14612 33532 -14548
rect 33468 -14692 33532 -14628
rect 33468 -14772 33532 -14708
rect 33468 -14852 33532 -14788
rect 33468 -14932 33532 -14868
rect 33468 -15012 33532 -14948
rect 33468 -15092 33532 -15028
rect 33468 -15172 33532 -15108
rect 33468 -15252 33532 -15188
rect 33468 -15332 33532 -15268
rect 33468 -15412 33532 -15348
rect 33468 -15492 33532 -15428
rect 33468 -15572 33532 -15508
rect 33468 -15652 33532 -15588
rect 33468 -15732 33532 -15668
rect 33468 -15812 33532 -15748
rect 39080 -10852 39144 -10788
rect 39080 -10932 39144 -10868
rect 39080 -11012 39144 -10948
rect 39080 -11092 39144 -11028
rect 39080 -11172 39144 -11108
rect 39080 -11252 39144 -11188
rect 39080 -11332 39144 -11268
rect 39080 -11412 39144 -11348
rect 39080 -11492 39144 -11428
rect 39080 -11572 39144 -11508
rect 39080 -11652 39144 -11588
rect 39080 -11732 39144 -11668
rect 39080 -11812 39144 -11748
rect 39080 -11892 39144 -11828
rect 39080 -11972 39144 -11908
rect 39080 -12052 39144 -11988
rect 39080 -12132 39144 -12068
rect 39080 -12212 39144 -12148
rect 39080 -12292 39144 -12228
rect 39080 -12372 39144 -12308
rect 39080 -12452 39144 -12388
rect 39080 -12532 39144 -12468
rect 39080 -12612 39144 -12548
rect 39080 -12692 39144 -12628
rect 39080 -12772 39144 -12708
rect 39080 -12852 39144 -12788
rect 39080 -12932 39144 -12868
rect 39080 -13012 39144 -12948
rect 39080 -13092 39144 -13028
rect 39080 -13172 39144 -13108
rect 39080 -13252 39144 -13188
rect 39080 -13332 39144 -13268
rect 39080 -13412 39144 -13348
rect 39080 -13492 39144 -13428
rect 39080 -13572 39144 -13508
rect 39080 -13652 39144 -13588
rect 39080 -13732 39144 -13668
rect 39080 -13812 39144 -13748
rect 39080 -13892 39144 -13828
rect 39080 -13972 39144 -13908
rect 39080 -14052 39144 -13988
rect 39080 -14132 39144 -14068
rect 39080 -14212 39144 -14148
rect 39080 -14292 39144 -14228
rect 39080 -14372 39144 -14308
rect 39080 -14452 39144 -14388
rect 39080 -14532 39144 -14468
rect 39080 -14612 39144 -14548
rect 39080 -14692 39144 -14628
rect 39080 -14772 39144 -14708
rect 39080 -14852 39144 -14788
rect 39080 -14932 39144 -14868
rect 39080 -15012 39144 -14948
rect 39080 -15092 39144 -15028
rect 39080 -15172 39144 -15108
rect 39080 -15252 39144 -15188
rect 39080 -15332 39144 -15268
rect 39080 -15412 39144 -15348
rect 39080 -15492 39144 -15428
rect 39080 -15572 39144 -15508
rect 39080 -15652 39144 -15588
rect 39080 -15732 39144 -15668
rect 39080 -15812 39144 -15748
rect -33876 -16172 -33812 -16108
rect -33876 -16252 -33812 -16188
rect -33876 -16332 -33812 -16268
rect -33876 -16412 -33812 -16348
rect -33876 -16492 -33812 -16428
rect -33876 -16572 -33812 -16508
rect -33876 -16652 -33812 -16588
rect -33876 -16732 -33812 -16668
rect -33876 -16812 -33812 -16748
rect -33876 -16892 -33812 -16828
rect -33876 -16972 -33812 -16908
rect -33876 -17052 -33812 -16988
rect -33876 -17132 -33812 -17068
rect -33876 -17212 -33812 -17148
rect -33876 -17292 -33812 -17228
rect -33876 -17372 -33812 -17308
rect -33876 -17452 -33812 -17388
rect -33876 -17532 -33812 -17468
rect -33876 -17612 -33812 -17548
rect -33876 -17692 -33812 -17628
rect -33876 -17772 -33812 -17708
rect -33876 -17852 -33812 -17788
rect -33876 -17932 -33812 -17868
rect -33876 -18012 -33812 -17948
rect -33876 -18092 -33812 -18028
rect -33876 -18172 -33812 -18108
rect -33876 -18252 -33812 -18188
rect -33876 -18332 -33812 -18268
rect -33876 -18412 -33812 -18348
rect -33876 -18492 -33812 -18428
rect -33876 -18572 -33812 -18508
rect -33876 -18652 -33812 -18588
rect -33876 -18732 -33812 -18668
rect -33876 -18812 -33812 -18748
rect -33876 -18892 -33812 -18828
rect -33876 -18972 -33812 -18908
rect -33876 -19052 -33812 -18988
rect -33876 -19132 -33812 -19068
rect -33876 -19212 -33812 -19148
rect -33876 -19292 -33812 -19228
rect -33876 -19372 -33812 -19308
rect -33876 -19452 -33812 -19388
rect -33876 -19532 -33812 -19468
rect -33876 -19612 -33812 -19548
rect -33876 -19692 -33812 -19628
rect -33876 -19772 -33812 -19708
rect -33876 -19852 -33812 -19788
rect -33876 -19932 -33812 -19868
rect -33876 -20012 -33812 -19948
rect -33876 -20092 -33812 -20028
rect -33876 -20172 -33812 -20108
rect -33876 -20252 -33812 -20188
rect -33876 -20332 -33812 -20268
rect -33876 -20412 -33812 -20348
rect -33876 -20492 -33812 -20428
rect -33876 -20572 -33812 -20508
rect -33876 -20652 -33812 -20588
rect -33876 -20732 -33812 -20668
rect -33876 -20812 -33812 -20748
rect -33876 -20892 -33812 -20828
rect -33876 -20972 -33812 -20908
rect -33876 -21052 -33812 -20988
rect -33876 -21132 -33812 -21068
rect -28264 -16172 -28200 -16108
rect -28264 -16252 -28200 -16188
rect -28264 -16332 -28200 -16268
rect -28264 -16412 -28200 -16348
rect -28264 -16492 -28200 -16428
rect -28264 -16572 -28200 -16508
rect -28264 -16652 -28200 -16588
rect -28264 -16732 -28200 -16668
rect -28264 -16812 -28200 -16748
rect -28264 -16892 -28200 -16828
rect -28264 -16972 -28200 -16908
rect -28264 -17052 -28200 -16988
rect -28264 -17132 -28200 -17068
rect -28264 -17212 -28200 -17148
rect -28264 -17292 -28200 -17228
rect -28264 -17372 -28200 -17308
rect -28264 -17452 -28200 -17388
rect -28264 -17532 -28200 -17468
rect -28264 -17612 -28200 -17548
rect -28264 -17692 -28200 -17628
rect -28264 -17772 -28200 -17708
rect -28264 -17852 -28200 -17788
rect -28264 -17932 -28200 -17868
rect -28264 -18012 -28200 -17948
rect -28264 -18092 -28200 -18028
rect -28264 -18172 -28200 -18108
rect -28264 -18252 -28200 -18188
rect -28264 -18332 -28200 -18268
rect -28264 -18412 -28200 -18348
rect -28264 -18492 -28200 -18428
rect -28264 -18572 -28200 -18508
rect -28264 -18652 -28200 -18588
rect -28264 -18732 -28200 -18668
rect -28264 -18812 -28200 -18748
rect -28264 -18892 -28200 -18828
rect -28264 -18972 -28200 -18908
rect -28264 -19052 -28200 -18988
rect -28264 -19132 -28200 -19068
rect -28264 -19212 -28200 -19148
rect -28264 -19292 -28200 -19228
rect -28264 -19372 -28200 -19308
rect -28264 -19452 -28200 -19388
rect -28264 -19532 -28200 -19468
rect -28264 -19612 -28200 -19548
rect -28264 -19692 -28200 -19628
rect -28264 -19772 -28200 -19708
rect -28264 -19852 -28200 -19788
rect -28264 -19932 -28200 -19868
rect -28264 -20012 -28200 -19948
rect -28264 -20092 -28200 -20028
rect -28264 -20172 -28200 -20108
rect -28264 -20252 -28200 -20188
rect -28264 -20332 -28200 -20268
rect -28264 -20412 -28200 -20348
rect -28264 -20492 -28200 -20428
rect -28264 -20572 -28200 -20508
rect -28264 -20652 -28200 -20588
rect -28264 -20732 -28200 -20668
rect -28264 -20812 -28200 -20748
rect -28264 -20892 -28200 -20828
rect -28264 -20972 -28200 -20908
rect -28264 -21052 -28200 -20988
rect -28264 -21132 -28200 -21068
rect -22652 -16172 -22588 -16108
rect -22652 -16252 -22588 -16188
rect -22652 -16332 -22588 -16268
rect -22652 -16412 -22588 -16348
rect -22652 -16492 -22588 -16428
rect -22652 -16572 -22588 -16508
rect -22652 -16652 -22588 -16588
rect -22652 -16732 -22588 -16668
rect -22652 -16812 -22588 -16748
rect -22652 -16892 -22588 -16828
rect -22652 -16972 -22588 -16908
rect -22652 -17052 -22588 -16988
rect -22652 -17132 -22588 -17068
rect -22652 -17212 -22588 -17148
rect -22652 -17292 -22588 -17228
rect -22652 -17372 -22588 -17308
rect -22652 -17452 -22588 -17388
rect -22652 -17532 -22588 -17468
rect -22652 -17612 -22588 -17548
rect -22652 -17692 -22588 -17628
rect -22652 -17772 -22588 -17708
rect -22652 -17852 -22588 -17788
rect -22652 -17932 -22588 -17868
rect -22652 -18012 -22588 -17948
rect -22652 -18092 -22588 -18028
rect -22652 -18172 -22588 -18108
rect -22652 -18252 -22588 -18188
rect -22652 -18332 -22588 -18268
rect -22652 -18412 -22588 -18348
rect -22652 -18492 -22588 -18428
rect -22652 -18572 -22588 -18508
rect -22652 -18652 -22588 -18588
rect -22652 -18732 -22588 -18668
rect -22652 -18812 -22588 -18748
rect -22652 -18892 -22588 -18828
rect -22652 -18972 -22588 -18908
rect -22652 -19052 -22588 -18988
rect -22652 -19132 -22588 -19068
rect -22652 -19212 -22588 -19148
rect -22652 -19292 -22588 -19228
rect -22652 -19372 -22588 -19308
rect -22652 -19452 -22588 -19388
rect -22652 -19532 -22588 -19468
rect -22652 -19612 -22588 -19548
rect -22652 -19692 -22588 -19628
rect -22652 -19772 -22588 -19708
rect -22652 -19852 -22588 -19788
rect -22652 -19932 -22588 -19868
rect -22652 -20012 -22588 -19948
rect -22652 -20092 -22588 -20028
rect -22652 -20172 -22588 -20108
rect -22652 -20252 -22588 -20188
rect -22652 -20332 -22588 -20268
rect -22652 -20412 -22588 -20348
rect -22652 -20492 -22588 -20428
rect -22652 -20572 -22588 -20508
rect -22652 -20652 -22588 -20588
rect -22652 -20732 -22588 -20668
rect -22652 -20812 -22588 -20748
rect -22652 -20892 -22588 -20828
rect -22652 -20972 -22588 -20908
rect -22652 -21052 -22588 -20988
rect -22652 -21132 -22588 -21068
rect -17040 -16172 -16976 -16108
rect -17040 -16252 -16976 -16188
rect -17040 -16332 -16976 -16268
rect -17040 -16412 -16976 -16348
rect -17040 -16492 -16976 -16428
rect -17040 -16572 -16976 -16508
rect -17040 -16652 -16976 -16588
rect -17040 -16732 -16976 -16668
rect -17040 -16812 -16976 -16748
rect -17040 -16892 -16976 -16828
rect -17040 -16972 -16976 -16908
rect -17040 -17052 -16976 -16988
rect -17040 -17132 -16976 -17068
rect -17040 -17212 -16976 -17148
rect -17040 -17292 -16976 -17228
rect -17040 -17372 -16976 -17308
rect -17040 -17452 -16976 -17388
rect -17040 -17532 -16976 -17468
rect -17040 -17612 -16976 -17548
rect -17040 -17692 -16976 -17628
rect -17040 -17772 -16976 -17708
rect -17040 -17852 -16976 -17788
rect -17040 -17932 -16976 -17868
rect -17040 -18012 -16976 -17948
rect -17040 -18092 -16976 -18028
rect -17040 -18172 -16976 -18108
rect -17040 -18252 -16976 -18188
rect -17040 -18332 -16976 -18268
rect -17040 -18412 -16976 -18348
rect -17040 -18492 -16976 -18428
rect -17040 -18572 -16976 -18508
rect -17040 -18652 -16976 -18588
rect -17040 -18732 -16976 -18668
rect -17040 -18812 -16976 -18748
rect -17040 -18892 -16976 -18828
rect -17040 -18972 -16976 -18908
rect -17040 -19052 -16976 -18988
rect -17040 -19132 -16976 -19068
rect -17040 -19212 -16976 -19148
rect -17040 -19292 -16976 -19228
rect -17040 -19372 -16976 -19308
rect -17040 -19452 -16976 -19388
rect -17040 -19532 -16976 -19468
rect -17040 -19612 -16976 -19548
rect -17040 -19692 -16976 -19628
rect -17040 -19772 -16976 -19708
rect -17040 -19852 -16976 -19788
rect -17040 -19932 -16976 -19868
rect -17040 -20012 -16976 -19948
rect -17040 -20092 -16976 -20028
rect -17040 -20172 -16976 -20108
rect -17040 -20252 -16976 -20188
rect -17040 -20332 -16976 -20268
rect -17040 -20412 -16976 -20348
rect -17040 -20492 -16976 -20428
rect -17040 -20572 -16976 -20508
rect -17040 -20652 -16976 -20588
rect -17040 -20732 -16976 -20668
rect -17040 -20812 -16976 -20748
rect -17040 -20892 -16976 -20828
rect -17040 -20972 -16976 -20908
rect -17040 -21052 -16976 -20988
rect -17040 -21132 -16976 -21068
rect -11428 -16172 -11364 -16108
rect -11428 -16252 -11364 -16188
rect -11428 -16332 -11364 -16268
rect -11428 -16412 -11364 -16348
rect -11428 -16492 -11364 -16428
rect -11428 -16572 -11364 -16508
rect -11428 -16652 -11364 -16588
rect -11428 -16732 -11364 -16668
rect -11428 -16812 -11364 -16748
rect -11428 -16892 -11364 -16828
rect -11428 -16972 -11364 -16908
rect -11428 -17052 -11364 -16988
rect -11428 -17132 -11364 -17068
rect -11428 -17212 -11364 -17148
rect -11428 -17292 -11364 -17228
rect -11428 -17372 -11364 -17308
rect -11428 -17452 -11364 -17388
rect -11428 -17532 -11364 -17468
rect -11428 -17612 -11364 -17548
rect -11428 -17692 -11364 -17628
rect -11428 -17772 -11364 -17708
rect -11428 -17852 -11364 -17788
rect -11428 -17932 -11364 -17868
rect -11428 -18012 -11364 -17948
rect -11428 -18092 -11364 -18028
rect -11428 -18172 -11364 -18108
rect -11428 -18252 -11364 -18188
rect -11428 -18332 -11364 -18268
rect -11428 -18412 -11364 -18348
rect -11428 -18492 -11364 -18428
rect -11428 -18572 -11364 -18508
rect -11428 -18652 -11364 -18588
rect -11428 -18732 -11364 -18668
rect -11428 -18812 -11364 -18748
rect -11428 -18892 -11364 -18828
rect -11428 -18972 -11364 -18908
rect -11428 -19052 -11364 -18988
rect -11428 -19132 -11364 -19068
rect -11428 -19212 -11364 -19148
rect -11428 -19292 -11364 -19228
rect -11428 -19372 -11364 -19308
rect -11428 -19452 -11364 -19388
rect -11428 -19532 -11364 -19468
rect -11428 -19612 -11364 -19548
rect -11428 -19692 -11364 -19628
rect -11428 -19772 -11364 -19708
rect -11428 -19852 -11364 -19788
rect -11428 -19932 -11364 -19868
rect -11428 -20012 -11364 -19948
rect -11428 -20092 -11364 -20028
rect -11428 -20172 -11364 -20108
rect -11428 -20252 -11364 -20188
rect -11428 -20332 -11364 -20268
rect -11428 -20412 -11364 -20348
rect -11428 -20492 -11364 -20428
rect -11428 -20572 -11364 -20508
rect -11428 -20652 -11364 -20588
rect -11428 -20732 -11364 -20668
rect -11428 -20812 -11364 -20748
rect -11428 -20892 -11364 -20828
rect -11428 -20972 -11364 -20908
rect -11428 -21052 -11364 -20988
rect -11428 -21132 -11364 -21068
rect -5816 -16172 -5752 -16108
rect -5816 -16252 -5752 -16188
rect -5816 -16332 -5752 -16268
rect -5816 -16412 -5752 -16348
rect -5816 -16492 -5752 -16428
rect -5816 -16572 -5752 -16508
rect -5816 -16652 -5752 -16588
rect -5816 -16732 -5752 -16668
rect -5816 -16812 -5752 -16748
rect -5816 -16892 -5752 -16828
rect -5816 -16972 -5752 -16908
rect -5816 -17052 -5752 -16988
rect -5816 -17132 -5752 -17068
rect -5816 -17212 -5752 -17148
rect -5816 -17292 -5752 -17228
rect -5816 -17372 -5752 -17308
rect -5816 -17452 -5752 -17388
rect -5816 -17532 -5752 -17468
rect -5816 -17612 -5752 -17548
rect -5816 -17692 -5752 -17628
rect -5816 -17772 -5752 -17708
rect -5816 -17852 -5752 -17788
rect -5816 -17932 -5752 -17868
rect -5816 -18012 -5752 -17948
rect -5816 -18092 -5752 -18028
rect -5816 -18172 -5752 -18108
rect -5816 -18252 -5752 -18188
rect -5816 -18332 -5752 -18268
rect -5816 -18412 -5752 -18348
rect -5816 -18492 -5752 -18428
rect -5816 -18572 -5752 -18508
rect -5816 -18652 -5752 -18588
rect -5816 -18732 -5752 -18668
rect -5816 -18812 -5752 -18748
rect -5816 -18892 -5752 -18828
rect -5816 -18972 -5752 -18908
rect -5816 -19052 -5752 -18988
rect -5816 -19132 -5752 -19068
rect -5816 -19212 -5752 -19148
rect -5816 -19292 -5752 -19228
rect -5816 -19372 -5752 -19308
rect -5816 -19452 -5752 -19388
rect -5816 -19532 -5752 -19468
rect -5816 -19612 -5752 -19548
rect -5816 -19692 -5752 -19628
rect -5816 -19772 -5752 -19708
rect -5816 -19852 -5752 -19788
rect -5816 -19932 -5752 -19868
rect -5816 -20012 -5752 -19948
rect -5816 -20092 -5752 -20028
rect -5816 -20172 -5752 -20108
rect -5816 -20252 -5752 -20188
rect -5816 -20332 -5752 -20268
rect -5816 -20412 -5752 -20348
rect -5816 -20492 -5752 -20428
rect -5816 -20572 -5752 -20508
rect -5816 -20652 -5752 -20588
rect -5816 -20732 -5752 -20668
rect -5816 -20812 -5752 -20748
rect -5816 -20892 -5752 -20828
rect -5816 -20972 -5752 -20908
rect -5816 -21052 -5752 -20988
rect -5816 -21132 -5752 -21068
rect -204 -16172 -140 -16108
rect -204 -16252 -140 -16188
rect -204 -16332 -140 -16268
rect -204 -16412 -140 -16348
rect -204 -16492 -140 -16428
rect -204 -16572 -140 -16508
rect -204 -16652 -140 -16588
rect -204 -16732 -140 -16668
rect -204 -16812 -140 -16748
rect -204 -16892 -140 -16828
rect -204 -16972 -140 -16908
rect -204 -17052 -140 -16988
rect -204 -17132 -140 -17068
rect -204 -17212 -140 -17148
rect -204 -17292 -140 -17228
rect -204 -17372 -140 -17308
rect -204 -17452 -140 -17388
rect -204 -17532 -140 -17468
rect -204 -17612 -140 -17548
rect -204 -17692 -140 -17628
rect -204 -17772 -140 -17708
rect -204 -17852 -140 -17788
rect -204 -17932 -140 -17868
rect -204 -18012 -140 -17948
rect -204 -18092 -140 -18028
rect -204 -18172 -140 -18108
rect -204 -18252 -140 -18188
rect -204 -18332 -140 -18268
rect -204 -18412 -140 -18348
rect -204 -18492 -140 -18428
rect -204 -18572 -140 -18508
rect -204 -18652 -140 -18588
rect -204 -18732 -140 -18668
rect -204 -18812 -140 -18748
rect -204 -18892 -140 -18828
rect -204 -18972 -140 -18908
rect -204 -19052 -140 -18988
rect -204 -19132 -140 -19068
rect -204 -19212 -140 -19148
rect -204 -19292 -140 -19228
rect -204 -19372 -140 -19308
rect -204 -19452 -140 -19388
rect -204 -19532 -140 -19468
rect -204 -19612 -140 -19548
rect -204 -19692 -140 -19628
rect -204 -19772 -140 -19708
rect -204 -19852 -140 -19788
rect -204 -19932 -140 -19868
rect -204 -20012 -140 -19948
rect -204 -20092 -140 -20028
rect -204 -20172 -140 -20108
rect -204 -20252 -140 -20188
rect -204 -20332 -140 -20268
rect -204 -20412 -140 -20348
rect -204 -20492 -140 -20428
rect -204 -20572 -140 -20508
rect -204 -20652 -140 -20588
rect -204 -20732 -140 -20668
rect -204 -20812 -140 -20748
rect -204 -20892 -140 -20828
rect -204 -20972 -140 -20908
rect -204 -21052 -140 -20988
rect -204 -21132 -140 -21068
rect 5408 -16172 5472 -16108
rect 5408 -16252 5472 -16188
rect 5408 -16332 5472 -16268
rect 5408 -16412 5472 -16348
rect 5408 -16492 5472 -16428
rect 5408 -16572 5472 -16508
rect 5408 -16652 5472 -16588
rect 5408 -16732 5472 -16668
rect 5408 -16812 5472 -16748
rect 5408 -16892 5472 -16828
rect 5408 -16972 5472 -16908
rect 5408 -17052 5472 -16988
rect 5408 -17132 5472 -17068
rect 5408 -17212 5472 -17148
rect 5408 -17292 5472 -17228
rect 5408 -17372 5472 -17308
rect 5408 -17452 5472 -17388
rect 5408 -17532 5472 -17468
rect 5408 -17612 5472 -17548
rect 5408 -17692 5472 -17628
rect 5408 -17772 5472 -17708
rect 5408 -17852 5472 -17788
rect 5408 -17932 5472 -17868
rect 5408 -18012 5472 -17948
rect 5408 -18092 5472 -18028
rect 5408 -18172 5472 -18108
rect 5408 -18252 5472 -18188
rect 5408 -18332 5472 -18268
rect 5408 -18412 5472 -18348
rect 5408 -18492 5472 -18428
rect 5408 -18572 5472 -18508
rect 5408 -18652 5472 -18588
rect 5408 -18732 5472 -18668
rect 5408 -18812 5472 -18748
rect 5408 -18892 5472 -18828
rect 5408 -18972 5472 -18908
rect 5408 -19052 5472 -18988
rect 5408 -19132 5472 -19068
rect 5408 -19212 5472 -19148
rect 5408 -19292 5472 -19228
rect 5408 -19372 5472 -19308
rect 5408 -19452 5472 -19388
rect 5408 -19532 5472 -19468
rect 5408 -19612 5472 -19548
rect 5408 -19692 5472 -19628
rect 5408 -19772 5472 -19708
rect 5408 -19852 5472 -19788
rect 5408 -19932 5472 -19868
rect 5408 -20012 5472 -19948
rect 5408 -20092 5472 -20028
rect 5408 -20172 5472 -20108
rect 5408 -20252 5472 -20188
rect 5408 -20332 5472 -20268
rect 5408 -20412 5472 -20348
rect 5408 -20492 5472 -20428
rect 5408 -20572 5472 -20508
rect 5408 -20652 5472 -20588
rect 5408 -20732 5472 -20668
rect 5408 -20812 5472 -20748
rect 5408 -20892 5472 -20828
rect 5408 -20972 5472 -20908
rect 5408 -21052 5472 -20988
rect 5408 -21132 5472 -21068
rect 11020 -16172 11084 -16108
rect 11020 -16252 11084 -16188
rect 11020 -16332 11084 -16268
rect 11020 -16412 11084 -16348
rect 11020 -16492 11084 -16428
rect 11020 -16572 11084 -16508
rect 11020 -16652 11084 -16588
rect 11020 -16732 11084 -16668
rect 11020 -16812 11084 -16748
rect 11020 -16892 11084 -16828
rect 11020 -16972 11084 -16908
rect 11020 -17052 11084 -16988
rect 11020 -17132 11084 -17068
rect 11020 -17212 11084 -17148
rect 11020 -17292 11084 -17228
rect 11020 -17372 11084 -17308
rect 11020 -17452 11084 -17388
rect 11020 -17532 11084 -17468
rect 11020 -17612 11084 -17548
rect 11020 -17692 11084 -17628
rect 11020 -17772 11084 -17708
rect 11020 -17852 11084 -17788
rect 11020 -17932 11084 -17868
rect 11020 -18012 11084 -17948
rect 11020 -18092 11084 -18028
rect 11020 -18172 11084 -18108
rect 11020 -18252 11084 -18188
rect 11020 -18332 11084 -18268
rect 11020 -18412 11084 -18348
rect 11020 -18492 11084 -18428
rect 11020 -18572 11084 -18508
rect 11020 -18652 11084 -18588
rect 11020 -18732 11084 -18668
rect 11020 -18812 11084 -18748
rect 11020 -18892 11084 -18828
rect 11020 -18972 11084 -18908
rect 11020 -19052 11084 -18988
rect 11020 -19132 11084 -19068
rect 11020 -19212 11084 -19148
rect 11020 -19292 11084 -19228
rect 11020 -19372 11084 -19308
rect 11020 -19452 11084 -19388
rect 11020 -19532 11084 -19468
rect 11020 -19612 11084 -19548
rect 11020 -19692 11084 -19628
rect 11020 -19772 11084 -19708
rect 11020 -19852 11084 -19788
rect 11020 -19932 11084 -19868
rect 11020 -20012 11084 -19948
rect 11020 -20092 11084 -20028
rect 11020 -20172 11084 -20108
rect 11020 -20252 11084 -20188
rect 11020 -20332 11084 -20268
rect 11020 -20412 11084 -20348
rect 11020 -20492 11084 -20428
rect 11020 -20572 11084 -20508
rect 11020 -20652 11084 -20588
rect 11020 -20732 11084 -20668
rect 11020 -20812 11084 -20748
rect 11020 -20892 11084 -20828
rect 11020 -20972 11084 -20908
rect 11020 -21052 11084 -20988
rect 11020 -21132 11084 -21068
rect 16632 -16172 16696 -16108
rect 16632 -16252 16696 -16188
rect 16632 -16332 16696 -16268
rect 16632 -16412 16696 -16348
rect 16632 -16492 16696 -16428
rect 16632 -16572 16696 -16508
rect 16632 -16652 16696 -16588
rect 16632 -16732 16696 -16668
rect 16632 -16812 16696 -16748
rect 16632 -16892 16696 -16828
rect 16632 -16972 16696 -16908
rect 16632 -17052 16696 -16988
rect 16632 -17132 16696 -17068
rect 16632 -17212 16696 -17148
rect 16632 -17292 16696 -17228
rect 16632 -17372 16696 -17308
rect 16632 -17452 16696 -17388
rect 16632 -17532 16696 -17468
rect 16632 -17612 16696 -17548
rect 16632 -17692 16696 -17628
rect 16632 -17772 16696 -17708
rect 16632 -17852 16696 -17788
rect 16632 -17932 16696 -17868
rect 16632 -18012 16696 -17948
rect 16632 -18092 16696 -18028
rect 16632 -18172 16696 -18108
rect 16632 -18252 16696 -18188
rect 16632 -18332 16696 -18268
rect 16632 -18412 16696 -18348
rect 16632 -18492 16696 -18428
rect 16632 -18572 16696 -18508
rect 16632 -18652 16696 -18588
rect 16632 -18732 16696 -18668
rect 16632 -18812 16696 -18748
rect 16632 -18892 16696 -18828
rect 16632 -18972 16696 -18908
rect 16632 -19052 16696 -18988
rect 16632 -19132 16696 -19068
rect 16632 -19212 16696 -19148
rect 16632 -19292 16696 -19228
rect 16632 -19372 16696 -19308
rect 16632 -19452 16696 -19388
rect 16632 -19532 16696 -19468
rect 16632 -19612 16696 -19548
rect 16632 -19692 16696 -19628
rect 16632 -19772 16696 -19708
rect 16632 -19852 16696 -19788
rect 16632 -19932 16696 -19868
rect 16632 -20012 16696 -19948
rect 16632 -20092 16696 -20028
rect 16632 -20172 16696 -20108
rect 16632 -20252 16696 -20188
rect 16632 -20332 16696 -20268
rect 16632 -20412 16696 -20348
rect 16632 -20492 16696 -20428
rect 16632 -20572 16696 -20508
rect 16632 -20652 16696 -20588
rect 16632 -20732 16696 -20668
rect 16632 -20812 16696 -20748
rect 16632 -20892 16696 -20828
rect 16632 -20972 16696 -20908
rect 16632 -21052 16696 -20988
rect 16632 -21132 16696 -21068
rect 22244 -16172 22308 -16108
rect 22244 -16252 22308 -16188
rect 22244 -16332 22308 -16268
rect 22244 -16412 22308 -16348
rect 22244 -16492 22308 -16428
rect 22244 -16572 22308 -16508
rect 22244 -16652 22308 -16588
rect 22244 -16732 22308 -16668
rect 22244 -16812 22308 -16748
rect 22244 -16892 22308 -16828
rect 22244 -16972 22308 -16908
rect 22244 -17052 22308 -16988
rect 22244 -17132 22308 -17068
rect 22244 -17212 22308 -17148
rect 22244 -17292 22308 -17228
rect 22244 -17372 22308 -17308
rect 22244 -17452 22308 -17388
rect 22244 -17532 22308 -17468
rect 22244 -17612 22308 -17548
rect 22244 -17692 22308 -17628
rect 22244 -17772 22308 -17708
rect 22244 -17852 22308 -17788
rect 22244 -17932 22308 -17868
rect 22244 -18012 22308 -17948
rect 22244 -18092 22308 -18028
rect 22244 -18172 22308 -18108
rect 22244 -18252 22308 -18188
rect 22244 -18332 22308 -18268
rect 22244 -18412 22308 -18348
rect 22244 -18492 22308 -18428
rect 22244 -18572 22308 -18508
rect 22244 -18652 22308 -18588
rect 22244 -18732 22308 -18668
rect 22244 -18812 22308 -18748
rect 22244 -18892 22308 -18828
rect 22244 -18972 22308 -18908
rect 22244 -19052 22308 -18988
rect 22244 -19132 22308 -19068
rect 22244 -19212 22308 -19148
rect 22244 -19292 22308 -19228
rect 22244 -19372 22308 -19308
rect 22244 -19452 22308 -19388
rect 22244 -19532 22308 -19468
rect 22244 -19612 22308 -19548
rect 22244 -19692 22308 -19628
rect 22244 -19772 22308 -19708
rect 22244 -19852 22308 -19788
rect 22244 -19932 22308 -19868
rect 22244 -20012 22308 -19948
rect 22244 -20092 22308 -20028
rect 22244 -20172 22308 -20108
rect 22244 -20252 22308 -20188
rect 22244 -20332 22308 -20268
rect 22244 -20412 22308 -20348
rect 22244 -20492 22308 -20428
rect 22244 -20572 22308 -20508
rect 22244 -20652 22308 -20588
rect 22244 -20732 22308 -20668
rect 22244 -20812 22308 -20748
rect 22244 -20892 22308 -20828
rect 22244 -20972 22308 -20908
rect 22244 -21052 22308 -20988
rect 22244 -21132 22308 -21068
rect 27856 -16172 27920 -16108
rect 27856 -16252 27920 -16188
rect 27856 -16332 27920 -16268
rect 27856 -16412 27920 -16348
rect 27856 -16492 27920 -16428
rect 27856 -16572 27920 -16508
rect 27856 -16652 27920 -16588
rect 27856 -16732 27920 -16668
rect 27856 -16812 27920 -16748
rect 27856 -16892 27920 -16828
rect 27856 -16972 27920 -16908
rect 27856 -17052 27920 -16988
rect 27856 -17132 27920 -17068
rect 27856 -17212 27920 -17148
rect 27856 -17292 27920 -17228
rect 27856 -17372 27920 -17308
rect 27856 -17452 27920 -17388
rect 27856 -17532 27920 -17468
rect 27856 -17612 27920 -17548
rect 27856 -17692 27920 -17628
rect 27856 -17772 27920 -17708
rect 27856 -17852 27920 -17788
rect 27856 -17932 27920 -17868
rect 27856 -18012 27920 -17948
rect 27856 -18092 27920 -18028
rect 27856 -18172 27920 -18108
rect 27856 -18252 27920 -18188
rect 27856 -18332 27920 -18268
rect 27856 -18412 27920 -18348
rect 27856 -18492 27920 -18428
rect 27856 -18572 27920 -18508
rect 27856 -18652 27920 -18588
rect 27856 -18732 27920 -18668
rect 27856 -18812 27920 -18748
rect 27856 -18892 27920 -18828
rect 27856 -18972 27920 -18908
rect 27856 -19052 27920 -18988
rect 27856 -19132 27920 -19068
rect 27856 -19212 27920 -19148
rect 27856 -19292 27920 -19228
rect 27856 -19372 27920 -19308
rect 27856 -19452 27920 -19388
rect 27856 -19532 27920 -19468
rect 27856 -19612 27920 -19548
rect 27856 -19692 27920 -19628
rect 27856 -19772 27920 -19708
rect 27856 -19852 27920 -19788
rect 27856 -19932 27920 -19868
rect 27856 -20012 27920 -19948
rect 27856 -20092 27920 -20028
rect 27856 -20172 27920 -20108
rect 27856 -20252 27920 -20188
rect 27856 -20332 27920 -20268
rect 27856 -20412 27920 -20348
rect 27856 -20492 27920 -20428
rect 27856 -20572 27920 -20508
rect 27856 -20652 27920 -20588
rect 27856 -20732 27920 -20668
rect 27856 -20812 27920 -20748
rect 27856 -20892 27920 -20828
rect 27856 -20972 27920 -20908
rect 27856 -21052 27920 -20988
rect 27856 -21132 27920 -21068
rect 33468 -16172 33532 -16108
rect 33468 -16252 33532 -16188
rect 33468 -16332 33532 -16268
rect 33468 -16412 33532 -16348
rect 33468 -16492 33532 -16428
rect 33468 -16572 33532 -16508
rect 33468 -16652 33532 -16588
rect 33468 -16732 33532 -16668
rect 33468 -16812 33532 -16748
rect 33468 -16892 33532 -16828
rect 33468 -16972 33532 -16908
rect 33468 -17052 33532 -16988
rect 33468 -17132 33532 -17068
rect 33468 -17212 33532 -17148
rect 33468 -17292 33532 -17228
rect 33468 -17372 33532 -17308
rect 33468 -17452 33532 -17388
rect 33468 -17532 33532 -17468
rect 33468 -17612 33532 -17548
rect 33468 -17692 33532 -17628
rect 33468 -17772 33532 -17708
rect 33468 -17852 33532 -17788
rect 33468 -17932 33532 -17868
rect 33468 -18012 33532 -17948
rect 33468 -18092 33532 -18028
rect 33468 -18172 33532 -18108
rect 33468 -18252 33532 -18188
rect 33468 -18332 33532 -18268
rect 33468 -18412 33532 -18348
rect 33468 -18492 33532 -18428
rect 33468 -18572 33532 -18508
rect 33468 -18652 33532 -18588
rect 33468 -18732 33532 -18668
rect 33468 -18812 33532 -18748
rect 33468 -18892 33532 -18828
rect 33468 -18972 33532 -18908
rect 33468 -19052 33532 -18988
rect 33468 -19132 33532 -19068
rect 33468 -19212 33532 -19148
rect 33468 -19292 33532 -19228
rect 33468 -19372 33532 -19308
rect 33468 -19452 33532 -19388
rect 33468 -19532 33532 -19468
rect 33468 -19612 33532 -19548
rect 33468 -19692 33532 -19628
rect 33468 -19772 33532 -19708
rect 33468 -19852 33532 -19788
rect 33468 -19932 33532 -19868
rect 33468 -20012 33532 -19948
rect 33468 -20092 33532 -20028
rect 33468 -20172 33532 -20108
rect 33468 -20252 33532 -20188
rect 33468 -20332 33532 -20268
rect 33468 -20412 33532 -20348
rect 33468 -20492 33532 -20428
rect 33468 -20572 33532 -20508
rect 33468 -20652 33532 -20588
rect 33468 -20732 33532 -20668
rect 33468 -20812 33532 -20748
rect 33468 -20892 33532 -20828
rect 33468 -20972 33532 -20908
rect 33468 -21052 33532 -20988
rect 33468 -21132 33532 -21068
rect 39080 -16172 39144 -16108
rect 39080 -16252 39144 -16188
rect 39080 -16332 39144 -16268
rect 39080 -16412 39144 -16348
rect 39080 -16492 39144 -16428
rect 39080 -16572 39144 -16508
rect 39080 -16652 39144 -16588
rect 39080 -16732 39144 -16668
rect 39080 -16812 39144 -16748
rect 39080 -16892 39144 -16828
rect 39080 -16972 39144 -16908
rect 39080 -17052 39144 -16988
rect 39080 -17132 39144 -17068
rect 39080 -17212 39144 -17148
rect 39080 -17292 39144 -17228
rect 39080 -17372 39144 -17308
rect 39080 -17452 39144 -17388
rect 39080 -17532 39144 -17468
rect 39080 -17612 39144 -17548
rect 39080 -17692 39144 -17628
rect 39080 -17772 39144 -17708
rect 39080 -17852 39144 -17788
rect 39080 -17932 39144 -17868
rect 39080 -18012 39144 -17948
rect 39080 -18092 39144 -18028
rect 39080 -18172 39144 -18108
rect 39080 -18252 39144 -18188
rect 39080 -18332 39144 -18268
rect 39080 -18412 39144 -18348
rect 39080 -18492 39144 -18428
rect 39080 -18572 39144 -18508
rect 39080 -18652 39144 -18588
rect 39080 -18732 39144 -18668
rect 39080 -18812 39144 -18748
rect 39080 -18892 39144 -18828
rect 39080 -18972 39144 -18908
rect 39080 -19052 39144 -18988
rect 39080 -19132 39144 -19068
rect 39080 -19212 39144 -19148
rect 39080 -19292 39144 -19228
rect 39080 -19372 39144 -19308
rect 39080 -19452 39144 -19388
rect 39080 -19532 39144 -19468
rect 39080 -19612 39144 -19548
rect 39080 -19692 39144 -19628
rect 39080 -19772 39144 -19708
rect 39080 -19852 39144 -19788
rect 39080 -19932 39144 -19868
rect 39080 -20012 39144 -19948
rect 39080 -20092 39144 -20028
rect 39080 -20172 39144 -20108
rect 39080 -20252 39144 -20188
rect 39080 -20332 39144 -20268
rect 39080 -20412 39144 -20348
rect 39080 -20492 39144 -20428
rect 39080 -20572 39144 -20508
rect 39080 -20652 39144 -20588
rect 39080 -20732 39144 -20668
rect 39080 -20812 39144 -20748
rect 39080 -20892 39144 -20828
rect 39080 -20972 39144 -20908
rect 39080 -21052 39144 -20988
rect 39080 -21132 39144 -21068
rect -33876 -21492 -33812 -21428
rect -33876 -21572 -33812 -21508
rect -33876 -21652 -33812 -21588
rect -33876 -21732 -33812 -21668
rect -33876 -21812 -33812 -21748
rect -33876 -21892 -33812 -21828
rect -33876 -21972 -33812 -21908
rect -33876 -22052 -33812 -21988
rect -33876 -22132 -33812 -22068
rect -33876 -22212 -33812 -22148
rect -33876 -22292 -33812 -22228
rect -33876 -22372 -33812 -22308
rect -33876 -22452 -33812 -22388
rect -33876 -22532 -33812 -22468
rect -33876 -22612 -33812 -22548
rect -33876 -22692 -33812 -22628
rect -33876 -22772 -33812 -22708
rect -33876 -22852 -33812 -22788
rect -33876 -22932 -33812 -22868
rect -33876 -23012 -33812 -22948
rect -33876 -23092 -33812 -23028
rect -33876 -23172 -33812 -23108
rect -33876 -23252 -33812 -23188
rect -33876 -23332 -33812 -23268
rect -33876 -23412 -33812 -23348
rect -33876 -23492 -33812 -23428
rect -33876 -23572 -33812 -23508
rect -33876 -23652 -33812 -23588
rect -33876 -23732 -33812 -23668
rect -33876 -23812 -33812 -23748
rect -33876 -23892 -33812 -23828
rect -33876 -23972 -33812 -23908
rect -33876 -24052 -33812 -23988
rect -33876 -24132 -33812 -24068
rect -33876 -24212 -33812 -24148
rect -33876 -24292 -33812 -24228
rect -33876 -24372 -33812 -24308
rect -33876 -24452 -33812 -24388
rect -33876 -24532 -33812 -24468
rect -33876 -24612 -33812 -24548
rect -33876 -24692 -33812 -24628
rect -33876 -24772 -33812 -24708
rect -33876 -24852 -33812 -24788
rect -33876 -24932 -33812 -24868
rect -33876 -25012 -33812 -24948
rect -33876 -25092 -33812 -25028
rect -33876 -25172 -33812 -25108
rect -33876 -25252 -33812 -25188
rect -33876 -25332 -33812 -25268
rect -33876 -25412 -33812 -25348
rect -33876 -25492 -33812 -25428
rect -33876 -25572 -33812 -25508
rect -33876 -25652 -33812 -25588
rect -33876 -25732 -33812 -25668
rect -33876 -25812 -33812 -25748
rect -33876 -25892 -33812 -25828
rect -33876 -25972 -33812 -25908
rect -33876 -26052 -33812 -25988
rect -33876 -26132 -33812 -26068
rect -33876 -26212 -33812 -26148
rect -33876 -26292 -33812 -26228
rect -33876 -26372 -33812 -26308
rect -33876 -26452 -33812 -26388
rect -28264 -21492 -28200 -21428
rect -28264 -21572 -28200 -21508
rect -28264 -21652 -28200 -21588
rect -28264 -21732 -28200 -21668
rect -28264 -21812 -28200 -21748
rect -28264 -21892 -28200 -21828
rect -28264 -21972 -28200 -21908
rect -28264 -22052 -28200 -21988
rect -28264 -22132 -28200 -22068
rect -28264 -22212 -28200 -22148
rect -28264 -22292 -28200 -22228
rect -28264 -22372 -28200 -22308
rect -28264 -22452 -28200 -22388
rect -28264 -22532 -28200 -22468
rect -28264 -22612 -28200 -22548
rect -28264 -22692 -28200 -22628
rect -28264 -22772 -28200 -22708
rect -28264 -22852 -28200 -22788
rect -28264 -22932 -28200 -22868
rect -28264 -23012 -28200 -22948
rect -28264 -23092 -28200 -23028
rect -28264 -23172 -28200 -23108
rect -28264 -23252 -28200 -23188
rect -28264 -23332 -28200 -23268
rect -28264 -23412 -28200 -23348
rect -28264 -23492 -28200 -23428
rect -28264 -23572 -28200 -23508
rect -28264 -23652 -28200 -23588
rect -28264 -23732 -28200 -23668
rect -28264 -23812 -28200 -23748
rect -28264 -23892 -28200 -23828
rect -28264 -23972 -28200 -23908
rect -28264 -24052 -28200 -23988
rect -28264 -24132 -28200 -24068
rect -28264 -24212 -28200 -24148
rect -28264 -24292 -28200 -24228
rect -28264 -24372 -28200 -24308
rect -28264 -24452 -28200 -24388
rect -28264 -24532 -28200 -24468
rect -28264 -24612 -28200 -24548
rect -28264 -24692 -28200 -24628
rect -28264 -24772 -28200 -24708
rect -28264 -24852 -28200 -24788
rect -28264 -24932 -28200 -24868
rect -28264 -25012 -28200 -24948
rect -28264 -25092 -28200 -25028
rect -28264 -25172 -28200 -25108
rect -28264 -25252 -28200 -25188
rect -28264 -25332 -28200 -25268
rect -28264 -25412 -28200 -25348
rect -28264 -25492 -28200 -25428
rect -28264 -25572 -28200 -25508
rect -28264 -25652 -28200 -25588
rect -28264 -25732 -28200 -25668
rect -28264 -25812 -28200 -25748
rect -28264 -25892 -28200 -25828
rect -28264 -25972 -28200 -25908
rect -28264 -26052 -28200 -25988
rect -28264 -26132 -28200 -26068
rect -28264 -26212 -28200 -26148
rect -28264 -26292 -28200 -26228
rect -28264 -26372 -28200 -26308
rect -28264 -26452 -28200 -26388
rect -22652 -21492 -22588 -21428
rect -22652 -21572 -22588 -21508
rect -22652 -21652 -22588 -21588
rect -22652 -21732 -22588 -21668
rect -22652 -21812 -22588 -21748
rect -22652 -21892 -22588 -21828
rect -22652 -21972 -22588 -21908
rect -22652 -22052 -22588 -21988
rect -22652 -22132 -22588 -22068
rect -22652 -22212 -22588 -22148
rect -22652 -22292 -22588 -22228
rect -22652 -22372 -22588 -22308
rect -22652 -22452 -22588 -22388
rect -22652 -22532 -22588 -22468
rect -22652 -22612 -22588 -22548
rect -22652 -22692 -22588 -22628
rect -22652 -22772 -22588 -22708
rect -22652 -22852 -22588 -22788
rect -22652 -22932 -22588 -22868
rect -22652 -23012 -22588 -22948
rect -22652 -23092 -22588 -23028
rect -22652 -23172 -22588 -23108
rect -22652 -23252 -22588 -23188
rect -22652 -23332 -22588 -23268
rect -22652 -23412 -22588 -23348
rect -22652 -23492 -22588 -23428
rect -22652 -23572 -22588 -23508
rect -22652 -23652 -22588 -23588
rect -22652 -23732 -22588 -23668
rect -22652 -23812 -22588 -23748
rect -22652 -23892 -22588 -23828
rect -22652 -23972 -22588 -23908
rect -22652 -24052 -22588 -23988
rect -22652 -24132 -22588 -24068
rect -22652 -24212 -22588 -24148
rect -22652 -24292 -22588 -24228
rect -22652 -24372 -22588 -24308
rect -22652 -24452 -22588 -24388
rect -22652 -24532 -22588 -24468
rect -22652 -24612 -22588 -24548
rect -22652 -24692 -22588 -24628
rect -22652 -24772 -22588 -24708
rect -22652 -24852 -22588 -24788
rect -22652 -24932 -22588 -24868
rect -22652 -25012 -22588 -24948
rect -22652 -25092 -22588 -25028
rect -22652 -25172 -22588 -25108
rect -22652 -25252 -22588 -25188
rect -22652 -25332 -22588 -25268
rect -22652 -25412 -22588 -25348
rect -22652 -25492 -22588 -25428
rect -22652 -25572 -22588 -25508
rect -22652 -25652 -22588 -25588
rect -22652 -25732 -22588 -25668
rect -22652 -25812 -22588 -25748
rect -22652 -25892 -22588 -25828
rect -22652 -25972 -22588 -25908
rect -22652 -26052 -22588 -25988
rect -22652 -26132 -22588 -26068
rect -22652 -26212 -22588 -26148
rect -22652 -26292 -22588 -26228
rect -22652 -26372 -22588 -26308
rect -22652 -26452 -22588 -26388
rect -17040 -21492 -16976 -21428
rect -17040 -21572 -16976 -21508
rect -17040 -21652 -16976 -21588
rect -17040 -21732 -16976 -21668
rect -17040 -21812 -16976 -21748
rect -17040 -21892 -16976 -21828
rect -17040 -21972 -16976 -21908
rect -17040 -22052 -16976 -21988
rect -17040 -22132 -16976 -22068
rect -17040 -22212 -16976 -22148
rect -17040 -22292 -16976 -22228
rect -17040 -22372 -16976 -22308
rect -17040 -22452 -16976 -22388
rect -17040 -22532 -16976 -22468
rect -17040 -22612 -16976 -22548
rect -17040 -22692 -16976 -22628
rect -17040 -22772 -16976 -22708
rect -17040 -22852 -16976 -22788
rect -17040 -22932 -16976 -22868
rect -17040 -23012 -16976 -22948
rect -17040 -23092 -16976 -23028
rect -17040 -23172 -16976 -23108
rect -17040 -23252 -16976 -23188
rect -17040 -23332 -16976 -23268
rect -17040 -23412 -16976 -23348
rect -17040 -23492 -16976 -23428
rect -17040 -23572 -16976 -23508
rect -17040 -23652 -16976 -23588
rect -17040 -23732 -16976 -23668
rect -17040 -23812 -16976 -23748
rect -17040 -23892 -16976 -23828
rect -17040 -23972 -16976 -23908
rect -17040 -24052 -16976 -23988
rect -17040 -24132 -16976 -24068
rect -17040 -24212 -16976 -24148
rect -17040 -24292 -16976 -24228
rect -17040 -24372 -16976 -24308
rect -17040 -24452 -16976 -24388
rect -17040 -24532 -16976 -24468
rect -17040 -24612 -16976 -24548
rect -17040 -24692 -16976 -24628
rect -17040 -24772 -16976 -24708
rect -17040 -24852 -16976 -24788
rect -17040 -24932 -16976 -24868
rect -17040 -25012 -16976 -24948
rect -17040 -25092 -16976 -25028
rect -17040 -25172 -16976 -25108
rect -17040 -25252 -16976 -25188
rect -17040 -25332 -16976 -25268
rect -17040 -25412 -16976 -25348
rect -17040 -25492 -16976 -25428
rect -17040 -25572 -16976 -25508
rect -17040 -25652 -16976 -25588
rect -17040 -25732 -16976 -25668
rect -17040 -25812 -16976 -25748
rect -17040 -25892 -16976 -25828
rect -17040 -25972 -16976 -25908
rect -17040 -26052 -16976 -25988
rect -17040 -26132 -16976 -26068
rect -17040 -26212 -16976 -26148
rect -17040 -26292 -16976 -26228
rect -17040 -26372 -16976 -26308
rect -17040 -26452 -16976 -26388
rect -11428 -21492 -11364 -21428
rect -11428 -21572 -11364 -21508
rect -11428 -21652 -11364 -21588
rect -11428 -21732 -11364 -21668
rect -11428 -21812 -11364 -21748
rect -11428 -21892 -11364 -21828
rect -11428 -21972 -11364 -21908
rect -11428 -22052 -11364 -21988
rect -11428 -22132 -11364 -22068
rect -11428 -22212 -11364 -22148
rect -11428 -22292 -11364 -22228
rect -11428 -22372 -11364 -22308
rect -11428 -22452 -11364 -22388
rect -11428 -22532 -11364 -22468
rect -11428 -22612 -11364 -22548
rect -11428 -22692 -11364 -22628
rect -11428 -22772 -11364 -22708
rect -11428 -22852 -11364 -22788
rect -11428 -22932 -11364 -22868
rect -11428 -23012 -11364 -22948
rect -11428 -23092 -11364 -23028
rect -11428 -23172 -11364 -23108
rect -11428 -23252 -11364 -23188
rect -11428 -23332 -11364 -23268
rect -11428 -23412 -11364 -23348
rect -11428 -23492 -11364 -23428
rect -11428 -23572 -11364 -23508
rect -11428 -23652 -11364 -23588
rect -11428 -23732 -11364 -23668
rect -11428 -23812 -11364 -23748
rect -11428 -23892 -11364 -23828
rect -11428 -23972 -11364 -23908
rect -11428 -24052 -11364 -23988
rect -11428 -24132 -11364 -24068
rect -11428 -24212 -11364 -24148
rect -11428 -24292 -11364 -24228
rect -11428 -24372 -11364 -24308
rect -11428 -24452 -11364 -24388
rect -11428 -24532 -11364 -24468
rect -11428 -24612 -11364 -24548
rect -11428 -24692 -11364 -24628
rect -11428 -24772 -11364 -24708
rect -11428 -24852 -11364 -24788
rect -11428 -24932 -11364 -24868
rect -11428 -25012 -11364 -24948
rect -11428 -25092 -11364 -25028
rect -11428 -25172 -11364 -25108
rect -11428 -25252 -11364 -25188
rect -11428 -25332 -11364 -25268
rect -11428 -25412 -11364 -25348
rect -11428 -25492 -11364 -25428
rect -11428 -25572 -11364 -25508
rect -11428 -25652 -11364 -25588
rect -11428 -25732 -11364 -25668
rect -11428 -25812 -11364 -25748
rect -11428 -25892 -11364 -25828
rect -11428 -25972 -11364 -25908
rect -11428 -26052 -11364 -25988
rect -11428 -26132 -11364 -26068
rect -11428 -26212 -11364 -26148
rect -11428 -26292 -11364 -26228
rect -11428 -26372 -11364 -26308
rect -11428 -26452 -11364 -26388
rect -5816 -21492 -5752 -21428
rect -5816 -21572 -5752 -21508
rect -5816 -21652 -5752 -21588
rect -5816 -21732 -5752 -21668
rect -5816 -21812 -5752 -21748
rect -5816 -21892 -5752 -21828
rect -5816 -21972 -5752 -21908
rect -5816 -22052 -5752 -21988
rect -5816 -22132 -5752 -22068
rect -5816 -22212 -5752 -22148
rect -5816 -22292 -5752 -22228
rect -5816 -22372 -5752 -22308
rect -5816 -22452 -5752 -22388
rect -5816 -22532 -5752 -22468
rect -5816 -22612 -5752 -22548
rect -5816 -22692 -5752 -22628
rect -5816 -22772 -5752 -22708
rect -5816 -22852 -5752 -22788
rect -5816 -22932 -5752 -22868
rect -5816 -23012 -5752 -22948
rect -5816 -23092 -5752 -23028
rect -5816 -23172 -5752 -23108
rect -5816 -23252 -5752 -23188
rect -5816 -23332 -5752 -23268
rect -5816 -23412 -5752 -23348
rect -5816 -23492 -5752 -23428
rect -5816 -23572 -5752 -23508
rect -5816 -23652 -5752 -23588
rect -5816 -23732 -5752 -23668
rect -5816 -23812 -5752 -23748
rect -5816 -23892 -5752 -23828
rect -5816 -23972 -5752 -23908
rect -5816 -24052 -5752 -23988
rect -5816 -24132 -5752 -24068
rect -5816 -24212 -5752 -24148
rect -5816 -24292 -5752 -24228
rect -5816 -24372 -5752 -24308
rect -5816 -24452 -5752 -24388
rect -5816 -24532 -5752 -24468
rect -5816 -24612 -5752 -24548
rect -5816 -24692 -5752 -24628
rect -5816 -24772 -5752 -24708
rect -5816 -24852 -5752 -24788
rect -5816 -24932 -5752 -24868
rect -5816 -25012 -5752 -24948
rect -5816 -25092 -5752 -25028
rect -5816 -25172 -5752 -25108
rect -5816 -25252 -5752 -25188
rect -5816 -25332 -5752 -25268
rect -5816 -25412 -5752 -25348
rect -5816 -25492 -5752 -25428
rect -5816 -25572 -5752 -25508
rect -5816 -25652 -5752 -25588
rect -5816 -25732 -5752 -25668
rect -5816 -25812 -5752 -25748
rect -5816 -25892 -5752 -25828
rect -5816 -25972 -5752 -25908
rect -5816 -26052 -5752 -25988
rect -5816 -26132 -5752 -26068
rect -5816 -26212 -5752 -26148
rect -5816 -26292 -5752 -26228
rect -5816 -26372 -5752 -26308
rect -5816 -26452 -5752 -26388
rect -204 -21492 -140 -21428
rect -204 -21572 -140 -21508
rect -204 -21652 -140 -21588
rect -204 -21732 -140 -21668
rect -204 -21812 -140 -21748
rect -204 -21892 -140 -21828
rect -204 -21972 -140 -21908
rect -204 -22052 -140 -21988
rect -204 -22132 -140 -22068
rect -204 -22212 -140 -22148
rect -204 -22292 -140 -22228
rect -204 -22372 -140 -22308
rect -204 -22452 -140 -22388
rect -204 -22532 -140 -22468
rect -204 -22612 -140 -22548
rect -204 -22692 -140 -22628
rect -204 -22772 -140 -22708
rect -204 -22852 -140 -22788
rect -204 -22932 -140 -22868
rect -204 -23012 -140 -22948
rect -204 -23092 -140 -23028
rect -204 -23172 -140 -23108
rect -204 -23252 -140 -23188
rect -204 -23332 -140 -23268
rect -204 -23412 -140 -23348
rect -204 -23492 -140 -23428
rect -204 -23572 -140 -23508
rect -204 -23652 -140 -23588
rect -204 -23732 -140 -23668
rect -204 -23812 -140 -23748
rect -204 -23892 -140 -23828
rect -204 -23972 -140 -23908
rect -204 -24052 -140 -23988
rect -204 -24132 -140 -24068
rect -204 -24212 -140 -24148
rect -204 -24292 -140 -24228
rect -204 -24372 -140 -24308
rect -204 -24452 -140 -24388
rect -204 -24532 -140 -24468
rect -204 -24612 -140 -24548
rect -204 -24692 -140 -24628
rect -204 -24772 -140 -24708
rect -204 -24852 -140 -24788
rect -204 -24932 -140 -24868
rect -204 -25012 -140 -24948
rect -204 -25092 -140 -25028
rect -204 -25172 -140 -25108
rect -204 -25252 -140 -25188
rect -204 -25332 -140 -25268
rect -204 -25412 -140 -25348
rect -204 -25492 -140 -25428
rect -204 -25572 -140 -25508
rect -204 -25652 -140 -25588
rect -204 -25732 -140 -25668
rect -204 -25812 -140 -25748
rect -204 -25892 -140 -25828
rect -204 -25972 -140 -25908
rect -204 -26052 -140 -25988
rect -204 -26132 -140 -26068
rect -204 -26212 -140 -26148
rect -204 -26292 -140 -26228
rect -204 -26372 -140 -26308
rect -204 -26452 -140 -26388
rect 5408 -21492 5472 -21428
rect 5408 -21572 5472 -21508
rect 5408 -21652 5472 -21588
rect 5408 -21732 5472 -21668
rect 5408 -21812 5472 -21748
rect 5408 -21892 5472 -21828
rect 5408 -21972 5472 -21908
rect 5408 -22052 5472 -21988
rect 5408 -22132 5472 -22068
rect 5408 -22212 5472 -22148
rect 5408 -22292 5472 -22228
rect 5408 -22372 5472 -22308
rect 5408 -22452 5472 -22388
rect 5408 -22532 5472 -22468
rect 5408 -22612 5472 -22548
rect 5408 -22692 5472 -22628
rect 5408 -22772 5472 -22708
rect 5408 -22852 5472 -22788
rect 5408 -22932 5472 -22868
rect 5408 -23012 5472 -22948
rect 5408 -23092 5472 -23028
rect 5408 -23172 5472 -23108
rect 5408 -23252 5472 -23188
rect 5408 -23332 5472 -23268
rect 5408 -23412 5472 -23348
rect 5408 -23492 5472 -23428
rect 5408 -23572 5472 -23508
rect 5408 -23652 5472 -23588
rect 5408 -23732 5472 -23668
rect 5408 -23812 5472 -23748
rect 5408 -23892 5472 -23828
rect 5408 -23972 5472 -23908
rect 5408 -24052 5472 -23988
rect 5408 -24132 5472 -24068
rect 5408 -24212 5472 -24148
rect 5408 -24292 5472 -24228
rect 5408 -24372 5472 -24308
rect 5408 -24452 5472 -24388
rect 5408 -24532 5472 -24468
rect 5408 -24612 5472 -24548
rect 5408 -24692 5472 -24628
rect 5408 -24772 5472 -24708
rect 5408 -24852 5472 -24788
rect 5408 -24932 5472 -24868
rect 5408 -25012 5472 -24948
rect 5408 -25092 5472 -25028
rect 5408 -25172 5472 -25108
rect 5408 -25252 5472 -25188
rect 5408 -25332 5472 -25268
rect 5408 -25412 5472 -25348
rect 5408 -25492 5472 -25428
rect 5408 -25572 5472 -25508
rect 5408 -25652 5472 -25588
rect 5408 -25732 5472 -25668
rect 5408 -25812 5472 -25748
rect 5408 -25892 5472 -25828
rect 5408 -25972 5472 -25908
rect 5408 -26052 5472 -25988
rect 5408 -26132 5472 -26068
rect 5408 -26212 5472 -26148
rect 5408 -26292 5472 -26228
rect 5408 -26372 5472 -26308
rect 5408 -26452 5472 -26388
rect 11020 -21492 11084 -21428
rect 11020 -21572 11084 -21508
rect 11020 -21652 11084 -21588
rect 11020 -21732 11084 -21668
rect 11020 -21812 11084 -21748
rect 11020 -21892 11084 -21828
rect 11020 -21972 11084 -21908
rect 11020 -22052 11084 -21988
rect 11020 -22132 11084 -22068
rect 11020 -22212 11084 -22148
rect 11020 -22292 11084 -22228
rect 11020 -22372 11084 -22308
rect 11020 -22452 11084 -22388
rect 11020 -22532 11084 -22468
rect 11020 -22612 11084 -22548
rect 11020 -22692 11084 -22628
rect 11020 -22772 11084 -22708
rect 11020 -22852 11084 -22788
rect 11020 -22932 11084 -22868
rect 11020 -23012 11084 -22948
rect 11020 -23092 11084 -23028
rect 11020 -23172 11084 -23108
rect 11020 -23252 11084 -23188
rect 11020 -23332 11084 -23268
rect 11020 -23412 11084 -23348
rect 11020 -23492 11084 -23428
rect 11020 -23572 11084 -23508
rect 11020 -23652 11084 -23588
rect 11020 -23732 11084 -23668
rect 11020 -23812 11084 -23748
rect 11020 -23892 11084 -23828
rect 11020 -23972 11084 -23908
rect 11020 -24052 11084 -23988
rect 11020 -24132 11084 -24068
rect 11020 -24212 11084 -24148
rect 11020 -24292 11084 -24228
rect 11020 -24372 11084 -24308
rect 11020 -24452 11084 -24388
rect 11020 -24532 11084 -24468
rect 11020 -24612 11084 -24548
rect 11020 -24692 11084 -24628
rect 11020 -24772 11084 -24708
rect 11020 -24852 11084 -24788
rect 11020 -24932 11084 -24868
rect 11020 -25012 11084 -24948
rect 11020 -25092 11084 -25028
rect 11020 -25172 11084 -25108
rect 11020 -25252 11084 -25188
rect 11020 -25332 11084 -25268
rect 11020 -25412 11084 -25348
rect 11020 -25492 11084 -25428
rect 11020 -25572 11084 -25508
rect 11020 -25652 11084 -25588
rect 11020 -25732 11084 -25668
rect 11020 -25812 11084 -25748
rect 11020 -25892 11084 -25828
rect 11020 -25972 11084 -25908
rect 11020 -26052 11084 -25988
rect 11020 -26132 11084 -26068
rect 11020 -26212 11084 -26148
rect 11020 -26292 11084 -26228
rect 11020 -26372 11084 -26308
rect 11020 -26452 11084 -26388
rect 16632 -21492 16696 -21428
rect 16632 -21572 16696 -21508
rect 16632 -21652 16696 -21588
rect 16632 -21732 16696 -21668
rect 16632 -21812 16696 -21748
rect 16632 -21892 16696 -21828
rect 16632 -21972 16696 -21908
rect 16632 -22052 16696 -21988
rect 16632 -22132 16696 -22068
rect 16632 -22212 16696 -22148
rect 16632 -22292 16696 -22228
rect 16632 -22372 16696 -22308
rect 16632 -22452 16696 -22388
rect 16632 -22532 16696 -22468
rect 16632 -22612 16696 -22548
rect 16632 -22692 16696 -22628
rect 16632 -22772 16696 -22708
rect 16632 -22852 16696 -22788
rect 16632 -22932 16696 -22868
rect 16632 -23012 16696 -22948
rect 16632 -23092 16696 -23028
rect 16632 -23172 16696 -23108
rect 16632 -23252 16696 -23188
rect 16632 -23332 16696 -23268
rect 16632 -23412 16696 -23348
rect 16632 -23492 16696 -23428
rect 16632 -23572 16696 -23508
rect 16632 -23652 16696 -23588
rect 16632 -23732 16696 -23668
rect 16632 -23812 16696 -23748
rect 16632 -23892 16696 -23828
rect 16632 -23972 16696 -23908
rect 16632 -24052 16696 -23988
rect 16632 -24132 16696 -24068
rect 16632 -24212 16696 -24148
rect 16632 -24292 16696 -24228
rect 16632 -24372 16696 -24308
rect 16632 -24452 16696 -24388
rect 16632 -24532 16696 -24468
rect 16632 -24612 16696 -24548
rect 16632 -24692 16696 -24628
rect 16632 -24772 16696 -24708
rect 16632 -24852 16696 -24788
rect 16632 -24932 16696 -24868
rect 16632 -25012 16696 -24948
rect 16632 -25092 16696 -25028
rect 16632 -25172 16696 -25108
rect 16632 -25252 16696 -25188
rect 16632 -25332 16696 -25268
rect 16632 -25412 16696 -25348
rect 16632 -25492 16696 -25428
rect 16632 -25572 16696 -25508
rect 16632 -25652 16696 -25588
rect 16632 -25732 16696 -25668
rect 16632 -25812 16696 -25748
rect 16632 -25892 16696 -25828
rect 16632 -25972 16696 -25908
rect 16632 -26052 16696 -25988
rect 16632 -26132 16696 -26068
rect 16632 -26212 16696 -26148
rect 16632 -26292 16696 -26228
rect 16632 -26372 16696 -26308
rect 16632 -26452 16696 -26388
rect 22244 -21492 22308 -21428
rect 22244 -21572 22308 -21508
rect 22244 -21652 22308 -21588
rect 22244 -21732 22308 -21668
rect 22244 -21812 22308 -21748
rect 22244 -21892 22308 -21828
rect 22244 -21972 22308 -21908
rect 22244 -22052 22308 -21988
rect 22244 -22132 22308 -22068
rect 22244 -22212 22308 -22148
rect 22244 -22292 22308 -22228
rect 22244 -22372 22308 -22308
rect 22244 -22452 22308 -22388
rect 22244 -22532 22308 -22468
rect 22244 -22612 22308 -22548
rect 22244 -22692 22308 -22628
rect 22244 -22772 22308 -22708
rect 22244 -22852 22308 -22788
rect 22244 -22932 22308 -22868
rect 22244 -23012 22308 -22948
rect 22244 -23092 22308 -23028
rect 22244 -23172 22308 -23108
rect 22244 -23252 22308 -23188
rect 22244 -23332 22308 -23268
rect 22244 -23412 22308 -23348
rect 22244 -23492 22308 -23428
rect 22244 -23572 22308 -23508
rect 22244 -23652 22308 -23588
rect 22244 -23732 22308 -23668
rect 22244 -23812 22308 -23748
rect 22244 -23892 22308 -23828
rect 22244 -23972 22308 -23908
rect 22244 -24052 22308 -23988
rect 22244 -24132 22308 -24068
rect 22244 -24212 22308 -24148
rect 22244 -24292 22308 -24228
rect 22244 -24372 22308 -24308
rect 22244 -24452 22308 -24388
rect 22244 -24532 22308 -24468
rect 22244 -24612 22308 -24548
rect 22244 -24692 22308 -24628
rect 22244 -24772 22308 -24708
rect 22244 -24852 22308 -24788
rect 22244 -24932 22308 -24868
rect 22244 -25012 22308 -24948
rect 22244 -25092 22308 -25028
rect 22244 -25172 22308 -25108
rect 22244 -25252 22308 -25188
rect 22244 -25332 22308 -25268
rect 22244 -25412 22308 -25348
rect 22244 -25492 22308 -25428
rect 22244 -25572 22308 -25508
rect 22244 -25652 22308 -25588
rect 22244 -25732 22308 -25668
rect 22244 -25812 22308 -25748
rect 22244 -25892 22308 -25828
rect 22244 -25972 22308 -25908
rect 22244 -26052 22308 -25988
rect 22244 -26132 22308 -26068
rect 22244 -26212 22308 -26148
rect 22244 -26292 22308 -26228
rect 22244 -26372 22308 -26308
rect 22244 -26452 22308 -26388
rect 27856 -21492 27920 -21428
rect 27856 -21572 27920 -21508
rect 27856 -21652 27920 -21588
rect 27856 -21732 27920 -21668
rect 27856 -21812 27920 -21748
rect 27856 -21892 27920 -21828
rect 27856 -21972 27920 -21908
rect 27856 -22052 27920 -21988
rect 27856 -22132 27920 -22068
rect 27856 -22212 27920 -22148
rect 27856 -22292 27920 -22228
rect 27856 -22372 27920 -22308
rect 27856 -22452 27920 -22388
rect 27856 -22532 27920 -22468
rect 27856 -22612 27920 -22548
rect 27856 -22692 27920 -22628
rect 27856 -22772 27920 -22708
rect 27856 -22852 27920 -22788
rect 27856 -22932 27920 -22868
rect 27856 -23012 27920 -22948
rect 27856 -23092 27920 -23028
rect 27856 -23172 27920 -23108
rect 27856 -23252 27920 -23188
rect 27856 -23332 27920 -23268
rect 27856 -23412 27920 -23348
rect 27856 -23492 27920 -23428
rect 27856 -23572 27920 -23508
rect 27856 -23652 27920 -23588
rect 27856 -23732 27920 -23668
rect 27856 -23812 27920 -23748
rect 27856 -23892 27920 -23828
rect 27856 -23972 27920 -23908
rect 27856 -24052 27920 -23988
rect 27856 -24132 27920 -24068
rect 27856 -24212 27920 -24148
rect 27856 -24292 27920 -24228
rect 27856 -24372 27920 -24308
rect 27856 -24452 27920 -24388
rect 27856 -24532 27920 -24468
rect 27856 -24612 27920 -24548
rect 27856 -24692 27920 -24628
rect 27856 -24772 27920 -24708
rect 27856 -24852 27920 -24788
rect 27856 -24932 27920 -24868
rect 27856 -25012 27920 -24948
rect 27856 -25092 27920 -25028
rect 27856 -25172 27920 -25108
rect 27856 -25252 27920 -25188
rect 27856 -25332 27920 -25268
rect 27856 -25412 27920 -25348
rect 27856 -25492 27920 -25428
rect 27856 -25572 27920 -25508
rect 27856 -25652 27920 -25588
rect 27856 -25732 27920 -25668
rect 27856 -25812 27920 -25748
rect 27856 -25892 27920 -25828
rect 27856 -25972 27920 -25908
rect 27856 -26052 27920 -25988
rect 27856 -26132 27920 -26068
rect 27856 -26212 27920 -26148
rect 27856 -26292 27920 -26228
rect 27856 -26372 27920 -26308
rect 27856 -26452 27920 -26388
rect 33468 -21492 33532 -21428
rect 33468 -21572 33532 -21508
rect 33468 -21652 33532 -21588
rect 33468 -21732 33532 -21668
rect 33468 -21812 33532 -21748
rect 33468 -21892 33532 -21828
rect 33468 -21972 33532 -21908
rect 33468 -22052 33532 -21988
rect 33468 -22132 33532 -22068
rect 33468 -22212 33532 -22148
rect 33468 -22292 33532 -22228
rect 33468 -22372 33532 -22308
rect 33468 -22452 33532 -22388
rect 33468 -22532 33532 -22468
rect 33468 -22612 33532 -22548
rect 33468 -22692 33532 -22628
rect 33468 -22772 33532 -22708
rect 33468 -22852 33532 -22788
rect 33468 -22932 33532 -22868
rect 33468 -23012 33532 -22948
rect 33468 -23092 33532 -23028
rect 33468 -23172 33532 -23108
rect 33468 -23252 33532 -23188
rect 33468 -23332 33532 -23268
rect 33468 -23412 33532 -23348
rect 33468 -23492 33532 -23428
rect 33468 -23572 33532 -23508
rect 33468 -23652 33532 -23588
rect 33468 -23732 33532 -23668
rect 33468 -23812 33532 -23748
rect 33468 -23892 33532 -23828
rect 33468 -23972 33532 -23908
rect 33468 -24052 33532 -23988
rect 33468 -24132 33532 -24068
rect 33468 -24212 33532 -24148
rect 33468 -24292 33532 -24228
rect 33468 -24372 33532 -24308
rect 33468 -24452 33532 -24388
rect 33468 -24532 33532 -24468
rect 33468 -24612 33532 -24548
rect 33468 -24692 33532 -24628
rect 33468 -24772 33532 -24708
rect 33468 -24852 33532 -24788
rect 33468 -24932 33532 -24868
rect 33468 -25012 33532 -24948
rect 33468 -25092 33532 -25028
rect 33468 -25172 33532 -25108
rect 33468 -25252 33532 -25188
rect 33468 -25332 33532 -25268
rect 33468 -25412 33532 -25348
rect 33468 -25492 33532 -25428
rect 33468 -25572 33532 -25508
rect 33468 -25652 33532 -25588
rect 33468 -25732 33532 -25668
rect 33468 -25812 33532 -25748
rect 33468 -25892 33532 -25828
rect 33468 -25972 33532 -25908
rect 33468 -26052 33532 -25988
rect 33468 -26132 33532 -26068
rect 33468 -26212 33532 -26148
rect 33468 -26292 33532 -26228
rect 33468 -26372 33532 -26308
rect 33468 -26452 33532 -26388
rect 39080 -21492 39144 -21428
rect 39080 -21572 39144 -21508
rect 39080 -21652 39144 -21588
rect 39080 -21732 39144 -21668
rect 39080 -21812 39144 -21748
rect 39080 -21892 39144 -21828
rect 39080 -21972 39144 -21908
rect 39080 -22052 39144 -21988
rect 39080 -22132 39144 -22068
rect 39080 -22212 39144 -22148
rect 39080 -22292 39144 -22228
rect 39080 -22372 39144 -22308
rect 39080 -22452 39144 -22388
rect 39080 -22532 39144 -22468
rect 39080 -22612 39144 -22548
rect 39080 -22692 39144 -22628
rect 39080 -22772 39144 -22708
rect 39080 -22852 39144 -22788
rect 39080 -22932 39144 -22868
rect 39080 -23012 39144 -22948
rect 39080 -23092 39144 -23028
rect 39080 -23172 39144 -23108
rect 39080 -23252 39144 -23188
rect 39080 -23332 39144 -23268
rect 39080 -23412 39144 -23348
rect 39080 -23492 39144 -23428
rect 39080 -23572 39144 -23508
rect 39080 -23652 39144 -23588
rect 39080 -23732 39144 -23668
rect 39080 -23812 39144 -23748
rect 39080 -23892 39144 -23828
rect 39080 -23972 39144 -23908
rect 39080 -24052 39144 -23988
rect 39080 -24132 39144 -24068
rect 39080 -24212 39144 -24148
rect 39080 -24292 39144 -24228
rect 39080 -24372 39144 -24308
rect 39080 -24452 39144 -24388
rect 39080 -24532 39144 -24468
rect 39080 -24612 39144 -24548
rect 39080 -24692 39144 -24628
rect 39080 -24772 39144 -24708
rect 39080 -24852 39144 -24788
rect 39080 -24932 39144 -24868
rect 39080 -25012 39144 -24948
rect 39080 -25092 39144 -25028
rect 39080 -25172 39144 -25108
rect 39080 -25252 39144 -25188
rect 39080 -25332 39144 -25268
rect 39080 -25412 39144 -25348
rect 39080 -25492 39144 -25428
rect 39080 -25572 39144 -25508
rect 39080 -25652 39144 -25588
rect 39080 -25732 39144 -25668
rect 39080 -25812 39144 -25748
rect 39080 -25892 39144 -25828
rect 39080 -25972 39144 -25908
rect 39080 -26052 39144 -25988
rect 39080 -26132 39144 -26068
rect 39080 -26212 39144 -26148
rect 39080 -26292 39144 -26228
rect 39080 -26372 39144 -26308
rect 39080 -26452 39144 -26388
rect -33876 -26812 -33812 -26748
rect -33876 -26892 -33812 -26828
rect -33876 -26972 -33812 -26908
rect -33876 -27052 -33812 -26988
rect -33876 -27132 -33812 -27068
rect -33876 -27212 -33812 -27148
rect -33876 -27292 -33812 -27228
rect -33876 -27372 -33812 -27308
rect -33876 -27452 -33812 -27388
rect -33876 -27532 -33812 -27468
rect -33876 -27612 -33812 -27548
rect -33876 -27692 -33812 -27628
rect -33876 -27772 -33812 -27708
rect -33876 -27852 -33812 -27788
rect -33876 -27932 -33812 -27868
rect -33876 -28012 -33812 -27948
rect -33876 -28092 -33812 -28028
rect -33876 -28172 -33812 -28108
rect -33876 -28252 -33812 -28188
rect -33876 -28332 -33812 -28268
rect -33876 -28412 -33812 -28348
rect -33876 -28492 -33812 -28428
rect -33876 -28572 -33812 -28508
rect -33876 -28652 -33812 -28588
rect -33876 -28732 -33812 -28668
rect -33876 -28812 -33812 -28748
rect -33876 -28892 -33812 -28828
rect -33876 -28972 -33812 -28908
rect -33876 -29052 -33812 -28988
rect -33876 -29132 -33812 -29068
rect -33876 -29212 -33812 -29148
rect -33876 -29292 -33812 -29228
rect -33876 -29372 -33812 -29308
rect -33876 -29452 -33812 -29388
rect -33876 -29532 -33812 -29468
rect -33876 -29612 -33812 -29548
rect -33876 -29692 -33812 -29628
rect -33876 -29772 -33812 -29708
rect -33876 -29852 -33812 -29788
rect -33876 -29932 -33812 -29868
rect -33876 -30012 -33812 -29948
rect -33876 -30092 -33812 -30028
rect -33876 -30172 -33812 -30108
rect -33876 -30252 -33812 -30188
rect -33876 -30332 -33812 -30268
rect -33876 -30412 -33812 -30348
rect -33876 -30492 -33812 -30428
rect -33876 -30572 -33812 -30508
rect -33876 -30652 -33812 -30588
rect -33876 -30732 -33812 -30668
rect -33876 -30812 -33812 -30748
rect -33876 -30892 -33812 -30828
rect -33876 -30972 -33812 -30908
rect -33876 -31052 -33812 -30988
rect -33876 -31132 -33812 -31068
rect -33876 -31212 -33812 -31148
rect -33876 -31292 -33812 -31228
rect -33876 -31372 -33812 -31308
rect -33876 -31452 -33812 -31388
rect -33876 -31532 -33812 -31468
rect -33876 -31612 -33812 -31548
rect -33876 -31692 -33812 -31628
rect -33876 -31772 -33812 -31708
rect -28264 -26812 -28200 -26748
rect -28264 -26892 -28200 -26828
rect -28264 -26972 -28200 -26908
rect -28264 -27052 -28200 -26988
rect -28264 -27132 -28200 -27068
rect -28264 -27212 -28200 -27148
rect -28264 -27292 -28200 -27228
rect -28264 -27372 -28200 -27308
rect -28264 -27452 -28200 -27388
rect -28264 -27532 -28200 -27468
rect -28264 -27612 -28200 -27548
rect -28264 -27692 -28200 -27628
rect -28264 -27772 -28200 -27708
rect -28264 -27852 -28200 -27788
rect -28264 -27932 -28200 -27868
rect -28264 -28012 -28200 -27948
rect -28264 -28092 -28200 -28028
rect -28264 -28172 -28200 -28108
rect -28264 -28252 -28200 -28188
rect -28264 -28332 -28200 -28268
rect -28264 -28412 -28200 -28348
rect -28264 -28492 -28200 -28428
rect -28264 -28572 -28200 -28508
rect -28264 -28652 -28200 -28588
rect -28264 -28732 -28200 -28668
rect -28264 -28812 -28200 -28748
rect -28264 -28892 -28200 -28828
rect -28264 -28972 -28200 -28908
rect -28264 -29052 -28200 -28988
rect -28264 -29132 -28200 -29068
rect -28264 -29212 -28200 -29148
rect -28264 -29292 -28200 -29228
rect -28264 -29372 -28200 -29308
rect -28264 -29452 -28200 -29388
rect -28264 -29532 -28200 -29468
rect -28264 -29612 -28200 -29548
rect -28264 -29692 -28200 -29628
rect -28264 -29772 -28200 -29708
rect -28264 -29852 -28200 -29788
rect -28264 -29932 -28200 -29868
rect -28264 -30012 -28200 -29948
rect -28264 -30092 -28200 -30028
rect -28264 -30172 -28200 -30108
rect -28264 -30252 -28200 -30188
rect -28264 -30332 -28200 -30268
rect -28264 -30412 -28200 -30348
rect -28264 -30492 -28200 -30428
rect -28264 -30572 -28200 -30508
rect -28264 -30652 -28200 -30588
rect -28264 -30732 -28200 -30668
rect -28264 -30812 -28200 -30748
rect -28264 -30892 -28200 -30828
rect -28264 -30972 -28200 -30908
rect -28264 -31052 -28200 -30988
rect -28264 -31132 -28200 -31068
rect -28264 -31212 -28200 -31148
rect -28264 -31292 -28200 -31228
rect -28264 -31372 -28200 -31308
rect -28264 -31452 -28200 -31388
rect -28264 -31532 -28200 -31468
rect -28264 -31612 -28200 -31548
rect -28264 -31692 -28200 -31628
rect -28264 -31772 -28200 -31708
rect -22652 -26812 -22588 -26748
rect -22652 -26892 -22588 -26828
rect -22652 -26972 -22588 -26908
rect -22652 -27052 -22588 -26988
rect -22652 -27132 -22588 -27068
rect -22652 -27212 -22588 -27148
rect -22652 -27292 -22588 -27228
rect -22652 -27372 -22588 -27308
rect -22652 -27452 -22588 -27388
rect -22652 -27532 -22588 -27468
rect -22652 -27612 -22588 -27548
rect -22652 -27692 -22588 -27628
rect -22652 -27772 -22588 -27708
rect -22652 -27852 -22588 -27788
rect -22652 -27932 -22588 -27868
rect -22652 -28012 -22588 -27948
rect -22652 -28092 -22588 -28028
rect -22652 -28172 -22588 -28108
rect -22652 -28252 -22588 -28188
rect -22652 -28332 -22588 -28268
rect -22652 -28412 -22588 -28348
rect -22652 -28492 -22588 -28428
rect -22652 -28572 -22588 -28508
rect -22652 -28652 -22588 -28588
rect -22652 -28732 -22588 -28668
rect -22652 -28812 -22588 -28748
rect -22652 -28892 -22588 -28828
rect -22652 -28972 -22588 -28908
rect -22652 -29052 -22588 -28988
rect -22652 -29132 -22588 -29068
rect -22652 -29212 -22588 -29148
rect -22652 -29292 -22588 -29228
rect -22652 -29372 -22588 -29308
rect -22652 -29452 -22588 -29388
rect -22652 -29532 -22588 -29468
rect -22652 -29612 -22588 -29548
rect -22652 -29692 -22588 -29628
rect -22652 -29772 -22588 -29708
rect -22652 -29852 -22588 -29788
rect -22652 -29932 -22588 -29868
rect -22652 -30012 -22588 -29948
rect -22652 -30092 -22588 -30028
rect -22652 -30172 -22588 -30108
rect -22652 -30252 -22588 -30188
rect -22652 -30332 -22588 -30268
rect -22652 -30412 -22588 -30348
rect -22652 -30492 -22588 -30428
rect -22652 -30572 -22588 -30508
rect -22652 -30652 -22588 -30588
rect -22652 -30732 -22588 -30668
rect -22652 -30812 -22588 -30748
rect -22652 -30892 -22588 -30828
rect -22652 -30972 -22588 -30908
rect -22652 -31052 -22588 -30988
rect -22652 -31132 -22588 -31068
rect -22652 -31212 -22588 -31148
rect -22652 -31292 -22588 -31228
rect -22652 -31372 -22588 -31308
rect -22652 -31452 -22588 -31388
rect -22652 -31532 -22588 -31468
rect -22652 -31612 -22588 -31548
rect -22652 -31692 -22588 -31628
rect -22652 -31772 -22588 -31708
rect -17040 -26812 -16976 -26748
rect -17040 -26892 -16976 -26828
rect -17040 -26972 -16976 -26908
rect -17040 -27052 -16976 -26988
rect -17040 -27132 -16976 -27068
rect -17040 -27212 -16976 -27148
rect -17040 -27292 -16976 -27228
rect -17040 -27372 -16976 -27308
rect -17040 -27452 -16976 -27388
rect -17040 -27532 -16976 -27468
rect -17040 -27612 -16976 -27548
rect -17040 -27692 -16976 -27628
rect -17040 -27772 -16976 -27708
rect -17040 -27852 -16976 -27788
rect -17040 -27932 -16976 -27868
rect -17040 -28012 -16976 -27948
rect -17040 -28092 -16976 -28028
rect -17040 -28172 -16976 -28108
rect -17040 -28252 -16976 -28188
rect -17040 -28332 -16976 -28268
rect -17040 -28412 -16976 -28348
rect -17040 -28492 -16976 -28428
rect -17040 -28572 -16976 -28508
rect -17040 -28652 -16976 -28588
rect -17040 -28732 -16976 -28668
rect -17040 -28812 -16976 -28748
rect -17040 -28892 -16976 -28828
rect -17040 -28972 -16976 -28908
rect -17040 -29052 -16976 -28988
rect -17040 -29132 -16976 -29068
rect -17040 -29212 -16976 -29148
rect -17040 -29292 -16976 -29228
rect -17040 -29372 -16976 -29308
rect -17040 -29452 -16976 -29388
rect -17040 -29532 -16976 -29468
rect -17040 -29612 -16976 -29548
rect -17040 -29692 -16976 -29628
rect -17040 -29772 -16976 -29708
rect -17040 -29852 -16976 -29788
rect -17040 -29932 -16976 -29868
rect -17040 -30012 -16976 -29948
rect -17040 -30092 -16976 -30028
rect -17040 -30172 -16976 -30108
rect -17040 -30252 -16976 -30188
rect -17040 -30332 -16976 -30268
rect -17040 -30412 -16976 -30348
rect -17040 -30492 -16976 -30428
rect -17040 -30572 -16976 -30508
rect -17040 -30652 -16976 -30588
rect -17040 -30732 -16976 -30668
rect -17040 -30812 -16976 -30748
rect -17040 -30892 -16976 -30828
rect -17040 -30972 -16976 -30908
rect -17040 -31052 -16976 -30988
rect -17040 -31132 -16976 -31068
rect -17040 -31212 -16976 -31148
rect -17040 -31292 -16976 -31228
rect -17040 -31372 -16976 -31308
rect -17040 -31452 -16976 -31388
rect -17040 -31532 -16976 -31468
rect -17040 -31612 -16976 -31548
rect -17040 -31692 -16976 -31628
rect -17040 -31772 -16976 -31708
rect -11428 -26812 -11364 -26748
rect -11428 -26892 -11364 -26828
rect -11428 -26972 -11364 -26908
rect -11428 -27052 -11364 -26988
rect -11428 -27132 -11364 -27068
rect -11428 -27212 -11364 -27148
rect -11428 -27292 -11364 -27228
rect -11428 -27372 -11364 -27308
rect -11428 -27452 -11364 -27388
rect -11428 -27532 -11364 -27468
rect -11428 -27612 -11364 -27548
rect -11428 -27692 -11364 -27628
rect -11428 -27772 -11364 -27708
rect -11428 -27852 -11364 -27788
rect -11428 -27932 -11364 -27868
rect -11428 -28012 -11364 -27948
rect -11428 -28092 -11364 -28028
rect -11428 -28172 -11364 -28108
rect -11428 -28252 -11364 -28188
rect -11428 -28332 -11364 -28268
rect -11428 -28412 -11364 -28348
rect -11428 -28492 -11364 -28428
rect -11428 -28572 -11364 -28508
rect -11428 -28652 -11364 -28588
rect -11428 -28732 -11364 -28668
rect -11428 -28812 -11364 -28748
rect -11428 -28892 -11364 -28828
rect -11428 -28972 -11364 -28908
rect -11428 -29052 -11364 -28988
rect -11428 -29132 -11364 -29068
rect -11428 -29212 -11364 -29148
rect -11428 -29292 -11364 -29228
rect -11428 -29372 -11364 -29308
rect -11428 -29452 -11364 -29388
rect -11428 -29532 -11364 -29468
rect -11428 -29612 -11364 -29548
rect -11428 -29692 -11364 -29628
rect -11428 -29772 -11364 -29708
rect -11428 -29852 -11364 -29788
rect -11428 -29932 -11364 -29868
rect -11428 -30012 -11364 -29948
rect -11428 -30092 -11364 -30028
rect -11428 -30172 -11364 -30108
rect -11428 -30252 -11364 -30188
rect -11428 -30332 -11364 -30268
rect -11428 -30412 -11364 -30348
rect -11428 -30492 -11364 -30428
rect -11428 -30572 -11364 -30508
rect -11428 -30652 -11364 -30588
rect -11428 -30732 -11364 -30668
rect -11428 -30812 -11364 -30748
rect -11428 -30892 -11364 -30828
rect -11428 -30972 -11364 -30908
rect -11428 -31052 -11364 -30988
rect -11428 -31132 -11364 -31068
rect -11428 -31212 -11364 -31148
rect -11428 -31292 -11364 -31228
rect -11428 -31372 -11364 -31308
rect -11428 -31452 -11364 -31388
rect -11428 -31532 -11364 -31468
rect -11428 -31612 -11364 -31548
rect -11428 -31692 -11364 -31628
rect -11428 -31772 -11364 -31708
rect -5816 -26812 -5752 -26748
rect -5816 -26892 -5752 -26828
rect -5816 -26972 -5752 -26908
rect -5816 -27052 -5752 -26988
rect -5816 -27132 -5752 -27068
rect -5816 -27212 -5752 -27148
rect -5816 -27292 -5752 -27228
rect -5816 -27372 -5752 -27308
rect -5816 -27452 -5752 -27388
rect -5816 -27532 -5752 -27468
rect -5816 -27612 -5752 -27548
rect -5816 -27692 -5752 -27628
rect -5816 -27772 -5752 -27708
rect -5816 -27852 -5752 -27788
rect -5816 -27932 -5752 -27868
rect -5816 -28012 -5752 -27948
rect -5816 -28092 -5752 -28028
rect -5816 -28172 -5752 -28108
rect -5816 -28252 -5752 -28188
rect -5816 -28332 -5752 -28268
rect -5816 -28412 -5752 -28348
rect -5816 -28492 -5752 -28428
rect -5816 -28572 -5752 -28508
rect -5816 -28652 -5752 -28588
rect -5816 -28732 -5752 -28668
rect -5816 -28812 -5752 -28748
rect -5816 -28892 -5752 -28828
rect -5816 -28972 -5752 -28908
rect -5816 -29052 -5752 -28988
rect -5816 -29132 -5752 -29068
rect -5816 -29212 -5752 -29148
rect -5816 -29292 -5752 -29228
rect -5816 -29372 -5752 -29308
rect -5816 -29452 -5752 -29388
rect -5816 -29532 -5752 -29468
rect -5816 -29612 -5752 -29548
rect -5816 -29692 -5752 -29628
rect -5816 -29772 -5752 -29708
rect -5816 -29852 -5752 -29788
rect -5816 -29932 -5752 -29868
rect -5816 -30012 -5752 -29948
rect -5816 -30092 -5752 -30028
rect -5816 -30172 -5752 -30108
rect -5816 -30252 -5752 -30188
rect -5816 -30332 -5752 -30268
rect -5816 -30412 -5752 -30348
rect -5816 -30492 -5752 -30428
rect -5816 -30572 -5752 -30508
rect -5816 -30652 -5752 -30588
rect -5816 -30732 -5752 -30668
rect -5816 -30812 -5752 -30748
rect -5816 -30892 -5752 -30828
rect -5816 -30972 -5752 -30908
rect -5816 -31052 -5752 -30988
rect -5816 -31132 -5752 -31068
rect -5816 -31212 -5752 -31148
rect -5816 -31292 -5752 -31228
rect -5816 -31372 -5752 -31308
rect -5816 -31452 -5752 -31388
rect -5816 -31532 -5752 -31468
rect -5816 -31612 -5752 -31548
rect -5816 -31692 -5752 -31628
rect -5816 -31772 -5752 -31708
rect -204 -26812 -140 -26748
rect -204 -26892 -140 -26828
rect -204 -26972 -140 -26908
rect -204 -27052 -140 -26988
rect -204 -27132 -140 -27068
rect -204 -27212 -140 -27148
rect -204 -27292 -140 -27228
rect -204 -27372 -140 -27308
rect -204 -27452 -140 -27388
rect -204 -27532 -140 -27468
rect -204 -27612 -140 -27548
rect -204 -27692 -140 -27628
rect -204 -27772 -140 -27708
rect -204 -27852 -140 -27788
rect -204 -27932 -140 -27868
rect -204 -28012 -140 -27948
rect -204 -28092 -140 -28028
rect -204 -28172 -140 -28108
rect -204 -28252 -140 -28188
rect -204 -28332 -140 -28268
rect -204 -28412 -140 -28348
rect -204 -28492 -140 -28428
rect -204 -28572 -140 -28508
rect -204 -28652 -140 -28588
rect -204 -28732 -140 -28668
rect -204 -28812 -140 -28748
rect -204 -28892 -140 -28828
rect -204 -28972 -140 -28908
rect -204 -29052 -140 -28988
rect -204 -29132 -140 -29068
rect -204 -29212 -140 -29148
rect -204 -29292 -140 -29228
rect -204 -29372 -140 -29308
rect -204 -29452 -140 -29388
rect -204 -29532 -140 -29468
rect -204 -29612 -140 -29548
rect -204 -29692 -140 -29628
rect -204 -29772 -140 -29708
rect -204 -29852 -140 -29788
rect -204 -29932 -140 -29868
rect -204 -30012 -140 -29948
rect -204 -30092 -140 -30028
rect -204 -30172 -140 -30108
rect -204 -30252 -140 -30188
rect -204 -30332 -140 -30268
rect -204 -30412 -140 -30348
rect -204 -30492 -140 -30428
rect -204 -30572 -140 -30508
rect -204 -30652 -140 -30588
rect -204 -30732 -140 -30668
rect -204 -30812 -140 -30748
rect -204 -30892 -140 -30828
rect -204 -30972 -140 -30908
rect -204 -31052 -140 -30988
rect -204 -31132 -140 -31068
rect -204 -31212 -140 -31148
rect -204 -31292 -140 -31228
rect -204 -31372 -140 -31308
rect -204 -31452 -140 -31388
rect -204 -31532 -140 -31468
rect -204 -31612 -140 -31548
rect -204 -31692 -140 -31628
rect -204 -31772 -140 -31708
rect 5408 -26812 5472 -26748
rect 5408 -26892 5472 -26828
rect 5408 -26972 5472 -26908
rect 5408 -27052 5472 -26988
rect 5408 -27132 5472 -27068
rect 5408 -27212 5472 -27148
rect 5408 -27292 5472 -27228
rect 5408 -27372 5472 -27308
rect 5408 -27452 5472 -27388
rect 5408 -27532 5472 -27468
rect 5408 -27612 5472 -27548
rect 5408 -27692 5472 -27628
rect 5408 -27772 5472 -27708
rect 5408 -27852 5472 -27788
rect 5408 -27932 5472 -27868
rect 5408 -28012 5472 -27948
rect 5408 -28092 5472 -28028
rect 5408 -28172 5472 -28108
rect 5408 -28252 5472 -28188
rect 5408 -28332 5472 -28268
rect 5408 -28412 5472 -28348
rect 5408 -28492 5472 -28428
rect 5408 -28572 5472 -28508
rect 5408 -28652 5472 -28588
rect 5408 -28732 5472 -28668
rect 5408 -28812 5472 -28748
rect 5408 -28892 5472 -28828
rect 5408 -28972 5472 -28908
rect 5408 -29052 5472 -28988
rect 5408 -29132 5472 -29068
rect 5408 -29212 5472 -29148
rect 5408 -29292 5472 -29228
rect 5408 -29372 5472 -29308
rect 5408 -29452 5472 -29388
rect 5408 -29532 5472 -29468
rect 5408 -29612 5472 -29548
rect 5408 -29692 5472 -29628
rect 5408 -29772 5472 -29708
rect 5408 -29852 5472 -29788
rect 5408 -29932 5472 -29868
rect 5408 -30012 5472 -29948
rect 5408 -30092 5472 -30028
rect 5408 -30172 5472 -30108
rect 5408 -30252 5472 -30188
rect 5408 -30332 5472 -30268
rect 5408 -30412 5472 -30348
rect 5408 -30492 5472 -30428
rect 5408 -30572 5472 -30508
rect 5408 -30652 5472 -30588
rect 5408 -30732 5472 -30668
rect 5408 -30812 5472 -30748
rect 5408 -30892 5472 -30828
rect 5408 -30972 5472 -30908
rect 5408 -31052 5472 -30988
rect 5408 -31132 5472 -31068
rect 5408 -31212 5472 -31148
rect 5408 -31292 5472 -31228
rect 5408 -31372 5472 -31308
rect 5408 -31452 5472 -31388
rect 5408 -31532 5472 -31468
rect 5408 -31612 5472 -31548
rect 5408 -31692 5472 -31628
rect 5408 -31772 5472 -31708
rect 11020 -26812 11084 -26748
rect 11020 -26892 11084 -26828
rect 11020 -26972 11084 -26908
rect 11020 -27052 11084 -26988
rect 11020 -27132 11084 -27068
rect 11020 -27212 11084 -27148
rect 11020 -27292 11084 -27228
rect 11020 -27372 11084 -27308
rect 11020 -27452 11084 -27388
rect 11020 -27532 11084 -27468
rect 11020 -27612 11084 -27548
rect 11020 -27692 11084 -27628
rect 11020 -27772 11084 -27708
rect 11020 -27852 11084 -27788
rect 11020 -27932 11084 -27868
rect 11020 -28012 11084 -27948
rect 11020 -28092 11084 -28028
rect 11020 -28172 11084 -28108
rect 11020 -28252 11084 -28188
rect 11020 -28332 11084 -28268
rect 11020 -28412 11084 -28348
rect 11020 -28492 11084 -28428
rect 11020 -28572 11084 -28508
rect 11020 -28652 11084 -28588
rect 11020 -28732 11084 -28668
rect 11020 -28812 11084 -28748
rect 11020 -28892 11084 -28828
rect 11020 -28972 11084 -28908
rect 11020 -29052 11084 -28988
rect 11020 -29132 11084 -29068
rect 11020 -29212 11084 -29148
rect 11020 -29292 11084 -29228
rect 11020 -29372 11084 -29308
rect 11020 -29452 11084 -29388
rect 11020 -29532 11084 -29468
rect 11020 -29612 11084 -29548
rect 11020 -29692 11084 -29628
rect 11020 -29772 11084 -29708
rect 11020 -29852 11084 -29788
rect 11020 -29932 11084 -29868
rect 11020 -30012 11084 -29948
rect 11020 -30092 11084 -30028
rect 11020 -30172 11084 -30108
rect 11020 -30252 11084 -30188
rect 11020 -30332 11084 -30268
rect 11020 -30412 11084 -30348
rect 11020 -30492 11084 -30428
rect 11020 -30572 11084 -30508
rect 11020 -30652 11084 -30588
rect 11020 -30732 11084 -30668
rect 11020 -30812 11084 -30748
rect 11020 -30892 11084 -30828
rect 11020 -30972 11084 -30908
rect 11020 -31052 11084 -30988
rect 11020 -31132 11084 -31068
rect 11020 -31212 11084 -31148
rect 11020 -31292 11084 -31228
rect 11020 -31372 11084 -31308
rect 11020 -31452 11084 -31388
rect 11020 -31532 11084 -31468
rect 11020 -31612 11084 -31548
rect 11020 -31692 11084 -31628
rect 11020 -31772 11084 -31708
rect 16632 -26812 16696 -26748
rect 16632 -26892 16696 -26828
rect 16632 -26972 16696 -26908
rect 16632 -27052 16696 -26988
rect 16632 -27132 16696 -27068
rect 16632 -27212 16696 -27148
rect 16632 -27292 16696 -27228
rect 16632 -27372 16696 -27308
rect 16632 -27452 16696 -27388
rect 16632 -27532 16696 -27468
rect 16632 -27612 16696 -27548
rect 16632 -27692 16696 -27628
rect 16632 -27772 16696 -27708
rect 16632 -27852 16696 -27788
rect 16632 -27932 16696 -27868
rect 16632 -28012 16696 -27948
rect 16632 -28092 16696 -28028
rect 16632 -28172 16696 -28108
rect 16632 -28252 16696 -28188
rect 16632 -28332 16696 -28268
rect 16632 -28412 16696 -28348
rect 16632 -28492 16696 -28428
rect 16632 -28572 16696 -28508
rect 16632 -28652 16696 -28588
rect 16632 -28732 16696 -28668
rect 16632 -28812 16696 -28748
rect 16632 -28892 16696 -28828
rect 16632 -28972 16696 -28908
rect 16632 -29052 16696 -28988
rect 16632 -29132 16696 -29068
rect 16632 -29212 16696 -29148
rect 16632 -29292 16696 -29228
rect 16632 -29372 16696 -29308
rect 16632 -29452 16696 -29388
rect 16632 -29532 16696 -29468
rect 16632 -29612 16696 -29548
rect 16632 -29692 16696 -29628
rect 16632 -29772 16696 -29708
rect 16632 -29852 16696 -29788
rect 16632 -29932 16696 -29868
rect 16632 -30012 16696 -29948
rect 16632 -30092 16696 -30028
rect 16632 -30172 16696 -30108
rect 16632 -30252 16696 -30188
rect 16632 -30332 16696 -30268
rect 16632 -30412 16696 -30348
rect 16632 -30492 16696 -30428
rect 16632 -30572 16696 -30508
rect 16632 -30652 16696 -30588
rect 16632 -30732 16696 -30668
rect 16632 -30812 16696 -30748
rect 16632 -30892 16696 -30828
rect 16632 -30972 16696 -30908
rect 16632 -31052 16696 -30988
rect 16632 -31132 16696 -31068
rect 16632 -31212 16696 -31148
rect 16632 -31292 16696 -31228
rect 16632 -31372 16696 -31308
rect 16632 -31452 16696 -31388
rect 16632 -31532 16696 -31468
rect 16632 -31612 16696 -31548
rect 16632 -31692 16696 -31628
rect 16632 -31772 16696 -31708
rect 22244 -26812 22308 -26748
rect 22244 -26892 22308 -26828
rect 22244 -26972 22308 -26908
rect 22244 -27052 22308 -26988
rect 22244 -27132 22308 -27068
rect 22244 -27212 22308 -27148
rect 22244 -27292 22308 -27228
rect 22244 -27372 22308 -27308
rect 22244 -27452 22308 -27388
rect 22244 -27532 22308 -27468
rect 22244 -27612 22308 -27548
rect 22244 -27692 22308 -27628
rect 22244 -27772 22308 -27708
rect 22244 -27852 22308 -27788
rect 22244 -27932 22308 -27868
rect 22244 -28012 22308 -27948
rect 22244 -28092 22308 -28028
rect 22244 -28172 22308 -28108
rect 22244 -28252 22308 -28188
rect 22244 -28332 22308 -28268
rect 22244 -28412 22308 -28348
rect 22244 -28492 22308 -28428
rect 22244 -28572 22308 -28508
rect 22244 -28652 22308 -28588
rect 22244 -28732 22308 -28668
rect 22244 -28812 22308 -28748
rect 22244 -28892 22308 -28828
rect 22244 -28972 22308 -28908
rect 22244 -29052 22308 -28988
rect 22244 -29132 22308 -29068
rect 22244 -29212 22308 -29148
rect 22244 -29292 22308 -29228
rect 22244 -29372 22308 -29308
rect 22244 -29452 22308 -29388
rect 22244 -29532 22308 -29468
rect 22244 -29612 22308 -29548
rect 22244 -29692 22308 -29628
rect 22244 -29772 22308 -29708
rect 22244 -29852 22308 -29788
rect 22244 -29932 22308 -29868
rect 22244 -30012 22308 -29948
rect 22244 -30092 22308 -30028
rect 22244 -30172 22308 -30108
rect 22244 -30252 22308 -30188
rect 22244 -30332 22308 -30268
rect 22244 -30412 22308 -30348
rect 22244 -30492 22308 -30428
rect 22244 -30572 22308 -30508
rect 22244 -30652 22308 -30588
rect 22244 -30732 22308 -30668
rect 22244 -30812 22308 -30748
rect 22244 -30892 22308 -30828
rect 22244 -30972 22308 -30908
rect 22244 -31052 22308 -30988
rect 22244 -31132 22308 -31068
rect 22244 -31212 22308 -31148
rect 22244 -31292 22308 -31228
rect 22244 -31372 22308 -31308
rect 22244 -31452 22308 -31388
rect 22244 -31532 22308 -31468
rect 22244 -31612 22308 -31548
rect 22244 -31692 22308 -31628
rect 22244 -31772 22308 -31708
rect 27856 -26812 27920 -26748
rect 27856 -26892 27920 -26828
rect 27856 -26972 27920 -26908
rect 27856 -27052 27920 -26988
rect 27856 -27132 27920 -27068
rect 27856 -27212 27920 -27148
rect 27856 -27292 27920 -27228
rect 27856 -27372 27920 -27308
rect 27856 -27452 27920 -27388
rect 27856 -27532 27920 -27468
rect 27856 -27612 27920 -27548
rect 27856 -27692 27920 -27628
rect 27856 -27772 27920 -27708
rect 27856 -27852 27920 -27788
rect 27856 -27932 27920 -27868
rect 27856 -28012 27920 -27948
rect 27856 -28092 27920 -28028
rect 27856 -28172 27920 -28108
rect 27856 -28252 27920 -28188
rect 27856 -28332 27920 -28268
rect 27856 -28412 27920 -28348
rect 27856 -28492 27920 -28428
rect 27856 -28572 27920 -28508
rect 27856 -28652 27920 -28588
rect 27856 -28732 27920 -28668
rect 27856 -28812 27920 -28748
rect 27856 -28892 27920 -28828
rect 27856 -28972 27920 -28908
rect 27856 -29052 27920 -28988
rect 27856 -29132 27920 -29068
rect 27856 -29212 27920 -29148
rect 27856 -29292 27920 -29228
rect 27856 -29372 27920 -29308
rect 27856 -29452 27920 -29388
rect 27856 -29532 27920 -29468
rect 27856 -29612 27920 -29548
rect 27856 -29692 27920 -29628
rect 27856 -29772 27920 -29708
rect 27856 -29852 27920 -29788
rect 27856 -29932 27920 -29868
rect 27856 -30012 27920 -29948
rect 27856 -30092 27920 -30028
rect 27856 -30172 27920 -30108
rect 27856 -30252 27920 -30188
rect 27856 -30332 27920 -30268
rect 27856 -30412 27920 -30348
rect 27856 -30492 27920 -30428
rect 27856 -30572 27920 -30508
rect 27856 -30652 27920 -30588
rect 27856 -30732 27920 -30668
rect 27856 -30812 27920 -30748
rect 27856 -30892 27920 -30828
rect 27856 -30972 27920 -30908
rect 27856 -31052 27920 -30988
rect 27856 -31132 27920 -31068
rect 27856 -31212 27920 -31148
rect 27856 -31292 27920 -31228
rect 27856 -31372 27920 -31308
rect 27856 -31452 27920 -31388
rect 27856 -31532 27920 -31468
rect 27856 -31612 27920 -31548
rect 27856 -31692 27920 -31628
rect 27856 -31772 27920 -31708
rect 33468 -26812 33532 -26748
rect 33468 -26892 33532 -26828
rect 33468 -26972 33532 -26908
rect 33468 -27052 33532 -26988
rect 33468 -27132 33532 -27068
rect 33468 -27212 33532 -27148
rect 33468 -27292 33532 -27228
rect 33468 -27372 33532 -27308
rect 33468 -27452 33532 -27388
rect 33468 -27532 33532 -27468
rect 33468 -27612 33532 -27548
rect 33468 -27692 33532 -27628
rect 33468 -27772 33532 -27708
rect 33468 -27852 33532 -27788
rect 33468 -27932 33532 -27868
rect 33468 -28012 33532 -27948
rect 33468 -28092 33532 -28028
rect 33468 -28172 33532 -28108
rect 33468 -28252 33532 -28188
rect 33468 -28332 33532 -28268
rect 33468 -28412 33532 -28348
rect 33468 -28492 33532 -28428
rect 33468 -28572 33532 -28508
rect 33468 -28652 33532 -28588
rect 33468 -28732 33532 -28668
rect 33468 -28812 33532 -28748
rect 33468 -28892 33532 -28828
rect 33468 -28972 33532 -28908
rect 33468 -29052 33532 -28988
rect 33468 -29132 33532 -29068
rect 33468 -29212 33532 -29148
rect 33468 -29292 33532 -29228
rect 33468 -29372 33532 -29308
rect 33468 -29452 33532 -29388
rect 33468 -29532 33532 -29468
rect 33468 -29612 33532 -29548
rect 33468 -29692 33532 -29628
rect 33468 -29772 33532 -29708
rect 33468 -29852 33532 -29788
rect 33468 -29932 33532 -29868
rect 33468 -30012 33532 -29948
rect 33468 -30092 33532 -30028
rect 33468 -30172 33532 -30108
rect 33468 -30252 33532 -30188
rect 33468 -30332 33532 -30268
rect 33468 -30412 33532 -30348
rect 33468 -30492 33532 -30428
rect 33468 -30572 33532 -30508
rect 33468 -30652 33532 -30588
rect 33468 -30732 33532 -30668
rect 33468 -30812 33532 -30748
rect 33468 -30892 33532 -30828
rect 33468 -30972 33532 -30908
rect 33468 -31052 33532 -30988
rect 33468 -31132 33532 -31068
rect 33468 -31212 33532 -31148
rect 33468 -31292 33532 -31228
rect 33468 -31372 33532 -31308
rect 33468 -31452 33532 -31388
rect 33468 -31532 33532 -31468
rect 33468 -31612 33532 -31548
rect 33468 -31692 33532 -31628
rect 33468 -31772 33532 -31708
rect 39080 -26812 39144 -26748
rect 39080 -26892 39144 -26828
rect 39080 -26972 39144 -26908
rect 39080 -27052 39144 -26988
rect 39080 -27132 39144 -27068
rect 39080 -27212 39144 -27148
rect 39080 -27292 39144 -27228
rect 39080 -27372 39144 -27308
rect 39080 -27452 39144 -27388
rect 39080 -27532 39144 -27468
rect 39080 -27612 39144 -27548
rect 39080 -27692 39144 -27628
rect 39080 -27772 39144 -27708
rect 39080 -27852 39144 -27788
rect 39080 -27932 39144 -27868
rect 39080 -28012 39144 -27948
rect 39080 -28092 39144 -28028
rect 39080 -28172 39144 -28108
rect 39080 -28252 39144 -28188
rect 39080 -28332 39144 -28268
rect 39080 -28412 39144 -28348
rect 39080 -28492 39144 -28428
rect 39080 -28572 39144 -28508
rect 39080 -28652 39144 -28588
rect 39080 -28732 39144 -28668
rect 39080 -28812 39144 -28748
rect 39080 -28892 39144 -28828
rect 39080 -28972 39144 -28908
rect 39080 -29052 39144 -28988
rect 39080 -29132 39144 -29068
rect 39080 -29212 39144 -29148
rect 39080 -29292 39144 -29228
rect 39080 -29372 39144 -29308
rect 39080 -29452 39144 -29388
rect 39080 -29532 39144 -29468
rect 39080 -29612 39144 -29548
rect 39080 -29692 39144 -29628
rect 39080 -29772 39144 -29708
rect 39080 -29852 39144 -29788
rect 39080 -29932 39144 -29868
rect 39080 -30012 39144 -29948
rect 39080 -30092 39144 -30028
rect 39080 -30172 39144 -30108
rect 39080 -30252 39144 -30188
rect 39080 -30332 39144 -30268
rect 39080 -30412 39144 -30348
rect 39080 -30492 39144 -30428
rect 39080 -30572 39144 -30508
rect 39080 -30652 39144 -30588
rect 39080 -30732 39144 -30668
rect 39080 -30812 39144 -30748
rect 39080 -30892 39144 -30828
rect 39080 -30972 39144 -30908
rect 39080 -31052 39144 -30988
rect 39080 -31132 39144 -31068
rect 39080 -31212 39144 -31148
rect 39080 -31292 39144 -31228
rect 39080 -31372 39144 -31308
rect 39080 -31452 39144 -31388
rect 39080 -31532 39144 -31468
rect 39080 -31612 39144 -31548
rect 39080 -31692 39144 -31628
rect 39080 -31772 39144 -31708
rect -33876 -32132 -33812 -32068
rect -33876 -32212 -33812 -32148
rect -33876 -32292 -33812 -32228
rect -33876 -32372 -33812 -32308
rect -33876 -32452 -33812 -32388
rect -33876 -32532 -33812 -32468
rect -33876 -32612 -33812 -32548
rect -33876 -32692 -33812 -32628
rect -33876 -32772 -33812 -32708
rect -33876 -32852 -33812 -32788
rect -33876 -32932 -33812 -32868
rect -33876 -33012 -33812 -32948
rect -33876 -33092 -33812 -33028
rect -33876 -33172 -33812 -33108
rect -33876 -33252 -33812 -33188
rect -33876 -33332 -33812 -33268
rect -33876 -33412 -33812 -33348
rect -33876 -33492 -33812 -33428
rect -33876 -33572 -33812 -33508
rect -33876 -33652 -33812 -33588
rect -33876 -33732 -33812 -33668
rect -33876 -33812 -33812 -33748
rect -33876 -33892 -33812 -33828
rect -33876 -33972 -33812 -33908
rect -33876 -34052 -33812 -33988
rect -33876 -34132 -33812 -34068
rect -33876 -34212 -33812 -34148
rect -33876 -34292 -33812 -34228
rect -33876 -34372 -33812 -34308
rect -33876 -34452 -33812 -34388
rect -33876 -34532 -33812 -34468
rect -33876 -34612 -33812 -34548
rect -33876 -34692 -33812 -34628
rect -33876 -34772 -33812 -34708
rect -33876 -34852 -33812 -34788
rect -33876 -34932 -33812 -34868
rect -33876 -35012 -33812 -34948
rect -33876 -35092 -33812 -35028
rect -33876 -35172 -33812 -35108
rect -33876 -35252 -33812 -35188
rect -33876 -35332 -33812 -35268
rect -33876 -35412 -33812 -35348
rect -33876 -35492 -33812 -35428
rect -33876 -35572 -33812 -35508
rect -33876 -35652 -33812 -35588
rect -33876 -35732 -33812 -35668
rect -33876 -35812 -33812 -35748
rect -33876 -35892 -33812 -35828
rect -33876 -35972 -33812 -35908
rect -33876 -36052 -33812 -35988
rect -33876 -36132 -33812 -36068
rect -33876 -36212 -33812 -36148
rect -33876 -36292 -33812 -36228
rect -33876 -36372 -33812 -36308
rect -33876 -36452 -33812 -36388
rect -33876 -36532 -33812 -36468
rect -33876 -36612 -33812 -36548
rect -33876 -36692 -33812 -36628
rect -33876 -36772 -33812 -36708
rect -33876 -36852 -33812 -36788
rect -33876 -36932 -33812 -36868
rect -33876 -37012 -33812 -36948
rect -33876 -37092 -33812 -37028
rect -28264 -32132 -28200 -32068
rect -28264 -32212 -28200 -32148
rect -28264 -32292 -28200 -32228
rect -28264 -32372 -28200 -32308
rect -28264 -32452 -28200 -32388
rect -28264 -32532 -28200 -32468
rect -28264 -32612 -28200 -32548
rect -28264 -32692 -28200 -32628
rect -28264 -32772 -28200 -32708
rect -28264 -32852 -28200 -32788
rect -28264 -32932 -28200 -32868
rect -28264 -33012 -28200 -32948
rect -28264 -33092 -28200 -33028
rect -28264 -33172 -28200 -33108
rect -28264 -33252 -28200 -33188
rect -28264 -33332 -28200 -33268
rect -28264 -33412 -28200 -33348
rect -28264 -33492 -28200 -33428
rect -28264 -33572 -28200 -33508
rect -28264 -33652 -28200 -33588
rect -28264 -33732 -28200 -33668
rect -28264 -33812 -28200 -33748
rect -28264 -33892 -28200 -33828
rect -28264 -33972 -28200 -33908
rect -28264 -34052 -28200 -33988
rect -28264 -34132 -28200 -34068
rect -28264 -34212 -28200 -34148
rect -28264 -34292 -28200 -34228
rect -28264 -34372 -28200 -34308
rect -28264 -34452 -28200 -34388
rect -28264 -34532 -28200 -34468
rect -28264 -34612 -28200 -34548
rect -28264 -34692 -28200 -34628
rect -28264 -34772 -28200 -34708
rect -28264 -34852 -28200 -34788
rect -28264 -34932 -28200 -34868
rect -28264 -35012 -28200 -34948
rect -28264 -35092 -28200 -35028
rect -28264 -35172 -28200 -35108
rect -28264 -35252 -28200 -35188
rect -28264 -35332 -28200 -35268
rect -28264 -35412 -28200 -35348
rect -28264 -35492 -28200 -35428
rect -28264 -35572 -28200 -35508
rect -28264 -35652 -28200 -35588
rect -28264 -35732 -28200 -35668
rect -28264 -35812 -28200 -35748
rect -28264 -35892 -28200 -35828
rect -28264 -35972 -28200 -35908
rect -28264 -36052 -28200 -35988
rect -28264 -36132 -28200 -36068
rect -28264 -36212 -28200 -36148
rect -28264 -36292 -28200 -36228
rect -28264 -36372 -28200 -36308
rect -28264 -36452 -28200 -36388
rect -28264 -36532 -28200 -36468
rect -28264 -36612 -28200 -36548
rect -28264 -36692 -28200 -36628
rect -28264 -36772 -28200 -36708
rect -28264 -36852 -28200 -36788
rect -28264 -36932 -28200 -36868
rect -28264 -37012 -28200 -36948
rect -28264 -37092 -28200 -37028
rect -22652 -32132 -22588 -32068
rect -22652 -32212 -22588 -32148
rect -22652 -32292 -22588 -32228
rect -22652 -32372 -22588 -32308
rect -22652 -32452 -22588 -32388
rect -22652 -32532 -22588 -32468
rect -22652 -32612 -22588 -32548
rect -22652 -32692 -22588 -32628
rect -22652 -32772 -22588 -32708
rect -22652 -32852 -22588 -32788
rect -22652 -32932 -22588 -32868
rect -22652 -33012 -22588 -32948
rect -22652 -33092 -22588 -33028
rect -22652 -33172 -22588 -33108
rect -22652 -33252 -22588 -33188
rect -22652 -33332 -22588 -33268
rect -22652 -33412 -22588 -33348
rect -22652 -33492 -22588 -33428
rect -22652 -33572 -22588 -33508
rect -22652 -33652 -22588 -33588
rect -22652 -33732 -22588 -33668
rect -22652 -33812 -22588 -33748
rect -22652 -33892 -22588 -33828
rect -22652 -33972 -22588 -33908
rect -22652 -34052 -22588 -33988
rect -22652 -34132 -22588 -34068
rect -22652 -34212 -22588 -34148
rect -22652 -34292 -22588 -34228
rect -22652 -34372 -22588 -34308
rect -22652 -34452 -22588 -34388
rect -22652 -34532 -22588 -34468
rect -22652 -34612 -22588 -34548
rect -22652 -34692 -22588 -34628
rect -22652 -34772 -22588 -34708
rect -22652 -34852 -22588 -34788
rect -22652 -34932 -22588 -34868
rect -22652 -35012 -22588 -34948
rect -22652 -35092 -22588 -35028
rect -22652 -35172 -22588 -35108
rect -22652 -35252 -22588 -35188
rect -22652 -35332 -22588 -35268
rect -22652 -35412 -22588 -35348
rect -22652 -35492 -22588 -35428
rect -22652 -35572 -22588 -35508
rect -22652 -35652 -22588 -35588
rect -22652 -35732 -22588 -35668
rect -22652 -35812 -22588 -35748
rect -22652 -35892 -22588 -35828
rect -22652 -35972 -22588 -35908
rect -22652 -36052 -22588 -35988
rect -22652 -36132 -22588 -36068
rect -22652 -36212 -22588 -36148
rect -22652 -36292 -22588 -36228
rect -22652 -36372 -22588 -36308
rect -22652 -36452 -22588 -36388
rect -22652 -36532 -22588 -36468
rect -22652 -36612 -22588 -36548
rect -22652 -36692 -22588 -36628
rect -22652 -36772 -22588 -36708
rect -22652 -36852 -22588 -36788
rect -22652 -36932 -22588 -36868
rect -22652 -37012 -22588 -36948
rect -22652 -37092 -22588 -37028
rect -17040 -32132 -16976 -32068
rect -17040 -32212 -16976 -32148
rect -17040 -32292 -16976 -32228
rect -17040 -32372 -16976 -32308
rect -17040 -32452 -16976 -32388
rect -17040 -32532 -16976 -32468
rect -17040 -32612 -16976 -32548
rect -17040 -32692 -16976 -32628
rect -17040 -32772 -16976 -32708
rect -17040 -32852 -16976 -32788
rect -17040 -32932 -16976 -32868
rect -17040 -33012 -16976 -32948
rect -17040 -33092 -16976 -33028
rect -17040 -33172 -16976 -33108
rect -17040 -33252 -16976 -33188
rect -17040 -33332 -16976 -33268
rect -17040 -33412 -16976 -33348
rect -17040 -33492 -16976 -33428
rect -17040 -33572 -16976 -33508
rect -17040 -33652 -16976 -33588
rect -17040 -33732 -16976 -33668
rect -17040 -33812 -16976 -33748
rect -17040 -33892 -16976 -33828
rect -17040 -33972 -16976 -33908
rect -17040 -34052 -16976 -33988
rect -17040 -34132 -16976 -34068
rect -17040 -34212 -16976 -34148
rect -17040 -34292 -16976 -34228
rect -17040 -34372 -16976 -34308
rect -17040 -34452 -16976 -34388
rect -17040 -34532 -16976 -34468
rect -17040 -34612 -16976 -34548
rect -17040 -34692 -16976 -34628
rect -17040 -34772 -16976 -34708
rect -17040 -34852 -16976 -34788
rect -17040 -34932 -16976 -34868
rect -17040 -35012 -16976 -34948
rect -17040 -35092 -16976 -35028
rect -17040 -35172 -16976 -35108
rect -17040 -35252 -16976 -35188
rect -17040 -35332 -16976 -35268
rect -17040 -35412 -16976 -35348
rect -17040 -35492 -16976 -35428
rect -17040 -35572 -16976 -35508
rect -17040 -35652 -16976 -35588
rect -17040 -35732 -16976 -35668
rect -17040 -35812 -16976 -35748
rect -17040 -35892 -16976 -35828
rect -17040 -35972 -16976 -35908
rect -17040 -36052 -16976 -35988
rect -17040 -36132 -16976 -36068
rect -17040 -36212 -16976 -36148
rect -17040 -36292 -16976 -36228
rect -17040 -36372 -16976 -36308
rect -17040 -36452 -16976 -36388
rect -17040 -36532 -16976 -36468
rect -17040 -36612 -16976 -36548
rect -17040 -36692 -16976 -36628
rect -17040 -36772 -16976 -36708
rect -17040 -36852 -16976 -36788
rect -17040 -36932 -16976 -36868
rect -17040 -37012 -16976 -36948
rect -17040 -37092 -16976 -37028
rect -11428 -32132 -11364 -32068
rect -11428 -32212 -11364 -32148
rect -11428 -32292 -11364 -32228
rect -11428 -32372 -11364 -32308
rect -11428 -32452 -11364 -32388
rect -11428 -32532 -11364 -32468
rect -11428 -32612 -11364 -32548
rect -11428 -32692 -11364 -32628
rect -11428 -32772 -11364 -32708
rect -11428 -32852 -11364 -32788
rect -11428 -32932 -11364 -32868
rect -11428 -33012 -11364 -32948
rect -11428 -33092 -11364 -33028
rect -11428 -33172 -11364 -33108
rect -11428 -33252 -11364 -33188
rect -11428 -33332 -11364 -33268
rect -11428 -33412 -11364 -33348
rect -11428 -33492 -11364 -33428
rect -11428 -33572 -11364 -33508
rect -11428 -33652 -11364 -33588
rect -11428 -33732 -11364 -33668
rect -11428 -33812 -11364 -33748
rect -11428 -33892 -11364 -33828
rect -11428 -33972 -11364 -33908
rect -11428 -34052 -11364 -33988
rect -11428 -34132 -11364 -34068
rect -11428 -34212 -11364 -34148
rect -11428 -34292 -11364 -34228
rect -11428 -34372 -11364 -34308
rect -11428 -34452 -11364 -34388
rect -11428 -34532 -11364 -34468
rect -11428 -34612 -11364 -34548
rect -11428 -34692 -11364 -34628
rect -11428 -34772 -11364 -34708
rect -11428 -34852 -11364 -34788
rect -11428 -34932 -11364 -34868
rect -11428 -35012 -11364 -34948
rect -11428 -35092 -11364 -35028
rect -11428 -35172 -11364 -35108
rect -11428 -35252 -11364 -35188
rect -11428 -35332 -11364 -35268
rect -11428 -35412 -11364 -35348
rect -11428 -35492 -11364 -35428
rect -11428 -35572 -11364 -35508
rect -11428 -35652 -11364 -35588
rect -11428 -35732 -11364 -35668
rect -11428 -35812 -11364 -35748
rect -11428 -35892 -11364 -35828
rect -11428 -35972 -11364 -35908
rect -11428 -36052 -11364 -35988
rect -11428 -36132 -11364 -36068
rect -11428 -36212 -11364 -36148
rect -11428 -36292 -11364 -36228
rect -11428 -36372 -11364 -36308
rect -11428 -36452 -11364 -36388
rect -11428 -36532 -11364 -36468
rect -11428 -36612 -11364 -36548
rect -11428 -36692 -11364 -36628
rect -11428 -36772 -11364 -36708
rect -11428 -36852 -11364 -36788
rect -11428 -36932 -11364 -36868
rect -11428 -37012 -11364 -36948
rect -11428 -37092 -11364 -37028
rect -5816 -32132 -5752 -32068
rect -5816 -32212 -5752 -32148
rect -5816 -32292 -5752 -32228
rect -5816 -32372 -5752 -32308
rect -5816 -32452 -5752 -32388
rect -5816 -32532 -5752 -32468
rect -5816 -32612 -5752 -32548
rect -5816 -32692 -5752 -32628
rect -5816 -32772 -5752 -32708
rect -5816 -32852 -5752 -32788
rect -5816 -32932 -5752 -32868
rect -5816 -33012 -5752 -32948
rect -5816 -33092 -5752 -33028
rect -5816 -33172 -5752 -33108
rect -5816 -33252 -5752 -33188
rect -5816 -33332 -5752 -33268
rect -5816 -33412 -5752 -33348
rect -5816 -33492 -5752 -33428
rect -5816 -33572 -5752 -33508
rect -5816 -33652 -5752 -33588
rect -5816 -33732 -5752 -33668
rect -5816 -33812 -5752 -33748
rect -5816 -33892 -5752 -33828
rect -5816 -33972 -5752 -33908
rect -5816 -34052 -5752 -33988
rect -5816 -34132 -5752 -34068
rect -5816 -34212 -5752 -34148
rect -5816 -34292 -5752 -34228
rect -5816 -34372 -5752 -34308
rect -5816 -34452 -5752 -34388
rect -5816 -34532 -5752 -34468
rect -5816 -34612 -5752 -34548
rect -5816 -34692 -5752 -34628
rect -5816 -34772 -5752 -34708
rect -5816 -34852 -5752 -34788
rect -5816 -34932 -5752 -34868
rect -5816 -35012 -5752 -34948
rect -5816 -35092 -5752 -35028
rect -5816 -35172 -5752 -35108
rect -5816 -35252 -5752 -35188
rect -5816 -35332 -5752 -35268
rect -5816 -35412 -5752 -35348
rect -5816 -35492 -5752 -35428
rect -5816 -35572 -5752 -35508
rect -5816 -35652 -5752 -35588
rect -5816 -35732 -5752 -35668
rect -5816 -35812 -5752 -35748
rect -5816 -35892 -5752 -35828
rect -5816 -35972 -5752 -35908
rect -5816 -36052 -5752 -35988
rect -5816 -36132 -5752 -36068
rect -5816 -36212 -5752 -36148
rect -5816 -36292 -5752 -36228
rect -5816 -36372 -5752 -36308
rect -5816 -36452 -5752 -36388
rect -5816 -36532 -5752 -36468
rect -5816 -36612 -5752 -36548
rect -5816 -36692 -5752 -36628
rect -5816 -36772 -5752 -36708
rect -5816 -36852 -5752 -36788
rect -5816 -36932 -5752 -36868
rect -5816 -37012 -5752 -36948
rect -5816 -37092 -5752 -37028
rect -204 -32132 -140 -32068
rect -204 -32212 -140 -32148
rect -204 -32292 -140 -32228
rect -204 -32372 -140 -32308
rect -204 -32452 -140 -32388
rect -204 -32532 -140 -32468
rect -204 -32612 -140 -32548
rect -204 -32692 -140 -32628
rect -204 -32772 -140 -32708
rect -204 -32852 -140 -32788
rect -204 -32932 -140 -32868
rect -204 -33012 -140 -32948
rect -204 -33092 -140 -33028
rect -204 -33172 -140 -33108
rect -204 -33252 -140 -33188
rect -204 -33332 -140 -33268
rect -204 -33412 -140 -33348
rect -204 -33492 -140 -33428
rect -204 -33572 -140 -33508
rect -204 -33652 -140 -33588
rect -204 -33732 -140 -33668
rect -204 -33812 -140 -33748
rect -204 -33892 -140 -33828
rect -204 -33972 -140 -33908
rect -204 -34052 -140 -33988
rect -204 -34132 -140 -34068
rect -204 -34212 -140 -34148
rect -204 -34292 -140 -34228
rect -204 -34372 -140 -34308
rect -204 -34452 -140 -34388
rect -204 -34532 -140 -34468
rect -204 -34612 -140 -34548
rect -204 -34692 -140 -34628
rect -204 -34772 -140 -34708
rect -204 -34852 -140 -34788
rect -204 -34932 -140 -34868
rect -204 -35012 -140 -34948
rect -204 -35092 -140 -35028
rect -204 -35172 -140 -35108
rect -204 -35252 -140 -35188
rect -204 -35332 -140 -35268
rect -204 -35412 -140 -35348
rect -204 -35492 -140 -35428
rect -204 -35572 -140 -35508
rect -204 -35652 -140 -35588
rect -204 -35732 -140 -35668
rect -204 -35812 -140 -35748
rect -204 -35892 -140 -35828
rect -204 -35972 -140 -35908
rect -204 -36052 -140 -35988
rect -204 -36132 -140 -36068
rect -204 -36212 -140 -36148
rect -204 -36292 -140 -36228
rect -204 -36372 -140 -36308
rect -204 -36452 -140 -36388
rect -204 -36532 -140 -36468
rect -204 -36612 -140 -36548
rect -204 -36692 -140 -36628
rect -204 -36772 -140 -36708
rect -204 -36852 -140 -36788
rect -204 -36932 -140 -36868
rect -204 -37012 -140 -36948
rect -204 -37092 -140 -37028
rect 5408 -32132 5472 -32068
rect 5408 -32212 5472 -32148
rect 5408 -32292 5472 -32228
rect 5408 -32372 5472 -32308
rect 5408 -32452 5472 -32388
rect 5408 -32532 5472 -32468
rect 5408 -32612 5472 -32548
rect 5408 -32692 5472 -32628
rect 5408 -32772 5472 -32708
rect 5408 -32852 5472 -32788
rect 5408 -32932 5472 -32868
rect 5408 -33012 5472 -32948
rect 5408 -33092 5472 -33028
rect 5408 -33172 5472 -33108
rect 5408 -33252 5472 -33188
rect 5408 -33332 5472 -33268
rect 5408 -33412 5472 -33348
rect 5408 -33492 5472 -33428
rect 5408 -33572 5472 -33508
rect 5408 -33652 5472 -33588
rect 5408 -33732 5472 -33668
rect 5408 -33812 5472 -33748
rect 5408 -33892 5472 -33828
rect 5408 -33972 5472 -33908
rect 5408 -34052 5472 -33988
rect 5408 -34132 5472 -34068
rect 5408 -34212 5472 -34148
rect 5408 -34292 5472 -34228
rect 5408 -34372 5472 -34308
rect 5408 -34452 5472 -34388
rect 5408 -34532 5472 -34468
rect 5408 -34612 5472 -34548
rect 5408 -34692 5472 -34628
rect 5408 -34772 5472 -34708
rect 5408 -34852 5472 -34788
rect 5408 -34932 5472 -34868
rect 5408 -35012 5472 -34948
rect 5408 -35092 5472 -35028
rect 5408 -35172 5472 -35108
rect 5408 -35252 5472 -35188
rect 5408 -35332 5472 -35268
rect 5408 -35412 5472 -35348
rect 5408 -35492 5472 -35428
rect 5408 -35572 5472 -35508
rect 5408 -35652 5472 -35588
rect 5408 -35732 5472 -35668
rect 5408 -35812 5472 -35748
rect 5408 -35892 5472 -35828
rect 5408 -35972 5472 -35908
rect 5408 -36052 5472 -35988
rect 5408 -36132 5472 -36068
rect 5408 -36212 5472 -36148
rect 5408 -36292 5472 -36228
rect 5408 -36372 5472 -36308
rect 5408 -36452 5472 -36388
rect 5408 -36532 5472 -36468
rect 5408 -36612 5472 -36548
rect 5408 -36692 5472 -36628
rect 5408 -36772 5472 -36708
rect 5408 -36852 5472 -36788
rect 5408 -36932 5472 -36868
rect 5408 -37012 5472 -36948
rect 5408 -37092 5472 -37028
rect 11020 -32132 11084 -32068
rect 11020 -32212 11084 -32148
rect 11020 -32292 11084 -32228
rect 11020 -32372 11084 -32308
rect 11020 -32452 11084 -32388
rect 11020 -32532 11084 -32468
rect 11020 -32612 11084 -32548
rect 11020 -32692 11084 -32628
rect 11020 -32772 11084 -32708
rect 11020 -32852 11084 -32788
rect 11020 -32932 11084 -32868
rect 11020 -33012 11084 -32948
rect 11020 -33092 11084 -33028
rect 11020 -33172 11084 -33108
rect 11020 -33252 11084 -33188
rect 11020 -33332 11084 -33268
rect 11020 -33412 11084 -33348
rect 11020 -33492 11084 -33428
rect 11020 -33572 11084 -33508
rect 11020 -33652 11084 -33588
rect 11020 -33732 11084 -33668
rect 11020 -33812 11084 -33748
rect 11020 -33892 11084 -33828
rect 11020 -33972 11084 -33908
rect 11020 -34052 11084 -33988
rect 11020 -34132 11084 -34068
rect 11020 -34212 11084 -34148
rect 11020 -34292 11084 -34228
rect 11020 -34372 11084 -34308
rect 11020 -34452 11084 -34388
rect 11020 -34532 11084 -34468
rect 11020 -34612 11084 -34548
rect 11020 -34692 11084 -34628
rect 11020 -34772 11084 -34708
rect 11020 -34852 11084 -34788
rect 11020 -34932 11084 -34868
rect 11020 -35012 11084 -34948
rect 11020 -35092 11084 -35028
rect 11020 -35172 11084 -35108
rect 11020 -35252 11084 -35188
rect 11020 -35332 11084 -35268
rect 11020 -35412 11084 -35348
rect 11020 -35492 11084 -35428
rect 11020 -35572 11084 -35508
rect 11020 -35652 11084 -35588
rect 11020 -35732 11084 -35668
rect 11020 -35812 11084 -35748
rect 11020 -35892 11084 -35828
rect 11020 -35972 11084 -35908
rect 11020 -36052 11084 -35988
rect 11020 -36132 11084 -36068
rect 11020 -36212 11084 -36148
rect 11020 -36292 11084 -36228
rect 11020 -36372 11084 -36308
rect 11020 -36452 11084 -36388
rect 11020 -36532 11084 -36468
rect 11020 -36612 11084 -36548
rect 11020 -36692 11084 -36628
rect 11020 -36772 11084 -36708
rect 11020 -36852 11084 -36788
rect 11020 -36932 11084 -36868
rect 11020 -37012 11084 -36948
rect 11020 -37092 11084 -37028
rect 16632 -32132 16696 -32068
rect 16632 -32212 16696 -32148
rect 16632 -32292 16696 -32228
rect 16632 -32372 16696 -32308
rect 16632 -32452 16696 -32388
rect 16632 -32532 16696 -32468
rect 16632 -32612 16696 -32548
rect 16632 -32692 16696 -32628
rect 16632 -32772 16696 -32708
rect 16632 -32852 16696 -32788
rect 16632 -32932 16696 -32868
rect 16632 -33012 16696 -32948
rect 16632 -33092 16696 -33028
rect 16632 -33172 16696 -33108
rect 16632 -33252 16696 -33188
rect 16632 -33332 16696 -33268
rect 16632 -33412 16696 -33348
rect 16632 -33492 16696 -33428
rect 16632 -33572 16696 -33508
rect 16632 -33652 16696 -33588
rect 16632 -33732 16696 -33668
rect 16632 -33812 16696 -33748
rect 16632 -33892 16696 -33828
rect 16632 -33972 16696 -33908
rect 16632 -34052 16696 -33988
rect 16632 -34132 16696 -34068
rect 16632 -34212 16696 -34148
rect 16632 -34292 16696 -34228
rect 16632 -34372 16696 -34308
rect 16632 -34452 16696 -34388
rect 16632 -34532 16696 -34468
rect 16632 -34612 16696 -34548
rect 16632 -34692 16696 -34628
rect 16632 -34772 16696 -34708
rect 16632 -34852 16696 -34788
rect 16632 -34932 16696 -34868
rect 16632 -35012 16696 -34948
rect 16632 -35092 16696 -35028
rect 16632 -35172 16696 -35108
rect 16632 -35252 16696 -35188
rect 16632 -35332 16696 -35268
rect 16632 -35412 16696 -35348
rect 16632 -35492 16696 -35428
rect 16632 -35572 16696 -35508
rect 16632 -35652 16696 -35588
rect 16632 -35732 16696 -35668
rect 16632 -35812 16696 -35748
rect 16632 -35892 16696 -35828
rect 16632 -35972 16696 -35908
rect 16632 -36052 16696 -35988
rect 16632 -36132 16696 -36068
rect 16632 -36212 16696 -36148
rect 16632 -36292 16696 -36228
rect 16632 -36372 16696 -36308
rect 16632 -36452 16696 -36388
rect 16632 -36532 16696 -36468
rect 16632 -36612 16696 -36548
rect 16632 -36692 16696 -36628
rect 16632 -36772 16696 -36708
rect 16632 -36852 16696 -36788
rect 16632 -36932 16696 -36868
rect 16632 -37012 16696 -36948
rect 16632 -37092 16696 -37028
rect 22244 -32132 22308 -32068
rect 22244 -32212 22308 -32148
rect 22244 -32292 22308 -32228
rect 22244 -32372 22308 -32308
rect 22244 -32452 22308 -32388
rect 22244 -32532 22308 -32468
rect 22244 -32612 22308 -32548
rect 22244 -32692 22308 -32628
rect 22244 -32772 22308 -32708
rect 22244 -32852 22308 -32788
rect 22244 -32932 22308 -32868
rect 22244 -33012 22308 -32948
rect 22244 -33092 22308 -33028
rect 22244 -33172 22308 -33108
rect 22244 -33252 22308 -33188
rect 22244 -33332 22308 -33268
rect 22244 -33412 22308 -33348
rect 22244 -33492 22308 -33428
rect 22244 -33572 22308 -33508
rect 22244 -33652 22308 -33588
rect 22244 -33732 22308 -33668
rect 22244 -33812 22308 -33748
rect 22244 -33892 22308 -33828
rect 22244 -33972 22308 -33908
rect 22244 -34052 22308 -33988
rect 22244 -34132 22308 -34068
rect 22244 -34212 22308 -34148
rect 22244 -34292 22308 -34228
rect 22244 -34372 22308 -34308
rect 22244 -34452 22308 -34388
rect 22244 -34532 22308 -34468
rect 22244 -34612 22308 -34548
rect 22244 -34692 22308 -34628
rect 22244 -34772 22308 -34708
rect 22244 -34852 22308 -34788
rect 22244 -34932 22308 -34868
rect 22244 -35012 22308 -34948
rect 22244 -35092 22308 -35028
rect 22244 -35172 22308 -35108
rect 22244 -35252 22308 -35188
rect 22244 -35332 22308 -35268
rect 22244 -35412 22308 -35348
rect 22244 -35492 22308 -35428
rect 22244 -35572 22308 -35508
rect 22244 -35652 22308 -35588
rect 22244 -35732 22308 -35668
rect 22244 -35812 22308 -35748
rect 22244 -35892 22308 -35828
rect 22244 -35972 22308 -35908
rect 22244 -36052 22308 -35988
rect 22244 -36132 22308 -36068
rect 22244 -36212 22308 -36148
rect 22244 -36292 22308 -36228
rect 22244 -36372 22308 -36308
rect 22244 -36452 22308 -36388
rect 22244 -36532 22308 -36468
rect 22244 -36612 22308 -36548
rect 22244 -36692 22308 -36628
rect 22244 -36772 22308 -36708
rect 22244 -36852 22308 -36788
rect 22244 -36932 22308 -36868
rect 22244 -37012 22308 -36948
rect 22244 -37092 22308 -37028
rect 27856 -32132 27920 -32068
rect 27856 -32212 27920 -32148
rect 27856 -32292 27920 -32228
rect 27856 -32372 27920 -32308
rect 27856 -32452 27920 -32388
rect 27856 -32532 27920 -32468
rect 27856 -32612 27920 -32548
rect 27856 -32692 27920 -32628
rect 27856 -32772 27920 -32708
rect 27856 -32852 27920 -32788
rect 27856 -32932 27920 -32868
rect 27856 -33012 27920 -32948
rect 27856 -33092 27920 -33028
rect 27856 -33172 27920 -33108
rect 27856 -33252 27920 -33188
rect 27856 -33332 27920 -33268
rect 27856 -33412 27920 -33348
rect 27856 -33492 27920 -33428
rect 27856 -33572 27920 -33508
rect 27856 -33652 27920 -33588
rect 27856 -33732 27920 -33668
rect 27856 -33812 27920 -33748
rect 27856 -33892 27920 -33828
rect 27856 -33972 27920 -33908
rect 27856 -34052 27920 -33988
rect 27856 -34132 27920 -34068
rect 27856 -34212 27920 -34148
rect 27856 -34292 27920 -34228
rect 27856 -34372 27920 -34308
rect 27856 -34452 27920 -34388
rect 27856 -34532 27920 -34468
rect 27856 -34612 27920 -34548
rect 27856 -34692 27920 -34628
rect 27856 -34772 27920 -34708
rect 27856 -34852 27920 -34788
rect 27856 -34932 27920 -34868
rect 27856 -35012 27920 -34948
rect 27856 -35092 27920 -35028
rect 27856 -35172 27920 -35108
rect 27856 -35252 27920 -35188
rect 27856 -35332 27920 -35268
rect 27856 -35412 27920 -35348
rect 27856 -35492 27920 -35428
rect 27856 -35572 27920 -35508
rect 27856 -35652 27920 -35588
rect 27856 -35732 27920 -35668
rect 27856 -35812 27920 -35748
rect 27856 -35892 27920 -35828
rect 27856 -35972 27920 -35908
rect 27856 -36052 27920 -35988
rect 27856 -36132 27920 -36068
rect 27856 -36212 27920 -36148
rect 27856 -36292 27920 -36228
rect 27856 -36372 27920 -36308
rect 27856 -36452 27920 -36388
rect 27856 -36532 27920 -36468
rect 27856 -36612 27920 -36548
rect 27856 -36692 27920 -36628
rect 27856 -36772 27920 -36708
rect 27856 -36852 27920 -36788
rect 27856 -36932 27920 -36868
rect 27856 -37012 27920 -36948
rect 27856 -37092 27920 -37028
rect 33468 -32132 33532 -32068
rect 33468 -32212 33532 -32148
rect 33468 -32292 33532 -32228
rect 33468 -32372 33532 -32308
rect 33468 -32452 33532 -32388
rect 33468 -32532 33532 -32468
rect 33468 -32612 33532 -32548
rect 33468 -32692 33532 -32628
rect 33468 -32772 33532 -32708
rect 33468 -32852 33532 -32788
rect 33468 -32932 33532 -32868
rect 33468 -33012 33532 -32948
rect 33468 -33092 33532 -33028
rect 33468 -33172 33532 -33108
rect 33468 -33252 33532 -33188
rect 33468 -33332 33532 -33268
rect 33468 -33412 33532 -33348
rect 33468 -33492 33532 -33428
rect 33468 -33572 33532 -33508
rect 33468 -33652 33532 -33588
rect 33468 -33732 33532 -33668
rect 33468 -33812 33532 -33748
rect 33468 -33892 33532 -33828
rect 33468 -33972 33532 -33908
rect 33468 -34052 33532 -33988
rect 33468 -34132 33532 -34068
rect 33468 -34212 33532 -34148
rect 33468 -34292 33532 -34228
rect 33468 -34372 33532 -34308
rect 33468 -34452 33532 -34388
rect 33468 -34532 33532 -34468
rect 33468 -34612 33532 -34548
rect 33468 -34692 33532 -34628
rect 33468 -34772 33532 -34708
rect 33468 -34852 33532 -34788
rect 33468 -34932 33532 -34868
rect 33468 -35012 33532 -34948
rect 33468 -35092 33532 -35028
rect 33468 -35172 33532 -35108
rect 33468 -35252 33532 -35188
rect 33468 -35332 33532 -35268
rect 33468 -35412 33532 -35348
rect 33468 -35492 33532 -35428
rect 33468 -35572 33532 -35508
rect 33468 -35652 33532 -35588
rect 33468 -35732 33532 -35668
rect 33468 -35812 33532 -35748
rect 33468 -35892 33532 -35828
rect 33468 -35972 33532 -35908
rect 33468 -36052 33532 -35988
rect 33468 -36132 33532 -36068
rect 33468 -36212 33532 -36148
rect 33468 -36292 33532 -36228
rect 33468 -36372 33532 -36308
rect 33468 -36452 33532 -36388
rect 33468 -36532 33532 -36468
rect 33468 -36612 33532 -36548
rect 33468 -36692 33532 -36628
rect 33468 -36772 33532 -36708
rect 33468 -36852 33532 -36788
rect 33468 -36932 33532 -36868
rect 33468 -37012 33532 -36948
rect 33468 -37092 33532 -37028
rect 39080 -32132 39144 -32068
rect 39080 -32212 39144 -32148
rect 39080 -32292 39144 -32228
rect 39080 -32372 39144 -32308
rect 39080 -32452 39144 -32388
rect 39080 -32532 39144 -32468
rect 39080 -32612 39144 -32548
rect 39080 -32692 39144 -32628
rect 39080 -32772 39144 -32708
rect 39080 -32852 39144 -32788
rect 39080 -32932 39144 -32868
rect 39080 -33012 39144 -32948
rect 39080 -33092 39144 -33028
rect 39080 -33172 39144 -33108
rect 39080 -33252 39144 -33188
rect 39080 -33332 39144 -33268
rect 39080 -33412 39144 -33348
rect 39080 -33492 39144 -33428
rect 39080 -33572 39144 -33508
rect 39080 -33652 39144 -33588
rect 39080 -33732 39144 -33668
rect 39080 -33812 39144 -33748
rect 39080 -33892 39144 -33828
rect 39080 -33972 39144 -33908
rect 39080 -34052 39144 -33988
rect 39080 -34132 39144 -34068
rect 39080 -34212 39144 -34148
rect 39080 -34292 39144 -34228
rect 39080 -34372 39144 -34308
rect 39080 -34452 39144 -34388
rect 39080 -34532 39144 -34468
rect 39080 -34612 39144 -34548
rect 39080 -34692 39144 -34628
rect 39080 -34772 39144 -34708
rect 39080 -34852 39144 -34788
rect 39080 -34932 39144 -34868
rect 39080 -35012 39144 -34948
rect 39080 -35092 39144 -35028
rect 39080 -35172 39144 -35108
rect 39080 -35252 39144 -35188
rect 39080 -35332 39144 -35268
rect 39080 -35412 39144 -35348
rect 39080 -35492 39144 -35428
rect 39080 -35572 39144 -35508
rect 39080 -35652 39144 -35588
rect 39080 -35732 39144 -35668
rect 39080 -35812 39144 -35748
rect 39080 -35892 39144 -35828
rect 39080 -35972 39144 -35908
rect 39080 -36052 39144 -35988
rect 39080 -36132 39144 -36068
rect 39080 -36212 39144 -36148
rect 39080 -36292 39144 -36228
rect 39080 -36372 39144 -36308
rect 39080 -36452 39144 -36388
rect 39080 -36532 39144 -36468
rect 39080 -36612 39144 -36548
rect 39080 -36692 39144 -36628
rect 39080 -36772 39144 -36708
rect 39080 -36852 39144 -36788
rect 39080 -36932 39144 -36868
rect 39080 -37012 39144 -36948
rect 39080 -37092 39144 -37028
<< mimcap >>
rect -39124 37012 -34124 37080
rect -39124 32148 -39056 37012
rect -34192 32148 -34124 37012
rect -39124 32080 -34124 32148
rect -33512 37012 -28512 37080
rect -33512 32148 -33444 37012
rect -28580 32148 -28512 37012
rect -33512 32080 -28512 32148
rect -27900 37012 -22900 37080
rect -27900 32148 -27832 37012
rect -22968 32148 -22900 37012
rect -27900 32080 -22900 32148
rect -22288 37012 -17288 37080
rect -22288 32148 -22220 37012
rect -17356 32148 -17288 37012
rect -22288 32080 -17288 32148
rect -16676 37012 -11676 37080
rect -16676 32148 -16608 37012
rect -11744 32148 -11676 37012
rect -16676 32080 -11676 32148
rect -11064 37012 -6064 37080
rect -11064 32148 -10996 37012
rect -6132 32148 -6064 37012
rect -11064 32080 -6064 32148
rect -5452 37012 -452 37080
rect -5452 32148 -5384 37012
rect -520 32148 -452 37012
rect -5452 32080 -452 32148
rect 160 37012 5160 37080
rect 160 32148 228 37012
rect 5092 32148 5160 37012
rect 160 32080 5160 32148
rect 5772 37012 10772 37080
rect 5772 32148 5840 37012
rect 10704 32148 10772 37012
rect 5772 32080 10772 32148
rect 11384 37012 16384 37080
rect 11384 32148 11452 37012
rect 16316 32148 16384 37012
rect 11384 32080 16384 32148
rect 16996 37012 21996 37080
rect 16996 32148 17064 37012
rect 21928 32148 21996 37012
rect 16996 32080 21996 32148
rect 22608 37012 27608 37080
rect 22608 32148 22676 37012
rect 27540 32148 27608 37012
rect 22608 32080 27608 32148
rect 28220 37012 33220 37080
rect 28220 32148 28288 37012
rect 33152 32148 33220 37012
rect 28220 32080 33220 32148
rect 33832 37012 38832 37080
rect 33832 32148 33900 37012
rect 38764 32148 38832 37012
rect 33832 32080 38832 32148
rect -39124 31692 -34124 31760
rect -39124 26828 -39056 31692
rect -34192 26828 -34124 31692
rect -39124 26760 -34124 26828
rect -33512 31692 -28512 31760
rect -33512 26828 -33444 31692
rect -28580 26828 -28512 31692
rect -33512 26760 -28512 26828
rect -27900 31692 -22900 31760
rect -27900 26828 -27832 31692
rect -22968 26828 -22900 31692
rect -27900 26760 -22900 26828
rect -22288 31692 -17288 31760
rect -22288 26828 -22220 31692
rect -17356 26828 -17288 31692
rect -22288 26760 -17288 26828
rect -16676 31692 -11676 31760
rect -16676 26828 -16608 31692
rect -11744 26828 -11676 31692
rect -16676 26760 -11676 26828
rect -11064 31692 -6064 31760
rect -11064 26828 -10996 31692
rect -6132 26828 -6064 31692
rect -11064 26760 -6064 26828
rect -5452 31692 -452 31760
rect -5452 26828 -5384 31692
rect -520 26828 -452 31692
rect -5452 26760 -452 26828
rect 160 31692 5160 31760
rect 160 26828 228 31692
rect 5092 26828 5160 31692
rect 160 26760 5160 26828
rect 5772 31692 10772 31760
rect 5772 26828 5840 31692
rect 10704 26828 10772 31692
rect 5772 26760 10772 26828
rect 11384 31692 16384 31760
rect 11384 26828 11452 31692
rect 16316 26828 16384 31692
rect 11384 26760 16384 26828
rect 16996 31692 21996 31760
rect 16996 26828 17064 31692
rect 21928 26828 21996 31692
rect 16996 26760 21996 26828
rect 22608 31692 27608 31760
rect 22608 26828 22676 31692
rect 27540 26828 27608 31692
rect 22608 26760 27608 26828
rect 28220 31692 33220 31760
rect 28220 26828 28288 31692
rect 33152 26828 33220 31692
rect 28220 26760 33220 26828
rect 33832 31692 38832 31760
rect 33832 26828 33900 31692
rect 38764 26828 38832 31692
rect 33832 26760 38832 26828
rect -39124 26372 -34124 26440
rect -39124 21508 -39056 26372
rect -34192 21508 -34124 26372
rect -39124 21440 -34124 21508
rect -33512 26372 -28512 26440
rect -33512 21508 -33444 26372
rect -28580 21508 -28512 26372
rect -33512 21440 -28512 21508
rect -27900 26372 -22900 26440
rect -27900 21508 -27832 26372
rect -22968 21508 -22900 26372
rect -27900 21440 -22900 21508
rect -22288 26372 -17288 26440
rect -22288 21508 -22220 26372
rect -17356 21508 -17288 26372
rect -22288 21440 -17288 21508
rect -16676 26372 -11676 26440
rect -16676 21508 -16608 26372
rect -11744 21508 -11676 26372
rect -16676 21440 -11676 21508
rect -11064 26372 -6064 26440
rect -11064 21508 -10996 26372
rect -6132 21508 -6064 26372
rect -11064 21440 -6064 21508
rect -5452 26372 -452 26440
rect -5452 21508 -5384 26372
rect -520 21508 -452 26372
rect -5452 21440 -452 21508
rect 160 26372 5160 26440
rect 160 21508 228 26372
rect 5092 21508 5160 26372
rect 160 21440 5160 21508
rect 5772 26372 10772 26440
rect 5772 21508 5840 26372
rect 10704 21508 10772 26372
rect 5772 21440 10772 21508
rect 11384 26372 16384 26440
rect 11384 21508 11452 26372
rect 16316 21508 16384 26372
rect 11384 21440 16384 21508
rect 16996 26372 21996 26440
rect 16996 21508 17064 26372
rect 21928 21508 21996 26372
rect 16996 21440 21996 21508
rect 22608 26372 27608 26440
rect 22608 21508 22676 26372
rect 27540 21508 27608 26372
rect 22608 21440 27608 21508
rect 28220 26372 33220 26440
rect 28220 21508 28288 26372
rect 33152 21508 33220 26372
rect 28220 21440 33220 21508
rect 33832 26372 38832 26440
rect 33832 21508 33900 26372
rect 38764 21508 38832 26372
rect 33832 21440 38832 21508
rect -39124 21052 -34124 21120
rect -39124 16188 -39056 21052
rect -34192 16188 -34124 21052
rect -39124 16120 -34124 16188
rect -33512 21052 -28512 21120
rect -33512 16188 -33444 21052
rect -28580 16188 -28512 21052
rect -33512 16120 -28512 16188
rect -27900 21052 -22900 21120
rect -27900 16188 -27832 21052
rect -22968 16188 -22900 21052
rect -27900 16120 -22900 16188
rect -22288 21052 -17288 21120
rect -22288 16188 -22220 21052
rect -17356 16188 -17288 21052
rect -22288 16120 -17288 16188
rect -16676 21052 -11676 21120
rect -16676 16188 -16608 21052
rect -11744 16188 -11676 21052
rect -16676 16120 -11676 16188
rect -11064 21052 -6064 21120
rect -11064 16188 -10996 21052
rect -6132 16188 -6064 21052
rect -11064 16120 -6064 16188
rect -5452 21052 -452 21120
rect -5452 16188 -5384 21052
rect -520 16188 -452 21052
rect -5452 16120 -452 16188
rect 160 21052 5160 21120
rect 160 16188 228 21052
rect 5092 16188 5160 21052
rect 160 16120 5160 16188
rect 5772 21052 10772 21120
rect 5772 16188 5840 21052
rect 10704 16188 10772 21052
rect 5772 16120 10772 16188
rect 11384 21052 16384 21120
rect 11384 16188 11452 21052
rect 16316 16188 16384 21052
rect 11384 16120 16384 16188
rect 16996 21052 21996 21120
rect 16996 16188 17064 21052
rect 21928 16188 21996 21052
rect 16996 16120 21996 16188
rect 22608 21052 27608 21120
rect 22608 16188 22676 21052
rect 27540 16188 27608 21052
rect 22608 16120 27608 16188
rect 28220 21052 33220 21120
rect 28220 16188 28288 21052
rect 33152 16188 33220 21052
rect 28220 16120 33220 16188
rect 33832 21052 38832 21120
rect 33832 16188 33900 21052
rect 38764 16188 38832 21052
rect 33832 16120 38832 16188
rect -39124 15732 -34124 15800
rect -39124 10868 -39056 15732
rect -34192 10868 -34124 15732
rect -39124 10800 -34124 10868
rect -33512 15732 -28512 15800
rect -33512 10868 -33444 15732
rect -28580 10868 -28512 15732
rect -33512 10800 -28512 10868
rect -27900 15732 -22900 15800
rect -27900 10868 -27832 15732
rect -22968 10868 -22900 15732
rect -27900 10800 -22900 10868
rect -22288 15732 -17288 15800
rect -22288 10868 -22220 15732
rect -17356 10868 -17288 15732
rect -22288 10800 -17288 10868
rect -16676 15732 -11676 15800
rect -16676 10868 -16608 15732
rect -11744 10868 -11676 15732
rect -16676 10800 -11676 10868
rect -11064 15732 -6064 15800
rect -11064 10868 -10996 15732
rect -6132 10868 -6064 15732
rect -11064 10800 -6064 10868
rect -5452 15732 -452 15800
rect -5452 10868 -5384 15732
rect -520 10868 -452 15732
rect -5452 10800 -452 10868
rect 160 15732 5160 15800
rect 160 10868 228 15732
rect 5092 10868 5160 15732
rect 160 10800 5160 10868
rect 5772 15732 10772 15800
rect 5772 10868 5840 15732
rect 10704 10868 10772 15732
rect 5772 10800 10772 10868
rect 11384 15732 16384 15800
rect 11384 10868 11452 15732
rect 16316 10868 16384 15732
rect 11384 10800 16384 10868
rect 16996 15732 21996 15800
rect 16996 10868 17064 15732
rect 21928 10868 21996 15732
rect 16996 10800 21996 10868
rect 22608 15732 27608 15800
rect 22608 10868 22676 15732
rect 27540 10868 27608 15732
rect 22608 10800 27608 10868
rect 28220 15732 33220 15800
rect 28220 10868 28288 15732
rect 33152 10868 33220 15732
rect 28220 10800 33220 10868
rect 33832 15732 38832 15800
rect 33832 10868 33900 15732
rect 38764 10868 38832 15732
rect 33832 10800 38832 10868
rect -39124 10412 -34124 10480
rect -39124 5548 -39056 10412
rect -34192 5548 -34124 10412
rect -39124 5480 -34124 5548
rect -33512 10412 -28512 10480
rect -33512 5548 -33444 10412
rect -28580 5548 -28512 10412
rect -33512 5480 -28512 5548
rect -27900 10412 -22900 10480
rect -27900 5548 -27832 10412
rect -22968 5548 -22900 10412
rect -27900 5480 -22900 5548
rect -22288 10412 -17288 10480
rect -22288 5548 -22220 10412
rect -17356 5548 -17288 10412
rect -22288 5480 -17288 5548
rect -16676 10412 -11676 10480
rect -16676 5548 -16608 10412
rect -11744 5548 -11676 10412
rect -16676 5480 -11676 5548
rect -11064 10412 -6064 10480
rect -11064 5548 -10996 10412
rect -6132 5548 -6064 10412
rect -11064 5480 -6064 5548
rect -5452 10412 -452 10480
rect -5452 5548 -5384 10412
rect -520 5548 -452 10412
rect -5452 5480 -452 5548
rect 160 10412 5160 10480
rect 160 5548 228 10412
rect 5092 5548 5160 10412
rect 160 5480 5160 5548
rect 5772 10412 10772 10480
rect 5772 5548 5840 10412
rect 10704 5548 10772 10412
rect 5772 5480 10772 5548
rect 11384 10412 16384 10480
rect 11384 5548 11452 10412
rect 16316 5548 16384 10412
rect 11384 5480 16384 5548
rect 16996 10412 21996 10480
rect 16996 5548 17064 10412
rect 21928 5548 21996 10412
rect 16996 5480 21996 5548
rect 22608 10412 27608 10480
rect 22608 5548 22676 10412
rect 27540 5548 27608 10412
rect 22608 5480 27608 5548
rect 28220 10412 33220 10480
rect 28220 5548 28288 10412
rect 33152 5548 33220 10412
rect 28220 5480 33220 5548
rect 33832 10412 38832 10480
rect 33832 5548 33900 10412
rect 38764 5548 38832 10412
rect 33832 5480 38832 5548
rect -39124 5092 -34124 5160
rect -39124 228 -39056 5092
rect -34192 228 -34124 5092
rect -39124 160 -34124 228
rect -33512 5092 -28512 5160
rect -33512 228 -33444 5092
rect -28580 228 -28512 5092
rect -33512 160 -28512 228
rect -27900 5092 -22900 5160
rect -27900 228 -27832 5092
rect -22968 228 -22900 5092
rect -27900 160 -22900 228
rect -22288 5092 -17288 5160
rect -22288 228 -22220 5092
rect -17356 228 -17288 5092
rect -22288 160 -17288 228
rect -16676 5092 -11676 5160
rect -16676 228 -16608 5092
rect -11744 228 -11676 5092
rect -16676 160 -11676 228
rect -11064 5092 -6064 5160
rect -11064 228 -10996 5092
rect -6132 228 -6064 5092
rect -11064 160 -6064 228
rect -5452 5092 -452 5160
rect -5452 228 -5384 5092
rect -520 228 -452 5092
rect -5452 160 -452 228
rect 160 5092 5160 5160
rect 160 228 228 5092
rect 5092 228 5160 5092
rect 160 160 5160 228
rect 5772 5092 10772 5160
rect 5772 228 5840 5092
rect 10704 228 10772 5092
rect 5772 160 10772 228
rect 11384 5092 16384 5160
rect 11384 228 11452 5092
rect 16316 228 16384 5092
rect 11384 160 16384 228
rect 16996 5092 21996 5160
rect 16996 228 17064 5092
rect 21928 228 21996 5092
rect 16996 160 21996 228
rect 22608 5092 27608 5160
rect 22608 228 22676 5092
rect 27540 228 27608 5092
rect 22608 160 27608 228
rect 28220 5092 33220 5160
rect 28220 228 28288 5092
rect 33152 228 33220 5092
rect 28220 160 33220 228
rect 33832 5092 38832 5160
rect 33832 228 33900 5092
rect 38764 228 38832 5092
rect 33832 160 38832 228
rect -39124 -228 -34124 -160
rect -39124 -5092 -39056 -228
rect -34192 -5092 -34124 -228
rect -39124 -5160 -34124 -5092
rect -33512 -228 -28512 -160
rect -33512 -5092 -33444 -228
rect -28580 -5092 -28512 -228
rect -33512 -5160 -28512 -5092
rect -27900 -228 -22900 -160
rect -27900 -5092 -27832 -228
rect -22968 -5092 -22900 -228
rect -27900 -5160 -22900 -5092
rect -22288 -228 -17288 -160
rect -22288 -5092 -22220 -228
rect -17356 -5092 -17288 -228
rect -22288 -5160 -17288 -5092
rect -16676 -228 -11676 -160
rect -16676 -5092 -16608 -228
rect -11744 -5092 -11676 -228
rect -16676 -5160 -11676 -5092
rect -11064 -228 -6064 -160
rect -11064 -5092 -10996 -228
rect -6132 -5092 -6064 -228
rect -11064 -5160 -6064 -5092
rect -5452 -228 -452 -160
rect -5452 -5092 -5384 -228
rect -520 -5092 -452 -228
rect -5452 -5160 -452 -5092
rect 160 -228 5160 -160
rect 160 -5092 228 -228
rect 5092 -5092 5160 -228
rect 160 -5160 5160 -5092
rect 5772 -228 10772 -160
rect 5772 -5092 5840 -228
rect 10704 -5092 10772 -228
rect 5772 -5160 10772 -5092
rect 11384 -228 16384 -160
rect 11384 -5092 11452 -228
rect 16316 -5092 16384 -228
rect 11384 -5160 16384 -5092
rect 16996 -228 21996 -160
rect 16996 -5092 17064 -228
rect 21928 -5092 21996 -228
rect 16996 -5160 21996 -5092
rect 22608 -228 27608 -160
rect 22608 -5092 22676 -228
rect 27540 -5092 27608 -228
rect 22608 -5160 27608 -5092
rect 28220 -228 33220 -160
rect 28220 -5092 28288 -228
rect 33152 -5092 33220 -228
rect 28220 -5160 33220 -5092
rect 33832 -228 38832 -160
rect 33832 -5092 33900 -228
rect 38764 -5092 38832 -228
rect 33832 -5160 38832 -5092
rect -39124 -5548 -34124 -5480
rect -39124 -10412 -39056 -5548
rect -34192 -10412 -34124 -5548
rect -39124 -10480 -34124 -10412
rect -33512 -5548 -28512 -5480
rect -33512 -10412 -33444 -5548
rect -28580 -10412 -28512 -5548
rect -33512 -10480 -28512 -10412
rect -27900 -5548 -22900 -5480
rect -27900 -10412 -27832 -5548
rect -22968 -10412 -22900 -5548
rect -27900 -10480 -22900 -10412
rect -22288 -5548 -17288 -5480
rect -22288 -10412 -22220 -5548
rect -17356 -10412 -17288 -5548
rect -22288 -10480 -17288 -10412
rect -16676 -5548 -11676 -5480
rect -16676 -10412 -16608 -5548
rect -11744 -10412 -11676 -5548
rect -16676 -10480 -11676 -10412
rect -11064 -5548 -6064 -5480
rect -11064 -10412 -10996 -5548
rect -6132 -10412 -6064 -5548
rect -11064 -10480 -6064 -10412
rect -5452 -5548 -452 -5480
rect -5452 -10412 -5384 -5548
rect -520 -10412 -452 -5548
rect -5452 -10480 -452 -10412
rect 160 -5548 5160 -5480
rect 160 -10412 228 -5548
rect 5092 -10412 5160 -5548
rect 160 -10480 5160 -10412
rect 5772 -5548 10772 -5480
rect 5772 -10412 5840 -5548
rect 10704 -10412 10772 -5548
rect 5772 -10480 10772 -10412
rect 11384 -5548 16384 -5480
rect 11384 -10412 11452 -5548
rect 16316 -10412 16384 -5548
rect 11384 -10480 16384 -10412
rect 16996 -5548 21996 -5480
rect 16996 -10412 17064 -5548
rect 21928 -10412 21996 -5548
rect 16996 -10480 21996 -10412
rect 22608 -5548 27608 -5480
rect 22608 -10412 22676 -5548
rect 27540 -10412 27608 -5548
rect 22608 -10480 27608 -10412
rect 28220 -5548 33220 -5480
rect 28220 -10412 28288 -5548
rect 33152 -10412 33220 -5548
rect 28220 -10480 33220 -10412
rect 33832 -5548 38832 -5480
rect 33832 -10412 33900 -5548
rect 38764 -10412 38832 -5548
rect 33832 -10480 38832 -10412
rect -39124 -10868 -34124 -10800
rect -39124 -15732 -39056 -10868
rect -34192 -15732 -34124 -10868
rect -39124 -15800 -34124 -15732
rect -33512 -10868 -28512 -10800
rect -33512 -15732 -33444 -10868
rect -28580 -15732 -28512 -10868
rect -33512 -15800 -28512 -15732
rect -27900 -10868 -22900 -10800
rect -27900 -15732 -27832 -10868
rect -22968 -15732 -22900 -10868
rect -27900 -15800 -22900 -15732
rect -22288 -10868 -17288 -10800
rect -22288 -15732 -22220 -10868
rect -17356 -15732 -17288 -10868
rect -22288 -15800 -17288 -15732
rect -16676 -10868 -11676 -10800
rect -16676 -15732 -16608 -10868
rect -11744 -15732 -11676 -10868
rect -16676 -15800 -11676 -15732
rect -11064 -10868 -6064 -10800
rect -11064 -15732 -10996 -10868
rect -6132 -15732 -6064 -10868
rect -11064 -15800 -6064 -15732
rect -5452 -10868 -452 -10800
rect -5452 -15732 -5384 -10868
rect -520 -15732 -452 -10868
rect -5452 -15800 -452 -15732
rect 160 -10868 5160 -10800
rect 160 -15732 228 -10868
rect 5092 -15732 5160 -10868
rect 160 -15800 5160 -15732
rect 5772 -10868 10772 -10800
rect 5772 -15732 5840 -10868
rect 10704 -15732 10772 -10868
rect 5772 -15800 10772 -15732
rect 11384 -10868 16384 -10800
rect 11384 -15732 11452 -10868
rect 16316 -15732 16384 -10868
rect 11384 -15800 16384 -15732
rect 16996 -10868 21996 -10800
rect 16996 -15732 17064 -10868
rect 21928 -15732 21996 -10868
rect 16996 -15800 21996 -15732
rect 22608 -10868 27608 -10800
rect 22608 -15732 22676 -10868
rect 27540 -15732 27608 -10868
rect 22608 -15800 27608 -15732
rect 28220 -10868 33220 -10800
rect 28220 -15732 28288 -10868
rect 33152 -15732 33220 -10868
rect 28220 -15800 33220 -15732
rect 33832 -10868 38832 -10800
rect 33832 -15732 33900 -10868
rect 38764 -15732 38832 -10868
rect 33832 -15800 38832 -15732
rect -39124 -16188 -34124 -16120
rect -39124 -21052 -39056 -16188
rect -34192 -21052 -34124 -16188
rect -39124 -21120 -34124 -21052
rect -33512 -16188 -28512 -16120
rect -33512 -21052 -33444 -16188
rect -28580 -21052 -28512 -16188
rect -33512 -21120 -28512 -21052
rect -27900 -16188 -22900 -16120
rect -27900 -21052 -27832 -16188
rect -22968 -21052 -22900 -16188
rect -27900 -21120 -22900 -21052
rect -22288 -16188 -17288 -16120
rect -22288 -21052 -22220 -16188
rect -17356 -21052 -17288 -16188
rect -22288 -21120 -17288 -21052
rect -16676 -16188 -11676 -16120
rect -16676 -21052 -16608 -16188
rect -11744 -21052 -11676 -16188
rect -16676 -21120 -11676 -21052
rect -11064 -16188 -6064 -16120
rect -11064 -21052 -10996 -16188
rect -6132 -21052 -6064 -16188
rect -11064 -21120 -6064 -21052
rect -5452 -16188 -452 -16120
rect -5452 -21052 -5384 -16188
rect -520 -21052 -452 -16188
rect -5452 -21120 -452 -21052
rect 160 -16188 5160 -16120
rect 160 -21052 228 -16188
rect 5092 -21052 5160 -16188
rect 160 -21120 5160 -21052
rect 5772 -16188 10772 -16120
rect 5772 -21052 5840 -16188
rect 10704 -21052 10772 -16188
rect 5772 -21120 10772 -21052
rect 11384 -16188 16384 -16120
rect 11384 -21052 11452 -16188
rect 16316 -21052 16384 -16188
rect 11384 -21120 16384 -21052
rect 16996 -16188 21996 -16120
rect 16996 -21052 17064 -16188
rect 21928 -21052 21996 -16188
rect 16996 -21120 21996 -21052
rect 22608 -16188 27608 -16120
rect 22608 -21052 22676 -16188
rect 27540 -21052 27608 -16188
rect 22608 -21120 27608 -21052
rect 28220 -16188 33220 -16120
rect 28220 -21052 28288 -16188
rect 33152 -21052 33220 -16188
rect 28220 -21120 33220 -21052
rect 33832 -16188 38832 -16120
rect 33832 -21052 33900 -16188
rect 38764 -21052 38832 -16188
rect 33832 -21120 38832 -21052
rect -39124 -21508 -34124 -21440
rect -39124 -26372 -39056 -21508
rect -34192 -26372 -34124 -21508
rect -39124 -26440 -34124 -26372
rect -33512 -21508 -28512 -21440
rect -33512 -26372 -33444 -21508
rect -28580 -26372 -28512 -21508
rect -33512 -26440 -28512 -26372
rect -27900 -21508 -22900 -21440
rect -27900 -26372 -27832 -21508
rect -22968 -26372 -22900 -21508
rect -27900 -26440 -22900 -26372
rect -22288 -21508 -17288 -21440
rect -22288 -26372 -22220 -21508
rect -17356 -26372 -17288 -21508
rect -22288 -26440 -17288 -26372
rect -16676 -21508 -11676 -21440
rect -16676 -26372 -16608 -21508
rect -11744 -26372 -11676 -21508
rect -16676 -26440 -11676 -26372
rect -11064 -21508 -6064 -21440
rect -11064 -26372 -10996 -21508
rect -6132 -26372 -6064 -21508
rect -11064 -26440 -6064 -26372
rect -5452 -21508 -452 -21440
rect -5452 -26372 -5384 -21508
rect -520 -26372 -452 -21508
rect -5452 -26440 -452 -26372
rect 160 -21508 5160 -21440
rect 160 -26372 228 -21508
rect 5092 -26372 5160 -21508
rect 160 -26440 5160 -26372
rect 5772 -21508 10772 -21440
rect 5772 -26372 5840 -21508
rect 10704 -26372 10772 -21508
rect 5772 -26440 10772 -26372
rect 11384 -21508 16384 -21440
rect 11384 -26372 11452 -21508
rect 16316 -26372 16384 -21508
rect 11384 -26440 16384 -26372
rect 16996 -21508 21996 -21440
rect 16996 -26372 17064 -21508
rect 21928 -26372 21996 -21508
rect 16996 -26440 21996 -26372
rect 22608 -21508 27608 -21440
rect 22608 -26372 22676 -21508
rect 27540 -26372 27608 -21508
rect 22608 -26440 27608 -26372
rect 28220 -21508 33220 -21440
rect 28220 -26372 28288 -21508
rect 33152 -26372 33220 -21508
rect 28220 -26440 33220 -26372
rect 33832 -21508 38832 -21440
rect 33832 -26372 33900 -21508
rect 38764 -26372 38832 -21508
rect 33832 -26440 38832 -26372
rect -39124 -26828 -34124 -26760
rect -39124 -31692 -39056 -26828
rect -34192 -31692 -34124 -26828
rect -39124 -31760 -34124 -31692
rect -33512 -26828 -28512 -26760
rect -33512 -31692 -33444 -26828
rect -28580 -31692 -28512 -26828
rect -33512 -31760 -28512 -31692
rect -27900 -26828 -22900 -26760
rect -27900 -31692 -27832 -26828
rect -22968 -31692 -22900 -26828
rect -27900 -31760 -22900 -31692
rect -22288 -26828 -17288 -26760
rect -22288 -31692 -22220 -26828
rect -17356 -31692 -17288 -26828
rect -22288 -31760 -17288 -31692
rect -16676 -26828 -11676 -26760
rect -16676 -31692 -16608 -26828
rect -11744 -31692 -11676 -26828
rect -16676 -31760 -11676 -31692
rect -11064 -26828 -6064 -26760
rect -11064 -31692 -10996 -26828
rect -6132 -31692 -6064 -26828
rect -11064 -31760 -6064 -31692
rect -5452 -26828 -452 -26760
rect -5452 -31692 -5384 -26828
rect -520 -31692 -452 -26828
rect -5452 -31760 -452 -31692
rect 160 -26828 5160 -26760
rect 160 -31692 228 -26828
rect 5092 -31692 5160 -26828
rect 160 -31760 5160 -31692
rect 5772 -26828 10772 -26760
rect 5772 -31692 5840 -26828
rect 10704 -31692 10772 -26828
rect 5772 -31760 10772 -31692
rect 11384 -26828 16384 -26760
rect 11384 -31692 11452 -26828
rect 16316 -31692 16384 -26828
rect 11384 -31760 16384 -31692
rect 16996 -26828 21996 -26760
rect 16996 -31692 17064 -26828
rect 21928 -31692 21996 -26828
rect 16996 -31760 21996 -31692
rect 22608 -26828 27608 -26760
rect 22608 -31692 22676 -26828
rect 27540 -31692 27608 -26828
rect 22608 -31760 27608 -31692
rect 28220 -26828 33220 -26760
rect 28220 -31692 28288 -26828
rect 33152 -31692 33220 -26828
rect 28220 -31760 33220 -31692
rect 33832 -26828 38832 -26760
rect 33832 -31692 33900 -26828
rect 38764 -31692 38832 -26828
rect 33832 -31760 38832 -31692
rect -39124 -32148 -34124 -32080
rect -39124 -37012 -39056 -32148
rect -34192 -37012 -34124 -32148
rect -39124 -37080 -34124 -37012
rect -33512 -32148 -28512 -32080
rect -33512 -37012 -33444 -32148
rect -28580 -37012 -28512 -32148
rect -33512 -37080 -28512 -37012
rect -27900 -32148 -22900 -32080
rect -27900 -37012 -27832 -32148
rect -22968 -37012 -22900 -32148
rect -27900 -37080 -22900 -37012
rect -22288 -32148 -17288 -32080
rect -22288 -37012 -22220 -32148
rect -17356 -37012 -17288 -32148
rect -22288 -37080 -17288 -37012
rect -16676 -32148 -11676 -32080
rect -16676 -37012 -16608 -32148
rect -11744 -37012 -11676 -32148
rect -16676 -37080 -11676 -37012
rect -11064 -32148 -6064 -32080
rect -11064 -37012 -10996 -32148
rect -6132 -37012 -6064 -32148
rect -11064 -37080 -6064 -37012
rect -5452 -32148 -452 -32080
rect -5452 -37012 -5384 -32148
rect -520 -37012 -452 -32148
rect -5452 -37080 -452 -37012
rect 160 -32148 5160 -32080
rect 160 -37012 228 -32148
rect 5092 -37012 5160 -32148
rect 160 -37080 5160 -37012
rect 5772 -32148 10772 -32080
rect 5772 -37012 5840 -32148
rect 10704 -37012 10772 -32148
rect 5772 -37080 10772 -37012
rect 11384 -32148 16384 -32080
rect 11384 -37012 11452 -32148
rect 16316 -37012 16384 -32148
rect 11384 -37080 16384 -37012
rect 16996 -32148 21996 -32080
rect 16996 -37012 17064 -32148
rect 21928 -37012 21996 -32148
rect 16996 -37080 21996 -37012
rect 22608 -32148 27608 -32080
rect 22608 -37012 22676 -32148
rect 27540 -37012 27608 -32148
rect 22608 -37080 27608 -37012
rect 28220 -32148 33220 -32080
rect 28220 -37012 28288 -32148
rect 33152 -37012 33220 -32148
rect 28220 -37080 33220 -37012
rect 33832 -32148 38832 -32080
rect 33832 -37012 33900 -32148
rect 38764 -37012 38832 -32148
rect 33832 -37080 38832 -37012
<< mimcapcontact >>
rect -39056 32148 -34192 37012
rect -33444 32148 -28580 37012
rect -27832 32148 -22968 37012
rect -22220 32148 -17356 37012
rect -16608 32148 -11744 37012
rect -10996 32148 -6132 37012
rect -5384 32148 -520 37012
rect 228 32148 5092 37012
rect 5840 32148 10704 37012
rect 11452 32148 16316 37012
rect 17064 32148 21928 37012
rect 22676 32148 27540 37012
rect 28288 32148 33152 37012
rect 33900 32148 38764 37012
rect -39056 26828 -34192 31692
rect -33444 26828 -28580 31692
rect -27832 26828 -22968 31692
rect -22220 26828 -17356 31692
rect -16608 26828 -11744 31692
rect -10996 26828 -6132 31692
rect -5384 26828 -520 31692
rect 228 26828 5092 31692
rect 5840 26828 10704 31692
rect 11452 26828 16316 31692
rect 17064 26828 21928 31692
rect 22676 26828 27540 31692
rect 28288 26828 33152 31692
rect 33900 26828 38764 31692
rect -39056 21508 -34192 26372
rect -33444 21508 -28580 26372
rect -27832 21508 -22968 26372
rect -22220 21508 -17356 26372
rect -16608 21508 -11744 26372
rect -10996 21508 -6132 26372
rect -5384 21508 -520 26372
rect 228 21508 5092 26372
rect 5840 21508 10704 26372
rect 11452 21508 16316 26372
rect 17064 21508 21928 26372
rect 22676 21508 27540 26372
rect 28288 21508 33152 26372
rect 33900 21508 38764 26372
rect -39056 16188 -34192 21052
rect -33444 16188 -28580 21052
rect -27832 16188 -22968 21052
rect -22220 16188 -17356 21052
rect -16608 16188 -11744 21052
rect -10996 16188 -6132 21052
rect -5384 16188 -520 21052
rect 228 16188 5092 21052
rect 5840 16188 10704 21052
rect 11452 16188 16316 21052
rect 17064 16188 21928 21052
rect 22676 16188 27540 21052
rect 28288 16188 33152 21052
rect 33900 16188 38764 21052
rect -39056 10868 -34192 15732
rect -33444 10868 -28580 15732
rect -27832 10868 -22968 15732
rect -22220 10868 -17356 15732
rect -16608 10868 -11744 15732
rect -10996 10868 -6132 15732
rect -5384 10868 -520 15732
rect 228 10868 5092 15732
rect 5840 10868 10704 15732
rect 11452 10868 16316 15732
rect 17064 10868 21928 15732
rect 22676 10868 27540 15732
rect 28288 10868 33152 15732
rect 33900 10868 38764 15732
rect -39056 5548 -34192 10412
rect -33444 5548 -28580 10412
rect -27832 5548 -22968 10412
rect -22220 5548 -17356 10412
rect -16608 5548 -11744 10412
rect -10996 5548 -6132 10412
rect -5384 5548 -520 10412
rect 228 5548 5092 10412
rect 5840 5548 10704 10412
rect 11452 5548 16316 10412
rect 17064 5548 21928 10412
rect 22676 5548 27540 10412
rect 28288 5548 33152 10412
rect 33900 5548 38764 10412
rect -39056 228 -34192 5092
rect -33444 228 -28580 5092
rect -27832 228 -22968 5092
rect -22220 228 -17356 5092
rect -16608 228 -11744 5092
rect -10996 228 -6132 5092
rect -5384 228 -520 5092
rect 228 228 5092 5092
rect 5840 228 10704 5092
rect 11452 228 16316 5092
rect 17064 228 21928 5092
rect 22676 228 27540 5092
rect 28288 228 33152 5092
rect 33900 228 38764 5092
rect -39056 -5092 -34192 -228
rect -33444 -5092 -28580 -228
rect -27832 -5092 -22968 -228
rect -22220 -5092 -17356 -228
rect -16608 -5092 -11744 -228
rect -10996 -5092 -6132 -228
rect -5384 -5092 -520 -228
rect 228 -5092 5092 -228
rect 5840 -5092 10704 -228
rect 11452 -5092 16316 -228
rect 17064 -5092 21928 -228
rect 22676 -5092 27540 -228
rect 28288 -5092 33152 -228
rect 33900 -5092 38764 -228
rect -39056 -10412 -34192 -5548
rect -33444 -10412 -28580 -5548
rect -27832 -10412 -22968 -5548
rect -22220 -10412 -17356 -5548
rect -16608 -10412 -11744 -5548
rect -10996 -10412 -6132 -5548
rect -5384 -10412 -520 -5548
rect 228 -10412 5092 -5548
rect 5840 -10412 10704 -5548
rect 11452 -10412 16316 -5548
rect 17064 -10412 21928 -5548
rect 22676 -10412 27540 -5548
rect 28288 -10412 33152 -5548
rect 33900 -10412 38764 -5548
rect -39056 -15732 -34192 -10868
rect -33444 -15732 -28580 -10868
rect -27832 -15732 -22968 -10868
rect -22220 -15732 -17356 -10868
rect -16608 -15732 -11744 -10868
rect -10996 -15732 -6132 -10868
rect -5384 -15732 -520 -10868
rect 228 -15732 5092 -10868
rect 5840 -15732 10704 -10868
rect 11452 -15732 16316 -10868
rect 17064 -15732 21928 -10868
rect 22676 -15732 27540 -10868
rect 28288 -15732 33152 -10868
rect 33900 -15732 38764 -10868
rect -39056 -21052 -34192 -16188
rect -33444 -21052 -28580 -16188
rect -27832 -21052 -22968 -16188
rect -22220 -21052 -17356 -16188
rect -16608 -21052 -11744 -16188
rect -10996 -21052 -6132 -16188
rect -5384 -21052 -520 -16188
rect 228 -21052 5092 -16188
rect 5840 -21052 10704 -16188
rect 11452 -21052 16316 -16188
rect 17064 -21052 21928 -16188
rect 22676 -21052 27540 -16188
rect 28288 -21052 33152 -16188
rect 33900 -21052 38764 -16188
rect -39056 -26372 -34192 -21508
rect -33444 -26372 -28580 -21508
rect -27832 -26372 -22968 -21508
rect -22220 -26372 -17356 -21508
rect -16608 -26372 -11744 -21508
rect -10996 -26372 -6132 -21508
rect -5384 -26372 -520 -21508
rect 228 -26372 5092 -21508
rect 5840 -26372 10704 -21508
rect 11452 -26372 16316 -21508
rect 17064 -26372 21928 -21508
rect 22676 -26372 27540 -21508
rect 28288 -26372 33152 -21508
rect 33900 -26372 38764 -21508
rect -39056 -31692 -34192 -26828
rect -33444 -31692 -28580 -26828
rect -27832 -31692 -22968 -26828
rect -22220 -31692 -17356 -26828
rect -16608 -31692 -11744 -26828
rect -10996 -31692 -6132 -26828
rect -5384 -31692 -520 -26828
rect 228 -31692 5092 -26828
rect 5840 -31692 10704 -26828
rect 11452 -31692 16316 -26828
rect 17064 -31692 21928 -26828
rect 22676 -31692 27540 -26828
rect 28288 -31692 33152 -26828
rect 33900 -31692 38764 -26828
rect -39056 -37012 -34192 -32148
rect -33444 -37012 -28580 -32148
rect -27832 -37012 -22968 -32148
rect -22220 -37012 -17356 -32148
rect -16608 -37012 -11744 -32148
rect -10996 -37012 -6132 -32148
rect -5384 -37012 -520 -32148
rect 228 -37012 5092 -32148
rect 5840 -37012 10704 -32148
rect 11452 -37012 16316 -32148
rect 17064 -37012 21928 -32148
rect 22676 -37012 27540 -32148
rect 28288 -37012 33152 -32148
rect 33900 -37012 38764 -32148
<< metal4 >>
rect -36676 37041 -36572 37240
rect -33896 37092 -33792 37240
rect -39085 37012 -34163 37041
rect -39085 32148 -39056 37012
rect -34192 32148 -34163 37012
rect -39085 32119 -34163 32148
rect -33896 37028 -33876 37092
rect -33812 37028 -33792 37092
rect -31064 37041 -30960 37240
rect -28284 37092 -28180 37240
rect -33896 37012 -33792 37028
rect -33896 36948 -33876 37012
rect -33812 36948 -33792 37012
rect -33896 36932 -33792 36948
rect -33896 36868 -33876 36932
rect -33812 36868 -33792 36932
rect -33896 36852 -33792 36868
rect -33896 36788 -33876 36852
rect -33812 36788 -33792 36852
rect -33896 36772 -33792 36788
rect -33896 36708 -33876 36772
rect -33812 36708 -33792 36772
rect -33896 36692 -33792 36708
rect -33896 36628 -33876 36692
rect -33812 36628 -33792 36692
rect -33896 36612 -33792 36628
rect -33896 36548 -33876 36612
rect -33812 36548 -33792 36612
rect -33896 36532 -33792 36548
rect -33896 36468 -33876 36532
rect -33812 36468 -33792 36532
rect -33896 36452 -33792 36468
rect -33896 36388 -33876 36452
rect -33812 36388 -33792 36452
rect -33896 36372 -33792 36388
rect -33896 36308 -33876 36372
rect -33812 36308 -33792 36372
rect -33896 36292 -33792 36308
rect -33896 36228 -33876 36292
rect -33812 36228 -33792 36292
rect -33896 36212 -33792 36228
rect -33896 36148 -33876 36212
rect -33812 36148 -33792 36212
rect -33896 36132 -33792 36148
rect -33896 36068 -33876 36132
rect -33812 36068 -33792 36132
rect -33896 36052 -33792 36068
rect -33896 35988 -33876 36052
rect -33812 35988 -33792 36052
rect -33896 35972 -33792 35988
rect -33896 35908 -33876 35972
rect -33812 35908 -33792 35972
rect -33896 35892 -33792 35908
rect -33896 35828 -33876 35892
rect -33812 35828 -33792 35892
rect -33896 35812 -33792 35828
rect -33896 35748 -33876 35812
rect -33812 35748 -33792 35812
rect -33896 35732 -33792 35748
rect -33896 35668 -33876 35732
rect -33812 35668 -33792 35732
rect -33896 35652 -33792 35668
rect -33896 35588 -33876 35652
rect -33812 35588 -33792 35652
rect -33896 35572 -33792 35588
rect -33896 35508 -33876 35572
rect -33812 35508 -33792 35572
rect -33896 35492 -33792 35508
rect -33896 35428 -33876 35492
rect -33812 35428 -33792 35492
rect -33896 35412 -33792 35428
rect -33896 35348 -33876 35412
rect -33812 35348 -33792 35412
rect -33896 35332 -33792 35348
rect -33896 35268 -33876 35332
rect -33812 35268 -33792 35332
rect -33896 35252 -33792 35268
rect -33896 35188 -33876 35252
rect -33812 35188 -33792 35252
rect -33896 35172 -33792 35188
rect -33896 35108 -33876 35172
rect -33812 35108 -33792 35172
rect -33896 35092 -33792 35108
rect -33896 35028 -33876 35092
rect -33812 35028 -33792 35092
rect -33896 35012 -33792 35028
rect -33896 34948 -33876 35012
rect -33812 34948 -33792 35012
rect -33896 34932 -33792 34948
rect -33896 34868 -33876 34932
rect -33812 34868 -33792 34932
rect -33896 34852 -33792 34868
rect -33896 34788 -33876 34852
rect -33812 34788 -33792 34852
rect -33896 34772 -33792 34788
rect -33896 34708 -33876 34772
rect -33812 34708 -33792 34772
rect -33896 34692 -33792 34708
rect -33896 34628 -33876 34692
rect -33812 34628 -33792 34692
rect -33896 34612 -33792 34628
rect -33896 34548 -33876 34612
rect -33812 34548 -33792 34612
rect -33896 34532 -33792 34548
rect -33896 34468 -33876 34532
rect -33812 34468 -33792 34532
rect -33896 34452 -33792 34468
rect -33896 34388 -33876 34452
rect -33812 34388 -33792 34452
rect -33896 34372 -33792 34388
rect -33896 34308 -33876 34372
rect -33812 34308 -33792 34372
rect -33896 34292 -33792 34308
rect -33896 34228 -33876 34292
rect -33812 34228 -33792 34292
rect -33896 34212 -33792 34228
rect -33896 34148 -33876 34212
rect -33812 34148 -33792 34212
rect -33896 34132 -33792 34148
rect -33896 34068 -33876 34132
rect -33812 34068 -33792 34132
rect -33896 34052 -33792 34068
rect -33896 33988 -33876 34052
rect -33812 33988 -33792 34052
rect -33896 33972 -33792 33988
rect -33896 33908 -33876 33972
rect -33812 33908 -33792 33972
rect -33896 33892 -33792 33908
rect -33896 33828 -33876 33892
rect -33812 33828 -33792 33892
rect -33896 33812 -33792 33828
rect -33896 33748 -33876 33812
rect -33812 33748 -33792 33812
rect -33896 33732 -33792 33748
rect -33896 33668 -33876 33732
rect -33812 33668 -33792 33732
rect -33896 33652 -33792 33668
rect -33896 33588 -33876 33652
rect -33812 33588 -33792 33652
rect -33896 33572 -33792 33588
rect -33896 33508 -33876 33572
rect -33812 33508 -33792 33572
rect -33896 33492 -33792 33508
rect -33896 33428 -33876 33492
rect -33812 33428 -33792 33492
rect -33896 33412 -33792 33428
rect -33896 33348 -33876 33412
rect -33812 33348 -33792 33412
rect -33896 33332 -33792 33348
rect -33896 33268 -33876 33332
rect -33812 33268 -33792 33332
rect -33896 33252 -33792 33268
rect -33896 33188 -33876 33252
rect -33812 33188 -33792 33252
rect -33896 33172 -33792 33188
rect -33896 33108 -33876 33172
rect -33812 33108 -33792 33172
rect -33896 33092 -33792 33108
rect -33896 33028 -33876 33092
rect -33812 33028 -33792 33092
rect -33896 33012 -33792 33028
rect -33896 32948 -33876 33012
rect -33812 32948 -33792 33012
rect -33896 32932 -33792 32948
rect -33896 32868 -33876 32932
rect -33812 32868 -33792 32932
rect -33896 32852 -33792 32868
rect -33896 32788 -33876 32852
rect -33812 32788 -33792 32852
rect -33896 32772 -33792 32788
rect -33896 32708 -33876 32772
rect -33812 32708 -33792 32772
rect -33896 32692 -33792 32708
rect -33896 32628 -33876 32692
rect -33812 32628 -33792 32692
rect -33896 32612 -33792 32628
rect -33896 32548 -33876 32612
rect -33812 32548 -33792 32612
rect -33896 32532 -33792 32548
rect -33896 32468 -33876 32532
rect -33812 32468 -33792 32532
rect -33896 32452 -33792 32468
rect -33896 32388 -33876 32452
rect -33812 32388 -33792 32452
rect -33896 32372 -33792 32388
rect -33896 32308 -33876 32372
rect -33812 32308 -33792 32372
rect -33896 32292 -33792 32308
rect -33896 32228 -33876 32292
rect -33812 32228 -33792 32292
rect -33896 32212 -33792 32228
rect -33896 32148 -33876 32212
rect -33812 32148 -33792 32212
rect -33896 32132 -33792 32148
rect -36676 31721 -36572 32119
rect -33896 32068 -33876 32132
rect -33812 32068 -33792 32132
rect -33473 37012 -28551 37041
rect -33473 32148 -33444 37012
rect -28580 32148 -28551 37012
rect -33473 32119 -28551 32148
rect -28284 37028 -28264 37092
rect -28200 37028 -28180 37092
rect -25452 37041 -25348 37240
rect -22672 37092 -22568 37240
rect -28284 37012 -28180 37028
rect -28284 36948 -28264 37012
rect -28200 36948 -28180 37012
rect -28284 36932 -28180 36948
rect -28284 36868 -28264 36932
rect -28200 36868 -28180 36932
rect -28284 36852 -28180 36868
rect -28284 36788 -28264 36852
rect -28200 36788 -28180 36852
rect -28284 36772 -28180 36788
rect -28284 36708 -28264 36772
rect -28200 36708 -28180 36772
rect -28284 36692 -28180 36708
rect -28284 36628 -28264 36692
rect -28200 36628 -28180 36692
rect -28284 36612 -28180 36628
rect -28284 36548 -28264 36612
rect -28200 36548 -28180 36612
rect -28284 36532 -28180 36548
rect -28284 36468 -28264 36532
rect -28200 36468 -28180 36532
rect -28284 36452 -28180 36468
rect -28284 36388 -28264 36452
rect -28200 36388 -28180 36452
rect -28284 36372 -28180 36388
rect -28284 36308 -28264 36372
rect -28200 36308 -28180 36372
rect -28284 36292 -28180 36308
rect -28284 36228 -28264 36292
rect -28200 36228 -28180 36292
rect -28284 36212 -28180 36228
rect -28284 36148 -28264 36212
rect -28200 36148 -28180 36212
rect -28284 36132 -28180 36148
rect -28284 36068 -28264 36132
rect -28200 36068 -28180 36132
rect -28284 36052 -28180 36068
rect -28284 35988 -28264 36052
rect -28200 35988 -28180 36052
rect -28284 35972 -28180 35988
rect -28284 35908 -28264 35972
rect -28200 35908 -28180 35972
rect -28284 35892 -28180 35908
rect -28284 35828 -28264 35892
rect -28200 35828 -28180 35892
rect -28284 35812 -28180 35828
rect -28284 35748 -28264 35812
rect -28200 35748 -28180 35812
rect -28284 35732 -28180 35748
rect -28284 35668 -28264 35732
rect -28200 35668 -28180 35732
rect -28284 35652 -28180 35668
rect -28284 35588 -28264 35652
rect -28200 35588 -28180 35652
rect -28284 35572 -28180 35588
rect -28284 35508 -28264 35572
rect -28200 35508 -28180 35572
rect -28284 35492 -28180 35508
rect -28284 35428 -28264 35492
rect -28200 35428 -28180 35492
rect -28284 35412 -28180 35428
rect -28284 35348 -28264 35412
rect -28200 35348 -28180 35412
rect -28284 35332 -28180 35348
rect -28284 35268 -28264 35332
rect -28200 35268 -28180 35332
rect -28284 35252 -28180 35268
rect -28284 35188 -28264 35252
rect -28200 35188 -28180 35252
rect -28284 35172 -28180 35188
rect -28284 35108 -28264 35172
rect -28200 35108 -28180 35172
rect -28284 35092 -28180 35108
rect -28284 35028 -28264 35092
rect -28200 35028 -28180 35092
rect -28284 35012 -28180 35028
rect -28284 34948 -28264 35012
rect -28200 34948 -28180 35012
rect -28284 34932 -28180 34948
rect -28284 34868 -28264 34932
rect -28200 34868 -28180 34932
rect -28284 34852 -28180 34868
rect -28284 34788 -28264 34852
rect -28200 34788 -28180 34852
rect -28284 34772 -28180 34788
rect -28284 34708 -28264 34772
rect -28200 34708 -28180 34772
rect -28284 34692 -28180 34708
rect -28284 34628 -28264 34692
rect -28200 34628 -28180 34692
rect -28284 34612 -28180 34628
rect -28284 34548 -28264 34612
rect -28200 34548 -28180 34612
rect -28284 34532 -28180 34548
rect -28284 34468 -28264 34532
rect -28200 34468 -28180 34532
rect -28284 34452 -28180 34468
rect -28284 34388 -28264 34452
rect -28200 34388 -28180 34452
rect -28284 34372 -28180 34388
rect -28284 34308 -28264 34372
rect -28200 34308 -28180 34372
rect -28284 34292 -28180 34308
rect -28284 34228 -28264 34292
rect -28200 34228 -28180 34292
rect -28284 34212 -28180 34228
rect -28284 34148 -28264 34212
rect -28200 34148 -28180 34212
rect -28284 34132 -28180 34148
rect -28284 34068 -28264 34132
rect -28200 34068 -28180 34132
rect -28284 34052 -28180 34068
rect -28284 33988 -28264 34052
rect -28200 33988 -28180 34052
rect -28284 33972 -28180 33988
rect -28284 33908 -28264 33972
rect -28200 33908 -28180 33972
rect -28284 33892 -28180 33908
rect -28284 33828 -28264 33892
rect -28200 33828 -28180 33892
rect -28284 33812 -28180 33828
rect -28284 33748 -28264 33812
rect -28200 33748 -28180 33812
rect -28284 33732 -28180 33748
rect -28284 33668 -28264 33732
rect -28200 33668 -28180 33732
rect -28284 33652 -28180 33668
rect -28284 33588 -28264 33652
rect -28200 33588 -28180 33652
rect -28284 33572 -28180 33588
rect -28284 33508 -28264 33572
rect -28200 33508 -28180 33572
rect -28284 33492 -28180 33508
rect -28284 33428 -28264 33492
rect -28200 33428 -28180 33492
rect -28284 33412 -28180 33428
rect -28284 33348 -28264 33412
rect -28200 33348 -28180 33412
rect -28284 33332 -28180 33348
rect -28284 33268 -28264 33332
rect -28200 33268 -28180 33332
rect -28284 33252 -28180 33268
rect -28284 33188 -28264 33252
rect -28200 33188 -28180 33252
rect -28284 33172 -28180 33188
rect -28284 33108 -28264 33172
rect -28200 33108 -28180 33172
rect -28284 33092 -28180 33108
rect -28284 33028 -28264 33092
rect -28200 33028 -28180 33092
rect -28284 33012 -28180 33028
rect -28284 32948 -28264 33012
rect -28200 32948 -28180 33012
rect -28284 32932 -28180 32948
rect -28284 32868 -28264 32932
rect -28200 32868 -28180 32932
rect -28284 32852 -28180 32868
rect -28284 32788 -28264 32852
rect -28200 32788 -28180 32852
rect -28284 32772 -28180 32788
rect -28284 32708 -28264 32772
rect -28200 32708 -28180 32772
rect -28284 32692 -28180 32708
rect -28284 32628 -28264 32692
rect -28200 32628 -28180 32692
rect -28284 32612 -28180 32628
rect -28284 32548 -28264 32612
rect -28200 32548 -28180 32612
rect -28284 32532 -28180 32548
rect -28284 32468 -28264 32532
rect -28200 32468 -28180 32532
rect -28284 32452 -28180 32468
rect -28284 32388 -28264 32452
rect -28200 32388 -28180 32452
rect -28284 32372 -28180 32388
rect -28284 32308 -28264 32372
rect -28200 32308 -28180 32372
rect -28284 32292 -28180 32308
rect -28284 32228 -28264 32292
rect -28200 32228 -28180 32292
rect -28284 32212 -28180 32228
rect -28284 32148 -28264 32212
rect -28200 32148 -28180 32212
rect -28284 32132 -28180 32148
rect -33896 31772 -33792 32068
rect -39085 31692 -34163 31721
rect -39085 26828 -39056 31692
rect -34192 26828 -34163 31692
rect -39085 26799 -34163 26828
rect -33896 31708 -33876 31772
rect -33812 31708 -33792 31772
rect -31064 31721 -30960 32119
rect -28284 32068 -28264 32132
rect -28200 32068 -28180 32132
rect -27861 37012 -22939 37041
rect -27861 32148 -27832 37012
rect -22968 32148 -22939 37012
rect -27861 32119 -22939 32148
rect -22672 37028 -22652 37092
rect -22588 37028 -22568 37092
rect -19840 37041 -19736 37240
rect -17060 37092 -16956 37240
rect -22672 37012 -22568 37028
rect -22672 36948 -22652 37012
rect -22588 36948 -22568 37012
rect -22672 36932 -22568 36948
rect -22672 36868 -22652 36932
rect -22588 36868 -22568 36932
rect -22672 36852 -22568 36868
rect -22672 36788 -22652 36852
rect -22588 36788 -22568 36852
rect -22672 36772 -22568 36788
rect -22672 36708 -22652 36772
rect -22588 36708 -22568 36772
rect -22672 36692 -22568 36708
rect -22672 36628 -22652 36692
rect -22588 36628 -22568 36692
rect -22672 36612 -22568 36628
rect -22672 36548 -22652 36612
rect -22588 36548 -22568 36612
rect -22672 36532 -22568 36548
rect -22672 36468 -22652 36532
rect -22588 36468 -22568 36532
rect -22672 36452 -22568 36468
rect -22672 36388 -22652 36452
rect -22588 36388 -22568 36452
rect -22672 36372 -22568 36388
rect -22672 36308 -22652 36372
rect -22588 36308 -22568 36372
rect -22672 36292 -22568 36308
rect -22672 36228 -22652 36292
rect -22588 36228 -22568 36292
rect -22672 36212 -22568 36228
rect -22672 36148 -22652 36212
rect -22588 36148 -22568 36212
rect -22672 36132 -22568 36148
rect -22672 36068 -22652 36132
rect -22588 36068 -22568 36132
rect -22672 36052 -22568 36068
rect -22672 35988 -22652 36052
rect -22588 35988 -22568 36052
rect -22672 35972 -22568 35988
rect -22672 35908 -22652 35972
rect -22588 35908 -22568 35972
rect -22672 35892 -22568 35908
rect -22672 35828 -22652 35892
rect -22588 35828 -22568 35892
rect -22672 35812 -22568 35828
rect -22672 35748 -22652 35812
rect -22588 35748 -22568 35812
rect -22672 35732 -22568 35748
rect -22672 35668 -22652 35732
rect -22588 35668 -22568 35732
rect -22672 35652 -22568 35668
rect -22672 35588 -22652 35652
rect -22588 35588 -22568 35652
rect -22672 35572 -22568 35588
rect -22672 35508 -22652 35572
rect -22588 35508 -22568 35572
rect -22672 35492 -22568 35508
rect -22672 35428 -22652 35492
rect -22588 35428 -22568 35492
rect -22672 35412 -22568 35428
rect -22672 35348 -22652 35412
rect -22588 35348 -22568 35412
rect -22672 35332 -22568 35348
rect -22672 35268 -22652 35332
rect -22588 35268 -22568 35332
rect -22672 35252 -22568 35268
rect -22672 35188 -22652 35252
rect -22588 35188 -22568 35252
rect -22672 35172 -22568 35188
rect -22672 35108 -22652 35172
rect -22588 35108 -22568 35172
rect -22672 35092 -22568 35108
rect -22672 35028 -22652 35092
rect -22588 35028 -22568 35092
rect -22672 35012 -22568 35028
rect -22672 34948 -22652 35012
rect -22588 34948 -22568 35012
rect -22672 34932 -22568 34948
rect -22672 34868 -22652 34932
rect -22588 34868 -22568 34932
rect -22672 34852 -22568 34868
rect -22672 34788 -22652 34852
rect -22588 34788 -22568 34852
rect -22672 34772 -22568 34788
rect -22672 34708 -22652 34772
rect -22588 34708 -22568 34772
rect -22672 34692 -22568 34708
rect -22672 34628 -22652 34692
rect -22588 34628 -22568 34692
rect -22672 34612 -22568 34628
rect -22672 34548 -22652 34612
rect -22588 34548 -22568 34612
rect -22672 34532 -22568 34548
rect -22672 34468 -22652 34532
rect -22588 34468 -22568 34532
rect -22672 34452 -22568 34468
rect -22672 34388 -22652 34452
rect -22588 34388 -22568 34452
rect -22672 34372 -22568 34388
rect -22672 34308 -22652 34372
rect -22588 34308 -22568 34372
rect -22672 34292 -22568 34308
rect -22672 34228 -22652 34292
rect -22588 34228 -22568 34292
rect -22672 34212 -22568 34228
rect -22672 34148 -22652 34212
rect -22588 34148 -22568 34212
rect -22672 34132 -22568 34148
rect -22672 34068 -22652 34132
rect -22588 34068 -22568 34132
rect -22672 34052 -22568 34068
rect -22672 33988 -22652 34052
rect -22588 33988 -22568 34052
rect -22672 33972 -22568 33988
rect -22672 33908 -22652 33972
rect -22588 33908 -22568 33972
rect -22672 33892 -22568 33908
rect -22672 33828 -22652 33892
rect -22588 33828 -22568 33892
rect -22672 33812 -22568 33828
rect -22672 33748 -22652 33812
rect -22588 33748 -22568 33812
rect -22672 33732 -22568 33748
rect -22672 33668 -22652 33732
rect -22588 33668 -22568 33732
rect -22672 33652 -22568 33668
rect -22672 33588 -22652 33652
rect -22588 33588 -22568 33652
rect -22672 33572 -22568 33588
rect -22672 33508 -22652 33572
rect -22588 33508 -22568 33572
rect -22672 33492 -22568 33508
rect -22672 33428 -22652 33492
rect -22588 33428 -22568 33492
rect -22672 33412 -22568 33428
rect -22672 33348 -22652 33412
rect -22588 33348 -22568 33412
rect -22672 33332 -22568 33348
rect -22672 33268 -22652 33332
rect -22588 33268 -22568 33332
rect -22672 33252 -22568 33268
rect -22672 33188 -22652 33252
rect -22588 33188 -22568 33252
rect -22672 33172 -22568 33188
rect -22672 33108 -22652 33172
rect -22588 33108 -22568 33172
rect -22672 33092 -22568 33108
rect -22672 33028 -22652 33092
rect -22588 33028 -22568 33092
rect -22672 33012 -22568 33028
rect -22672 32948 -22652 33012
rect -22588 32948 -22568 33012
rect -22672 32932 -22568 32948
rect -22672 32868 -22652 32932
rect -22588 32868 -22568 32932
rect -22672 32852 -22568 32868
rect -22672 32788 -22652 32852
rect -22588 32788 -22568 32852
rect -22672 32772 -22568 32788
rect -22672 32708 -22652 32772
rect -22588 32708 -22568 32772
rect -22672 32692 -22568 32708
rect -22672 32628 -22652 32692
rect -22588 32628 -22568 32692
rect -22672 32612 -22568 32628
rect -22672 32548 -22652 32612
rect -22588 32548 -22568 32612
rect -22672 32532 -22568 32548
rect -22672 32468 -22652 32532
rect -22588 32468 -22568 32532
rect -22672 32452 -22568 32468
rect -22672 32388 -22652 32452
rect -22588 32388 -22568 32452
rect -22672 32372 -22568 32388
rect -22672 32308 -22652 32372
rect -22588 32308 -22568 32372
rect -22672 32292 -22568 32308
rect -22672 32228 -22652 32292
rect -22588 32228 -22568 32292
rect -22672 32212 -22568 32228
rect -22672 32148 -22652 32212
rect -22588 32148 -22568 32212
rect -22672 32132 -22568 32148
rect -28284 31772 -28180 32068
rect -33896 31692 -33792 31708
rect -33896 31628 -33876 31692
rect -33812 31628 -33792 31692
rect -33896 31612 -33792 31628
rect -33896 31548 -33876 31612
rect -33812 31548 -33792 31612
rect -33896 31532 -33792 31548
rect -33896 31468 -33876 31532
rect -33812 31468 -33792 31532
rect -33896 31452 -33792 31468
rect -33896 31388 -33876 31452
rect -33812 31388 -33792 31452
rect -33896 31372 -33792 31388
rect -33896 31308 -33876 31372
rect -33812 31308 -33792 31372
rect -33896 31292 -33792 31308
rect -33896 31228 -33876 31292
rect -33812 31228 -33792 31292
rect -33896 31212 -33792 31228
rect -33896 31148 -33876 31212
rect -33812 31148 -33792 31212
rect -33896 31132 -33792 31148
rect -33896 31068 -33876 31132
rect -33812 31068 -33792 31132
rect -33896 31052 -33792 31068
rect -33896 30988 -33876 31052
rect -33812 30988 -33792 31052
rect -33896 30972 -33792 30988
rect -33896 30908 -33876 30972
rect -33812 30908 -33792 30972
rect -33896 30892 -33792 30908
rect -33896 30828 -33876 30892
rect -33812 30828 -33792 30892
rect -33896 30812 -33792 30828
rect -33896 30748 -33876 30812
rect -33812 30748 -33792 30812
rect -33896 30732 -33792 30748
rect -33896 30668 -33876 30732
rect -33812 30668 -33792 30732
rect -33896 30652 -33792 30668
rect -33896 30588 -33876 30652
rect -33812 30588 -33792 30652
rect -33896 30572 -33792 30588
rect -33896 30508 -33876 30572
rect -33812 30508 -33792 30572
rect -33896 30492 -33792 30508
rect -33896 30428 -33876 30492
rect -33812 30428 -33792 30492
rect -33896 30412 -33792 30428
rect -33896 30348 -33876 30412
rect -33812 30348 -33792 30412
rect -33896 30332 -33792 30348
rect -33896 30268 -33876 30332
rect -33812 30268 -33792 30332
rect -33896 30252 -33792 30268
rect -33896 30188 -33876 30252
rect -33812 30188 -33792 30252
rect -33896 30172 -33792 30188
rect -33896 30108 -33876 30172
rect -33812 30108 -33792 30172
rect -33896 30092 -33792 30108
rect -33896 30028 -33876 30092
rect -33812 30028 -33792 30092
rect -33896 30012 -33792 30028
rect -33896 29948 -33876 30012
rect -33812 29948 -33792 30012
rect -33896 29932 -33792 29948
rect -33896 29868 -33876 29932
rect -33812 29868 -33792 29932
rect -33896 29852 -33792 29868
rect -33896 29788 -33876 29852
rect -33812 29788 -33792 29852
rect -33896 29772 -33792 29788
rect -33896 29708 -33876 29772
rect -33812 29708 -33792 29772
rect -33896 29692 -33792 29708
rect -33896 29628 -33876 29692
rect -33812 29628 -33792 29692
rect -33896 29612 -33792 29628
rect -33896 29548 -33876 29612
rect -33812 29548 -33792 29612
rect -33896 29532 -33792 29548
rect -33896 29468 -33876 29532
rect -33812 29468 -33792 29532
rect -33896 29452 -33792 29468
rect -33896 29388 -33876 29452
rect -33812 29388 -33792 29452
rect -33896 29372 -33792 29388
rect -33896 29308 -33876 29372
rect -33812 29308 -33792 29372
rect -33896 29292 -33792 29308
rect -33896 29228 -33876 29292
rect -33812 29228 -33792 29292
rect -33896 29212 -33792 29228
rect -33896 29148 -33876 29212
rect -33812 29148 -33792 29212
rect -33896 29132 -33792 29148
rect -33896 29068 -33876 29132
rect -33812 29068 -33792 29132
rect -33896 29052 -33792 29068
rect -33896 28988 -33876 29052
rect -33812 28988 -33792 29052
rect -33896 28972 -33792 28988
rect -33896 28908 -33876 28972
rect -33812 28908 -33792 28972
rect -33896 28892 -33792 28908
rect -33896 28828 -33876 28892
rect -33812 28828 -33792 28892
rect -33896 28812 -33792 28828
rect -33896 28748 -33876 28812
rect -33812 28748 -33792 28812
rect -33896 28732 -33792 28748
rect -33896 28668 -33876 28732
rect -33812 28668 -33792 28732
rect -33896 28652 -33792 28668
rect -33896 28588 -33876 28652
rect -33812 28588 -33792 28652
rect -33896 28572 -33792 28588
rect -33896 28508 -33876 28572
rect -33812 28508 -33792 28572
rect -33896 28492 -33792 28508
rect -33896 28428 -33876 28492
rect -33812 28428 -33792 28492
rect -33896 28412 -33792 28428
rect -33896 28348 -33876 28412
rect -33812 28348 -33792 28412
rect -33896 28332 -33792 28348
rect -33896 28268 -33876 28332
rect -33812 28268 -33792 28332
rect -33896 28252 -33792 28268
rect -33896 28188 -33876 28252
rect -33812 28188 -33792 28252
rect -33896 28172 -33792 28188
rect -33896 28108 -33876 28172
rect -33812 28108 -33792 28172
rect -33896 28092 -33792 28108
rect -33896 28028 -33876 28092
rect -33812 28028 -33792 28092
rect -33896 28012 -33792 28028
rect -33896 27948 -33876 28012
rect -33812 27948 -33792 28012
rect -33896 27932 -33792 27948
rect -33896 27868 -33876 27932
rect -33812 27868 -33792 27932
rect -33896 27852 -33792 27868
rect -33896 27788 -33876 27852
rect -33812 27788 -33792 27852
rect -33896 27772 -33792 27788
rect -33896 27708 -33876 27772
rect -33812 27708 -33792 27772
rect -33896 27692 -33792 27708
rect -33896 27628 -33876 27692
rect -33812 27628 -33792 27692
rect -33896 27612 -33792 27628
rect -33896 27548 -33876 27612
rect -33812 27548 -33792 27612
rect -33896 27532 -33792 27548
rect -33896 27468 -33876 27532
rect -33812 27468 -33792 27532
rect -33896 27452 -33792 27468
rect -33896 27388 -33876 27452
rect -33812 27388 -33792 27452
rect -33896 27372 -33792 27388
rect -33896 27308 -33876 27372
rect -33812 27308 -33792 27372
rect -33896 27292 -33792 27308
rect -33896 27228 -33876 27292
rect -33812 27228 -33792 27292
rect -33896 27212 -33792 27228
rect -33896 27148 -33876 27212
rect -33812 27148 -33792 27212
rect -33896 27132 -33792 27148
rect -33896 27068 -33876 27132
rect -33812 27068 -33792 27132
rect -33896 27052 -33792 27068
rect -33896 26988 -33876 27052
rect -33812 26988 -33792 27052
rect -33896 26972 -33792 26988
rect -33896 26908 -33876 26972
rect -33812 26908 -33792 26972
rect -33896 26892 -33792 26908
rect -33896 26828 -33876 26892
rect -33812 26828 -33792 26892
rect -33896 26812 -33792 26828
rect -36676 26401 -36572 26799
rect -33896 26748 -33876 26812
rect -33812 26748 -33792 26812
rect -33473 31692 -28551 31721
rect -33473 26828 -33444 31692
rect -28580 26828 -28551 31692
rect -33473 26799 -28551 26828
rect -28284 31708 -28264 31772
rect -28200 31708 -28180 31772
rect -25452 31721 -25348 32119
rect -22672 32068 -22652 32132
rect -22588 32068 -22568 32132
rect -22249 37012 -17327 37041
rect -22249 32148 -22220 37012
rect -17356 32148 -17327 37012
rect -22249 32119 -17327 32148
rect -17060 37028 -17040 37092
rect -16976 37028 -16956 37092
rect -14228 37041 -14124 37240
rect -11448 37092 -11344 37240
rect -17060 37012 -16956 37028
rect -17060 36948 -17040 37012
rect -16976 36948 -16956 37012
rect -17060 36932 -16956 36948
rect -17060 36868 -17040 36932
rect -16976 36868 -16956 36932
rect -17060 36852 -16956 36868
rect -17060 36788 -17040 36852
rect -16976 36788 -16956 36852
rect -17060 36772 -16956 36788
rect -17060 36708 -17040 36772
rect -16976 36708 -16956 36772
rect -17060 36692 -16956 36708
rect -17060 36628 -17040 36692
rect -16976 36628 -16956 36692
rect -17060 36612 -16956 36628
rect -17060 36548 -17040 36612
rect -16976 36548 -16956 36612
rect -17060 36532 -16956 36548
rect -17060 36468 -17040 36532
rect -16976 36468 -16956 36532
rect -17060 36452 -16956 36468
rect -17060 36388 -17040 36452
rect -16976 36388 -16956 36452
rect -17060 36372 -16956 36388
rect -17060 36308 -17040 36372
rect -16976 36308 -16956 36372
rect -17060 36292 -16956 36308
rect -17060 36228 -17040 36292
rect -16976 36228 -16956 36292
rect -17060 36212 -16956 36228
rect -17060 36148 -17040 36212
rect -16976 36148 -16956 36212
rect -17060 36132 -16956 36148
rect -17060 36068 -17040 36132
rect -16976 36068 -16956 36132
rect -17060 36052 -16956 36068
rect -17060 35988 -17040 36052
rect -16976 35988 -16956 36052
rect -17060 35972 -16956 35988
rect -17060 35908 -17040 35972
rect -16976 35908 -16956 35972
rect -17060 35892 -16956 35908
rect -17060 35828 -17040 35892
rect -16976 35828 -16956 35892
rect -17060 35812 -16956 35828
rect -17060 35748 -17040 35812
rect -16976 35748 -16956 35812
rect -17060 35732 -16956 35748
rect -17060 35668 -17040 35732
rect -16976 35668 -16956 35732
rect -17060 35652 -16956 35668
rect -17060 35588 -17040 35652
rect -16976 35588 -16956 35652
rect -17060 35572 -16956 35588
rect -17060 35508 -17040 35572
rect -16976 35508 -16956 35572
rect -17060 35492 -16956 35508
rect -17060 35428 -17040 35492
rect -16976 35428 -16956 35492
rect -17060 35412 -16956 35428
rect -17060 35348 -17040 35412
rect -16976 35348 -16956 35412
rect -17060 35332 -16956 35348
rect -17060 35268 -17040 35332
rect -16976 35268 -16956 35332
rect -17060 35252 -16956 35268
rect -17060 35188 -17040 35252
rect -16976 35188 -16956 35252
rect -17060 35172 -16956 35188
rect -17060 35108 -17040 35172
rect -16976 35108 -16956 35172
rect -17060 35092 -16956 35108
rect -17060 35028 -17040 35092
rect -16976 35028 -16956 35092
rect -17060 35012 -16956 35028
rect -17060 34948 -17040 35012
rect -16976 34948 -16956 35012
rect -17060 34932 -16956 34948
rect -17060 34868 -17040 34932
rect -16976 34868 -16956 34932
rect -17060 34852 -16956 34868
rect -17060 34788 -17040 34852
rect -16976 34788 -16956 34852
rect -17060 34772 -16956 34788
rect -17060 34708 -17040 34772
rect -16976 34708 -16956 34772
rect -17060 34692 -16956 34708
rect -17060 34628 -17040 34692
rect -16976 34628 -16956 34692
rect -17060 34612 -16956 34628
rect -17060 34548 -17040 34612
rect -16976 34548 -16956 34612
rect -17060 34532 -16956 34548
rect -17060 34468 -17040 34532
rect -16976 34468 -16956 34532
rect -17060 34452 -16956 34468
rect -17060 34388 -17040 34452
rect -16976 34388 -16956 34452
rect -17060 34372 -16956 34388
rect -17060 34308 -17040 34372
rect -16976 34308 -16956 34372
rect -17060 34292 -16956 34308
rect -17060 34228 -17040 34292
rect -16976 34228 -16956 34292
rect -17060 34212 -16956 34228
rect -17060 34148 -17040 34212
rect -16976 34148 -16956 34212
rect -17060 34132 -16956 34148
rect -17060 34068 -17040 34132
rect -16976 34068 -16956 34132
rect -17060 34052 -16956 34068
rect -17060 33988 -17040 34052
rect -16976 33988 -16956 34052
rect -17060 33972 -16956 33988
rect -17060 33908 -17040 33972
rect -16976 33908 -16956 33972
rect -17060 33892 -16956 33908
rect -17060 33828 -17040 33892
rect -16976 33828 -16956 33892
rect -17060 33812 -16956 33828
rect -17060 33748 -17040 33812
rect -16976 33748 -16956 33812
rect -17060 33732 -16956 33748
rect -17060 33668 -17040 33732
rect -16976 33668 -16956 33732
rect -17060 33652 -16956 33668
rect -17060 33588 -17040 33652
rect -16976 33588 -16956 33652
rect -17060 33572 -16956 33588
rect -17060 33508 -17040 33572
rect -16976 33508 -16956 33572
rect -17060 33492 -16956 33508
rect -17060 33428 -17040 33492
rect -16976 33428 -16956 33492
rect -17060 33412 -16956 33428
rect -17060 33348 -17040 33412
rect -16976 33348 -16956 33412
rect -17060 33332 -16956 33348
rect -17060 33268 -17040 33332
rect -16976 33268 -16956 33332
rect -17060 33252 -16956 33268
rect -17060 33188 -17040 33252
rect -16976 33188 -16956 33252
rect -17060 33172 -16956 33188
rect -17060 33108 -17040 33172
rect -16976 33108 -16956 33172
rect -17060 33092 -16956 33108
rect -17060 33028 -17040 33092
rect -16976 33028 -16956 33092
rect -17060 33012 -16956 33028
rect -17060 32948 -17040 33012
rect -16976 32948 -16956 33012
rect -17060 32932 -16956 32948
rect -17060 32868 -17040 32932
rect -16976 32868 -16956 32932
rect -17060 32852 -16956 32868
rect -17060 32788 -17040 32852
rect -16976 32788 -16956 32852
rect -17060 32772 -16956 32788
rect -17060 32708 -17040 32772
rect -16976 32708 -16956 32772
rect -17060 32692 -16956 32708
rect -17060 32628 -17040 32692
rect -16976 32628 -16956 32692
rect -17060 32612 -16956 32628
rect -17060 32548 -17040 32612
rect -16976 32548 -16956 32612
rect -17060 32532 -16956 32548
rect -17060 32468 -17040 32532
rect -16976 32468 -16956 32532
rect -17060 32452 -16956 32468
rect -17060 32388 -17040 32452
rect -16976 32388 -16956 32452
rect -17060 32372 -16956 32388
rect -17060 32308 -17040 32372
rect -16976 32308 -16956 32372
rect -17060 32292 -16956 32308
rect -17060 32228 -17040 32292
rect -16976 32228 -16956 32292
rect -17060 32212 -16956 32228
rect -17060 32148 -17040 32212
rect -16976 32148 -16956 32212
rect -17060 32132 -16956 32148
rect -22672 31772 -22568 32068
rect -28284 31692 -28180 31708
rect -28284 31628 -28264 31692
rect -28200 31628 -28180 31692
rect -28284 31612 -28180 31628
rect -28284 31548 -28264 31612
rect -28200 31548 -28180 31612
rect -28284 31532 -28180 31548
rect -28284 31468 -28264 31532
rect -28200 31468 -28180 31532
rect -28284 31452 -28180 31468
rect -28284 31388 -28264 31452
rect -28200 31388 -28180 31452
rect -28284 31372 -28180 31388
rect -28284 31308 -28264 31372
rect -28200 31308 -28180 31372
rect -28284 31292 -28180 31308
rect -28284 31228 -28264 31292
rect -28200 31228 -28180 31292
rect -28284 31212 -28180 31228
rect -28284 31148 -28264 31212
rect -28200 31148 -28180 31212
rect -28284 31132 -28180 31148
rect -28284 31068 -28264 31132
rect -28200 31068 -28180 31132
rect -28284 31052 -28180 31068
rect -28284 30988 -28264 31052
rect -28200 30988 -28180 31052
rect -28284 30972 -28180 30988
rect -28284 30908 -28264 30972
rect -28200 30908 -28180 30972
rect -28284 30892 -28180 30908
rect -28284 30828 -28264 30892
rect -28200 30828 -28180 30892
rect -28284 30812 -28180 30828
rect -28284 30748 -28264 30812
rect -28200 30748 -28180 30812
rect -28284 30732 -28180 30748
rect -28284 30668 -28264 30732
rect -28200 30668 -28180 30732
rect -28284 30652 -28180 30668
rect -28284 30588 -28264 30652
rect -28200 30588 -28180 30652
rect -28284 30572 -28180 30588
rect -28284 30508 -28264 30572
rect -28200 30508 -28180 30572
rect -28284 30492 -28180 30508
rect -28284 30428 -28264 30492
rect -28200 30428 -28180 30492
rect -28284 30412 -28180 30428
rect -28284 30348 -28264 30412
rect -28200 30348 -28180 30412
rect -28284 30332 -28180 30348
rect -28284 30268 -28264 30332
rect -28200 30268 -28180 30332
rect -28284 30252 -28180 30268
rect -28284 30188 -28264 30252
rect -28200 30188 -28180 30252
rect -28284 30172 -28180 30188
rect -28284 30108 -28264 30172
rect -28200 30108 -28180 30172
rect -28284 30092 -28180 30108
rect -28284 30028 -28264 30092
rect -28200 30028 -28180 30092
rect -28284 30012 -28180 30028
rect -28284 29948 -28264 30012
rect -28200 29948 -28180 30012
rect -28284 29932 -28180 29948
rect -28284 29868 -28264 29932
rect -28200 29868 -28180 29932
rect -28284 29852 -28180 29868
rect -28284 29788 -28264 29852
rect -28200 29788 -28180 29852
rect -28284 29772 -28180 29788
rect -28284 29708 -28264 29772
rect -28200 29708 -28180 29772
rect -28284 29692 -28180 29708
rect -28284 29628 -28264 29692
rect -28200 29628 -28180 29692
rect -28284 29612 -28180 29628
rect -28284 29548 -28264 29612
rect -28200 29548 -28180 29612
rect -28284 29532 -28180 29548
rect -28284 29468 -28264 29532
rect -28200 29468 -28180 29532
rect -28284 29452 -28180 29468
rect -28284 29388 -28264 29452
rect -28200 29388 -28180 29452
rect -28284 29372 -28180 29388
rect -28284 29308 -28264 29372
rect -28200 29308 -28180 29372
rect -28284 29292 -28180 29308
rect -28284 29228 -28264 29292
rect -28200 29228 -28180 29292
rect -28284 29212 -28180 29228
rect -28284 29148 -28264 29212
rect -28200 29148 -28180 29212
rect -28284 29132 -28180 29148
rect -28284 29068 -28264 29132
rect -28200 29068 -28180 29132
rect -28284 29052 -28180 29068
rect -28284 28988 -28264 29052
rect -28200 28988 -28180 29052
rect -28284 28972 -28180 28988
rect -28284 28908 -28264 28972
rect -28200 28908 -28180 28972
rect -28284 28892 -28180 28908
rect -28284 28828 -28264 28892
rect -28200 28828 -28180 28892
rect -28284 28812 -28180 28828
rect -28284 28748 -28264 28812
rect -28200 28748 -28180 28812
rect -28284 28732 -28180 28748
rect -28284 28668 -28264 28732
rect -28200 28668 -28180 28732
rect -28284 28652 -28180 28668
rect -28284 28588 -28264 28652
rect -28200 28588 -28180 28652
rect -28284 28572 -28180 28588
rect -28284 28508 -28264 28572
rect -28200 28508 -28180 28572
rect -28284 28492 -28180 28508
rect -28284 28428 -28264 28492
rect -28200 28428 -28180 28492
rect -28284 28412 -28180 28428
rect -28284 28348 -28264 28412
rect -28200 28348 -28180 28412
rect -28284 28332 -28180 28348
rect -28284 28268 -28264 28332
rect -28200 28268 -28180 28332
rect -28284 28252 -28180 28268
rect -28284 28188 -28264 28252
rect -28200 28188 -28180 28252
rect -28284 28172 -28180 28188
rect -28284 28108 -28264 28172
rect -28200 28108 -28180 28172
rect -28284 28092 -28180 28108
rect -28284 28028 -28264 28092
rect -28200 28028 -28180 28092
rect -28284 28012 -28180 28028
rect -28284 27948 -28264 28012
rect -28200 27948 -28180 28012
rect -28284 27932 -28180 27948
rect -28284 27868 -28264 27932
rect -28200 27868 -28180 27932
rect -28284 27852 -28180 27868
rect -28284 27788 -28264 27852
rect -28200 27788 -28180 27852
rect -28284 27772 -28180 27788
rect -28284 27708 -28264 27772
rect -28200 27708 -28180 27772
rect -28284 27692 -28180 27708
rect -28284 27628 -28264 27692
rect -28200 27628 -28180 27692
rect -28284 27612 -28180 27628
rect -28284 27548 -28264 27612
rect -28200 27548 -28180 27612
rect -28284 27532 -28180 27548
rect -28284 27468 -28264 27532
rect -28200 27468 -28180 27532
rect -28284 27452 -28180 27468
rect -28284 27388 -28264 27452
rect -28200 27388 -28180 27452
rect -28284 27372 -28180 27388
rect -28284 27308 -28264 27372
rect -28200 27308 -28180 27372
rect -28284 27292 -28180 27308
rect -28284 27228 -28264 27292
rect -28200 27228 -28180 27292
rect -28284 27212 -28180 27228
rect -28284 27148 -28264 27212
rect -28200 27148 -28180 27212
rect -28284 27132 -28180 27148
rect -28284 27068 -28264 27132
rect -28200 27068 -28180 27132
rect -28284 27052 -28180 27068
rect -28284 26988 -28264 27052
rect -28200 26988 -28180 27052
rect -28284 26972 -28180 26988
rect -28284 26908 -28264 26972
rect -28200 26908 -28180 26972
rect -28284 26892 -28180 26908
rect -28284 26828 -28264 26892
rect -28200 26828 -28180 26892
rect -28284 26812 -28180 26828
rect -33896 26452 -33792 26748
rect -39085 26372 -34163 26401
rect -39085 21508 -39056 26372
rect -34192 21508 -34163 26372
rect -39085 21479 -34163 21508
rect -33896 26388 -33876 26452
rect -33812 26388 -33792 26452
rect -31064 26401 -30960 26799
rect -28284 26748 -28264 26812
rect -28200 26748 -28180 26812
rect -27861 31692 -22939 31721
rect -27861 26828 -27832 31692
rect -22968 26828 -22939 31692
rect -27861 26799 -22939 26828
rect -22672 31708 -22652 31772
rect -22588 31708 -22568 31772
rect -19840 31721 -19736 32119
rect -17060 32068 -17040 32132
rect -16976 32068 -16956 32132
rect -16637 37012 -11715 37041
rect -16637 32148 -16608 37012
rect -11744 32148 -11715 37012
rect -16637 32119 -11715 32148
rect -11448 37028 -11428 37092
rect -11364 37028 -11344 37092
rect -8616 37041 -8512 37240
rect -5836 37092 -5732 37240
rect -11448 37012 -11344 37028
rect -11448 36948 -11428 37012
rect -11364 36948 -11344 37012
rect -11448 36932 -11344 36948
rect -11448 36868 -11428 36932
rect -11364 36868 -11344 36932
rect -11448 36852 -11344 36868
rect -11448 36788 -11428 36852
rect -11364 36788 -11344 36852
rect -11448 36772 -11344 36788
rect -11448 36708 -11428 36772
rect -11364 36708 -11344 36772
rect -11448 36692 -11344 36708
rect -11448 36628 -11428 36692
rect -11364 36628 -11344 36692
rect -11448 36612 -11344 36628
rect -11448 36548 -11428 36612
rect -11364 36548 -11344 36612
rect -11448 36532 -11344 36548
rect -11448 36468 -11428 36532
rect -11364 36468 -11344 36532
rect -11448 36452 -11344 36468
rect -11448 36388 -11428 36452
rect -11364 36388 -11344 36452
rect -11448 36372 -11344 36388
rect -11448 36308 -11428 36372
rect -11364 36308 -11344 36372
rect -11448 36292 -11344 36308
rect -11448 36228 -11428 36292
rect -11364 36228 -11344 36292
rect -11448 36212 -11344 36228
rect -11448 36148 -11428 36212
rect -11364 36148 -11344 36212
rect -11448 36132 -11344 36148
rect -11448 36068 -11428 36132
rect -11364 36068 -11344 36132
rect -11448 36052 -11344 36068
rect -11448 35988 -11428 36052
rect -11364 35988 -11344 36052
rect -11448 35972 -11344 35988
rect -11448 35908 -11428 35972
rect -11364 35908 -11344 35972
rect -11448 35892 -11344 35908
rect -11448 35828 -11428 35892
rect -11364 35828 -11344 35892
rect -11448 35812 -11344 35828
rect -11448 35748 -11428 35812
rect -11364 35748 -11344 35812
rect -11448 35732 -11344 35748
rect -11448 35668 -11428 35732
rect -11364 35668 -11344 35732
rect -11448 35652 -11344 35668
rect -11448 35588 -11428 35652
rect -11364 35588 -11344 35652
rect -11448 35572 -11344 35588
rect -11448 35508 -11428 35572
rect -11364 35508 -11344 35572
rect -11448 35492 -11344 35508
rect -11448 35428 -11428 35492
rect -11364 35428 -11344 35492
rect -11448 35412 -11344 35428
rect -11448 35348 -11428 35412
rect -11364 35348 -11344 35412
rect -11448 35332 -11344 35348
rect -11448 35268 -11428 35332
rect -11364 35268 -11344 35332
rect -11448 35252 -11344 35268
rect -11448 35188 -11428 35252
rect -11364 35188 -11344 35252
rect -11448 35172 -11344 35188
rect -11448 35108 -11428 35172
rect -11364 35108 -11344 35172
rect -11448 35092 -11344 35108
rect -11448 35028 -11428 35092
rect -11364 35028 -11344 35092
rect -11448 35012 -11344 35028
rect -11448 34948 -11428 35012
rect -11364 34948 -11344 35012
rect -11448 34932 -11344 34948
rect -11448 34868 -11428 34932
rect -11364 34868 -11344 34932
rect -11448 34852 -11344 34868
rect -11448 34788 -11428 34852
rect -11364 34788 -11344 34852
rect -11448 34772 -11344 34788
rect -11448 34708 -11428 34772
rect -11364 34708 -11344 34772
rect -11448 34692 -11344 34708
rect -11448 34628 -11428 34692
rect -11364 34628 -11344 34692
rect -11448 34612 -11344 34628
rect -11448 34548 -11428 34612
rect -11364 34548 -11344 34612
rect -11448 34532 -11344 34548
rect -11448 34468 -11428 34532
rect -11364 34468 -11344 34532
rect -11448 34452 -11344 34468
rect -11448 34388 -11428 34452
rect -11364 34388 -11344 34452
rect -11448 34372 -11344 34388
rect -11448 34308 -11428 34372
rect -11364 34308 -11344 34372
rect -11448 34292 -11344 34308
rect -11448 34228 -11428 34292
rect -11364 34228 -11344 34292
rect -11448 34212 -11344 34228
rect -11448 34148 -11428 34212
rect -11364 34148 -11344 34212
rect -11448 34132 -11344 34148
rect -11448 34068 -11428 34132
rect -11364 34068 -11344 34132
rect -11448 34052 -11344 34068
rect -11448 33988 -11428 34052
rect -11364 33988 -11344 34052
rect -11448 33972 -11344 33988
rect -11448 33908 -11428 33972
rect -11364 33908 -11344 33972
rect -11448 33892 -11344 33908
rect -11448 33828 -11428 33892
rect -11364 33828 -11344 33892
rect -11448 33812 -11344 33828
rect -11448 33748 -11428 33812
rect -11364 33748 -11344 33812
rect -11448 33732 -11344 33748
rect -11448 33668 -11428 33732
rect -11364 33668 -11344 33732
rect -11448 33652 -11344 33668
rect -11448 33588 -11428 33652
rect -11364 33588 -11344 33652
rect -11448 33572 -11344 33588
rect -11448 33508 -11428 33572
rect -11364 33508 -11344 33572
rect -11448 33492 -11344 33508
rect -11448 33428 -11428 33492
rect -11364 33428 -11344 33492
rect -11448 33412 -11344 33428
rect -11448 33348 -11428 33412
rect -11364 33348 -11344 33412
rect -11448 33332 -11344 33348
rect -11448 33268 -11428 33332
rect -11364 33268 -11344 33332
rect -11448 33252 -11344 33268
rect -11448 33188 -11428 33252
rect -11364 33188 -11344 33252
rect -11448 33172 -11344 33188
rect -11448 33108 -11428 33172
rect -11364 33108 -11344 33172
rect -11448 33092 -11344 33108
rect -11448 33028 -11428 33092
rect -11364 33028 -11344 33092
rect -11448 33012 -11344 33028
rect -11448 32948 -11428 33012
rect -11364 32948 -11344 33012
rect -11448 32932 -11344 32948
rect -11448 32868 -11428 32932
rect -11364 32868 -11344 32932
rect -11448 32852 -11344 32868
rect -11448 32788 -11428 32852
rect -11364 32788 -11344 32852
rect -11448 32772 -11344 32788
rect -11448 32708 -11428 32772
rect -11364 32708 -11344 32772
rect -11448 32692 -11344 32708
rect -11448 32628 -11428 32692
rect -11364 32628 -11344 32692
rect -11448 32612 -11344 32628
rect -11448 32548 -11428 32612
rect -11364 32548 -11344 32612
rect -11448 32532 -11344 32548
rect -11448 32468 -11428 32532
rect -11364 32468 -11344 32532
rect -11448 32452 -11344 32468
rect -11448 32388 -11428 32452
rect -11364 32388 -11344 32452
rect -11448 32372 -11344 32388
rect -11448 32308 -11428 32372
rect -11364 32308 -11344 32372
rect -11448 32292 -11344 32308
rect -11448 32228 -11428 32292
rect -11364 32228 -11344 32292
rect -11448 32212 -11344 32228
rect -11448 32148 -11428 32212
rect -11364 32148 -11344 32212
rect -11448 32132 -11344 32148
rect -17060 31772 -16956 32068
rect -22672 31692 -22568 31708
rect -22672 31628 -22652 31692
rect -22588 31628 -22568 31692
rect -22672 31612 -22568 31628
rect -22672 31548 -22652 31612
rect -22588 31548 -22568 31612
rect -22672 31532 -22568 31548
rect -22672 31468 -22652 31532
rect -22588 31468 -22568 31532
rect -22672 31452 -22568 31468
rect -22672 31388 -22652 31452
rect -22588 31388 -22568 31452
rect -22672 31372 -22568 31388
rect -22672 31308 -22652 31372
rect -22588 31308 -22568 31372
rect -22672 31292 -22568 31308
rect -22672 31228 -22652 31292
rect -22588 31228 -22568 31292
rect -22672 31212 -22568 31228
rect -22672 31148 -22652 31212
rect -22588 31148 -22568 31212
rect -22672 31132 -22568 31148
rect -22672 31068 -22652 31132
rect -22588 31068 -22568 31132
rect -22672 31052 -22568 31068
rect -22672 30988 -22652 31052
rect -22588 30988 -22568 31052
rect -22672 30972 -22568 30988
rect -22672 30908 -22652 30972
rect -22588 30908 -22568 30972
rect -22672 30892 -22568 30908
rect -22672 30828 -22652 30892
rect -22588 30828 -22568 30892
rect -22672 30812 -22568 30828
rect -22672 30748 -22652 30812
rect -22588 30748 -22568 30812
rect -22672 30732 -22568 30748
rect -22672 30668 -22652 30732
rect -22588 30668 -22568 30732
rect -22672 30652 -22568 30668
rect -22672 30588 -22652 30652
rect -22588 30588 -22568 30652
rect -22672 30572 -22568 30588
rect -22672 30508 -22652 30572
rect -22588 30508 -22568 30572
rect -22672 30492 -22568 30508
rect -22672 30428 -22652 30492
rect -22588 30428 -22568 30492
rect -22672 30412 -22568 30428
rect -22672 30348 -22652 30412
rect -22588 30348 -22568 30412
rect -22672 30332 -22568 30348
rect -22672 30268 -22652 30332
rect -22588 30268 -22568 30332
rect -22672 30252 -22568 30268
rect -22672 30188 -22652 30252
rect -22588 30188 -22568 30252
rect -22672 30172 -22568 30188
rect -22672 30108 -22652 30172
rect -22588 30108 -22568 30172
rect -22672 30092 -22568 30108
rect -22672 30028 -22652 30092
rect -22588 30028 -22568 30092
rect -22672 30012 -22568 30028
rect -22672 29948 -22652 30012
rect -22588 29948 -22568 30012
rect -22672 29932 -22568 29948
rect -22672 29868 -22652 29932
rect -22588 29868 -22568 29932
rect -22672 29852 -22568 29868
rect -22672 29788 -22652 29852
rect -22588 29788 -22568 29852
rect -22672 29772 -22568 29788
rect -22672 29708 -22652 29772
rect -22588 29708 -22568 29772
rect -22672 29692 -22568 29708
rect -22672 29628 -22652 29692
rect -22588 29628 -22568 29692
rect -22672 29612 -22568 29628
rect -22672 29548 -22652 29612
rect -22588 29548 -22568 29612
rect -22672 29532 -22568 29548
rect -22672 29468 -22652 29532
rect -22588 29468 -22568 29532
rect -22672 29452 -22568 29468
rect -22672 29388 -22652 29452
rect -22588 29388 -22568 29452
rect -22672 29372 -22568 29388
rect -22672 29308 -22652 29372
rect -22588 29308 -22568 29372
rect -22672 29292 -22568 29308
rect -22672 29228 -22652 29292
rect -22588 29228 -22568 29292
rect -22672 29212 -22568 29228
rect -22672 29148 -22652 29212
rect -22588 29148 -22568 29212
rect -22672 29132 -22568 29148
rect -22672 29068 -22652 29132
rect -22588 29068 -22568 29132
rect -22672 29052 -22568 29068
rect -22672 28988 -22652 29052
rect -22588 28988 -22568 29052
rect -22672 28972 -22568 28988
rect -22672 28908 -22652 28972
rect -22588 28908 -22568 28972
rect -22672 28892 -22568 28908
rect -22672 28828 -22652 28892
rect -22588 28828 -22568 28892
rect -22672 28812 -22568 28828
rect -22672 28748 -22652 28812
rect -22588 28748 -22568 28812
rect -22672 28732 -22568 28748
rect -22672 28668 -22652 28732
rect -22588 28668 -22568 28732
rect -22672 28652 -22568 28668
rect -22672 28588 -22652 28652
rect -22588 28588 -22568 28652
rect -22672 28572 -22568 28588
rect -22672 28508 -22652 28572
rect -22588 28508 -22568 28572
rect -22672 28492 -22568 28508
rect -22672 28428 -22652 28492
rect -22588 28428 -22568 28492
rect -22672 28412 -22568 28428
rect -22672 28348 -22652 28412
rect -22588 28348 -22568 28412
rect -22672 28332 -22568 28348
rect -22672 28268 -22652 28332
rect -22588 28268 -22568 28332
rect -22672 28252 -22568 28268
rect -22672 28188 -22652 28252
rect -22588 28188 -22568 28252
rect -22672 28172 -22568 28188
rect -22672 28108 -22652 28172
rect -22588 28108 -22568 28172
rect -22672 28092 -22568 28108
rect -22672 28028 -22652 28092
rect -22588 28028 -22568 28092
rect -22672 28012 -22568 28028
rect -22672 27948 -22652 28012
rect -22588 27948 -22568 28012
rect -22672 27932 -22568 27948
rect -22672 27868 -22652 27932
rect -22588 27868 -22568 27932
rect -22672 27852 -22568 27868
rect -22672 27788 -22652 27852
rect -22588 27788 -22568 27852
rect -22672 27772 -22568 27788
rect -22672 27708 -22652 27772
rect -22588 27708 -22568 27772
rect -22672 27692 -22568 27708
rect -22672 27628 -22652 27692
rect -22588 27628 -22568 27692
rect -22672 27612 -22568 27628
rect -22672 27548 -22652 27612
rect -22588 27548 -22568 27612
rect -22672 27532 -22568 27548
rect -22672 27468 -22652 27532
rect -22588 27468 -22568 27532
rect -22672 27452 -22568 27468
rect -22672 27388 -22652 27452
rect -22588 27388 -22568 27452
rect -22672 27372 -22568 27388
rect -22672 27308 -22652 27372
rect -22588 27308 -22568 27372
rect -22672 27292 -22568 27308
rect -22672 27228 -22652 27292
rect -22588 27228 -22568 27292
rect -22672 27212 -22568 27228
rect -22672 27148 -22652 27212
rect -22588 27148 -22568 27212
rect -22672 27132 -22568 27148
rect -22672 27068 -22652 27132
rect -22588 27068 -22568 27132
rect -22672 27052 -22568 27068
rect -22672 26988 -22652 27052
rect -22588 26988 -22568 27052
rect -22672 26972 -22568 26988
rect -22672 26908 -22652 26972
rect -22588 26908 -22568 26972
rect -22672 26892 -22568 26908
rect -22672 26828 -22652 26892
rect -22588 26828 -22568 26892
rect -22672 26812 -22568 26828
rect -28284 26452 -28180 26748
rect -33896 26372 -33792 26388
rect -33896 26308 -33876 26372
rect -33812 26308 -33792 26372
rect -33896 26292 -33792 26308
rect -33896 26228 -33876 26292
rect -33812 26228 -33792 26292
rect -33896 26212 -33792 26228
rect -33896 26148 -33876 26212
rect -33812 26148 -33792 26212
rect -33896 26132 -33792 26148
rect -33896 26068 -33876 26132
rect -33812 26068 -33792 26132
rect -33896 26052 -33792 26068
rect -33896 25988 -33876 26052
rect -33812 25988 -33792 26052
rect -33896 25972 -33792 25988
rect -33896 25908 -33876 25972
rect -33812 25908 -33792 25972
rect -33896 25892 -33792 25908
rect -33896 25828 -33876 25892
rect -33812 25828 -33792 25892
rect -33896 25812 -33792 25828
rect -33896 25748 -33876 25812
rect -33812 25748 -33792 25812
rect -33896 25732 -33792 25748
rect -33896 25668 -33876 25732
rect -33812 25668 -33792 25732
rect -33896 25652 -33792 25668
rect -33896 25588 -33876 25652
rect -33812 25588 -33792 25652
rect -33896 25572 -33792 25588
rect -33896 25508 -33876 25572
rect -33812 25508 -33792 25572
rect -33896 25492 -33792 25508
rect -33896 25428 -33876 25492
rect -33812 25428 -33792 25492
rect -33896 25412 -33792 25428
rect -33896 25348 -33876 25412
rect -33812 25348 -33792 25412
rect -33896 25332 -33792 25348
rect -33896 25268 -33876 25332
rect -33812 25268 -33792 25332
rect -33896 25252 -33792 25268
rect -33896 25188 -33876 25252
rect -33812 25188 -33792 25252
rect -33896 25172 -33792 25188
rect -33896 25108 -33876 25172
rect -33812 25108 -33792 25172
rect -33896 25092 -33792 25108
rect -33896 25028 -33876 25092
rect -33812 25028 -33792 25092
rect -33896 25012 -33792 25028
rect -33896 24948 -33876 25012
rect -33812 24948 -33792 25012
rect -33896 24932 -33792 24948
rect -33896 24868 -33876 24932
rect -33812 24868 -33792 24932
rect -33896 24852 -33792 24868
rect -33896 24788 -33876 24852
rect -33812 24788 -33792 24852
rect -33896 24772 -33792 24788
rect -33896 24708 -33876 24772
rect -33812 24708 -33792 24772
rect -33896 24692 -33792 24708
rect -33896 24628 -33876 24692
rect -33812 24628 -33792 24692
rect -33896 24612 -33792 24628
rect -33896 24548 -33876 24612
rect -33812 24548 -33792 24612
rect -33896 24532 -33792 24548
rect -33896 24468 -33876 24532
rect -33812 24468 -33792 24532
rect -33896 24452 -33792 24468
rect -33896 24388 -33876 24452
rect -33812 24388 -33792 24452
rect -33896 24372 -33792 24388
rect -33896 24308 -33876 24372
rect -33812 24308 -33792 24372
rect -33896 24292 -33792 24308
rect -33896 24228 -33876 24292
rect -33812 24228 -33792 24292
rect -33896 24212 -33792 24228
rect -33896 24148 -33876 24212
rect -33812 24148 -33792 24212
rect -33896 24132 -33792 24148
rect -33896 24068 -33876 24132
rect -33812 24068 -33792 24132
rect -33896 24052 -33792 24068
rect -33896 23988 -33876 24052
rect -33812 23988 -33792 24052
rect -33896 23972 -33792 23988
rect -33896 23908 -33876 23972
rect -33812 23908 -33792 23972
rect -33896 23892 -33792 23908
rect -33896 23828 -33876 23892
rect -33812 23828 -33792 23892
rect -33896 23812 -33792 23828
rect -33896 23748 -33876 23812
rect -33812 23748 -33792 23812
rect -33896 23732 -33792 23748
rect -33896 23668 -33876 23732
rect -33812 23668 -33792 23732
rect -33896 23652 -33792 23668
rect -33896 23588 -33876 23652
rect -33812 23588 -33792 23652
rect -33896 23572 -33792 23588
rect -33896 23508 -33876 23572
rect -33812 23508 -33792 23572
rect -33896 23492 -33792 23508
rect -33896 23428 -33876 23492
rect -33812 23428 -33792 23492
rect -33896 23412 -33792 23428
rect -33896 23348 -33876 23412
rect -33812 23348 -33792 23412
rect -33896 23332 -33792 23348
rect -33896 23268 -33876 23332
rect -33812 23268 -33792 23332
rect -33896 23252 -33792 23268
rect -33896 23188 -33876 23252
rect -33812 23188 -33792 23252
rect -33896 23172 -33792 23188
rect -33896 23108 -33876 23172
rect -33812 23108 -33792 23172
rect -33896 23092 -33792 23108
rect -33896 23028 -33876 23092
rect -33812 23028 -33792 23092
rect -33896 23012 -33792 23028
rect -33896 22948 -33876 23012
rect -33812 22948 -33792 23012
rect -33896 22932 -33792 22948
rect -33896 22868 -33876 22932
rect -33812 22868 -33792 22932
rect -33896 22852 -33792 22868
rect -33896 22788 -33876 22852
rect -33812 22788 -33792 22852
rect -33896 22772 -33792 22788
rect -33896 22708 -33876 22772
rect -33812 22708 -33792 22772
rect -33896 22692 -33792 22708
rect -33896 22628 -33876 22692
rect -33812 22628 -33792 22692
rect -33896 22612 -33792 22628
rect -33896 22548 -33876 22612
rect -33812 22548 -33792 22612
rect -33896 22532 -33792 22548
rect -33896 22468 -33876 22532
rect -33812 22468 -33792 22532
rect -33896 22452 -33792 22468
rect -33896 22388 -33876 22452
rect -33812 22388 -33792 22452
rect -33896 22372 -33792 22388
rect -33896 22308 -33876 22372
rect -33812 22308 -33792 22372
rect -33896 22292 -33792 22308
rect -33896 22228 -33876 22292
rect -33812 22228 -33792 22292
rect -33896 22212 -33792 22228
rect -33896 22148 -33876 22212
rect -33812 22148 -33792 22212
rect -33896 22132 -33792 22148
rect -33896 22068 -33876 22132
rect -33812 22068 -33792 22132
rect -33896 22052 -33792 22068
rect -33896 21988 -33876 22052
rect -33812 21988 -33792 22052
rect -33896 21972 -33792 21988
rect -33896 21908 -33876 21972
rect -33812 21908 -33792 21972
rect -33896 21892 -33792 21908
rect -33896 21828 -33876 21892
rect -33812 21828 -33792 21892
rect -33896 21812 -33792 21828
rect -33896 21748 -33876 21812
rect -33812 21748 -33792 21812
rect -33896 21732 -33792 21748
rect -33896 21668 -33876 21732
rect -33812 21668 -33792 21732
rect -33896 21652 -33792 21668
rect -33896 21588 -33876 21652
rect -33812 21588 -33792 21652
rect -33896 21572 -33792 21588
rect -33896 21508 -33876 21572
rect -33812 21508 -33792 21572
rect -33896 21492 -33792 21508
rect -36676 21081 -36572 21479
rect -33896 21428 -33876 21492
rect -33812 21428 -33792 21492
rect -33473 26372 -28551 26401
rect -33473 21508 -33444 26372
rect -28580 21508 -28551 26372
rect -33473 21479 -28551 21508
rect -28284 26388 -28264 26452
rect -28200 26388 -28180 26452
rect -25452 26401 -25348 26799
rect -22672 26748 -22652 26812
rect -22588 26748 -22568 26812
rect -22249 31692 -17327 31721
rect -22249 26828 -22220 31692
rect -17356 26828 -17327 31692
rect -22249 26799 -17327 26828
rect -17060 31708 -17040 31772
rect -16976 31708 -16956 31772
rect -14228 31721 -14124 32119
rect -11448 32068 -11428 32132
rect -11364 32068 -11344 32132
rect -11025 37012 -6103 37041
rect -11025 32148 -10996 37012
rect -6132 32148 -6103 37012
rect -11025 32119 -6103 32148
rect -5836 37028 -5816 37092
rect -5752 37028 -5732 37092
rect -3004 37041 -2900 37240
rect -224 37092 -120 37240
rect -5836 37012 -5732 37028
rect -5836 36948 -5816 37012
rect -5752 36948 -5732 37012
rect -5836 36932 -5732 36948
rect -5836 36868 -5816 36932
rect -5752 36868 -5732 36932
rect -5836 36852 -5732 36868
rect -5836 36788 -5816 36852
rect -5752 36788 -5732 36852
rect -5836 36772 -5732 36788
rect -5836 36708 -5816 36772
rect -5752 36708 -5732 36772
rect -5836 36692 -5732 36708
rect -5836 36628 -5816 36692
rect -5752 36628 -5732 36692
rect -5836 36612 -5732 36628
rect -5836 36548 -5816 36612
rect -5752 36548 -5732 36612
rect -5836 36532 -5732 36548
rect -5836 36468 -5816 36532
rect -5752 36468 -5732 36532
rect -5836 36452 -5732 36468
rect -5836 36388 -5816 36452
rect -5752 36388 -5732 36452
rect -5836 36372 -5732 36388
rect -5836 36308 -5816 36372
rect -5752 36308 -5732 36372
rect -5836 36292 -5732 36308
rect -5836 36228 -5816 36292
rect -5752 36228 -5732 36292
rect -5836 36212 -5732 36228
rect -5836 36148 -5816 36212
rect -5752 36148 -5732 36212
rect -5836 36132 -5732 36148
rect -5836 36068 -5816 36132
rect -5752 36068 -5732 36132
rect -5836 36052 -5732 36068
rect -5836 35988 -5816 36052
rect -5752 35988 -5732 36052
rect -5836 35972 -5732 35988
rect -5836 35908 -5816 35972
rect -5752 35908 -5732 35972
rect -5836 35892 -5732 35908
rect -5836 35828 -5816 35892
rect -5752 35828 -5732 35892
rect -5836 35812 -5732 35828
rect -5836 35748 -5816 35812
rect -5752 35748 -5732 35812
rect -5836 35732 -5732 35748
rect -5836 35668 -5816 35732
rect -5752 35668 -5732 35732
rect -5836 35652 -5732 35668
rect -5836 35588 -5816 35652
rect -5752 35588 -5732 35652
rect -5836 35572 -5732 35588
rect -5836 35508 -5816 35572
rect -5752 35508 -5732 35572
rect -5836 35492 -5732 35508
rect -5836 35428 -5816 35492
rect -5752 35428 -5732 35492
rect -5836 35412 -5732 35428
rect -5836 35348 -5816 35412
rect -5752 35348 -5732 35412
rect -5836 35332 -5732 35348
rect -5836 35268 -5816 35332
rect -5752 35268 -5732 35332
rect -5836 35252 -5732 35268
rect -5836 35188 -5816 35252
rect -5752 35188 -5732 35252
rect -5836 35172 -5732 35188
rect -5836 35108 -5816 35172
rect -5752 35108 -5732 35172
rect -5836 35092 -5732 35108
rect -5836 35028 -5816 35092
rect -5752 35028 -5732 35092
rect -5836 35012 -5732 35028
rect -5836 34948 -5816 35012
rect -5752 34948 -5732 35012
rect -5836 34932 -5732 34948
rect -5836 34868 -5816 34932
rect -5752 34868 -5732 34932
rect -5836 34852 -5732 34868
rect -5836 34788 -5816 34852
rect -5752 34788 -5732 34852
rect -5836 34772 -5732 34788
rect -5836 34708 -5816 34772
rect -5752 34708 -5732 34772
rect -5836 34692 -5732 34708
rect -5836 34628 -5816 34692
rect -5752 34628 -5732 34692
rect -5836 34612 -5732 34628
rect -5836 34548 -5816 34612
rect -5752 34548 -5732 34612
rect -5836 34532 -5732 34548
rect -5836 34468 -5816 34532
rect -5752 34468 -5732 34532
rect -5836 34452 -5732 34468
rect -5836 34388 -5816 34452
rect -5752 34388 -5732 34452
rect -5836 34372 -5732 34388
rect -5836 34308 -5816 34372
rect -5752 34308 -5732 34372
rect -5836 34292 -5732 34308
rect -5836 34228 -5816 34292
rect -5752 34228 -5732 34292
rect -5836 34212 -5732 34228
rect -5836 34148 -5816 34212
rect -5752 34148 -5732 34212
rect -5836 34132 -5732 34148
rect -5836 34068 -5816 34132
rect -5752 34068 -5732 34132
rect -5836 34052 -5732 34068
rect -5836 33988 -5816 34052
rect -5752 33988 -5732 34052
rect -5836 33972 -5732 33988
rect -5836 33908 -5816 33972
rect -5752 33908 -5732 33972
rect -5836 33892 -5732 33908
rect -5836 33828 -5816 33892
rect -5752 33828 -5732 33892
rect -5836 33812 -5732 33828
rect -5836 33748 -5816 33812
rect -5752 33748 -5732 33812
rect -5836 33732 -5732 33748
rect -5836 33668 -5816 33732
rect -5752 33668 -5732 33732
rect -5836 33652 -5732 33668
rect -5836 33588 -5816 33652
rect -5752 33588 -5732 33652
rect -5836 33572 -5732 33588
rect -5836 33508 -5816 33572
rect -5752 33508 -5732 33572
rect -5836 33492 -5732 33508
rect -5836 33428 -5816 33492
rect -5752 33428 -5732 33492
rect -5836 33412 -5732 33428
rect -5836 33348 -5816 33412
rect -5752 33348 -5732 33412
rect -5836 33332 -5732 33348
rect -5836 33268 -5816 33332
rect -5752 33268 -5732 33332
rect -5836 33252 -5732 33268
rect -5836 33188 -5816 33252
rect -5752 33188 -5732 33252
rect -5836 33172 -5732 33188
rect -5836 33108 -5816 33172
rect -5752 33108 -5732 33172
rect -5836 33092 -5732 33108
rect -5836 33028 -5816 33092
rect -5752 33028 -5732 33092
rect -5836 33012 -5732 33028
rect -5836 32948 -5816 33012
rect -5752 32948 -5732 33012
rect -5836 32932 -5732 32948
rect -5836 32868 -5816 32932
rect -5752 32868 -5732 32932
rect -5836 32852 -5732 32868
rect -5836 32788 -5816 32852
rect -5752 32788 -5732 32852
rect -5836 32772 -5732 32788
rect -5836 32708 -5816 32772
rect -5752 32708 -5732 32772
rect -5836 32692 -5732 32708
rect -5836 32628 -5816 32692
rect -5752 32628 -5732 32692
rect -5836 32612 -5732 32628
rect -5836 32548 -5816 32612
rect -5752 32548 -5732 32612
rect -5836 32532 -5732 32548
rect -5836 32468 -5816 32532
rect -5752 32468 -5732 32532
rect -5836 32452 -5732 32468
rect -5836 32388 -5816 32452
rect -5752 32388 -5732 32452
rect -5836 32372 -5732 32388
rect -5836 32308 -5816 32372
rect -5752 32308 -5732 32372
rect -5836 32292 -5732 32308
rect -5836 32228 -5816 32292
rect -5752 32228 -5732 32292
rect -5836 32212 -5732 32228
rect -5836 32148 -5816 32212
rect -5752 32148 -5732 32212
rect -5836 32132 -5732 32148
rect -11448 31772 -11344 32068
rect -17060 31692 -16956 31708
rect -17060 31628 -17040 31692
rect -16976 31628 -16956 31692
rect -17060 31612 -16956 31628
rect -17060 31548 -17040 31612
rect -16976 31548 -16956 31612
rect -17060 31532 -16956 31548
rect -17060 31468 -17040 31532
rect -16976 31468 -16956 31532
rect -17060 31452 -16956 31468
rect -17060 31388 -17040 31452
rect -16976 31388 -16956 31452
rect -17060 31372 -16956 31388
rect -17060 31308 -17040 31372
rect -16976 31308 -16956 31372
rect -17060 31292 -16956 31308
rect -17060 31228 -17040 31292
rect -16976 31228 -16956 31292
rect -17060 31212 -16956 31228
rect -17060 31148 -17040 31212
rect -16976 31148 -16956 31212
rect -17060 31132 -16956 31148
rect -17060 31068 -17040 31132
rect -16976 31068 -16956 31132
rect -17060 31052 -16956 31068
rect -17060 30988 -17040 31052
rect -16976 30988 -16956 31052
rect -17060 30972 -16956 30988
rect -17060 30908 -17040 30972
rect -16976 30908 -16956 30972
rect -17060 30892 -16956 30908
rect -17060 30828 -17040 30892
rect -16976 30828 -16956 30892
rect -17060 30812 -16956 30828
rect -17060 30748 -17040 30812
rect -16976 30748 -16956 30812
rect -17060 30732 -16956 30748
rect -17060 30668 -17040 30732
rect -16976 30668 -16956 30732
rect -17060 30652 -16956 30668
rect -17060 30588 -17040 30652
rect -16976 30588 -16956 30652
rect -17060 30572 -16956 30588
rect -17060 30508 -17040 30572
rect -16976 30508 -16956 30572
rect -17060 30492 -16956 30508
rect -17060 30428 -17040 30492
rect -16976 30428 -16956 30492
rect -17060 30412 -16956 30428
rect -17060 30348 -17040 30412
rect -16976 30348 -16956 30412
rect -17060 30332 -16956 30348
rect -17060 30268 -17040 30332
rect -16976 30268 -16956 30332
rect -17060 30252 -16956 30268
rect -17060 30188 -17040 30252
rect -16976 30188 -16956 30252
rect -17060 30172 -16956 30188
rect -17060 30108 -17040 30172
rect -16976 30108 -16956 30172
rect -17060 30092 -16956 30108
rect -17060 30028 -17040 30092
rect -16976 30028 -16956 30092
rect -17060 30012 -16956 30028
rect -17060 29948 -17040 30012
rect -16976 29948 -16956 30012
rect -17060 29932 -16956 29948
rect -17060 29868 -17040 29932
rect -16976 29868 -16956 29932
rect -17060 29852 -16956 29868
rect -17060 29788 -17040 29852
rect -16976 29788 -16956 29852
rect -17060 29772 -16956 29788
rect -17060 29708 -17040 29772
rect -16976 29708 -16956 29772
rect -17060 29692 -16956 29708
rect -17060 29628 -17040 29692
rect -16976 29628 -16956 29692
rect -17060 29612 -16956 29628
rect -17060 29548 -17040 29612
rect -16976 29548 -16956 29612
rect -17060 29532 -16956 29548
rect -17060 29468 -17040 29532
rect -16976 29468 -16956 29532
rect -17060 29452 -16956 29468
rect -17060 29388 -17040 29452
rect -16976 29388 -16956 29452
rect -17060 29372 -16956 29388
rect -17060 29308 -17040 29372
rect -16976 29308 -16956 29372
rect -17060 29292 -16956 29308
rect -17060 29228 -17040 29292
rect -16976 29228 -16956 29292
rect -17060 29212 -16956 29228
rect -17060 29148 -17040 29212
rect -16976 29148 -16956 29212
rect -17060 29132 -16956 29148
rect -17060 29068 -17040 29132
rect -16976 29068 -16956 29132
rect -17060 29052 -16956 29068
rect -17060 28988 -17040 29052
rect -16976 28988 -16956 29052
rect -17060 28972 -16956 28988
rect -17060 28908 -17040 28972
rect -16976 28908 -16956 28972
rect -17060 28892 -16956 28908
rect -17060 28828 -17040 28892
rect -16976 28828 -16956 28892
rect -17060 28812 -16956 28828
rect -17060 28748 -17040 28812
rect -16976 28748 -16956 28812
rect -17060 28732 -16956 28748
rect -17060 28668 -17040 28732
rect -16976 28668 -16956 28732
rect -17060 28652 -16956 28668
rect -17060 28588 -17040 28652
rect -16976 28588 -16956 28652
rect -17060 28572 -16956 28588
rect -17060 28508 -17040 28572
rect -16976 28508 -16956 28572
rect -17060 28492 -16956 28508
rect -17060 28428 -17040 28492
rect -16976 28428 -16956 28492
rect -17060 28412 -16956 28428
rect -17060 28348 -17040 28412
rect -16976 28348 -16956 28412
rect -17060 28332 -16956 28348
rect -17060 28268 -17040 28332
rect -16976 28268 -16956 28332
rect -17060 28252 -16956 28268
rect -17060 28188 -17040 28252
rect -16976 28188 -16956 28252
rect -17060 28172 -16956 28188
rect -17060 28108 -17040 28172
rect -16976 28108 -16956 28172
rect -17060 28092 -16956 28108
rect -17060 28028 -17040 28092
rect -16976 28028 -16956 28092
rect -17060 28012 -16956 28028
rect -17060 27948 -17040 28012
rect -16976 27948 -16956 28012
rect -17060 27932 -16956 27948
rect -17060 27868 -17040 27932
rect -16976 27868 -16956 27932
rect -17060 27852 -16956 27868
rect -17060 27788 -17040 27852
rect -16976 27788 -16956 27852
rect -17060 27772 -16956 27788
rect -17060 27708 -17040 27772
rect -16976 27708 -16956 27772
rect -17060 27692 -16956 27708
rect -17060 27628 -17040 27692
rect -16976 27628 -16956 27692
rect -17060 27612 -16956 27628
rect -17060 27548 -17040 27612
rect -16976 27548 -16956 27612
rect -17060 27532 -16956 27548
rect -17060 27468 -17040 27532
rect -16976 27468 -16956 27532
rect -17060 27452 -16956 27468
rect -17060 27388 -17040 27452
rect -16976 27388 -16956 27452
rect -17060 27372 -16956 27388
rect -17060 27308 -17040 27372
rect -16976 27308 -16956 27372
rect -17060 27292 -16956 27308
rect -17060 27228 -17040 27292
rect -16976 27228 -16956 27292
rect -17060 27212 -16956 27228
rect -17060 27148 -17040 27212
rect -16976 27148 -16956 27212
rect -17060 27132 -16956 27148
rect -17060 27068 -17040 27132
rect -16976 27068 -16956 27132
rect -17060 27052 -16956 27068
rect -17060 26988 -17040 27052
rect -16976 26988 -16956 27052
rect -17060 26972 -16956 26988
rect -17060 26908 -17040 26972
rect -16976 26908 -16956 26972
rect -17060 26892 -16956 26908
rect -17060 26828 -17040 26892
rect -16976 26828 -16956 26892
rect -17060 26812 -16956 26828
rect -22672 26452 -22568 26748
rect -28284 26372 -28180 26388
rect -28284 26308 -28264 26372
rect -28200 26308 -28180 26372
rect -28284 26292 -28180 26308
rect -28284 26228 -28264 26292
rect -28200 26228 -28180 26292
rect -28284 26212 -28180 26228
rect -28284 26148 -28264 26212
rect -28200 26148 -28180 26212
rect -28284 26132 -28180 26148
rect -28284 26068 -28264 26132
rect -28200 26068 -28180 26132
rect -28284 26052 -28180 26068
rect -28284 25988 -28264 26052
rect -28200 25988 -28180 26052
rect -28284 25972 -28180 25988
rect -28284 25908 -28264 25972
rect -28200 25908 -28180 25972
rect -28284 25892 -28180 25908
rect -28284 25828 -28264 25892
rect -28200 25828 -28180 25892
rect -28284 25812 -28180 25828
rect -28284 25748 -28264 25812
rect -28200 25748 -28180 25812
rect -28284 25732 -28180 25748
rect -28284 25668 -28264 25732
rect -28200 25668 -28180 25732
rect -28284 25652 -28180 25668
rect -28284 25588 -28264 25652
rect -28200 25588 -28180 25652
rect -28284 25572 -28180 25588
rect -28284 25508 -28264 25572
rect -28200 25508 -28180 25572
rect -28284 25492 -28180 25508
rect -28284 25428 -28264 25492
rect -28200 25428 -28180 25492
rect -28284 25412 -28180 25428
rect -28284 25348 -28264 25412
rect -28200 25348 -28180 25412
rect -28284 25332 -28180 25348
rect -28284 25268 -28264 25332
rect -28200 25268 -28180 25332
rect -28284 25252 -28180 25268
rect -28284 25188 -28264 25252
rect -28200 25188 -28180 25252
rect -28284 25172 -28180 25188
rect -28284 25108 -28264 25172
rect -28200 25108 -28180 25172
rect -28284 25092 -28180 25108
rect -28284 25028 -28264 25092
rect -28200 25028 -28180 25092
rect -28284 25012 -28180 25028
rect -28284 24948 -28264 25012
rect -28200 24948 -28180 25012
rect -28284 24932 -28180 24948
rect -28284 24868 -28264 24932
rect -28200 24868 -28180 24932
rect -28284 24852 -28180 24868
rect -28284 24788 -28264 24852
rect -28200 24788 -28180 24852
rect -28284 24772 -28180 24788
rect -28284 24708 -28264 24772
rect -28200 24708 -28180 24772
rect -28284 24692 -28180 24708
rect -28284 24628 -28264 24692
rect -28200 24628 -28180 24692
rect -28284 24612 -28180 24628
rect -28284 24548 -28264 24612
rect -28200 24548 -28180 24612
rect -28284 24532 -28180 24548
rect -28284 24468 -28264 24532
rect -28200 24468 -28180 24532
rect -28284 24452 -28180 24468
rect -28284 24388 -28264 24452
rect -28200 24388 -28180 24452
rect -28284 24372 -28180 24388
rect -28284 24308 -28264 24372
rect -28200 24308 -28180 24372
rect -28284 24292 -28180 24308
rect -28284 24228 -28264 24292
rect -28200 24228 -28180 24292
rect -28284 24212 -28180 24228
rect -28284 24148 -28264 24212
rect -28200 24148 -28180 24212
rect -28284 24132 -28180 24148
rect -28284 24068 -28264 24132
rect -28200 24068 -28180 24132
rect -28284 24052 -28180 24068
rect -28284 23988 -28264 24052
rect -28200 23988 -28180 24052
rect -28284 23972 -28180 23988
rect -28284 23908 -28264 23972
rect -28200 23908 -28180 23972
rect -28284 23892 -28180 23908
rect -28284 23828 -28264 23892
rect -28200 23828 -28180 23892
rect -28284 23812 -28180 23828
rect -28284 23748 -28264 23812
rect -28200 23748 -28180 23812
rect -28284 23732 -28180 23748
rect -28284 23668 -28264 23732
rect -28200 23668 -28180 23732
rect -28284 23652 -28180 23668
rect -28284 23588 -28264 23652
rect -28200 23588 -28180 23652
rect -28284 23572 -28180 23588
rect -28284 23508 -28264 23572
rect -28200 23508 -28180 23572
rect -28284 23492 -28180 23508
rect -28284 23428 -28264 23492
rect -28200 23428 -28180 23492
rect -28284 23412 -28180 23428
rect -28284 23348 -28264 23412
rect -28200 23348 -28180 23412
rect -28284 23332 -28180 23348
rect -28284 23268 -28264 23332
rect -28200 23268 -28180 23332
rect -28284 23252 -28180 23268
rect -28284 23188 -28264 23252
rect -28200 23188 -28180 23252
rect -28284 23172 -28180 23188
rect -28284 23108 -28264 23172
rect -28200 23108 -28180 23172
rect -28284 23092 -28180 23108
rect -28284 23028 -28264 23092
rect -28200 23028 -28180 23092
rect -28284 23012 -28180 23028
rect -28284 22948 -28264 23012
rect -28200 22948 -28180 23012
rect -28284 22932 -28180 22948
rect -28284 22868 -28264 22932
rect -28200 22868 -28180 22932
rect -28284 22852 -28180 22868
rect -28284 22788 -28264 22852
rect -28200 22788 -28180 22852
rect -28284 22772 -28180 22788
rect -28284 22708 -28264 22772
rect -28200 22708 -28180 22772
rect -28284 22692 -28180 22708
rect -28284 22628 -28264 22692
rect -28200 22628 -28180 22692
rect -28284 22612 -28180 22628
rect -28284 22548 -28264 22612
rect -28200 22548 -28180 22612
rect -28284 22532 -28180 22548
rect -28284 22468 -28264 22532
rect -28200 22468 -28180 22532
rect -28284 22452 -28180 22468
rect -28284 22388 -28264 22452
rect -28200 22388 -28180 22452
rect -28284 22372 -28180 22388
rect -28284 22308 -28264 22372
rect -28200 22308 -28180 22372
rect -28284 22292 -28180 22308
rect -28284 22228 -28264 22292
rect -28200 22228 -28180 22292
rect -28284 22212 -28180 22228
rect -28284 22148 -28264 22212
rect -28200 22148 -28180 22212
rect -28284 22132 -28180 22148
rect -28284 22068 -28264 22132
rect -28200 22068 -28180 22132
rect -28284 22052 -28180 22068
rect -28284 21988 -28264 22052
rect -28200 21988 -28180 22052
rect -28284 21972 -28180 21988
rect -28284 21908 -28264 21972
rect -28200 21908 -28180 21972
rect -28284 21892 -28180 21908
rect -28284 21828 -28264 21892
rect -28200 21828 -28180 21892
rect -28284 21812 -28180 21828
rect -28284 21748 -28264 21812
rect -28200 21748 -28180 21812
rect -28284 21732 -28180 21748
rect -28284 21668 -28264 21732
rect -28200 21668 -28180 21732
rect -28284 21652 -28180 21668
rect -28284 21588 -28264 21652
rect -28200 21588 -28180 21652
rect -28284 21572 -28180 21588
rect -28284 21508 -28264 21572
rect -28200 21508 -28180 21572
rect -28284 21492 -28180 21508
rect -33896 21132 -33792 21428
rect -39085 21052 -34163 21081
rect -39085 16188 -39056 21052
rect -34192 16188 -34163 21052
rect -39085 16159 -34163 16188
rect -33896 21068 -33876 21132
rect -33812 21068 -33792 21132
rect -31064 21081 -30960 21479
rect -28284 21428 -28264 21492
rect -28200 21428 -28180 21492
rect -27861 26372 -22939 26401
rect -27861 21508 -27832 26372
rect -22968 21508 -22939 26372
rect -27861 21479 -22939 21508
rect -22672 26388 -22652 26452
rect -22588 26388 -22568 26452
rect -19840 26401 -19736 26799
rect -17060 26748 -17040 26812
rect -16976 26748 -16956 26812
rect -16637 31692 -11715 31721
rect -16637 26828 -16608 31692
rect -11744 26828 -11715 31692
rect -16637 26799 -11715 26828
rect -11448 31708 -11428 31772
rect -11364 31708 -11344 31772
rect -8616 31721 -8512 32119
rect -5836 32068 -5816 32132
rect -5752 32068 -5732 32132
rect -5413 37012 -491 37041
rect -5413 32148 -5384 37012
rect -520 32148 -491 37012
rect -5413 32119 -491 32148
rect -224 37028 -204 37092
rect -140 37028 -120 37092
rect 2608 37041 2712 37240
rect 5388 37092 5492 37240
rect -224 37012 -120 37028
rect -224 36948 -204 37012
rect -140 36948 -120 37012
rect -224 36932 -120 36948
rect -224 36868 -204 36932
rect -140 36868 -120 36932
rect -224 36852 -120 36868
rect -224 36788 -204 36852
rect -140 36788 -120 36852
rect -224 36772 -120 36788
rect -224 36708 -204 36772
rect -140 36708 -120 36772
rect -224 36692 -120 36708
rect -224 36628 -204 36692
rect -140 36628 -120 36692
rect -224 36612 -120 36628
rect -224 36548 -204 36612
rect -140 36548 -120 36612
rect -224 36532 -120 36548
rect -224 36468 -204 36532
rect -140 36468 -120 36532
rect -224 36452 -120 36468
rect -224 36388 -204 36452
rect -140 36388 -120 36452
rect -224 36372 -120 36388
rect -224 36308 -204 36372
rect -140 36308 -120 36372
rect -224 36292 -120 36308
rect -224 36228 -204 36292
rect -140 36228 -120 36292
rect -224 36212 -120 36228
rect -224 36148 -204 36212
rect -140 36148 -120 36212
rect -224 36132 -120 36148
rect -224 36068 -204 36132
rect -140 36068 -120 36132
rect -224 36052 -120 36068
rect -224 35988 -204 36052
rect -140 35988 -120 36052
rect -224 35972 -120 35988
rect -224 35908 -204 35972
rect -140 35908 -120 35972
rect -224 35892 -120 35908
rect -224 35828 -204 35892
rect -140 35828 -120 35892
rect -224 35812 -120 35828
rect -224 35748 -204 35812
rect -140 35748 -120 35812
rect -224 35732 -120 35748
rect -224 35668 -204 35732
rect -140 35668 -120 35732
rect -224 35652 -120 35668
rect -224 35588 -204 35652
rect -140 35588 -120 35652
rect -224 35572 -120 35588
rect -224 35508 -204 35572
rect -140 35508 -120 35572
rect -224 35492 -120 35508
rect -224 35428 -204 35492
rect -140 35428 -120 35492
rect -224 35412 -120 35428
rect -224 35348 -204 35412
rect -140 35348 -120 35412
rect -224 35332 -120 35348
rect -224 35268 -204 35332
rect -140 35268 -120 35332
rect -224 35252 -120 35268
rect -224 35188 -204 35252
rect -140 35188 -120 35252
rect -224 35172 -120 35188
rect -224 35108 -204 35172
rect -140 35108 -120 35172
rect -224 35092 -120 35108
rect -224 35028 -204 35092
rect -140 35028 -120 35092
rect -224 35012 -120 35028
rect -224 34948 -204 35012
rect -140 34948 -120 35012
rect -224 34932 -120 34948
rect -224 34868 -204 34932
rect -140 34868 -120 34932
rect -224 34852 -120 34868
rect -224 34788 -204 34852
rect -140 34788 -120 34852
rect -224 34772 -120 34788
rect -224 34708 -204 34772
rect -140 34708 -120 34772
rect -224 34692 -120 34708
rect -224 34628 -204 34692
rect -140 34628 -120 34692
rect -224 34612 -120 34628
rect -224 34548 -204 34612
rect -140 34548 -120 34612
rect -224 34532 -120 34548
rect -224 34468 -204 34532
rect -140 34468 -120 34532
rect -224 34452 -120 34468
rect -224 34388 -204 34452
rect -140 34388 -120 34452
rect -224 34372 -120 34388
rect -224 34308 -204 34372
rect -140 34308 -120 34372
rect -224 34292 -120 34308
rect -224 34228 -204 34292
rect -140 34228 -120 34292
rect -224 34212 -120 34228
rect -224 34148 -204 34212
rect -140 34148 -120 34212
rect -224 34132 -120 34148
rect -224 34068 -204 34132
rect -140 34068 -120 34132
rect -224 34052 -120 34068
rect -224 33988 -204 34052
rect -140 33988 -120 34052
rect -224 33972 -120 33988
rect -224 33908 -204 33972
rect -140 33908 -120 33972
rect -224 33892 -120 33908
rect -224 33828 -204 33892
rect -140 33828 -120 33892
rect -224 33812 -120 33828
rect -224 33748 -204 33812
rect -140 33748 -120 33812
rect -224 33732 -120 33748
rect -224 33668 -204 33732
rect -140 33668 -120 33732
rect -224 33652 -120 33668
rect -224 33588 -204 33652
rect -140 33588 -120 33652
rect -224 33572 -120 33588
rect -224 33508 -204 33572
rect -140 33508 -120 33572
rect -224 33492 -120 33508
rect -224 33428 -204 33492
rect -140 33428 -120 33492
rect -224 33412 -120 33428
rect -224 33348 -204 33412
rect -140 33348 -120 33412
rect -224 33332 -120 33348
rect -224 33268 -204 33332
rect -140 33268 -120 33332
rect -224 33252 -120 33268
rect -224 33188 -204 33252
rect -140 33188 -120 33252
rect -224 33172 -120 33188
rect -224 33108 -204 33172
rect -140 33108 -120 33172
rect -224 33092 -120 33108
rect -224 33028 -204 33092
rect -140 33028 -120 33092
rect -224 33012 -120 33028
rect -224 32948 -204 33012
rect -140 32948 -120 33012
rect -224 32932 -120 32948
rect -224 32868 -204 32932
rect -140 32868 -120 32932
rect -224 32852 -120 32868
rect -224 32788 -204 32852
rect -140 32788 -120 32852
rect -224 32772 -120 32788
rect -224 32708 -204 32772
rect -140 32708 -120 32772
rect -224 32692 -120 32708
rect -224 32628 -204 32692
rect -140 32628 -120 32692
rect -224 32612 -120 32628
rect -224 32548 -204 32612
rect -140 32548 -120 32612
rect -224 32532 -120 32548
rect -224 32468 -204 32532
rect -140 32468 -120 32532
rect -224 32452 -120 32468
rect -224 32388 -204 32452
rect -140 32388 -120 32452
rect -224 32372 -120 32388
rect -224 32308 -204 32372
rect -140 32308 -120 32372
rect -224 32292 -120 32308
rect -224 32228 -204 32292
rect -140 32228 -120 32292
rect -224 32212 -120 32228
rect -224 32148 -204 32212
rect -140 32148 -120 32212
rect -224 32132 -120 32148
rect -5836 31772 -5732 32068
rect -11448 31692 -11344 31708
rect -11448 31628 -11428 31692
rect -11364 31628 -11344 31692
rect -11448 31612 -11344 31628
rect -11448 31548 -11428 31612
rect -11364 31548 -11344 31612
rect -11448 31532 -11344 31548
rect -11448 31468 -11428 31532
rect -11364 31468 -11344 31532
rect -11448 31452 -11344 31468
rect -11448 31388 -11428 31452
rect -11364 31388 -11344 31452
rect -11448 31372 -11344 31388
rect -11448 31308 -11428 31372
rect -11364 31308 -11344 31372
rect -11448 31292 -11344 31308
rect -11448 31228 -11428 31292
rect -11364 31228 -11344 31292
rect -11448 31212 -11344 31228
rect -11448 31148 -11428 31212
rect -11364 31148 -11344 31212
rect -11448 31132 -11344 31148
rect -11448 31068 -11428 31132
rect -11364 31068 -11344 31132
rect -11448 31052 -11344 31068
rect -11448 30988 -11428 31052
rect -11364 30988 -11344 31052
rect -11448 30972 -11344 30988
rect -11448 30908 -11428 30972
rect -11364 30908 -11344 30972
rect -11448 30892 -11344 30908
rect -11448 30828 -11428 30892
rect -11364 30828 -11344 30892
rect -11448 30812 -11344 30828
rect -11448 30748 -11428 30812
rect -11364 30748 -11344 30812
rect -11448 30732 -11344 30748
rect -11448 30668 -11428 30732
rect -11364 30668 -11344 30732
rect -11448 30652 -11344 30668
rect -11448 30588 -11428 30652
rect -11364 30588 -11344 30652
rect -11448 30572 -11344 30588
rect -11448 30508 -11428 30572
rect -11364 30508 -11344 30572
rect -11448 30492 -11344 30508
rect -11448 30428 -11428 30492
rect -11364 30428 -11344 30492
rect -11448 30412 -11344 30428
rect -11448 30348 -11428 30412
rect -11364 30348 -11344 30412
rect -11448 30332 -11344 30348
rect -11448 30268 -11428 30332
rect -11364 30268 -11344 30332
rect -11448 30252 -11344 30268
rect -11448 30188 -11428 30252
rect -11364 30188 -11344 30252
rect -11448 30172 -11344 30188
rect -11448 30108 -11428 30172
rect -11364 30108 -11344 30172
rect -11448 30092 -11344 30108
rect -11448 30028 -11428 30092
rect -11364 30028 -11344 30092
rect -11448 30012 -11344 30028
rect -11448 29948 -11428 30012
rect -11364 29948 -11344 30012
rect -11448 29932 -11344 29948
rect -11448 29868 -11428 29932
rect -11364 29868 -11344 29932
rect -11448 29852 -11344 29868
rect -11448 29788 -11428 29852
rect -11364 29788 -11344 29852
rect -11448 29772 -11344 29788
rect -11448 29708 -11428 29772
rect -11364 29708 -11344 29772
rect -11448 29692 -11344 29708
rect -11448 29628 -11428 29692
rect -11364 29628 -11344 29692
rect -11448 29612 -11344 29628
rect -11448 29548 -11428 29612
rect -11364 29548 -11344 29612
rect -11448 29532 -11344 29548
rect -11448 29468 -11428 29532
rect -11364 29468 -11344 29532
rect -11448 29452 -11344 29468
rect -11448 29388 -11428 29452
rect -11364 29388 -11344 29452
rect -11448 29372 -11344 29388
rect -11448 29308 -11428 29372
rect -11364 29308 -11344 29372
rect -11448 29292 -11344 29308
rect -11448 29228 -11428 29292
rect -11364 29228 -11344 29292
rect -11448 29212 -11344 29228
rect -11448 29148 -11428 29212
rect -11364 29148 -11344 29212
rect -11448 29132 -11344 29148
rect -11448 29068 -11428 29132
rect -11364 29068 -11344 29132
rect -11448 29052 -11344 29068
rect -11448 28988 -11428 29052
rect -11364 28988 -11344 29052
rect -11448 28972 -11344 28988
rect -11448 28908 -11428 28972
rect -11364 28908 -11344 28972
rect -11448 28892 -11344 28908
rect -11448 28828 -11428 28892
rect -11364 28828 -11344 28892
rect -11448 28812 -11344 28828
rect -11448 28748 -11428 28812
rect -11364 28748 -11344 28812
rect -11448 28732 -11344 28748
rect -11448 28668 -11428 28732
rect -11364 28668 -11344 28732
rect -11448 28652 -11344 28668
rect -11448 28588 -11428 28652
rect -11364 28588 -11344 28652
rect -11448 28572 -11344 28588
rect -11448 28508 -11428 28572
rect -11364 28508 -11344 28572
rect -11448 28492 -11344 28508
rect -11448 28428 -11428 28492
rect -11364 28428 -11344 28492
rect -11448 28412 -11344 28428
rect -11448 28348 -11428 28412
rect -11364 28348 -11344 28412
rect -11448 28332 -11344 28348
rect -11448 28268 -11428 28332
rect -11364 28268 -11344 28332
rect -11448 28252 -11344 28268
rect -11448 28188 -11428 28252
rect -11364 28188 -11344 28252
rect -11448 28172 -11344 28188
rect -11448 28108 -11428 28172
rect -11364 28108 -11344 28172
rect -11448 28092 -11344 28108
rect -11448 28028 -11428 28092
rect -11364 28028 -11344 28092
rect -11448 28012 -11344 28028
rect -11448 27948 -11428 28012
rect -11364 27948 -11344 28012
rect -11448 27932 -11344 27948
rect -11448 27868 -11428 27932
rect -11364 27868 -11344 27932
rect -11448 27852 -11344 27868
rect -11448 27788 -11428 27852
rect -11364 27788 -11344 27852
rect -11448 27772 -11344 27788
rect -11448 27708 -11428 27772
rect -11364 27708 -11344 27772
rect -11448 27692 -11344 27708
rect -11448 27628 -11428 27692
rect -11364 27628 -11344 27692
rect -11448 27612 -11344 27628
rect -11448 27548 -11428 27612
rect -11364 27548 -11344 27612
rect -11448 27532 -11344 27548
rect -11448 27468 -11428 27532
rect -11364 27468 -11344 27532
rect -11448 27452 -11344 27468
rect -11448 27388 -11428 27452
rect -11364 27388 -11344 27452
rect -11448 27372 -11344 27388
rect -11448 27308 -11428 27372
rect -11364 27308 -11344 27372
rect -11448 27292 -11344 27308
rect -11448 27228 -11428 27292
rect -11364 27228 -11344 27292
rect -11448 27212 -11344 27228
rect -11448 27148 -11428 27212
rect -11364 27148 -11344 27212
rect -11448 27132 -11344 27148
rect -11448 27068 -11428 27132
rect -11364 27068 -11344 27132
rect -11448 27052 -11344 27068
rect -11448 26988 -11428 27052
rect -11364 26988 -11344 27052
rect -11448 26972 -11344 26988
rect -11448 26908 -11428 26972
rect -11364 26908 -11344 26972
rect -11448 26892 -11344 26908
rect -11448 26828 -11428 26892
rect -11364 26828 -11344 26892
rect -11448 26812 -11344 26828
rect -17060 26452 -16956 26748
rect -22672 26372 -22568 26388
rect -22672 26308 -22652 26372
rect -22588 26308 -22568 26372
rect -22672 26292 -22568 26308
rect -22672 26228 -22652 26292
rect -22588 26228 -22568 26292
rect -22672 26212 -22568 26228
rect -22672 26148 -22652 26212
rect -22588 26148 -22568 26212
rect -22672 26132 -22568 26148
rect -22672 26068 -22652 26132
rect -22588 26068 -22568 26132
rect -22672 26052 -22568 26068
rect -22672 25988 -22652 26052
rect -22588 25988 -22568 26052
rect -22672 25972 -22568 25988
rect -22672 25908 -22652 25972
rect -22588 25908 -22568 25972
rect -22672 25892 -22568 25908
rect -22672 25828 -22652 25892
rect -22588 25828 -22568 25892
rect -22672 25812 -22568 25828
rect -22672 25748 -22652 25812
rect -22588 25748 -22568 25812
rect -22672 25732 -22568 25748
rect -22672 25668 -22652 25732
rect -22588 25668 -22568 25732
rect -22672 25652 -22568 25668
rect -22672 25588 -22652 25652
rect -22588 25588 -22568 25652
rect -22672 25572 -22568 25588
rect -22672 25508 -22652 25572
rect -22588 25508 -22568 25572
rect -22672 25492 -22568 25508
rect -22672 25428 -22652 25492
rect -22588 25428 -22568 25492
rect -22672 25412 -22568 25428
rect -22672 25348 -22652 25412
rect -22588 25348 -22568 25412
rect -22672 25332 -22568 25348
rect -22672 25268 -22652 25332
rect -22588 25268 -22568 25332
rect -22672 25252 -22568 25268
rect -22672 25188 -22652 25252
rect -22588 25188 -22568 25252
rect -22672 25172 -22568 25188
rect -22672 25108 -22652 25172
rect -22588 25108 -22568 25172
rect -22672 25092 -22568 25108
rect -22672 25028 -22652 25092
rect -22588 25028 -22568 25092
rect -22672 25012 -22568 25028
rect -22672 24948 -22652 25012
rect -22588 24948 -22568 25012
rect -22672 24932 -22568 24948
rect -22672 24868 -22652 24932
rect -22588 24868 -22568 24932
rect -22672 24852 -22568 24868
rect -22672 24788 -22652 24852
rect -22588 24788 -22568 24852
rect -22672 24772 -22568 24788
rect -22672 24708 -22652 24772
rect -22588 24708 -22568 24772
rect -22672 24692 -22568 24708
rect -22672 24628 -22652 24692
rect -22588 24628 -22568 24692
rect -22672 24612 -22568 24628
rect -22672 24548 -22652 24612
rect -22588 24548 -22568 24612
rect -22672 24532 -22568 24548
rect -22672 24468 -22652 24532
rect -22588 24468 -22568 24532
rect -22672 24452 -22568 24468
rect -22672 24388 -22652 24452
rect -22588 24388 -22568 24452
rect -22672 24372 -22568 24388
rect -22672 24308 -22652 24372
rect -22588 24308 -22568 24372
rect -22672 24292 -22568 24308
rect -22672 24228 -22652 24292
rect -22588 24228 -22568 24292
rect -22672 24212 -22568 24228
rect -22672 24148 -22652 24212
rect -22588 24148 -22568 24212
rect -22672 24132 -22568 24148
rect -22672 24068 -22652 24132
rect -22588 24068 -22568 24132
rect -22672 24052 -22568 24068
rect -22672 23988 -22652 24052
rect -22588 23988 -22568 24052
rect -22672 23972 -22568 23988
rect -22672 23908 -22652 23972
rect -22588 23908 -22568 23972
rect -22672 23892 -22568 23908
rect -22672 23828 -22652 23892
rect -22588 23828 -22568 23892
rect -22672 23812 -22568 23828
rect -22672 23748 -22652 23812
rect -22588 23748 -22568 23812
rect -22672 23732 -22568 23748
rect -22672 23668 -22652 23732
rect -22588 23668 -22568 23732
rect -22672 23652 -22568 23668
rect -22672 23588 -22652 23652
rect -22588 23588 -22568 23652
rect -22672 23572 -22568 23588
rect -22672 23508 -22652 23572
rect -22588 23508 -22568 23572
rect -22672 23492 -22568 23508
rect -22672 23428 -22652 23492
rect -22588 23428 -22568 23492
rect -22672 23412 -22568 23428
rect -22672 23348 -22652 23412
rect -22588 23348 -22568 23412
rect -22672 23332 -22568 23348
rect -22672 23268 -22652 23332
rect -22588 23268 -22568 23332
rect -22672 23252 -22568 23268
rect -22672 23188 -22652 23252
rect -22588 23188 -22568 23252
rect -22672 23172 -22568 23188
rect -22672 23108 -22652 23172
rect -22588 23108 -22568 23172
rect -22672 23092 -22568 23108
rect -22672 23028 -22652 23092
rect -22588 23028 -22568 23092
rect -22672 23012 -22568 23028
rect -22672 22948 -22652 23012
rect -22588 22948 -22568 23012
rect -22672 22932 -22568 22948
rect -22672 22868 -22652 22932
rect -22588 22868 -22568 22932
rect -22672 22852 -22568 22868
rect -22672 22788 -22652 22852
rect -22588 22788 -22568 22852
rect -22672 22772 -22568 22788
rect -22672 22708 -22652 22772
rect -22588 22708 -22568 22772
rect -22672 22692 -22568 22708
rect -22672 22628 -22652 22692
rect -22588 22628 -22568 22692
rect -22672 22612 -22568 22628
rect -22672 22548 -22652 22612
rect -22588 22548 -22568 22612
rect -22672 22532 -22568 22548
rect -22672 22468 -22652 22532
rect -22588 22468 -22568 22532
rect -22672 22452 -22568 22468
rect -22672 22388 -22652 22452
rect -22588 22388 -22568 22452
rect -22672 22372 -22568 22388
rect -22672 22308 -22652 22372
rect -22588 22308 -22568 22372
rect -22672 22292 -22568 22308
rect -22672 22228 -22652 22292
rect -22588 22228 -22568 22292
rect -22672 22212 -22568 22228
rect -22672 22148 -22652 22212
rect -22588 22148 -22568 22212
rect -22672 22132 -22568 22148
rect -22672 22068 -22652 22132
rect -22588 22068 -22568 22132
rect -22672 22052 -22568 22068
rect -22672 21988 -22652 22052
rect -22588 21988 -22568 22052
rect -22672 21972 -22568 21988
rect -22672 21908 -22652 21972
rect -22588 21908 -22568 21972
rect -22672 21892 -22568 21908
rect -22672 21828 -22652 21892
rect -22588 21828 -22568 21892
rect -22672 21812 -22568 21828
rect -22672 21748 -22652 21812
rect -22588 21748 -22568 21812
rect -22672 21732 -22568 21748
rect -22672 21668 -22652 21732
rect -22588 21668 -22568 21732
rect -22672 21652 -22568 21668
rect -22672 21588 -22652 21652
rect -22588 21588 -22568 21652
rect -22672 21572 -22568 21588
rect -22672 21508 -22652 21572
rect -22588 21508 -22568 21572
rect -22672 21492 -22568 21508
rect -28284 21132 -28180 21428
rect -33896 21052 -33792 21068
rect -33896 20988 -33876 21052
rect -33812 20988 -33792 21052
rect -33896 20972 -33792 20988
rect -33896 20908 -33876 20972
rect -33812 20908 -33792 20972
rect -33896 20892 -33792 20908
rect -33896 20828 -33876 20892
rect -33812 20828 -33792 20892
rect -33896 20812 -33792 20828
rect -33896 20748 -33876 20812
rect -33812 20748 -33792 20812
rect -33896 20732 -33792 20748
rect -33896 20668 -33876 20732
rect -33812 20668 -33792 20732
rect -33896 20652 -33792 20668
rect -33896 20588 -33876 20652
rect -33812 20588 -33792 20652
rect -33896 20572 -33792 20588
rect -33896 20508 -33876 20572
rect -33812 20508 -33792 20572
rect -33896 20492 -33792 20508
rect -33896 20428 -33876 20492
rect -33812 20428 -33792 20492
rect -33896 20412 -33792 20428
rect -33896 20348 -33876 20412
rect -33812 20348 -33792 20412
rect -33896 20332 -33792 20348
rect -33896 20268 -33876 20332
rect -33812 20268 -33792 20332
rect -33896 20252 -33792 20268
rect -33896 20188 -33876 20252
rect -33812 20188 -33792 20252
rect -33896 20172 -33792 20188
rect -33896 20108 -33876 20172
rect -33812 20108 -33792 20172
rect -33896 20092 -33792 20108
rect -33896 20028 -33876 20092
rect -33812 20028 -33792 20092
rect -33896 20012 -33792 20028
rect -33896 19948 -33876 20012
rect -33812 19948 -33792 20012
rect -33896 19932 -33792 19948
rect -33896 19868 -33876 19932
rect -33812 19868 -33792 19932
rect -33896 19852 -33792 19868
rect -33896 19788 -33876 19852
rect -33812 19788 -33792 19852
rect -33896 19772 -33792 19788
rect -33896 19708 -33876 19772
rect -33812 19708 -33792 19772
rect -33896 19692 -33792 19708
rect -33896 19628 -33876 19692
rect -33812 19628 -33792 19692
rect -33896 19612 -33792 19628
rect -33896 19548 -33876 19612
rect -33812 19548 -33792 19612
rect -33896 19532 -33792 19548
rect -33896 19468 -33876 19532
rect -33812 19468 -33792 19532
rect -33896 19452 -33792 19468
rect -33896 19388 -33876 19452
rect -33812 19388 -33792 19452
rect -33896 19372 -33792 19388
rect -33896 19308 -33876 19372
rect -33812 19308 -33792 19372
rect -33896 19292 -33792 19308
rect -33896 19228 -33876 19292
rect -33812 19228 -33792 19292
rect -33896 19212 -33792 19228
rect -33896 19148 -33876 19212
rect -33812 19148 -33792 19212
rect -33896 19132 -33792 19148
rect -33896 19068 -33876 19132
rect -33812 19068 -33792 19132
rect -33896 19052 -33792 19068
rect -33896 18988 -33876 19052
rect -33812 18988 -33792 19052
rect -33896 18972 -33792 18988
rect -33896 18908 -33876 18972
rect -33812 18908 -33792 18972
rect -33896 18892 -33792 18908
rect -33896 18828 -33876 18892
rect -33812 18828 -33792 18892
rect -33896 18812 -33792 18828
rect -33896 18748 -33876 18812
rect -33812 18748 -33792 18812
rect -33896 18732 -33792 18748
rect -33896 18668 -33876 18732
rect -33812 18668 -33792 18732
rect -33896 18652 -33792 18668
rect -33896 18588 -33876 18652
rect -33812 18588 -33792 18652
rect -33896 18572 -33792 18588
rect -33896 18508 -33876 18572
rect -33812 18508 -33792 18572
rect -33896 18492 -33792 18508
rect -33896 18428 -33876 18492
rect -33812 18428 -33792 18492
rect -33896 18412 -33792 18428
rect -33896 18348 -33876 18412
rect -33812 18348 -33792 18412
rect -33896 18332 -33792 18348
rect -33896 18268 -33876 18332
rect -33812 18268 -33792 18332
rect -33896 18252 -33792 18268
rect -33896 18188 -33876 18252
rect -33812 18188 -33792 18252
rect -33896 18172 -33792 18188
rect -33896 18108 -33876 18172
rect -33812 18108 -33792 18172
rect -33896 18092 -33792 18108
rect -33896 18028 -33876 18092
rect -33812 18028 -33792 18092
rect -33896 18012 -33792 18028
rect -33896 17948 -33876 18012
rect -33812 17948 -33792 18012
rect -33896 17932 -33792 17948
rect -33896 17868 -33876 17932
rect -33812 17868 -33792 17932
rect -33896 17852 -33792 17868
rect -33896 17788 -33876 17852
rect -33812 17788 -33792 17852
rect -33896 17772 -33792 17788
rect -33896 17708 -33876 17772
rect -33812 17708 -33792 17772
rect -33896 17692 -33792 17708
rect -33896 17628 -33876 17692
rect -33812 17628 -33792 17692
rect -33896 17612 -33792 17628
rect -33896 17548 -33876 17612
rect -33812 17548 -33792 17612
rect -33896 17532 -33792 17548
rect -33896 17468 -33876 17532
rect -33812 17468 -33792 17532
rect -33896 17452 -33792 17468
rect -33896 17388 -33876 17452
rect -33812 17388 -33792 17452
rect -33896 17372 -33792 17388
rect -33896 17308 -33876 17372
rect -33812 17308 -33792 17372
rect -33896 17292 -33792 17308
rect -33896 17228 -33876 17292
rect -33812 17228 -33792 17292
rect -33896 17212 -33792 17228
rect -33896 17148 -33876 17212
rect -33812 17148 -33792 17212
rect -33896 17132 -33792 17148
rect -33896 17068 -33876 17132
rect -33812 17068 -33792 17132
rect -33896 17052 -33792 17068
rect -33896 16988 -33876 17052
rect -33812 16988 -33792 17052
rect -33896 16972 -33792 16988
rect -33896 16908 -33876 16972
rect -33812 16908 -33792 16972
rect -33896 16892 -33792 16908
rect -33896 16828 -33876 16892
rect -33812 16828 -33792 16892
rect -33896 16812 -33792 16828
rect -33896 16748 -33876 16812
rect -33812 16748 -33792 16812
rect -33896 16732 -33792 16748
rect -33896 16668 -33876 16732
rect -33812 16668 -33792 16732
rect -33896 16652 -33792 16668
rect -33896 16588 -33876 16652
rect -33812 16588 -33792 16652
rect -33896 16572 -33792 16588
rect -33896 16508 -33876 16572
rect -33812 16508 -33792 16572
rect -33896 16492 -33792 16508
rect -33896 16428 -33876 16492
rect -33812 16428 -33792 16492
rect -33896 16412 -33792 16428
rect -33896 16348 -33876 16412
rect -33812 16348 -33792 16412
rect -33896 16332 -33792 16348
rect -33896 16268 -33876 16332
rect -33812 16268 -33792 16332
rect -33896 16252 -33792 16268
rect -33896 16188 -33876 16252
rect -33812 16188 -33792 16252
rect -33896 16172 -33792 16188
rect -36676 15761 -36572 16159
rect -33896 16108 -33876 16172
rect -33812 16108 -33792 16172
rect -33473 21052 -28551 21081
rect -33473 16188 -33444 21052
rect -28580 16188 -28551 21052
rect -33473 16159 -28551 16188
rect -28284 21068 -28264 21132
rect -28200 21068 -28180 21132
rect -25452 21081 -25348 21479
rect -22672 21428 -22652 21492
rect -22588 21428 -22568 21492
rect -22249 26372 -17327 26401
rect -22249 21508 -22220 26372
rect -17356 21508 -17327 26372
rect -22249 21479 -17327 21508
rect -17060 26388 -17040 26452
rect -16976 26388 -16956 26452
rect -14228 26401 -14124 26799
rect -11448 26748 -11428 26812
rect -11364 26748 -11344 26812
rect -11025 31692 -6103 31721
rect -11025 26828 -10996 31692
rect -6132 26828 -6103 31692
rect -11025 26799 -6103 26828
rect -5836 31708 -5816 31772
rect -5752 31708 -5732 31772
rect -3004 31721 -2900 32119
rect -224 32068 -204 32132
rect -140 32068 -120 32132
rect 199 37012 5121 37041
rect 199 32148 228 37012
rect 5092 32148 5121 37012
rect 199 32119 5121 32148
rect 5388 37028 5408 37092
rect 5472 37028 5492 37092
rect 8220 37041 8324 37240
rect 11000 37092 11104 37240
rect 5388 37012 5492 37028
rect 5388 36948 5408 37012
rect 5472 36948 5492 37012
rect 5388 36932 5492 36948
rect 5388 36868 5408 36932
rect 5472 36868 5492 36932
rect 5388 36852 5492 36868
rect 5388 36788 5408 36852
rect 5472 36788 5492 36852
rect 5388 36772 5492 36788
rect 5388 36708 5408 36772
rect 5472 36708 5492 36772
rect 5388 36692 5492 36708
rect 5388 36628 5408 36692
rect 5472 36628 5492 36692
rect 5388 36612 5492 36628
rect 5388 36548 5408 36612
rect 5472 36548 5492 36612
rect 5388 36532 5492 36548
rect 5388 36468 5408 36532
rect 5472 36468 5492 36532
rect 5388 36452 5492 36468
rect 5388 36388 5408 36452
rect 5472 36388 5492 36452
rect 5388 36372 5492 36388
rect 5388 36308 5408 36372
rect 5472 36308 5492 36372
rect 5388 36292 5492 36308
rect 5388 36228 5408 36292
rect 5472 36228 5492 36292
rect 5388 36212 5492 36228
rect 5388 36148 5408 36212
rect 5472 36148 5492 36212
rect 5388 36132 5492 36148
rect 5388 36068 5408 36132
rect 5472 36068 5492 36132
rect 5388 36052 5492 36068
rect 5388 35988 5408 36052
rect 5472 35988 5492 36052
rect 5388 35972 5492 35988
rect 5388 35908 5408 35972
rect 5472 35908 5492 35972
rect 5388 35892 5492 35908
rect 5388 35828 5408 35892
rect 5472 35828 5492 35892
rect 5388 35812 5492 35828
rect 5388 35748 5408 35812
rect 5472 35748 5492 35812
rect 5388 35732 5492 35748
rect 5388 35668 5408 35732
rect 5472 35668 5492 35732
rect 5388 35652 5492 35668
rect 5388 35588 5408 35652
rect 5472 35588 5492 35652
rect 5388 35572 5492 35588
rect 5388 35508 5408 35572
rect 5472 35508 5492 35572
rect 5388 35492 5492 35508
rect 5388 35428 5408 35492
rect 5472 35428 5492 35492
rect 5388 35412 5492 35428
rect 5388 35348 5408 35412
rect 5472 35348 5492 35412
rect 5388 35332 5492 35348
rect 5388 35268 5408 35332
rect 5472 35268 5492 35332
rect 5388 35252 5492 35268
rect 5388 35188 5408 35252
rect 5472 35188 5492 35252
rect 5388 35172 5492 35188
rect 5388 35108 5408 35172
rect 5472 35108 5492 35172
rect 5388 35092 5492 35108
rect 5388 35028 5408 35092
rect 5472 35028 5492 35092
rect 5388 35012 5492 35028
rect 5388 34948 5408 35012
rect 5472 34948 5492 35012
rect 5388 34932 5492 34948
rect 5388 34868 5408 34932
rect 5472 34868 5492 34932
rect 5388 34852 5492 34868
rect 5388 34788 5408 34852
rect 5472 34788 5492 34852
rect 5388 34772 5492 34788
rect 5388 34708 5408 34772
rect 5472 34708 5492 34772
rect 5388 34692 5492 34708
rect 5388 34628 5408 34692
rect 5472 34628 5492 34692
rect 5388 34612 5492 34628
rect 5388 34548 5408 34612
rect 5472 34548 5492 34612
rect 5388 34532 5492 34548
rect 5388 34468 5408 34532
rect 5472 34468 5492 34532
rect 5388 34452 5492 34468
rect 5388 34388 5408 34452
rect 5472 34388 5492 34452
rect 5388 34372 5492 34388
rect 5388 34308 5408 34372
rect 5472 34308 5492 34372
rect 5388 34292 5492 34308
rect 5388 34228 5408 34292
rect 5472 34228 5492 34292
rect 5388 34212 5492 34228
rect 5388 34148 5408 34212
rect 5472 34148 5492 34212
rect 5388 34132 5492 34148
rect 5388 34068 5408 34132
rect 5472 34068 5492 34132
rect 5388 34052 5492 34068
rect 5388 33988 5408 34052
rect 5472 33988 5492 34052
rect 5388 33972 5492 33988
rect 5388 33908 5408 33972
rect 5472 33908 5492 33972
rect 5388 33892 5492 33908
rect 5388 33828 5408 33892
rect 5472 33828 5492 33892
rect 5388 33812 5492 33828
rect 5388 33748 5408 33812
rect 5472 33748 5492 33812
rect 5388 33732 5492 33748
rect 5388 33668 5408 33732
rect 5472 33668 5492 33732
rect 5388 33652 5492 33668
rect 5388 33588 5408 33652
rect 5472 33588 5492 33652
rect 5388 33572 5492 33588
rect 5388 33508 5408 33572
rect 5472 33508 5492 33572
rect 5388 33492 5492 33508
rect 5388 33428 5408 33492
rect 5472 33428 5492 33492
rect 5388 33412 5492 33428
rect 5388 33348 5408 33412
rect 5472 33348 5492 33412
rect 5388 33332 5492 33348
rect 5388 33268 5408 33332
rect 5472 33268 5492 33332
rect 5388 33252 5492 33268
rect 5388 33188 5408 33252
rect 5472 33188 5492 33252
rect 5388 33172 5492 33188
rect 5388 33108 5408 33172
rect 5472 33108 5492 33172
rect 5388 33092 5492 33108
rect 5388 33028 5408 33092
rect 5472 33028 5492 33092
rect 5388 33012 5492 33028
rect 5388 32948 5408 33012
rect 5472 32948 5492 33012
rect 5388 32932 5492 32948
rect 5388 32868 5408 32932
rect 5472 32868 5492 32932
rect 5388 32852 5492 32868
rect 5388 32788 5408 32852
rect 5472 32788 5492 32852
rect 5388 32772 5492 32788
rect 5388 32708 5408 32772
rect 5472 32708 5492 32772
rect 5388 32692 5492 32708
rect 5388 32628 5408 32692
rect 5472 32628 5492 32692
rect 5388 32612 5492 32628
rect 5388 32548 5408 32612
rect 5472 32548 5492 32612
rect 5388 32532 5492 32548
rect 5388 32468 5408 32532
rect 5472 32468 5492 32532
rect 5388 32452 5492 32468
rect 5388 32388 5408 32452
rect 5472 32388 5492 32452
rect 5388 32372 5492 32388
rect 5388 32308 5408 32372
rect 5472 32308 5492 32372
rect 5388 32292 5492 32308
rect 5388 32228 5408 32292
rect 5472 32228 5492 32292
rect 5388 32212 5492 32228
rect 5388 32148 5408 32212
rect 5472 32148 5492 32212
rect 5388 32132 5492 32148
rect -224 31772 -120 32068
rect -5836 31692 -5732 31708
rect -5836 31628 -5816 31692
rect -5752 31628 -5732 31692
rect -5836 31612 -5732 31628
rect -5836 31548 -5816 31612
rect -5752 31548 -5732 31612
rect -5836 31532 -5732 31548
rect -5836 31468 -5816 31532
rect -5752 31468 -5732 31532
rect -5836 31452 -5732 31468
rect -5836 31388 -5816 31452
rect -5752 31388 -5732 31452
rect -5836 31372 -5732 31388
rect -5836 31308 -5816 31372
rect -5752 31308 -5732 31372
rect -5836 31292 -5732 31308
rect -5836 31228 -5816 31292
rect -5752 31228 -5732 31292
rect -5836 31212 -5732 31228
rect -5836 31148 -5816 31212
rect -5752 31148 -5732 31212
rect -5836 31132 -5732 31148
rect -5836 31068 -5816 31132
rect -5752 31068 -5732 31132
rect -5836 31052 -5732 31068
rect -5836 30988 -5816 31052
rect -5752 30988 -5732 31052
rect -5836 30972 -5732 30988
rect -5836 30908 -5816 30972
rect -5752 30908 -5732 30972
rect -5836 30892 -5732 30908
rect -5836 30828 -5816 30892
rect -5752 30828 -5732 30892
rect -5836 30812 -5732 30828
rect -5836 30748 -5816 30812
rect -5752 30748 -5732 30812
rect -5836 30732 -5732 30748
rect -5836 30668 -5816 30732
rect -5752 30668 -5732 30732
rect -5836 30652 -5732 30668
rect -5836 30588 -5816 30652
rect -5752 30588 -5732 30652
rect -5836 30572 -5732 30588
rect -5836 30508 -5816 30572
rect -5752 30508 -5732 30572
rect -5836 30492 -5732 30508
rect -5836 30428 -5816 30492
rect -5752 30428 -5732 30492
rect -5836 30412 -5732 30428
rect -5836 30348 -5816 30412
rect -5752 30348 -5732 30412
rect -5836 30332 -5732 30348
rect -5836 30268 -5816 30332
rect -5752 30268 -5732 30332
rect -5836 30252 -5732 30268
rect -5836 30188 -5816 30252
rect -5752 30188 -5732 30252
rect -5836 30172 -5732 30188
rect -5836 30108 -5816 30172
rect -5752 30108 -5732 30172
rect -5836 30092 -5732 30108
rect -5836 30028 -5816 30092
rect -5752 30028 -5732 30092
rect -5836 30012 -5732 30028
rect -5836 29948 -5816 30012
rect -5752 29948 -5732 30012
rect -5836 29932 -5732 29948
rect -5836 29868 -5816 29932
rect -5752 29868 -5732 29932
rect -5836 29852 -5732 29868
rect -5836 29788 -5816 29852
rect -5752 29788 -5732 29852
rect -5836 29772 -5732 29788
rect -5836 29708 -5816 29772
rect -5752 29708 -5732 29772
rect -5836 29692 -5732 29708
rect -5836 29628 -5816 29692
rect -5752 29628 -5732 29692
rect -5836 29612 -5732 29628
rect -5836 29548 -5816 29612
rect -5752 29548 -5732 29612
rect -5836 29532 -5732 29548
rect -5836 29468 -5816 29532
rect -5752 29468 -5732 29532
rect -5836 29452 -5732 29468
rect -5836 29388 -5816 29452
rect -5752 29388 -5732 29452
rect -5836 29372 -5732 29388
rect -5836 29308 -5816 29372
rect -5752 29308 -5732 29372
rect -5836 29292 -5732 29308
rect -5836 29228 -5816 29292
rect -5752 29228 -5732 29292
rect -5836 29212 -5732 29228
rect -5836 29148 -5816 29212
rect -5752 29148 -5732 29212
rect -5836 29132 -5732 29148
rect -5836 29068 -5816 29132
rect -5752 29068 -5732 29132
rect -5836 29052 -5732 29068
rect -5836 28988 -5816 29052
rect -5752 28988 -5732 29052
rect -5836 28972 -5732 28988
rect -5836 28908 -5816 28972
rect -5752 28908 -5732 28972
rect -5836 28892 -5732 28908
rect -5836 28828 -5816 28892
rect -5752 28828 -5732 28892
rect -5836 28812 -5732 28828
rect -5836 28748 -5816 28812
rect -5752 28748 -5732 28812
rect -5836 28732 -5732 28748
rect -5836 28668 -5816 28732
rect -5752 28668 -5732 28732
rect -5836 28652 -5732 28668
rect -5836 28588 -5816 28652
rect -5752 28588 -5732 28652
rect -5836 28572 -5732 28588
rect -5836 28508 -5816 28572
rect -5752 28508 -5732 28572
rect -5836 28492 -5732 28508
rect -5836 28428 -5816 28492
rect -5752 28428 -5732 28492
rect -5836 28412 -5732 28428
rect -5836 28348 -5816 28412
rect -5752 28348 -5732 28412
rect -5836 28332 -5732 28348
rect -5836 28268 -5816 28332
rect -5752 28268 -5732 28332
rect -5836 28252 -5732 28268
rect -5836 28188 -5816 28252
rect -5752 28188 -5732 28252
rect -5836 28172 -5732 28188
rect -5836 28108 -5816 28172
rect -5752 28108 -5732 28172
rect -5836 28092 -5732 28108
rect -5836 28028 -5816 28092
rect -5752 28028 -5732 28092
rect -5836 28012 -5732 28028
rect -5836 27948 -5816 28012
rect -5752 27948 -5732 28012
rect -5836 27932 -5732 27948
rect -5836 27868 -5816 27932
rect -5752 27868 -5732 27932
rect -5836 27852 -5732 27868
rect -5836 27788 -5816 27852
rect -5752 27788 -5732 27852
rect -5836 27772 -5732 27788
rect -5836 27708 -5816 27772
rect -5752 27708 -5732 27772
rect -5836 27692 -5732 27708
rect -5836 27628 -5816 27692
rect -5752 27628 -5732 27692
rect -5836 27612 -5732 27628
rect -5836 27548 -5816 27612
rect -5752 27548 -5732 27612
rect -5836 27532 -5732 27548
rect -5836 27468 -5816 27532
rect -5752 27468 -5732 27532
rect -5836 27452 -5732 27468
rect -5836 27388 -5816 27452
rect -5752 27388 -5732 27452
rect -5836 27372 -5732 27388
rect -5836 27308 -5816 27372
rect -5752 27308 -5732 27372
rect -5836 27292 -5732 27308
rect -5836 27228 -5816 27292
rect -5752 27228 -5732 27292
rect -5836 27212 -5732 27228
rect -5836 27148 -5816 27212
rect -5752 27148 -5732 27212
rect -5836 27132 -5732 27148
rect -5836 27068 -5816 27132
rect -5752 27068 -5732 27132
rect -5836 27052 -5732 27068
rect -5836 26988 -5816 27052
rect -5752 26988 -5732 27052
rect -5836 26972 -5732 26988
rect -5836 26908 -5816 26972
rect -5752 26908 -5732 26972
rect -5836 26892 -5732 26908
rect -5836 26828 -5816 26892
rect -5752 26828 -5732 26892
rect -5836 26812 -5732 26828
rect -11448 26452 -11344 26748
rect -17060 26372 -16956 26388
rect -17060 26308 -17040 26372
rect -16976 26308 -16956 26372
rect -17060 26292 -16956 26308
rect -17060 26228 -17040 26292
rect -16976 26228 -16956 26292
rect -17060 26212 -16956 26228
rect -17060 26148 -17040 26212
rect -16976 26148 -16956 26212
rect -17060 26132 -16956 26148
rect -17060 26068 -17040 26132
rect -16976 26068 -16956 26132
rect -17060 26052 -16956 26068
rect -17060 25988 -17040 26052
rect -16976 25988 -16956 26052
rect -17060 25972 -16956 25988
rect -17060 25908 -17040 25972
rect -16976 25908 -16956 25972
rect -17060 25892 -16956 25908
rect -17060 25828 -17040 25892
rect -16976 25828 -16956 25892
rect -17060 25812 -16956 25828
rect -17060 25748 -17040 25812
rect -16976 25748 -16956 25812
rect -17060 25732 -16956 25748
rect -17060 25668 -17040 25732
rect -16976 25668 -16956 25732
rect -17060 25652 -16956 25668
rect -17060 25588 -17040 25652
rect -16976 25588 -16956 25652
rect -17060 25572 -16956 25588
rect -17060 25508 -17040 25572
rect -16976 25508 -16956 25572
rect -17060 25492 -16956 25508
rect -17060 25428 -17040 25492
rect -16976 25428 -16956 25492
rect -17060 25412 -16956 25428
rect -17060 25348 -17040 25412
rect -16976 25348 -16956 25412
rect -17060 25332 -16956 25348
rect -17060 25268 -17040 25332
rect -16976 25268 -16956 25332
rect -17060 25252 -16956 25268
rect -17060 25188 -17040 25252
rect -16976 25188 -16956 25252
rect -17060 25172 -16956 25188
rect -17060 25108 -17040 25172
rect -16976 25108 -16956 25172
rect -17060 25092 -16956 25108
rect -17060 25028 -17040 25092
rect -16976 25028 -16956 25092
rect -17060 25012 -16956 25028
rect -17060 24948 -17040 25012
rect -16976 24948 -16956 25012
rect -17060 24932 -16956 24948
rect -17060 24868 -17040 24932
rect -16976 24868 -16956 24932
rect -17060 24852 -16956 24868
rect -17060 24788 -17040 24852
rect -16976 24788 -16956 24852
rect -17060 24772 -16956 24788
rect -17060 24708 -17040 24772
rect -16976 24708 -16956 24772
rect -17060 24692 -16956 24708
rect -17060 24628 -17040 24692
rect -16976 24628 -16956 24692
rect -17060 24612 -16956 24628
rect -17060 24548 -17040 24612
rect -16976 24548 -16956 24612
rect -17060 24532 -16956 24548
rect -17060 24468 -17040 24532
rect -16976 24468 -16956 24532
rect -17060 24452 -16956 24468
rect -17060 24388 -17040 24452
rect -16976 24388 -16956 24452
rect -17060 24372 -16956 24388
rect -17060 24308 -17040 24372
rect -16976 24308 -16956 24372
rect -17060 24292 -16956 24308
rect -17060 24228 -17040 24292
rect -16976 24228 -16956 24292
rect -17060 24212 -16956 24228
rect -17060 24148 -17040 24212
rect -16976 24148 -16956 24212
rect -17060 24132 -16956 24148
rect -17060 24068 -17040 24132
rect -16976 24068 -16956 24132
rect -17060 24052 -16956 24068
rect -17060 23988 -17040 24052
rect -16976 23988 -16956 24052
rect -17060 23972 -16956 23988
rect -17060 23908 -17040 23972
rect -16976 23908 -16956 23972
rect -17060 23892 -16956 23908
rect -17060 23828 -17040 23892
rect -16976 23828 -16956 23892
rect -17060 23812 -16956 23828
rect -17060 23748 -17040 23812
rect -16976 23748 -16956 23812
rect -17060 23732 -16956 23748
rect -17060 23668 -17040 23732
rect -16976 23668 -16956 23732
rect -17060 23652 -16956 23668
rect -17060 23588 -17040 23652
rect -16976 23588 -16956 23652
rect -17060 23572 -16956 23588
rect -17060 23508 -17040 23572
rect -16976 23508 -16956 23572
rect -17060 23492 -16956 23508
rect -17060 23428 -17040 23492
rect -16976 23428 -16956 23492
rect -17060 23412 -16956 23428
rect -17060 23348 -17040 23412
rect -16976 23348 -16956 23412
rect -17060 23332 -16956 23348
rect -17060 23268 -17040 23332
rect -16976 23268 -16956 23332
rect -17060 23252 -16956 23268
rect -17060 23188 -17040 23252
rect -16976 23188 -16956 23252
rect -17060 23172 -16956 23188
rect -17060 23108 -17040 23172
rect -16976 23108 -16956 23172
rect -17060 23092 -16956 23108
rect -17060 23028 -17040 23092
rect -16976 23028 -16956 23092
rect -17060 23012 -16956 23028
rect -17060 22948 -17040 23012
rect -16976 22948 -16956 23012
rect -17060 22932 -16956 22948
rect -17060 22868 -17040 22932
rect -16976 22868 -16956 22932
rect -17060 22852 -16956 22868
rect -17060 22788 -17040 22852
rect -16976 22788 -16956 22852
rect -17060 22772 -16956 22788
rect -17060 22708 -17040 22772
rect -16976 22708 -16956 22772
rect -17060 22692 -16956 22708
rect -17060 22628 -17040 22692
rect -16976 22628 -16956 22692
rect -17060 22612 -16956 22628
rect -17060 22548 -17040 22612
rect -16976 22548 -16956 22612
rect -17060 22532 -16956 22548
rect -17060 22468 -17040 22532
rect -16976 22468 -16956 22532
rect -17060 22452 -16956 22468
rect -17060 22388 -17040 22452
rect -16976 22388 -16956 22452
rect -17060 22372 -16956 22388
rect -17060 22308 -17040 22372
rect -16976 22308 -16956 22372
rect -17060 22292 -16956 22308
rect -17060 22228 -17040 22292
rect -16976 22228 -16956 22292
rect -17060 22212 -16956 22228
rect -17060 22148 -17040 22212
rect -16976 22148 -16956 22212
rect -17060 22132 -16956 22148
rect -17060 22068 -17040 22132
rect -16976 22068 -16956 22132
rect -17060 22052 -16956 22068
rect -17060 21988 -17040 22052
rect -16976 21988 -16956 22052
rect -17060 21972 -16956 21988
rect -17060 21908 -17040 21972
rect -16976 21908 -16956 21972
rect -17060 21892 -16956 21908
rect -17060 21828 -17040 21892
rect -16976 21828 -16956 21892
rect -17060 21812 -16956 21828
rect -17060 21748 -17040 21812
rect -16976 21748 -16956 21812
rect -17060 21732 -16956 21748
rect -17060 21668 -17040 21732
rect -16976 21668 -16956 21732
rect -17060 21652 -16956 21668
rect -17060 21588 -17040 21652
rect -16976 21588 -16956 21652
rect -17060 21572 -16956 21588
rect -17060 21508 -17040 21572
rect -16976 21508 -16956 21572
rect -17060 21492 -16956 21508
rect -22672 21132 -22568 21428
rect -28284 21052 -28180 21068
rect -28284 20988 -28264 21052
rect -28200 20988 -28180 21052
rect -28284 20972 -28180 20988
rect -28284 20908 -28264 20972
rect -28200 20908 -28180 20972
rect -28284 20892 -28180 20908
rect -28284 20828 -28264 20892
rect -28200 20828 -28180 20892
rect -28284 20812 -28180 20828
rect -28284 20748 -28264 20812
rect -28200 20748 -28180 20812
rect -28284 20732 -28180 20748
rect -28284 20668 -28264 20732
rect -28200 20668 -28180 20732
rect -28284 20652 -28180 20668
rect -28284 20588 -28264 20652
rect -28200 20588 -28180 20652
rect -28284 20572 -28180 20588
rect -28284 20508 -28264 20572
rect -28200 20508 -28180 20572
rect -28284 20492 -28180 20508
rect -28284 20428 -28264 20492
rect -28200 20428 -28180 20492
rect -28284 20412 -28180 20428
rect -28284 20348 -28264 20412
rect -28200 20348 -28180 20412
rect -28284 20332 -28180 20348
rect -28284 20268 -28264 20332
rect -28200 20268 -28180 20332
rect -28284 20252 -28180 20268
rect -28284 20188 -28264 20252
rect -28200 20188 -28180 20252
rect -28284 20172 -28180 20188
rect -28284 20108 -28264 20172
rect -28200 20108 -28180 20172
rect -28284 20092 -28180 20108
rect -28284 20028 -28264 20092
rect -28200 20028 -28180 20092
rect -28284 20012 -28180 20028
rect -28284 19948 -28264 20012
rect -28200 19948 -28180 20012
rect -28284 19932 -28180 19948
rect -28284 19868 -28264 19932
rect -28200 19868 -28180 19932
rect -28284 19852 -28180 19868
rect -28284 19788 -28264 19852
rect -28200 19788 -28180 19852
rect -28284 19772 -28180 19788
rect -28284 19708 -28264 19772
rect -28200 19708 -28180 19772
rect -28284 19692 -28180 19708
rect -28284 19628 -28264 19692
rect -28200 19628 -28180 19692
rect -28284 19612 -28180 19628
rect -28284 19548 -28264 19612
rect -28200 19548 -28180 19612
rect -28284 19532 -28180 19548
rect -28284 19468 -28264 19532
rect -28200 19468 -28180 19532
rect -28284 19452 -28180 19468
rect -28284 19388 -28264 19452
rect -28200 19388 -28180 19452
rect -28284 19372 -28180 19388
rect -28284 19308 -28264 19372
rect -28200 19308 -28180 19372
rect -28284 19292 -28180 19308
rect -28284 19228 -28264 19292
rect -28200 19228 -28180 19292
rect -28284 19212 -28180 19228
rect -28284 19148 -28264 19212
rect -28200 19148 -28180 19212
rect -28284 19132 -28180 19148
rect -28284 19068 -28264 19132
rect -28200 19068 -28180 19132
rect -28284 19052 -28180 19068
rect -28284 18988 -28264 19052
rect -28200 18988 -28180 19052
rect -28284 18972 -28180 18988
rect -28284 18908 -28264 18972
rect -28200 18908 -28180 18972
rect -28284 18892 -28180 18908
rect -28284 18828 -28264 18892
rect -28200 18828 -28180 18892
rect -28284 18812 -28180 18828
rect -28284 18748 -28264 18812
rect -28200 18748 -28180 18812
rect -28284 18732 -28180 18748
rect -28284 18668 -28264 18732
rect -28200 18668 -28180 18732
rect -28284 18652 -28180 18668
rect -28284 18588 -28264 18652
rect -28200 18588 -28180 18652
rect -28284 18572 -28180 18588
rect -28284 18508 -28264 18572
rect -28200 18508 -28180 18572
rect -28284 18492 -28180 18508
rect -28284 18428 -28264 18492
rect -28200 18428 -28180 18492
rect -28284 18412 -28180 18428
rect -28284 18348 -28264 18412
rect -28200 18348 -28180 18412
rect -28284 18332 -28180 18348
rect -28284 18268 -28264 18332
rect -28200 18268 -28180 18332
rect -28284 18252 -28180 18268
rect -28284 18188 -28264 18252
rect -28200 18188 -28180 18252
rect -28284 18172 -28180 18188
rect -28284 18108 -28264 18172
rect -28200 18108 -28180 18172
rect -28284 18092 -28180 18108
rect -28284 18028 -28264 18092
rect -28200 18028 -28180 18092
rect -28284 18012 -28180 18028
rect -28284 17948 -28264 18012
rect -28200 17948 -28180 18012
rect -28284 17932 -28180 17948
rect -28284 17868 -28264 17932
rect -28200 17868 -28180 17932
rect -28284 17852 -28180 17868
rect -28284 17788 -28264 17852
rect -28200 17788 -28180 17852
rect -28284 17772 -28180 17788
rect -28284 17708 -28264 17772
rect -28200 17708 -28180 17772
rect -28284 17692 -28180 17708
rect -28284 17628 -28264 17692
rect -28200 17628 -28180 17692
rect -28284 17612 -28180 17628
rect -28284 17548 -28264 17612
rect -28200 17548 -28180 17612
rect -28284 17532 -28180 17548
rect -28284 17468 -28264 17532
rect -28200 17468 -28180 17532
rect -28284 17452 -28180 17468
rect -28284 17388 -28264 17452
rect -28200 17388 -28180 17452
rect -28284 17372 -28180 17388
rect -28284 17308 -28264 17372
rect -28200 17308 -28180 17372
rect -28284 17292 -28180 17308
rect -28284 17228 -28264 17292
rect -28200 17228 -28180 17292
rect -28284 17212 -28180 17228
rect -28284 17148 -28264 17212
rect -28200 17148 -28180 17212
rect -28284 17132 -28180 17148
rect -28284 17068 -28264 17132
rect -28200 17068 -28180 17132
rect -28284 17052 -28180 17068
rect -28284 16988 -28264 17052
rect -28200 16988 -28180 17052
rect -28284 16972 -28180 16988
rect -28284 16908 -28264 16972
rect -28200 16908 -28180 16972
rect -28284 16892 -28180 16908
rect -28284 16828 -28264 16892
rect -28200 16828 -28180 16892
rect -28284 16812 -28180 16828
rect -28284 16748 -28264 16812
rect -28200 16748 -28180 16812
rect -28284 16732 -28180 16748
rect -28284 16668 -28264 16732
rect -28200 16668 -28180 16732
rect -28284 16652 -28180 16668
rect -28284 16588 -28264 16652
rect -28200 16588 -28180 16652
rect -28284 16572 -28180 16588
rect -28284 16508 -28264 16572
rect -28200 16508 -28180 16572
rect -28284 16492 -28180 16508
rect -28284 16428 -28264 16492
rect -28200 16428 -28180 16492
rect -28284 16412 -28180 16428
rect -28284 16348 -28264 16412
rect -28200 16348 -28180 16412
rect -28284 16332 -28180 16348
rect -28284 16268 -28264 16332
rect -28200 16268 -28180 16332
rect -28284 16252 -28180 16268
rect -28284 16188 -28264 16252
rect -28200 16188 -28180 16252
rect -28284 16172 -28180 16188
rect -33896 15812 -33792 16108
rect -39085 15732 -34163 15761
rect -39085 10868 -39056 15732
rect -34192 10868 -34163 15732
rect -39085 10839 -34163 10868
rect -33896 15748 -33876 15812
rect -33812 15748 -33792 15812
rect -31064 15761 -30960 16159
rect -28284 16108 -28264 16172
rect -28200 16108 -28180 16172
rect -27861 21052 -22939 21081
rect -27861 16188 -27832 21052
rect -22968 16188 -22939 21052
rect -27861 16159 -22939 16188
rect -22672 21068 -22652 21132
rect -22588 21068 -22568 21132
rect -19840 21081 -19736 21479
rect -17060 21428 -17040 21492
rect -16976 21428 -16956 21492
rect -16637 26372 -11715 26401
rect -16637 21508 -16608 26372
rect -11744 21508 -11715 26372
rect -16637 21479 -11715 21508
rect -11448 26388 -11428 26452
rect -11364 26388 -11344 26452
rect -8616 26401 -8512 26799
rect -5836 26748 -5816 26812
rect -5752 26748 -5732 26812
rect -5413 31692 -491 31721
rect -5413 26828 -5384 31692
rect -520 26828 -491 31692
rect -5413 26799 -491 26828
rect -224 31708 -204 31772
rect -140 31708 -120 31772
rect 2608 31721 2712 32119
rect 5388 32068 5408 32132
rect 5472 32068 5492 32132
rect 5811 37012 10733 37041
rect 5811 32148 5840 37012
rect 10704 32148 10733 37012
rect 5811 32119 10733 32148
rect 11000 37028 11020 37092
rect 11084 37028 11104 37092
rect 13832 37041 13936 37240
rect 16612 37092 16716 37240
rect 11000 37012 11104 37028
rect 11000 36948 11020 37012
rect 11084 36948 11104 37012
rect 11000 36932 11104 36948
rect 11000 36868 11020 36932
rect 11084 36868 11104 36932
rect 11000 36852 11104 36868
rect 11000 36788 11020 36852
rect 11084 36788 11104 36852
rect 11000 36772 11104 36788
rect 11000 36708 11020 36772
rect 11084 36708 11104 36772
rect 11000 36692 11104 36708
rect 11000 36628 11020 36692
rect 11084 36628 11104 36692
rect 11000 36612 11104 36628
rect 11000 36548 11020 36612
rect 11084 36548 11104 36612
rect 11000 36532 11104 36548
rect 11000 36468 11020 36532
rect 11084 36468 11104 36532
rect 11000 36452 11104 36468
rect 11000 36388 11020 36452
rect 11084 36388 11104 36452
rect 11000 36372 11104 36388
rect 11000 36308 11020 36372
rect 11084 36308 11104 36372
rect 11000 36292 11104 36308
rect 11000 36228 11020 36292
rect 11084 36228 11104 36292
rect 11000 36212 11104 36228
rect 11000 36148 11020 36212
rect 11084 36148 11104 36212
rect 11000 36132 11104 36148
rect 11000 36068 11020 36132
rect 11084 36068 11104 36132
rect 11000 36052 11104 36068
rect 11000 35988 11020 36052
rect 11084 35988 11104 36052
rect 11000 35972 11104 35988
rect 11000 35908 11020 35972
rect 11084 35908 11104 35972
rect 11000 35892 11104 35908
rect 11000 35828 11020 35892
rect 11084 35828 11104 35892
rect 11000 35812 11104 35828
rect 11000 35748 11020 35812
rect 11084 35748 11104 35812
rect 11000 35732 11104 35748
rect 11000 35668 11020 35732
rect 11084 35668 11104 35732
rect 11000 35652 11104 35668
rect 11000 35588 11020 35652
rect 11084 35588 11104 35652
rect 11000 35572 11104 35588
rect 11000 35508 11020 35572
rect 11084 35508 11104 35572
rect 11000 35492 11104 35508
rect 11000 35428 11020 35492
rect 11084 35428 11104 35492
rect 11000 35412 11104 35428
rect 11000 35348 11020 35412
rect 11084 35348 11104 35412
rect 11000 35332 11104 35348
rect 11000 35268 11020 35332
rect 11084 35268 11104 35332
rect 11000 35252 11104 35268
rect 11000 35188 11020 35252
rect 11084 35188 11104 35252
rect 11000 35172 11104 35188
rect 11000 35108 11020 35172
rect 11084 35108 11104 35172
rect 11000 35092 11104 35108
rect 11000 35028 11020 35092
rect 11084 35028 11104 35092
rect 11000 35012 11104 35028
rect 11000 34948 11020 35012
rect 11084 34948 11104 35012
rect 11000 34932 11104 34948
rect 11000 34868 11020 34932
rect 11084 34868 11104 34932
rect 11000 34852 11104 34868
rect 11000 34788 11020 34852
rect 11084 34788 11104 34852
rect 11000 34772 11104 34788
rect 11000 34708 11020 34772
rect 11084 34708 11104 34772
rect 11000 34692 11104 34708
rect 11000 34628 11020 34692
rect 11084 34628 11104 34692
rect 11000 34612 11104 34628
rect 11000 34548 11020 34612
rect 11084 34548 11104 34612
rect 11000 34532 11104 34548
rect 11000 34468 11020 34532
rect 11084 34468 11104 34532
rect 11000 34452 11104 34468
rect 11000 34388 11020 34452
rect 11084 34388 11104 34452
rect 11000 34372 11104 34388
rect 11000 34308 11020 34372
rect 11084 34308 11104 34372
rect 11000 34292 11104 34308
rect 11000 34228 11020 34292
rect 11084 34228 11104 34292
rect 11000 34212 11104 34228
rect 11000 34148 11020 34212
rect 11084 34148 11104 34212
rect 11000 34132 11104 34148
rect 11000 34068 11020 34132
rect 11084 34068 11104 34132
rect 11000 34052 11104 34068
rect 11000 33988 11020 34052
rect 11084 33988 11104 34052
rect 11000 33972 11104 33988
rect 11000 33908 11020 33972
rect 11084 33908 11104 33972
rect 11000 33892 11104 33908
rect 11000 33828 11020 33892
rect 11084 33828 11104 33892
rect 11000 33812 11104 33828
rect 11000 33748 11020 33812
rect 11084 33748 11104 33812
rect 11000 33732 11104 33748
rect 11000 33668 11020 33732
rect 11084 33668 11104 33732
rect 11000 33652 11104 33668
rect 11000 33588 11020 33652
rect 11084 33588 11104 33652
rect 11000 33572 11104 33588
rect 11000 33508 11020 33572
rect 11084 33508 11104 33572
rect 11000 33492 11104 33508
rect 11000 33428 11020 33492
rect 11084 33428 11104 33492
rect 11000 33412 11104 33428
rect 11000 33348 11020 33412
rect 11084 33348 11104 33412
rect 11000 33332 11104 33348
rect 11000 33268 11020 33332
rect 11084 33268 11104 33332
rect 11000 33252 11104 33268
rect 11000 33188 11020 33252
rect 11084 33188 11104 33252
rect 11000 33172 11104 33188
rect 11000 33108 11020 33172
rect 11084 33108 11104 33172
rect 11000 33092 11104 33108
rect 11000 33028 11020 33092
rect 11084 33028 11104 33092
rect 11000 33012 11104 33028
rect 11000 32948 11020 33012
rect 11084 32948 11104 33012
rect 11000 32932 11104 32948
rect 11000 32868 11020 32932
rect 11084 32868 11104 32932
rect 11000 32852 11104 32868
rect 11000 32788 11020 32852
rect 11084 32788 11104 32852
rect 11000 32772 11104 32788
rect 11000 32708 11020 32772
rect 11084 32708 11104 32772
rect 11000 32692 11104 32708
rect 11000 32628 11020 32692
rect 11084 32628 11104 32692
rect 11000 32612 11104 32628
rect 11000 32548 11020 32612
rect 11084 32548 11104 32612
rect 11000 32532 11104 32548
rect 11000 32468 11020 32532
rect 11084 32468 11104 32532
rect 11000 32452 11104 32468
rect 11000 32388 11020 32452
rect 11084 32388 11104 32452
rect 11000 32372 11104 32388
rect 11000 32308 11020 32372
rect 11084 32308 11104 32372
rect 11000 32292 11104 32308
rect 11000 32228 11020 32292
rect 11084 32228 11104 32292
rect 11000 32212 11104 32228
rect 11000 32148 11020 32212
rect 11084 32148 11104 32212
rect 11000 32132 11104 32148
rect 5388 31772 5492 32068
rect -224 31692 -120 31708
rect -224 31628 -204 31692
rect -140 31628 -120 31692
rect -224 31612 -120 31628
rect -224 31548 -204 31612
rect -140 31548 -120 31612
rect -224 31532 -120 31548
rect -224 31468 -204 31532
rect -140 31468 -120 31532
rect -224 31452 -120 31468
rect -224 31388 -204 31452
rect -140 31388 -120 31452
rect -224 31372 -120 31388
rect -224 31308 -204 31372
rect -140 31308 -120 31372
rect -224 31292 -120 31308
rect -224 31228 -204 31292
rect -140 31228 -120 31292
rect -224 31212 -120 31228
rect -224 31148 -204 31212
rect -140 31148 -120 31212
rect -224 31132 -120 31148
rect -224 31068 -204 31132
rect -140 31068 -120 31132
rect -224 31052 -120 31068
rect -224 30988 -204 31052
rect -140 30988 -120 31052
rect -224 30972 -120 30988
rect -224 30908 -204 30972
rect -140 30908 -120 30972
rect -224 30892 -120 30908
rect -224 30828 -204 30892
rect -140 30828 -120 30892
rect -224 30812 -120 30828
rect -224 30748 -204 30812
rect -140 30748 -120 30812
rect -224 30732 -120 30748
rect -224 30668 -204 30732
rect -140 30668 -120 30732
rect -224 30652 -120 30668
rect -224 30588 -204 30652
rect -140 30588 -120 30652
rect -224 30572 -120 30588
rect -224 30508 -204 30572
rect -140 30508 -120 30572
rect -224 30492 -120 30508
rect -224 30428 -204 30492
rect -140 30428 -120 30492
rect -224 30412 -120 30428
rect -224 30348 -204 30412
rect -140 30348 -120 30412
rect -224 30332 -120 30348
rect -224 30268 -204 30332
rect -140 30268 -120 30332
rect -224 30252 -120 30268
rect -224 30188 -204 30252
rect -140 30188 -120 30252
rect -224 30172 -120 30188
rect -224 30108 -204 30172
rect -140 30108 -120 30172
rect -224 30092 -120 30108
rect -224 30028 -204 30092
rect -140 30028 -120 30092
rect -224 30012 -120 30028
rect -224 29948 -204 30012
rect -140 29948 -120 30012
rect -224 29932 -120 29948
rect -224 29868 -204 29932
rect -140 29868 -120 29932
rect -224 29852 -120 29868
rect -224 29788 -204 29852
rect -140 29788 -120 29852
rect -224 29772 -120 29788
rect -224 29708 -204 29772
rect -140 29708 -120 29772
rect -224 29692 -120 29708
rect -224 29628 -204 29692
rect -140 29628 -120 29692
rect -224 29612 -120 29628
rect -224 29548 -204 29612
rect -140 29548 -120 29612
rect -224 29532 -120 29548
rect -224 29468 -204 29532
rect -140 29468 -120 29532
rect -224 29452 -120 29468
rect -224 29388 -204 29452
rect -140 29388 -120 29452
rect -224 29372 -120 29388
rect -224 29308 -204 29372
rect -140 29308 -120 29372
rect -224 29292 -120 29308
rect -224 29228 -204 29292
rect -140 29228 -120 29292
rect -224 29212 -120 29228
rect -224 29148 -204 29212
rect -140 29148 -120 29212
rect -224 29132 -120 29148
rect -224 29068 -204 29132
rect -140 29068 -120 29132
rect -224 29052 -120 29068
rect -224 28988 -204 29052
rect -140 28988 -120 29052
rect -224 28972 -120 28988
rect -224 28908 -204 28972
rect -140 28908 -120 28972
rect -224 28892 -120 28908
rect -224 28828 -204 28892
rect -140 28828 -120 28892
rect -224 28812 -120 28828
rect -224 28748 -204 28812
rect -140 28748 -120 28812
rect -224 28732 -120 28748
rect -224 28668 -204 28732
rect -140 28668 -120 28732
rect -224 28652 -120 28668
rect -224 28588 -204 28652
rect -140 28588 -120 28652
rect -224 28572 -120 28588
rect -224 28508 -204 28572
rect -140 28508 -120 28572
rect -224 28492 -120 28508
rect -224 28428 -204 28492
rect -140 28428 -120 28492
rect -224 28412 -120 28428
rect -224 28348 -204 28412
rect -140 28348 -120 28412
rect -224 28332 -120 28348
rect -224 28268 -204 28332
rect -140 28268 -120 28332
rect -224 28252 -120 28268
rect -224 28188 -204 28252
rect -140 28188 -120 28252
rect -224 28172 -120 28188
rect -224 28108 -204 28172
rect -140 28108 -120 28172
rect -224 28092 -120 28108
rect -224 28028 -204 28092
rect -140 28028 -120 28092
rect -224 28012 -120 28028
rect -224 27948 -204 28012
rect -140 27948 -120 28012
rect -224 27932 -120 27948
rect -224 27868 -204 27932
rect -140 27868 -120 27932
rect -224 27852 -120 27868
rect -224 27788 -204 27852
rect -140 27788 -120 27852
rect -224 27772 -120 27788
rect -224 27708 -204 27772
rect -140 27708 -120 27772
rect -224 27692 -120 27708
rect -224 27628 -204 27692
rect -140 27628 -120 27692
rect -224 27612 -120 27628
rect -224 27548 -204 27612
rect -140 27548 -120 27612
rect -224 27532 -120 27548
rect -224 27468 -204 27532
rect -140 27468 -120 27532
rect -224 27452 -120 27468
rect -224 27388 -204 27452
rect -140 27388 -120 27452
rect -224 27372 -120 27388
rect -224 27308 -204 27372
rect -140 27308 -120 27372
rect -224 27292 -120 27308
rect -224 27228 -204 27292
rect -140 27228 -120 27292
rect -224 27212 -120 27228
rect -224 27148 -204 27212
rect -140 27148 -120 27212
rect -224 27132 -120 27148
rect -224 27068 -204 27132
rect -140 27068 -120 27132
rect -224 27052 -120 27068
rect -224 26988 -204 27052
rect -140 26988 -120 27052
rect -224 26972 -120 26988
rect -224 26908 -204 26972
rect -140 26908 -120 26972
rect -224 26892 -120 26908
rect -224 26828 -204 26892
rect -140 26828 -120 26892
rect -224 26812 -120 26828
rect -5836 26452 -5732 26748
rect -11448 26372 -11344 26388
rect -11448 26308 -11428 26372
rect -11364 26308 -11344 26372
rect -11448 26292 -11344 26308
rect -11448 26228 -11428 26292
rect -11364 26228 -11344 26292
rect -11448 26212 -11344 26228
rect -11448 26148 -11428 26212
rect -11364 26148 -11344 26212
rect -11448 26132 -11344 26148
rect -11448 26068 -11428 26132
rect -11364 26068 -11344 26132
rect -11448 26052 -11344 26068
rect -11448 25988 -11428 26052
rect -11364 25988 -11344 26052
rect -11448 25972 -11344 25988
rect -11448 25908 -11428 25972
rect -11364 25908 -11344 25972
rect -11448 25892 -11344 25908
rect -11448 25828 -11428 25892
rect -11364 25828 -11344 25892
rect -11448 25812 -11344 25828
rect -11448 25748 -11428 25812
rect -11364 25748 -11344 25812
rect -11448 25732 -11344 25748
rect -11448 25668 -11428 25732
rect -11364 25668 -11344 25732
rect -11448 25652 -11344 25668
rect -11448 25588 -11428 25652
rect -11364 25588 -11344 25652
rect -11448 25572 -11344 25588
rect -11448 25508 -11428 25572
rect -11364 25508 -11344 25572
rect -11448 25492 -11344 25508
rect -11448 25428 -11428 25492
rect -11364 25428 -11344 25492
rect -11448 25412 -11344 25428
rect -11448 25348 -11428 25412
rect -11364 25348 -11344 25412
rect -11448 25332 -11344 25348
rect -11448 25268 -11428 25332
rect -11364 25268 -11344 25332
rect -11448 25252 -11344 25268
rect -11448 25188 -11428 25252
rect -11364 25188 -11344 25252
rect -11448 25172 -11344 25188
rect -11448 25108 -11428 25172
rect -11364 25108 -11344 25172
rect -11448 25092 -11344 25108
rect -11448 25028 -11428 25092
rect -11364 25028 -11344 25092
rect -11448 25012 -11344 25028
rect -11448 24948 -11428 25012
rect -11364 24948 -11344 25012
rect -11448 24932 -11344 24948
rect -11448 24868 -11428 24932
rect -11364 24868 -11344 24932
rect -11448 24852 -11344 24868
rect -11448 24788 -11428 24852
rect -11364 24788 -11344 24852
rect -11448 24772 -11344 24788
rect -11448 24708 -11428 24772
rect -11364 24708 -11344 24772
rect -11448 24692 -11344 24708
rect -11448 24628 -11428 24692
rect -11364 24628 -11344 24692
rect -11448 24612 -11344 24628
rect -11448 24548 -11428 24612
rect -11364 24548 -11344 24612
rect -11448 24532 -11344 24548
rect -11448 24468 -11428 24532
rect -11364 24468 -11344 24532
rect -11448 24452 -11344 24468
rect -11448 24388 -11428 24452
rect -11364 24388 -11344 24452
rect -11448 24372 -11344 24388
rect -11448 24308 -11428 24372
rect -11364 24308 -11344 24372
rect -11448 24292 -11344 24308
rect -11448 24228 -11428 24292
rect -11364 24228 -11344 24292
rect -11448 24212 -11344 24228
rect -11448 24148 -11428 24212
rect -11364 24148 -11344 24212
rect -11448 24132 -11344 24148
rect -11448 24068 -11428 24132
rect -11364 24068 -11344 24132
rect -11448 24052 -11344 24068
rect -11448 23988 -11428 24052
rect -11364 23988 -11344 24052
rect -11448 23972 -11344 23988
rect -11448 23908 -11428 23972
rect -11364 23908 -11344 23972
rect -11448 23892 -11344 23908
rect -11448 23828 -11428 23892
rect -11364 23828 -11344 23892
rect -11448 23812 -11344 23828
rect -11448 23748 -11428 23812
rect -11364 23748 -11344 23812
rect -11448 23732 -11344 23748
rect -11448 23668 -11428 23732
rect -11364 23668 -11344 23732
rect -11448 23652 -11344 23668
rect -11448 23588 -11428 23652
rect -11364 23588 -11344 23652
rect -11448 23572 -11344 23588
rect -11448 23508 -11428 23572
rect -11364 23508 -11344 23572
rect -11448 23492 -11344 23508
rect -11448 23428 -11428 23492
rect -11364 23428 -11344 23492
rect -11448 23412 -11344 23428
rect -11448 23348 -11428 23412
rect -11364 23348 -11344 23412
rect -11448 23332 -11344 23348
rect -11448 23268 -11428 23332
rect -11364 23268 -11344 23332
rect -11448 23252 -11344 23268
rect -11448 23188 -11428 23252
rect -11364 23188 -11344 23252
rect -11448 23172 -11344 23188
rect -11448 23108 -11428 23172
rect -11364 23108 -11344 23172
rect -11448 23092 -11344 23108
rect -11448 23028 -11428 23092
rect -11364 23028 -11344 23092
rect -11448 23012 -11344 23028
rect -11448 22948 -11428 23012
rect -11364 22948 -11344 23012
rect -11448 22932 -11344 22948
rect -11448 22868 -11428 22932
rect -11364 22868 -11344 22932
rect -11448 22852 -11344 22868
rect -11448 22788 -11428 22852
rect -11364 22788 -11344 22852
rect -11448 22772 -11344 22788
rect -11448 22708 -11428 22772
rect -11364 22708 -11344 22772
rect -11448 22692 -11344 22708
rect -11448 22628 -11428 22692
rect -11364 22628 -11344 22692
rect -11448 22612 -11344 22628
rect -11448 22548 -11428 22612
rect -11364 22548 -11344 22612
rect -11448 22532 -11344 22548
rect -11448 22468 -11428 22532
rect -11364 22468 -11344 22532
rect -11448 22452 -11344 22468
rect -11448 22388 -11428 22452
rect -11364 22388 -11344 22452
rect -11448 22372 -11344 22388
rect -11448 22308 -11428 22372
rect -11364 22308 -11344 22372
rect -11448 22292 -11344 22308
rect -11448 22228 -11428 22292
rect -11364 22228 -11344 22292
rect -11448 22212 -11344 22228
rect -11448 22148 -11428 22212
rect -11364 22148 -11344 22212
rect -11448 22132 -11344 22148
rect -11448 22068 -11428 22132
rect -11364 22068 -11344 22132
rect -11448 22052 -11344 22068
rect -11448 21988 -11428 22052
rect -11364 21988 -11344 22052
rect -11448 21972 -11344 21988
rect -11448 21908 -11428 21972
rect -11364 21908 -11344 21972
rect -11448 21892 -11344 21908
rect -11448 21828 -11428 21892
rect -11364 21828 -11344 21892
rect -11448 21812 -11344 21828
rect -11448 21748 -11428 21812
rect -11364 21748 -11344 21812
rect -11448 21732 -11344 21748
rect -11448 21668 -11428 21732
rect -11364 21668 -11344 21732
rect -11448 21652 -11344 21668
rect -11448 21588 -11428 21652
rect -11364 21588 -11344 21652
rect -11448 21572 -11344 21588
rect -11448 21508 -11428 21572
rect -11364 21508 -11344 21572
rect -11448 21492 -11344 21508
rect -17060 21132 -16956 21428
rect -22672 21052 -22568 21068
rect -22672 20988 -22652 21052
rect -22588 20988 -22568 21052
rect -22672 20972 -22568 20988
rect -22672 20908 -22652 20972
rect -22588 20908 -22568 20972
rect -22672 20892 -22568 20908
rect -22672 20828 -22652 20892
rect -22588 20828 -22568 20892
rect -22672 20812 -22568 20828
rect -22672 20748 -22652 20812
rect -22588 20748 -22568 20812
rect -22672 20732 -22568 20748
rect -22672 20668 -22652 20732
rect -22588 20668 -22568 20732
rect -22672 20652 -22568 20668
rect -22672 20588 -22652 20652
rect -22588 20588 -22568 20652
rect -22672 20572 -22568 20588
rect -22672 20508 -22652 20572
rect -22588 20508 -22568 20572
rect -22672 20492 -22568 20508
rect -22672 20428 -22652 20492
rect -22588 20428 -22568 20492
rect -22672 20412 -22568 20428
rect -22672 20348 -22652 20412
rect -22588 20348 -22568 20412
rect -22672 20332 -22568 20348
rect -22672 20268 -22652 20332
rect -22588 20268 -22568 20332
rect -22672 20252 -22568 20268
rect -22672 20188 -22652 20252
rect -22588 20188 -22568 20252
rect -22672 20172 -22568 20188
rect -22672 20108 -22652 20172
rect -22588 20108 -22568 20172
rect -22672 20092 -22568 20108
rect -22672 20028 -22652 20092
rect -22588 20028 -22568 20092
rect -22672 20012 -22568 20028
rect -22672 19948 -22652 20012
rect -22588 19948 -22568 20012
rect -22672 19932 -22568 19948
rect -22672 19868 -22652 19932
rect -22588 19868 -22568 19932
rect -22672 19852 -22568 19868
rect -22672 19788 -22652 19852
rect -22588 19788 -22568 19852
rect -22672 19772 -22568 19788
rect -22672 19708 -22652 19772
rect -22588 19708 -22568 19772
rect -22672 19692 -22568 19708
rect -22672 19628 -22652 19692
rect -22588 19628 -22568 19692
rect -22672 19612 -22568 19628
rect -22672 19548 -22652 19612
rect -22588 19548 -22568 19612
rect -22672 19532 -22568 19548
rect -22672 19468 -22652 19532
rect -22588 19468 -22568 19532
rect -22672 19452 -22568 19468
rect -22672 19388 -22652 19452
rect -22588 19388 -22568 19452
rect -22672 19372 -22568 19388
rect -22672 19308 -22652 19372
rect -22588 19308 -22568 19372
rect -22672 19292 -22568 19308
rect -22672 19228 -22652 19292
rect -22588 19228 -22568 19292
rect -22672 19212 -22568 19228
rect -22672 19148 -22652 19212
rect -22588 19148 -22568 19212
rect -22672 19132 -22568 19148
rect -22672 19068 -22652 19132
rect -22588 19068 -22568 19132
rect -22672 19052 -22568 19068
rect -22672 18988 -22652 19052
rect -22588 18988 -22568 19052
rect -22672 18972 -22568 18988
rect -22672 18908 -22652 18972
rect -22588 18908 -22568 18972
rect -22672 18892 -22568 18908
rect -22672 18828 -22652 18892
rect -22588 18828 -22568 18892
rect -22672 18812 -22568 18828
rect -22672 18748 -22652 18812
rect -22588 18748 -22568 18812
rect -22672 18732 -22568 18748
rect -22672 18668 -22652 18732
rect -22588 18668 -22568 18732
rect -22672 18652 -22568 18668
rect -22672 18588 -22652 18652
rect -22588 18588 -22568 18652
rect -22672 18572 -22568 18588
rect -22672 18508 -22652 18572
rect -22588 18508 -22568 18572
rect -22672 18492 -22568 18508
rect -22672 18428 -22652 18492
rect -22588 18428 -22568 18492
rect -22672 18412 -22568 18428
rect -22672 18348 -22652 18412
rect -22588 18348 -22568 18412
rect -22672 18332 -22568 18348
rect -22672 18268 -22652 18332
rect -22588 18268 -22568 18332
rect -22672 18252 -22568 18268
rect -22672 18188 -22652 18252
rect -22588 18188 -22568 18252
rect -22672 18172 -22568 18188
rect -22672 18108 -22652 18172
rect -22588 18108 -22568 18172
rect -22672 18092 -22568 18108
rect -22672 18028 -22652 18092
rect -22588 18028 -22568 18092
rect -22672 18012 -22568 18028
rect -22672 17948 -22652 18012
rect -22588 17948 -22568 18012
rect -22672 17932 -22568 17948
rect -22672 17868 -22652 17932
rect -22588 17868 -22568 17932
rect -22672 17852 -22568 17868
rect -22672 17788 -22652 17852
rect -22588 17788 -22568 17852
rect -22672 17772 -22568 17788
rect -22672 17708 -22652 17772
rect -22588 17708 -22568 17772
rect -22672 17692 -22568 17708
rect -22672 17628 -22652 17692
rect -22588 17628 -22568 17692
rect -22672 17612 -22568 17628
rect -22672 17548 -22652 17612
rect -22588 17548 -22568 17612
rect -22672 17532 -22568 17548
rect -22672 17468 -22652 17532
rect -22588 17468 -22568 17532
rect -22672 17452 -22568 17468
rect -22672 17388 -22652 17452
rect -22588 17388 -22568 17452
rect -22672 17372 -22568 17388
rect -22672 17308 -22652 17372
rect -22588 17308 -22568 17372
rect -22672 17292 -22568 17308
rect -22672 17228 -22652 17292
rect -22588 17228 -22568 17292
rect -22672 17212 -22568 17228
rect -22672 17148 -22652 17212
rect -22588 17148 -22568 17212
rect -22672 17132 -22568 17148
rect -22672 17068 -22652 17132
rect -22588 17068 -22568 17132
rect -22672 17052 -22568 17068
rect -22672 16988 -22652 17052
rect -22588 16988 -22568 17052
rect -22672 16972 -22568 16988
rect -22672 16908 -22652 16972
rect -22588 16908 -22568 16972
rect -22672 16892 -22568 16908
rect -22672 16828 -22652 16892
rect -22588 16828 -22568 16892
rect -22672 16812 -22568 16828
rect -22672 16748 -22652 16812
rect -22588 16748 -22568 16812
rect -22672 16732 -22568 16748
rect -22672 16668 -22652 16732
rect -22588 16668 -22568 16732
rect -22672 16652 -22568 16668
rect -22672 16588 -22652 16652
rect -22588 16588 -22568 16652
rect -22672 16572 -22568 16588
rect -22672 16508 -22652 16572
rect -22588 16508 -22568 16572
rect -22672 16492 -22568 16508
rect -22672 16428 -22652 16492
rect -22588 16428 -22568 16492
rect -22672 16412 -22568 16428
rect -22672 16348 -22652 16412
rect -22588 16348 -22568 16412
rect -22672 16332 -22568 16348
rect -22672 16268 -22652 16332
rect -22588 16268 -22568 16332
rect -22672 16252 -22568 16268
rect -22672 16188 -22652 16252
rect -22588 16188 -22568 16252
rect -22672 16172 -22568 16188
rect -28284 15812 -28180 16108
rect -33896 15732 -33792 15748
rect -33896 15668 -33876 15732
rect -33812 15668 -33792 15732
rect -33896 15652 -33792 15668
rect -33896 15588 -33876 15652
rect -33812 15588 -33792 15652
rect -33896 15572 -33792 15588
rect -33896 15508 -33876 15572
rect -33812 15508 -33792 15572
rect -33896 15492 -33792 15508
rect -33896 15428 -33876 15492
rect -33812 15428 -33792 15492
rect -33896 15412 -33792 15428
rect -33896 15348 -33876 15412
rect -33812 15348 -33792 15412
rect -33896 15332 -33792 15348
rect -33896 15268 -33876 15332
rect -33812 15268 -33792 15332
rect -33896 15252 -33792 15268
rect -33896 15188 -33876 15252
rect -33812 15188 -33792 15252
rect -33896 15172 -33792 15188
rect -33896 15108 -33876 15172
rect -33812 15108 -33792 15172
rect -33896 15092 -33792 15108
rect -33896 15028 -33876 15092
rect -33812 15028 -33792 15092
rect -33896 15012 -33792 15028
rect -33896 14948 -33876 15012
rect -33812 14948 -33792 15012
rect -33896 14932 -33792 14948
rect -33896 14868 -33876 14932
rect -33812 14868 -33792 14932
rect -33896 14852 -33792 14868
rect -33896 14788 -33876 14852
rect -33812 14788 -33792 14852
rect -33896 14772 -33792 14788
rect -33896 14708 -33876 14772
rect -33812 14708 -33792 14772
rect -33896 14692 -33792 14708
rect -33896 14628 -33876 14692
rect -33812 14628 -33792 14692
rect -33896 14612 -33792 14628
rect -33896 14548 -33876 14612
rect -33812 14548 -33792 14612
rect -33896 14532 -33792 14548
rect -33896 14468 -33876 14532
rect -33812 14468 -33792 14532
rect -33896 14452 -33792 14468
rect -33896 14388 -33876 14452
rect -33812 14388 -33792 14452
rect -33896 14372 -33792 14388
rect -33896 14308 -33876 14372
rect -33812 14308 -33792 14372
rect -33896 14292 -33792 14308
rect -33896 14228 -33876 14292
rect -33812 14228 -33792 14292
rect -33896 14212 -33792 14228
rect -33896 14148 -33876 14212
rect -33812 14148 -33792 14212
rect -33896 14132 -33792 14148
rect -33896 14068 -33876 14132
rect -33812 14068 -33792 14132
rect -33896 14052 -33792 14068
rect -33896 13988 -33876 14052
rect -33812 13988 -33792 14052
rect -33896 13972 -33792 13988
rect -33896 13908 -33876 13972
rect -33812 13908 -33792 13972
rect -33896 13892 -33792 13908
rect -33896 13828 -33876 13892
rect -33812 13828 -33792 13892
rect -33896 13812 -33792 13828
rect -33896 13748 -33876 13812
rect -33812 13748 -33792 13812
rect -33896 13732 -33792 13748
rect -33896 13668 -33876 13732
rect -33812 13668 -33792 13732
rect -33896 13652 -33792 13668
rect -33896 13588 -33876 13652
rect -33812 13588 -33792 13652
rect -33896 13572 -33792 13588
rect -33896 13508 -33876 13572
rect -33812 13508 -33792 13572
rect -33896 13492 -33792 13508
rect -33896 13428 -33876 13492
rect -33812 13428 -33792 13492
rect -33896 13412 -33792 13428
rect -33896 13348 -33876 13412
rect -33812 13348 -33792 13412
rect -33896 13332 -33792 13348
rect -33896 13268 -33876 13332
rect -33812 13268 -33792 13332
rect -33896 13252 -33792 13268
rect -33896 13188 -33876 13252
rect -33812 13188 -33792 13252
rect -33896 13172 -33792 13188
rect -33896 13108 -33876 13172
rect -33812 13108 -33792 13172
rect -33896 13092 -33792 13108
rect -33896 13028 -33876 13092
rect -33812 13028 -33792 13092
rect -33896 13012 -33792 13028
rect -33896 12948 -33876 13012
rect -33812 12948 -33792 13012
rect -33896 12932 -33792 12948
rect -33896 12868 -33876 12932
rect -33812 12868 -33792 12932
rect -33896 12852 -33792 12868
rect -33896 12788 -33876 12852
rect -33812 12788 -33792 12852
rect -33896 12772 -33792 12788
rect -33896 12708 -33876 12772
rect -33812 12708 -33792 12772
rect -33896 12692 -33792 12708
rect -33896 12628 -33876 12692
rect -33812 12628 -33792 12692
rect -33896 12612 -33792 12628
rect -33896 12548 -33876 12612
rect -33812 12548 -33792 12612
rect -33896 12532 -33792 12548
rect -33896 12468 -33876 12532
rect -33812 12468 -33792 12532
rect -33896 12452 -33792 12468
rect -33896 12388 -33876 12452
rect -33812 12388 -33792 12452
rect -33896 12372 -33792 12388
rect -33896 12308 -33876 12372
rect -33812 12308 -33792 12372
rect -33896 12292 -33792 12308
rect -33896 12228 -33876 12292
rect -33812 12228 -33792 12292
rect -33896 12212 -33792 12228
rect -33896 12148 -33876 12212
rect -33812 12148 -33792 12212
rect -33896 12132 -33792 12148
rect -33896 12068 -33876 12132
rect -33812 12068 -33792 12132
rect -33896 12052 -33792 12068
rect -33896 11988 -33876 12052
rect -33812 11988 -33792 12052
rect -33896 11972 -33792 11988
rect -33896 11908 -33876 11972
rect -33812 11908 -33792 11972
rect -33896 11892 -33792 11908
rect -33896 11828 -33876 11892
rect -33812 11828 -33792 11892
rect -33896 11812 -33792 11828
rect -33896 11748 -33876 11812
rect -33812 11748 -33792 11812
rect -33896 11732 -33792 11748
rect -33896 11668 -33876 11732
rect -33812 11668 -33792 11732
rect -33896 11652 -33792 11668
rect -33896 11588 -33876 11652
rect -33812 11588 -33792 11652
rect -33896 11572 -33792 11588
rect -33896 11508 -33876 11572
rect -33812 11508 -33792 11572
rect -33896 11492 -33792 11508
rect -33896 11428 -33876 11492
rect -33812 11428 -33792 11492
rect -33896 11412 -33792 11428
rect -33896 11348 -33876 11412
rect -33812 11348 -33792 11412
rect -33896 11332 -33792 11348
rect -33896 11268 -33876 11332
rect -33812 11268 -33792 11332
rect -33896 11252 -33792 11268
rect -33896 11188 -33876 11252
rect -33812 11188 -33792 11252
rect -33896 11172 -33792 11188
rect -33896 11108 -33876 11172
rect -33812 11108 -33792 11172
rect -33896 11092 -33792 11108
rect -33896 11028 -33876 11092
rect -33812 11028 -33792 11092
rect -33896 11012 -33792 11028
rect -33896 10948 -33876 11012
rect -33812 10948 -33792 11012
rect -33896 10932 -33792 10948
rect -33896 10868 -33876 10932
rect -33812 10868 -33792 10932
rect -33896 10852 -33792 10868
rect -36676 10441 -36572 10839
rect -33896 10788 -33876 10852
rect -33812 10788 -33792 10852
rect -33473 15732 -28551 15761
rect -33473 10868 -33444 15732
rect -28580 10868 -28551 15732
rect -33473 10839 -28551 10868
rect -28284 15748 -28264 15812
rect -28200 15748 -28180 15812
rect -25452 15761 -25348 16159
rect -22672 16108 -22652 16172
rect -22588 16108 -22568 16172
rect -22249 21052 -17327 21081
rect -22249 16188 -22220 21052
rect -17356 16188 -17327 21052
rect -22249 16159 -17327 16188
rect -17060 21068 -17040 21132
rect -16976 21068 -16956 21132
rect -14228 21081 -14124 21479
rect -11448 21428 -11428 21492
rect -11364 21428 -11344 21492
rect -11025 26372 -6103 26401
rect -11025 21508 -10996 26372
rect -6132 21508 -6103 26372
rect -11025 21479 -6103 21508
rect -5836 26388 -5816 26452
rect -5752 26388 -5732 26452
rect -3004 26401 -2900 26799
rect -224 26748 -204 26812
rect -140 26748 -120 26812
rect 199 31692 5121 31721
rect 199 26828 228 31692
rect 5092 26828 5121 31692
rect 199 26799 5121 26828
rect 5388 31708 5408 31772
rect 5472 31708 5492 31772
rect 8220 31721 8324 32119
rect 11000 32068 11020 32132
rect 11084 32068 11104 32132
rect 11423 37012 16345 37041
rect 11423 32148 11452 37012
rect 16316 32148 16345 37012
rect 11423 32119 16345 32148
rect 16612 37028 16632 37092
rect 16696 37028 16716 37092
rect 19444 37041 19548 37240
rect 22224 37092 22328 37240
rect 16612 37012 16716 37028
rect 16612 36948 16632 37012
rect 16696 36948 16716 37012
rect 16612 36932 16716 36948
rect 16612 36868 16632 36932
rect 16696 36868 16716 36932
rect 16612 36852 16716 36868
rect 16612 36788 16632 36852
rect 16696 36788 16716 36852
rect 16612 36772 16716 36788
rect 16612 36708 16632 36772
rect 16696 36708 16716 36772
rect 16612 36692 16716 36708
rect 16612 36628 16632 36692
rect 16696 36628 16716 36692
rect 16612 36612 16716 36628
rect 16612 36548 16632 36612
rect 16696 36548 16716 36612
rect 16612 36532 16716 36548
rect 16612 36468 16632 36532
rect 16696 36468 16716 36532
rect 16612 36452 16716 36468
rect 16612 36388 16632 36452
rect 16696 36388 16716 36452
rect 16612 36372 16716 36388
rect 16612 36308 16632 36372
rect 16696 36308 16716 36372
rect 16612 36292 16716 36308
rect 16612 36228 16632 36292
rect 16696 36228 16716 36292
rect 16612 36212 16716 36228
rect 16612 36148 16632 36212
rect 16696 36148 16716 36212
rect 16612 36132 16716 36148
rect 16612 36068 16632 36132
rect 16696 36068 16716 36132
rect 16612 36052 16716 36068
rect 16612 35988 16632 36052
rect 16696 35988 16716 36052
rect 16612 35972 16716 35988
rect 16612 35908 16632 35972
rect 16696 35908 16716 35972
rect 16612 35892 16716 35908
rect 16612 35828 16632 35892
rect 16696 35828 16716 35892
rect 16612 35812 16716 35828
rect 16612 35748 16632 35812
rect 16696 35748 16716 35812
rect 16612 35732 16716 35748
rect 16612 35668 16632 35732
rect 16696 35668 16716 35732
rect 16612 35652 16716 35668
rect 16612 35588 16632 35652
rect 16696 35588 16716 35652
rect 16612 35572 16716 35588
rect 16612 35508 16632 35572
rect 16696 35508 16716 35572
rect 16612 35492 16716 35508
rect 16612 35428 16632 35492
rect 16696 35428 16716 35492
rect 16612 35412 16716 35428
rect 16612 35348 16632 35412
rect 16696 35348 16716 35412
rect 16612 35332 16716 35348
rect 16612 35268 16632 35332
rect 16696 35268 16716 35332
rect 16612 35252 16716 35268
rect 16612 35188 16632 35252
rect 16696 35188 16716 35252
rect 16612 35172 16716 35188
rect 16612 35108 16632 35172
rect 16696 35108 16716 35172
rect 16612 35092 16716 35108
rect 16612 35028 16632 35092
rect 16696 35028 16716 35092
rect 16612 35012 16716 35028
rect 16612 34948 16632 35012
rect 16696 34948 16716 35012
rect 16612 34932 16716 34948
rect 16612 34868 16632 34932
rect 16696 34868 16716 34932
rect 16612 34852 16716 34868
rect 16612 34788 16632 34852
rect 16696 34788 16716 34852
rect 16612 34772 16716 34788
rect 16612 34708 16632 34772
rect 16696 34708 16716 34772
rect 16612 34692 16716 34708
rect 16612 34628 16632 34692
rect 16696 34628 16716 34692
rect 16612 34612 16716 34628
rect 16612 34548 16632 34612
rect 16696 34548 16716 34612
rect 16612 34532 16716 34548
rect 16612 34468 16632 34532
rect 16696 34468 16716 34532
rect 16612 34452 16716 34468
rect 16612 34388 16632 34452
rect 16696 34388 16716 34452
rect 16612 34372 16716 34388
rect 16612 34308 16632 34372
rect 16696 34308 16716 34372
rect 16612 34292 16716 34308
rect 16612 34228 16632 34292
rect 16696 34228 16716 34292
rect 16612 34212 16716 34228
rect 16612 34148 16632 34212
rect 16696 34148 16716 34212
rect 16612 34132 16716 34148
rect 16612 34068 16632 34132
rect 16696 34068 16716 34132
rect 16612 34052 16716 34068
rect 16612 33988 16632 34052
rect 16696 33988 16716 34052
rect 16612 33972 16716 33988
rect 16612 33908 16632 33972
rect 16696 33908 16716 33972
rect 16612 33892 16716 33908
rect 16612 33828 16632 33892
rect 16696 33828 16716 33892
rect 16612 33812 16716 33828
rect 16612 33748 16632 33812
rect 16696 33748 16716 33812
rect 16612 33732 16716 33748
rect 16612 33668 16632 33732
rect 16696 33668 16716 33732
rect 16612 33652 16716 33668
rect 16612 33588 16632 33652
rect 16696 33588 16716 33652
rect 16612 33572 16716 33588
rect 16612 33508 16632 33572
rect 16696 33508 16716 33572
rect 16612 33492 16716 33508
rect 16612 33428 16632 33492
rect 16696 33428 16716 33492
rect 16612 33412 16716 33428
rect 16612 33348 16632 33412
rect 16696 33348 16716 33412
rect 16612 33332 16716 33348
rect 16612 33268 16632 33332
rect 16696 33268 16716 33332
rect 16612 33252 16716 33268
rect 16612 33188 16632 33252
rect 16696 33188 16716 33252
rect 16612 33172 16716 33188
rect 16612 33108 16632 33172
rect 16696 33108 16716 33172
rect 16612 33092 16716 33108
rect 16612 33028 16632 33092
rect 16696 33028 16716 33092
rect 16612 33012 16716 33028
rect 16612 32948 16632 33012
rect 16696 32948 16716 33012
rect 16612 32932 16716 32948
rect 16612 32868 16632 32932
rect 16696 32868 16716 32932
rect 16612 32852 16716 32868
rect 16612 32788 16632 32852
rect 16696 32788 16716 32852
rect 16612 32772 16716 32788
rect 16612 32708 16632 32772
rect 16696 32708 16716 32772
rect 16612 32692 16716 32708
rect 16612 32628 16632 32692
rect 16696 32628 16716 32692
rect 16612 32612 16716 32628
rect 16612 32548 16632 32612
rect 16696 32548 16716 32612
rect 16612 32532 16716 32548
rect 16612 32468 16632 32532
rect 16696 32468 16716 32532
rect 16612 32452 16716 32468
rect 16612 32388 16632 32452
rect 16696 32388 16716 32452
rect 16612 32372 16716 32388
rect 16612 32308 16632 32372
rect 16696 32308 16716 32372
rect 16612 32292 16716 32308
rect 16612 32228 16632 32292
rect 16696 32228 16716 32292
rect 16612 32212 16716 32228
rect 16612 32148 16632 32212
rect 16696 32148 16716 32212
rect 16612 32132 16716 32148
rect 11000 31772 11104 32068
rect 5388 31692 5492 31708
rect 5388 31628 5408 31692
rect 5472 31628 5492 31692
rect 5388 31612 5492 31628
rect 5388 31548 5408 31612
rect 5472 31548 5492 31612
rect 5388 31532 5492 31548
rect 5388 31468 5408 31532
rect 5472 31468 5492 31532
rect 5388 31452 5492 31468
rect 5388 31388 5408 31452
rect 5472 31388 5492 31452
rect 5388 31372 5492 31388
rect 5388 31308 5408 31372
rect 5472 31308 5492 31372
rect 5388 31292 5492 31308
rect 5388 31228 5408 31292
rect 5472 31228 5492 31292
rect 5388 31212 5492 31228
rect 5388 31148 5408 31212
rect 5472 31148 5492 31212
rect 5388 31132 5492 31148
rect 5388 31068 5408 31132
rect 5472 31068 5492 31132
rect 5388 31052 5492 31068
rect 5388 30988 5408 31052
rect 5472 30988 5492 31052
rect 5388 30972 5492 30988
rect 5388 30908 5408 30972
rect 5472 30908 5492 30972
rect 5388 30892 5492 30908
rect 5388 30828 5408 30892
rect 5472 30828 5492 30892
rect 5388 30812 5492 30828
rect 5388 30748 5408 30812
rect 5472 30748 5492 30812
rect 5388 30732 5492 30748
rect 5388 30668 5408 30732
rect 5472 30668 5492 30732
rect 5388 30652 5492 30668
rect 5388 30588 5408 30652
rect 5472 30588 5492 30652
rect 5388 30572 5492 30588
rect 5388 30508 5408 30572
rect 5472 30508 5492 30572
rect 5388 30492 5492 30508
rect 5388 30428 5408 30492
rect 5472 30428 5492 30492
rect 5388 30412 5492 30428
rect 5388 30348 5408 30412
rect 5472 30348 5492 30412
rect 5388 30332 5492 30348
rect 5388 30268 5408 30332
rect 5472 30268 5492 30332
rect 5388 30252 5492 30268
rect 5388 30188 5408 30252
rect 5472 30188 5492 30252
rect 5388 30172 5492 30188
rect 5388 30108 5408 30172
rect 5472 30108 5492 30172
rect 5388 30092 5492 30108
rect 5388 30028 5408 30092
rect 5472 30028 5492 30092
rect 5388 30012 5492 30028
rect 5388 29948 5408 30012
rect 5472 29948 5492 30012
rect 5388 29932 5492 29948
rect 5388 29868 5408 29932
rect 5472 29868 5492 29932
rect 5388 29852 5492 29868
rect 5388 29788 5408 29852
rect 5472 29788 5492 29852
rect 5388 29772 5492 29788
rect 5388 29708 5408 29772
rect 5472 29708 5492 29772
rect 5388 29692 5492 29708
rect 5388 29628 5408 29692
rect 5472 29628 5492 29692
rect 5388 29612 5492 29628
rect 5388 29548 5408 29612
rect 5472 29548 5492 29612
rect 5388 29532 5492 29548
rect 5388 29468 5408 29532
rect 5472 29468 5492 29532
rect 5388 29452 5492 29468
rect 5388 29388 5408 29452
rect 5472 29388 5492 29452
rect 5388 29372 5492 29388
rect 5388 29308 5408 29372
rect 5472 29308 5492 29372
rect 5388 29292 5492 29308
rect 5388 29228 5408 29292
rect 5472 29228 5492 29292
rect 5388 29212 5492 29228
rect 5388 29148 5408 29212
rect 5472 29148 5492 29212
rect 5388 29132 5492 29148
rect 5388 29068 5408 29132
rect 5472 29068 5492 29132
rect 5388 29052 5492 29068
rect 5388 28988 5408 29052
rect 5472 28988 5492 29052
rect 5388 28972 5492 28988
rect 5388 28908 5408 28972
rect 5472 28908 5492 28972
rect 5388 28892 5492 28908
rect 5388 28828 5408 28892
rect 5472 28828 5492 28892
rect 5388 28812 5492 28828
rect 5388 28748 5408 28812
rect 5472 28748 5492 28812
rect 5388 28732 5492 28748
rect 5388 28668 5408 28732
rect 5472 28668 5492 28732
rect 5388 28652 5492 28668
rect 5388 28588 5408 28652
rect 5472 28588 5492 28652
rect 5388 28572 5492 28588
rect 5388 28508 5408 28572
rect 5472 28508 5492 28572
rect 5388 28492 5492 28508
rect 5388 28428 5408 28492
rect 5472 28428 5492 28492
rect 5388 28412 5492 28428
rect 5388 28348 5408 28412
rect 5472 28348 5492 28412
rect 5388 28332 5492 28348
rect 5388 28268 5408 28332
rect 5472 28268 5492 28332
rect 5388 28252 5492 28268
rect 5388 28188 5408 28252
rect 5472 28188 5492 28252
rect 5388 28172 5492 28188
rect 5388 28108 5408 28172
rect 5472 28108 5492 28172
rect 5388 28092 5492 28108
rect 5388 28028 5408 28092
rect 5472 28028 5492 28092
rect 5388 28012 5492 28028
rect 5388 27948 5408 28012
rect 5472 27948 5492 28012
rect 5388 27932 5492 27948
rect 5388 27868 5408 27932
rect 5472 27868 5492 27932
rect 5388 27852 5492 27868
rect 5388 27788 5408 27852
rect 5472 27788 5492 27852
rect 5388 27772 5492 27788
rect 5388 27708 5408 27772
rect 5472 27708 5492 27772
rect 5388 27692 5492 27708
rect 5388 27628 5408 27692
rect 5472 27628 5492 27692
rect 5388 27612 5492 27628
rect 5388 27548 5408 27612
rect 5472 27548 5492 27612
rect 5388 27532 5492 27548
rect 5388 27468 5408 27532
rect 5472 27468 5492 27532
rect 5388 27452 5492 27468
rect 5388 27388 5408 27452
rect 5472 27388 5492 27452
rect 5388 27372 5492 27388
rect 5388 27308 5408 27372
rect 5472 27308 5492 27372
rect 5388 27292 5492 27308
rect 5388 27228 5408 27292
rect 5472 27228 5492 27292
rect 5388 27212 5492 27228
rect 5388 27148 5408 27212
rect 5472 27148 5492 27212
rect 5388 27132 5492 27148
rect 5388 27068 5408 27132
rect 5472 27068 5492 27132
rect 5388 27052 5492 27068
rect 5388 26988 5408 27052
rect 5472 26988 5492 27052
rect 5388 26972 5492 26988
rect 5388 26908 5408 26972
rect 5472 26908 5492 26972
rect 5388 26892 5492 26908
rect 5388 26828 5408 26892
rect 5472 26828 5492 26892
rect 5388 26812 5492 26828
rect -224 26452 -120 26748
rect -5836 26372 -5732 26388
rect -5836 26308 -5816 26372
rect -5752 26308 -5732 26372
rect -5836 26292 -5732 26308
rect -5836 26228 -5816 26292
rect -5752 26228 -5732 26292
rect -5836 26212 -5732 26228
rect -5836 26148 -5816 26212
rect -5752 26148 -5732 26212
rect -5836 26132 -5732 26148
rect -5836 26068 -5816 26132
rect -5752 26068 -5732 26132
rect -5836 26052 -5732 26068
rect -5836 25988 -5816 26052
rect -5752 25988 -5732 26052
rect -5836 25972 -5732 25988
rect -5836 25908 -5816 25972
rect -5752 25908 -5732 25972
rect -5836 25892 -5732 25908
rect -5836 25828 -5816 25892
rect -5752 25828 -5732 25892
rect -5836 25812 -5732 25828
rect -5836 25748 -5816 25812
rect -5752 25748 -5732 25812
rect -5836 25732 -5732 25748
rect -5836 25668 -5816 25732
rect -5752 25668 -5732 25732
rect -5836 25652 -5732 25668
rect -5836 25588 -5816 25652
rect -5752 25588 -5732 25652
rect -5836 25572 -5732 25588
rect -5836 25508 -5816 25572
rect -5752 25508 -5732 25572
rect -5836 25492 -5732 25508
rect -5836 25428 -5816 25492
rect -5752 25428 -5732 25492
rect -5836 25412 -5732 25428
rect -5836 25348 -5816 25412
rect -5752 25348 -5732 25412
rect -5836 25332 -5732 25348
rect -5836 25268 -5816 25332
rect -5752 25268 -5732 25332
rect -5836 25252 -5732 25268
rect -5836 25188 -5816 25252
rect -5752 25188 -5732 25252
rect -5836 25172 -5732 25188
rect -5836 25108 -5816 25172
rect -5752 25108 -5732 25172
rect -5836 25092 -5732 25108
rect -5836 25028 -5816 25092
rect -5752 25028 -5732 25092
rect -5836 25012 -5732 25028
rect -5836 24948 -5816 25012
rect -5752 24948 -5732 25012
rect -5836 24932 -5732 24948
rect -5836 24868 -5816 24932
rect -5752 24868 -5732 24932
rect -5836 24852 -5732 24868
rect -5836 24788 -5816 24852
rect -5752 24788 -5732 24852
rect -5836 24772 -5732 24788
rect -5836 24708 -5816 24772
rect -5752 24708 -5732 24772
rect -5836 24692 -5732 24708
rect -5836 24628 -5816 24692
rect -5752 24628 -5732 24692
rect -5836 24612 -5732 24628
rect -5836 24548 -5816 24612
rect -5752 24548 -5732 24612
rect -5836 24532 -5732 24548
rect -5836 24468 -5816 24532
rect -5752 24468 -5732 24532
rect -5836 24452 -5732 24468
rect -5836 24388 -5816 24452
rect -5752 24388 -5732 24452
rect -5836 24372 -5732 24388
rect -5836 24308 -5816 24372
rect -5752 24308 -5732 24372
rect -5836 24292 -5732 24308
rect -5836 24228 -5816 24292
rect -5752 24228 -5732 24292
rect -5836 24212 -5732 24228
rect -5836 24148 -5816 24212
rect -5752 24148 -5732 24212
rect -5836 24132 -5732 24148
rect -5836 24068 -5816 24132
rect -5752 24068 -5732 24132
rect -5836 24052 -5732 24068
rect -5836 23988 -5816 24052
rect -5752 23988 -5732 24052
rect -5836 23972 -5732 23988
rect -5836 23908 -5816 23972
rect -5752 23908 -5732 23972
rect -5836 23892 -5732 23908
rect -5836 23828 -5816 23892
rect -5752 23828 -5732 23892
rect -5836 23812 -5732 23828
rect -5836 23748 -5816 23812
rect -5752 23748 -5732 23812
rect -5836 23732 -5732 23748
rect -5836 23668 -5816 23732
rect -5752 23668 -5732 23732
rect -5836 23652 -5732 23668
rect -5836 23588 -5816 23652
rect -5752 23588 -5732 23652
rect -5836 23572 -5732 23588
rect -5836 23508 -5816 23572
rect -5752 23508 -5732 23572
rect -5836 23492 -5732 23508
rect -5836 23428 -5816 23492
rect -5752 23428 -5732 23492
rect -5836 23412 -5732 23428
rect -5836 23348 -5816 23412
rect -5752 23348 -5732 23412
rect -5836 23332 -5732 23348
rect -5836 23268 -5816 23332
rect -5752 23268 -5732 23332
rect -5836 23252 -5732 23268
rect -5836 23188 -5816 23252
rect -5752 23188 -5732 23252
rect -5836 23172 -5732 23188
rect -5836 23108 -5816 23172
rect -5752 23108 -5732 23172
rect -5836 23092 -5732 23108
rect -5836 23028 -5816 23092
rect -5752 23028 -5732 23092
rect -5836 23012 -5732 23028
rect -5836 22948 -5816 23012
rect -5752 22948 -5732 23012
rect -5836 22932 -5732 22948
rect -5836 22868 -5816 22932
rect -5752 22868 -5732 22932
rect -5836 22852 -5732 22868
rect -5836 22788 -5816 22852
rect -5752 22788 -5732 22852
rect -5836 22772 -5732 22788
rect -5836 22708 -5816 22772
rect -5752 22708 -5732 22772
rect -5836 22692 -5732 22708
rect -5836 22628 -5816 22692
rect -5752 22628 -5732 22692
rect -5836 22612 -5732 22628
rect -5836 22548 -5816 22612
rect -5752 22548 -5732 22612
rect -5836 22532 -5732 22548
rect -5836 22468 -5816 22532
rect -5752 22468 -5732 22532
rect -5836 22452 -5732 22468
rect -5836 22388 -5816 22452
rect -5752 22388 -5732 22452
rect -5836 22372 -5732 22388
rect -5836 22308 -5816 22372
rect -5752 22308 -5732 22372
rect -5836 22292 -5732 22308
rect -5836 22228 -5816 22292
rect -5752 22228 -5732 22292
rect -5836 22212 -5732 22228
rect -5836 22148 -5816 22212
rect -5752 22148 -5732 22212
rect -5836 22132 -5732 22148
rect -5836 22068 -5816 22132
rect -5752 22068 -5732 22132
rect -5836 22052 -5732 22068
rect -5836 21988 -5816 22052
rect -5752 21988 -5732 22052
rect -5836 21972 -5732 21988
rect -5836 21908 -5816 21972
rect -5752 21908 -5732 21972
rect -5836 21892 -5732 21908
rect -5836 21828 -5816 21892
rect -5752 21828 -5732 21892
rect -5836 21812 -5732 21828
rect -5836 21748 -5816 21812
rect -5752 21748 -5732 21812
rect -5836 21732 -5732 21748
rect -5836 21668 -5816 21732
rect -5752 21668 -5732 21732
rect -5836 21652 -5732 21668
rect -5836 21588 -5816 21652
rect -5752 21588 -5732 21652
rect -5836 21572 -5732 21588
rect -5836 21508 -5816 21572
rect -5752 21508 -5732 21572
rect -5836 21492 -5732 21508
rect -11448 21132 -11344 21428
rect -17060 21052 -16956 21068
rect -17060 20988 -17040 21052
rect -16976 20988 -16956 21052
rect -17060 20972 -16956 20988
rect -17060 20908 -17040 20972
rect -16976 20908 -16956 20972
rect -17060 20892 -16956 20908
rect -17060 20828 -17040 20892
rect -16976 20828 -16956 20892
rect -17060 20812 -16956 20828
rect -17060 20748 -17040 20812
rect -16976 20748 -16956 20812
rect -17060 20732 -16956 20748
rect -17060 20668 -17040 20732
rect -16976 20668 -16956 20732
rect -17060 20652 -16956 20668
rect -17060 20588 -17040 20652
rect -16976 20588 -16956 20652
rect -17060 20572 -16956 20588
rect -17060 20508 -17040 20572
rect -16976 20508 -16956 20572
rect -17060 20492 -16956 20508
rect -17060 20428 -17040 20492
rect -16976 20428 -16956 20492
rect -17060 20412 -16956 20428
rect -17060 20348 -17040 20412
rect -16976 20348 -16956 20412
rect -17060 20332 -16956 20348
rect -17060 20268 -17040 20332
rect -16976 20268 -16956 20332
rect -17060 20252 -16956 20268
rect -17060 20188 -17040 20252
rect -16976 20188 -16956 20252
rect -17060 20172 -16956 20188
rect -17060 20108 -17040 20172
rect -16976 20108 -16956 20172
rect -17060 20092 -16956 20108
rect -17060 20028 -17040 20092
rect -16976 20028 -16956 20092
rect -17060 20012 -16956 20028
rect -17060 19948 -17040 20012
rect -16976 19948 -16956 20012
rect -17060 19932 -16956 19948
rect -17060 19868 -17040 19932
rect -16976 19868 -16956 19932
rect -17060 19852 -16956 19868
rect -17060 19788 -17040 19852
rect -16976 19788 -16956 19852
rect -17060 19772 -16956 19788
rect -17060 19708 -17040 19772
rect -16976 19708 -16956 19772
rect -17060 19692 -16956 19708
rect -17060 19628 -17040 19692
rect -16976 19628 -16956 19692
rect -17060 19612 -16956 19628
rect -17060 19548 -17040 19612
rect -16976 19548 -16956 19612
rect -17060 19532 -16956 19548
rect -17060 19468 -17040 19532
rect -16976 19468 -16956 19532
rect -17060 19452 -16956 19468
rect -17060 19388 -17040 19452
rect -16976 19388 -16956 19452
rect -17060 19372 -16956 19388
rect -17060 19308 -17040 19372
rect -16976 19308 -16956 19372
rect -17060 19292 -16956 19308
rect -17060 19228 -17040 19292
rect -16976 19228 -16956 19292
rect -17060 19212 -16956 19228
rect -17060 19148 -17040 19212
rect -16976 19148 -16956 19212
rect -17060 19132 -16956 19148
rect -17060 19068 -17040 19132
rect -16976 19068 -16956 19132
rect -17060 19052 -16956 19068
rect -17060 18988 -17040 19052
rect -16976 18988 -16956 19052
rect -17060 18972 -16956 18988
rect -17060 18908 -17040 18972
rect -16976 18908 -16956 18972
rect -17060 18892 -16956 18908
rect -17060 18828 -17040 18892
rect -16976 18828 -16956 18892
rect -17060 18812 -16956 18828
rect -17060 18748 -17040 18812
rect -16976 18748 -16956 18812
rect -17060 18732 -16956 18748
rect -17060 18668 -17040 18732
rect -16976 18668 -16956 18732
rect -17060 18652 -16956 18668
rect -17060 18588 -17040 18652
rect -16976 18588 -16956 18652
rect -17060 18572 -16956 18588
rect -17060 18508 -17040 18572
rect -16976 18508 -16956 18572
rect -17060 18492 -16956 18508
rect -17060 18428 -17040 18492
rect -16976 18428 -16956 18492
rect -17060 18412 -16956 18428
rect -17060 18348 -17040 18412
rect -16976 18348 -16956 18412
rect -17060 18332 -16956 18348
rect -17060 18268 -17040 18332
rect -16976 18268 -16956 18332
rect -17060 18252 -16956 18268
rect -17060 18188 -17040 18252
rect -16976 18188 -16956 18252
rect -17060 18172 -16956 18188
rect -17060 18108 -17040 18172
rect -16976 18108 -16956 18172
rect -17060 18092 -16956 18108
rect -17060 18028 -17040 18092
rect -16976 18028 -16956 18092
rect -17060 18012 -16956 18028
rect -17060 17948 -17040 18012
rect -16976 17948 -16956 18012
rect -17060 17932 -16956 17948
rect -17060 17868 -17040 17932
rect -16976 17868 -16956 17932
rect -17060 17852 -16956 17868
rect -17060 17788 -17040 17852
rect -16976 17788 -16956 17852
rect -17060 17772 -16956 17788
rect -17060 17708 -17040 17772
rect -16976 17708 -16956 17772
rect -17060 17692 -16956 17708
rect -17060 17628 -17040 17692
rect -16976 17628 -16956 17692
rect -17060 17612 -16956 17628
rect -17060 17548 -17040 17612
rect -16976 17548 -16956 17612
rect -17060 17532 -16956 17548
rect -17060 17468 -17040 17532
rect -16976 17468 -16956 17532
rect -17060 17452 -16956 17468
rect -17060 17388 -17040 17452
rect -16976 17388 -16956 17452
rect -17060 17372 -16956 17388
rect -17060 17308 -17040 17372
rect -16976 17308 -16956 17372
rect -17060 17292 -16956 17308
rect -17060 17228 -17040 17292
rect -16976 17228 -16956 17292
rect -17060 17212 -16956 17228
rect -17060 17148 -17040 17212
rect -16976 17148 -16956 17212
rect -17060 17132 -16956 17148
rect -17060 17068 -17040 17132
rect -16976 17068 -16956 17132
rect -17060 17052 -16956 17068
rect -17060 16988 -17040 17052
rect -16976 16988 -16956 17052
rect -17060 16972 -16956 16988
rect -17060 16908 -17040 16972
rect -16976 16908 -16956 16972
rect -17060 16892 -16956 16908
rect -17060 16828 -17040 16892
rect -16976 16828 -16956 16892
rect -17060 16812 -16956 16828
rect -17060 16748 -17040 16812
rect -16976 16748 -16956 16812
rect -17060 16732 -16956 16748
rect -17060 16668 -17040 16732
rect -16976 16668 -16956 16732
rect -17060 16652 -16956 16668
rect -17060 16588 -17040 16652
rect -16976 16588 -16956 16652
rect -17060 16572 -16956 16588
rect -17060 16508 -17040 16572
rect -16976 16508 -16956 16572
rect -17060 16492 -16956 16508
rect -17060 16428 -17040 16492
rect -16976 16428 -16956 16492
rect -17060 16412 -16956 16428
rect -17060 16348 -17040 16412
rect -16976 16348 -16956 16412
rect -17060 16332 -16956 16348
rect -17060 16268 -17040 16332
rect -16976 16268 -16956 16332
rect -17060 16252 -16956 16268
rect -17060 16188 -17040 16252
rect -16976 16188 -16956 16252
rect -17060 16172 -16956 16188
rect -22672 15812 -22568 16108
rect -28284 15732 -28180 15748
rect -28284 15668 -28264 15732
rect -28200 15668 -28180 15732
rect -28284 15652 -28180 15668
rect -28284 15588 -28264 15652
rect -28200 15588 -28180 15652
rect -28284 15572 -28180 15588
rect -28284 15508 -28264 15572
rect -28200 15508 -28180 15572
rect -28284 15492 -28180 15508
rect -28284 15428 -28264 15492
rect -28200 15428 -28180 15492
rect -28284 15412 -28180 15428
rect -28284 15348 -28264 15412
rect -28200 15348 -28180 15412
rect -28284 15332 -28180 15348
rect -28284 15268 -28264 15332
rect -28200 15268 -28180 15332
rect -28284 15252 -28180 15268
rect -28284 15188 -28264 15252
rect -28200 15188 -28180 15252
rect -28284 15172 -28180 15188
rect -28284 15108 -28264 15172
rect -28200 15108 -28180 15172
rect -28284 15092 -28180 15108
rect -28284 15028 -28264 15092
rect -28200 15028 -28180 15092
rect -28284 15012 -28180 15028
rect -28284 14948 -28264 15012
rect -28200 14948 -28180 15012
rect -28284 14932 -28180 14948
rect -28284 14868 -28264 14932
rect -28200 14868 -28180 14932
rect -28284 14852 -28180 14868
rect -28284 14788 -28264 14852
rect -28200 14788 -28180 14852
rect -28284 14772 -28180 14788
rect -28284 14708 -28264 14772
rect -28200 14708 -28180 14772
rect -28284 14692 -28180 14708
rect -28284 14628 -28264 14692
rect -28200 14628 -28180 14692
rect -28284 14612 -28180 14628
rect -28284 14548 -28264 14612
rect -28200 14548 -28180 14612
rect -28284 14532 -28180 14548
rect -28284 14468 -28264 14532
rect -28200 14468 -28180 14532
rect -28284 14452 -28180 14468
rect -28284 14388 -28264 14452
rect -28200 14388 -28180 14452
rect -28284 14372 -28180 14388
rect -28284 14308 -28264 14372
rect -28200 14308 -28180 14372
rect -28284 14292 -28180 14308
rect -28284 14228 -28264 14292
rect -28200 14228 -28180 14292
rect -28284 14212 -28180 14228
rect -28284 14148 -28264 14212
rect -28200 14148 -28180 14212
rect -28284 14132 -28180 14148
rect -28284 14068 -28264 14132
rect -28200 14068 -28180 14132
rect -28284 14052 -28180 14068
rect -28284 13988 -28264 14052
rect -28200 13988 -28180 14052
rect -28284 13972 -28180 13988
rect -28284 13908 -28264 13972
rect -28200 13908 -28180 13972
rect -28284 13892 -28180 13908
rect -28284 13828 -28264 13892
rect -28200 13828 -28180 13892
rect -28284 13812 -28180 13828
rect -28284 13748 -28264 13812
rect -28200 13748 -28180 13812
rect -28284 13732 -28180 13748
rect -28284 13668 -28264 13732
rect -28200 13668 -28180 13732
rect -28284 13652 -28180 13668
rect -28284 13588 -28264 13652
rect -28200 13588 -28180 13652
rect -28284 13572 -28180 13588
rect -28284 13508 -28264 13572
rect -28200 13508 -28180 13572
rect -28284 13492 -28180 13508
rect -28284 13428 -28264 13492
rect -28200 13428 -28180 13492
rect -28284 13412 -28180 13428
rect -28284 13348 -28264 13412
rect -28200 13348 -28180 13412
rect -28284 13332 -28180 13348
rect -28284 13268 -28264 13332
rect -28200 13268 -28180 13332
rect -28284 13252 -28180 13268
rect -28284 13188 -28264 13252
rect -28200 13188 -28180 13252
rect -28284 13172 -28180 13188
rect -28284 13108 -28264 13172
rect -28200 13108 -28180 13172
rect -28284 13092 -28180 13108
rect -28284 13028 -28264 13092
rect -28200 13028 -28180 13092
rect -28284 13012 -28180 13028
rect -28284 12948 -28264 13012
rect -28200 12948 -28180 13012
rect -28284 12932 -28180 12948
rect -28284 12868 -28264 12932
rect -28200 12868 -28180 12932
rect -28284 12852 -28180 12868
rect -28284 12788 -28264 12852
rect -28200 12788 -28180 12852
rect -28284 12772 -28180 12788
rect -28284 12708 -28264 12772
rect -28200 12708 -28180 12772
rect -28284 12692 -28180 12708
rect -28284 12628 -28264 12692
rect -28200 12628 -28180 12692
rect -28284 12612 -28180 12628
rect -28284 12548 -28264 12612
rect -28200 12548 -28180 12612
rect -28284 12532 -28180 12548
rect -28284 12468 -28264 12532
rect -28200 12468 -28180 12532
rect -28284 12452 -28180 12468
rect -28284 12388 -28264 12452
rect -28200 12388 -28180 12452
rect -28284 12372 -28180 12388
rect -28284 12308 -28264 12372
rect -28200 12308 -28180 12372
rect -28284 12292 -28180 12308
rect -28284 12228 -28264 12292
rect -28200 12228 -28180 12292
rect -28284 12212 -28180 12228
rect -28284 12148 -28264 12212
rect -28200 12148 -28180 12212
rect -28284 12132 -28180 12148
rect -28284 12068 -28264 12132
rect -28200 12068 -28180 12132
rect -28284 12052 -28180 12068
rect -28284 11988 -28264 12052
rect -28200 11988 -28180 12052
rect -28284 11972 -28180 11988
rect -28284 11908 -28264 11972
rect -28200 11908 -28180 11972
rect -28284 11892 -28180 11908
rect -28284 11828 -28264 11892
rect -28200 11828 -28180 11892
rect -28284 11812 -28180 11828
rect -28284 11748 -28264 11812
rect -28200 11748 -28180 11812
rect -28284 11732 -28180 11748
rect -28284 11668 -28264 11732
rect -28200 11668 -28180 11732
rect -28284 11652 -28180 11668
rect -28284 11588 -28264 11652
rect -28200 11588 -28180 11652
rect -28284 11572 -28180 11588
rect -28284 11508 -28264 11572
rect -28200 11508 -28180 11572
rect -28284 11492 -28180 11508
rect -28284 11428 -28264 11492
rect -28200 11428 -28180 11492
rect -28284 11412 -28180 11428
rect -28284 11348 -28264 11412
rect -28200 11348 -28180 11412
rect -28284 11332 -28180 11348
rect -28284 11268 -28264 11332
rect -28200 11268 -28180 11332
rect -28284 11252 -28180 11268
rect -28284 11188 -28264 11252
rect -28200 11188 -28180 11252
rect -28284 11172 -28180 11188
rect -28284 11108 -28264 11172
rect -28200 11108 -28180 11172
rect -28284 11092 -28180 11108
rect -28284 11028 -28264 11092
rect -28200 11028 -28180 11092
rect -28284 11012 -28180 11028
rect -28284 10948 -28264 11012
rect -28200 10948 -28180 11012
rect -28284 10932 -28180 10948
rect -28284 10868 -28264 10932
rect -28200 10868 -28180 10932
rect -28284 10852 -28180 10868
rect -33896 10492 -33792 10788
rect -39085 10412 -34163 10441
rect -39085 5548 -39056 10412
rect -34192 5548 -34163 10412
rect -39085 5519 -34163 5548
rect -33896 10428 -33876 10492
rect -33812 10428 -33792 10492
rect -31064 10441 -30960 10839
rect -28284 10788 -28264 10852
rect -28200 10788 -28180 10852
rect -27861 15732 -22939 15761
rect -27861 10868 -27832 15732
rect -22968 10868 -22939 15732
rect -27861 10839 -22939 10868
rect -22672 15748 -22652 15812
rect -22588 15748 -22568 15812
rect -19840 15761 -19736 16159
rect -17060 16108 -17040 16172
rect -16976 16108 -16956 16172
rect -16637 21052 -11715 21081
rect -16637 16188 -16608 21052
rect -11744 16188 -11715 21052
rect -16637 16159 -11715 16188
rect -11448 21068 -11428 21132
rect -11364 21068 -11344 21132
rect -8616 21081 -8512 21479
rect -5836 21428 -5816 21492
rect -5752 21428 -5732 21492
rect -5413 26372 -491 26401
rect -5413 21508 -5384 26372
rect -520 21508 -491 26372
rect -5413 21479 -491 21508
rect -224 26388 -204 26452
rect -140 26388 -120 26452
rect 2608 26401 2712 26799
rect 5388 26748 5408 26812
rect 5472 26748 5492 26812
rect 5811 31692 10733 31721
rect 5811 26828 5840 31692
rect 10704 26828 10733 31692
rect 5811 26799 10733 26828
rect 11000 31708 11020 31772
rect 11084 31708 11104 31772
rect 13832 31721 13936 32119
rect 16612 32068 16632 32132
rect 16696 32068 16716 32132
rect 17035 37012 21957 37041
rect 17035 32148 17064 37012
rect 21928 32148 21957 37012
rect 17035 32119 21957 32148
rect 22224 37028 22244 37092
rect 22308 37028 22328 37092
rect 25056 37041 25160 37240
rect 27836 37092 27940 37240
rect 22224 37012 22328 37028
rect 22224 36948 22244 37012
rect 22308 36948 22328 37012
rect 22224 36932 22328 36948
rect 22224 36868 22244 36932
rect 22308 36868 22328 36932
rect 22224 36852 22328 36868
rect 22224 36788 22244 36852
rect 22308 36788 22328 36852
rect 22224 36772 22328 36788
rect 22224 36708 22244 36772
rect 22308 36708 22328 36772
rect 22224 36692 22328 36708
rect 22224 36628 22244 36692
rect 22308 36628 22328 36692
rect 22224 36612 22328 36628
rect 22224 36548 22244 36612
rect 22308 36548 22328 36612
rect 22224 36532 22328 36548
rect 22224 36468 22244 36532
rect 22308 36468 22328 36532
rect 22224 36452 22328 36468
rect 22224 36388 22244 36452
rect 22308 36388 22328 36452
rect 22224 36372 22328 36388
rect 22224 36308 22244 36372
rect 22308 36308 22328 36372
rect 22224 36292 22328 36308
rect 22224 36228 22244 36292
rect 22308 36228 22328 36292
rect 22224 36212 22328 36228
rect 22224 36148 22244 36212
rect 22308 36148 22328 36212
rect 22224 36132 22328 36148
rect 22224 36068 22244 36132
rect 22308 36068 22328 36132
rect 22224 36052 22328 36068
rect 22224 35988 22244 36052
rect 22308 35988 22328 36052
rect 22224 35972 22328 35988
rect 22224 35908 22244 35972
rect 22308 35908 22328 35972
rect 22224 35892 22328 35908
rect 22224 35828 22244 35892
rect 22308 35828 22328 35892
rect 22224 35812 22328 35828
rect 22224 35748 22244 35812
rect 22308 35748 22328 35812
rect 22224 35732 22328 35748
rect 22224 35668 22244 35732
rect 22308 35668 22328 35732
rect 22224 35652 22328 35668
rect 22224 35588 22244 35652
rect 22308 35588 22328 35652
rect 22224 35572 22328 35588
rect 22224 35508 22244 35572
rect 22308 35508 22328 35572
rect 22224 35492 22328 35508
rect 22224 35428 22244 35492
rect 22308 35428 22328 35492
rect 22224 35412 22328 35428
rect 22224 35348 22244 35412
rect 22308 35348 22328 35412
rect 22224 35332 22328 35348
rect 22224 35268 22244 35332
rect 22308 35268 22328 35332
rect 22224 35252 22328 35268
rect 22224 35188 22244 35252
rect 22308 35188 22328 35252
rect 22224 35172 22328 35188
rect 22224 35108 22244 35172
rect 22308 35108 22328 35172
rect 22224 35092 22328 35108
rect 22224 35028 22244 35092
rect 22308 35028 22328 35092
rect 22224 35012 22328 35028
rect 22224 34948 22244 35012
rect 22308 34948 22328 35012
rect 22224 34932 22328 34948
rect 22224 34868 22244 34932
rect 22308 34868 22328 34932
rect 22224 34852 22328 34868
rect 22224 34788 22244 34852
rect 22308 34788 22328 34852
rect 22224 34772 22328 34788
rect 22224 34708 22244 34772
rect 22308 34708 22328 34772
rect 22224 34692 22328 34708
rect 22224 34628 22244 34692
rect 22308 34628 22328 34692
rect 22224 34612 22328 34628
rect 22224 34548 22244 34612
rect 22308 34548 22328 34612
rect 22224 34532 22328 34548
rect 22224 34468 22244 34532
rect 22308 34468 22328 34532
rect 22224 34452 22328 34468
rect 22224 34388 22244 34452
rect 22308 34388 22328 34452
rect 22224 34372 22328 34388
rect 22224 34308 22244 34372
rect 22308 34308 22328 34372
rect 22224 34292 22328 34308
rect 22224 34228 22244 34292
rect 22308 34228 22328 34292
rect 22224 34212 22328 34228
rect 22224 34148 22244 34212
rect 22308 34148 22328 34212
rect 22224 34132 22328 34148
rect 22224 34068 22244 34132
rect 22308 34068 22328 34132
rect 22224 34052 22328 34068
rect 22224 33988 22244 34052
rect 22308 33988 22328 34052
rect 22224 33972 22328 33988
rect 22224 33908 22244 33972
rect 22308 33908 22328 33972
rect 22224 33892 22328 33908
rect 22224 33828 22244 33892
rect 22308 33828 22328 33892
rect 22224 33812 22328 33828
rect 22224 33748 22244 33812
rect 22308 33748 22328 33812
rect 22224 33732 22328 33748
rect 22224 33668 22244 33732
rect 22308 33668 22328 33732
rect 22224 33652 22328 33668
rect 22224 33588 22244 33652
rect 22308 33588 22328 33652
rect 22224 33572 22328 33588
rect 22224 33508 22244 33572
rect 22308 33508 22328 33572
rect 22224 33492 22328 33508
rect 22224 33428 22244 33492
rect 22308 33428 22328 33492
rect 22224 33412 22328 33428
rect 22224 33348 22244 33412
rect 22308 33348 22328 33412
rect 22224 33332 22328 33348
rect 22224 33268 22244 33332
rect 22308 33268 22328 33332
rect 22224 33252 22328 33268
rect 22224 33188 22244 33252
rect 22308 33188 22328 33252
rect 22224 33172 22328 33188
rect 22224 33108 22244 33172
rect 22308 33108 22328 33172
rect 22224 33092 22328 33108
rect 22224 33028 22244 33092
rect 22308 33028 22328 33092
rect 22224 33012 22328 33028
rect 22224 32948 22244 33012
rect 22308 32948 22328 33012
rect 22224 32932 22328 32948
rect 22224 32868 22244 32932
rect 22308 32868 22328 32932
rect 22224 32852 22328 32868
rect 22224 32788 22244 32852
rect 22308 32788 22328 32852
rect 22224 32772 22328 32788
rect 22224 32708 22244 32772
rect 22308 32708 22328 32772
rect 22224 32692 22328 32708
rect 22224 32628 22244 32692
rect 22308 32628 22328 32692
rect 22224 32612 22328 32628
rect 22224 32548 22244 32612
rect 22308 32548 22328 32612
rect 22224 32532 22328 32548
rect 22224 32468 22244 32532
rect 22308 32468 22328 32532
rect 22224 32452 22328 32468
rect 22224 32388 22244 32452
rect 22308 32388 22328 32452
rect 22224 32372 22328 32388
rect 22224 32308 22244 32372
rect 22308 32308 22328 32372
rect 22224 32292 22328 32308
rect 22224 32228 22244 32292
rect 22308 32228 22328 32292
rect 22224 32212 22328 32228
rect 22224 32148 22244 32212
rect 22308 32148 22328 32212
rect 22224 32132 22328 32148
rect 16612 31772 16716 32068
rect 11000 31692 11104 31708
rect 11000 31628 11020 31692
rect 11084 31628 11104 31692
rect 11000 31612 11104 31628
rect 11000 31548 11020 31612
rect 11084 31548 11104 31612
rect 11000 31532 11104 31548
rect 11000 31468 11020 31532
rect 11084 31468 11104 31532
rect 11000 31452 11104 31468
rect 11000 31388 11020 31452
rect 11084 31388 11104 31452
rect 11000 31372 11104 31388
rect 11000 31308 11020 31372
rect 11084 31308 11104 31372
rect 11000 31292 11104 31308
rect 11000 31228 11020 31292
rect 11084 31228 11104 31292
rect 11000 31212 11104 31228
rect 11000 31148 11020 31212
rect 11084 31148 11104 31212
rect 11000 31132 11104 31148
rect 11000 31068 11020 31132
rect 11084 31068 11104 31132
rect 11000 31052 11104 31068
rect 11000 30988 11020 31052
rect 11084 30988 11104 31052
rect 11000 30972 11104 30988
rect 11000 30908 11020 30972
rect 11084 30908 11104 30972
rect 11000 30892 11104 30908
rect 11000 30828 11020 30892
rect 11084 30828 11104 30892
rect 11000 30812 11104 30828
rect 11000 30748 11020 30812
rect 11084 30748 11104 30812
rect 11000 30732 11104 30748
rect 11000 30668 11020 30732
rect 11084 30668 11104 30732
rect 11000 30652 11104 30668
rect 11000 30588 11020 30652
rect 11084 30588 11104 30652
rect 11000 30572 11104 30588
rect 11000 30508 11020 30572
rect 11084 30508 11104 30572
rect 11000 30492 11104 30508
rect 11000 30428 11020 30492
rect 11084 30428 11104 30492
rect 11000 30412 11104 30428
rect 11000 30348 11020 30412
rect 11084 30348 11104 30412
rect 11000 30332 11104 30348
rect 11000 30268 11020 30332
rect 11084 30268 11104 30332
rect 11000 30252 11104 30268
rect 11000 30188 11020 30252
rect 11084 30188 11104 30252
rect 11000 30172 11104 30188
rect 11000 30108 11020 30172
rect 11084 30108 11104 30172
rect 11000 30092 11104 30108
rect 11000 30028 11020 30092
rect 11084 30028 11104 30092
rect 11000 30012 11104 30028
rect 11000 29948 11020 30012
rect 11084 29948 11104 30012
rect 11000 29932 11104 29948
rect 11000 29868 11020 29932
rect 11084 29868 11104 29932
rect 11000 29852 11104 29868
rect 11000 29788 11020 29852
rect 11084 29788 11104 29852
rect 11000 29772 11104 29788
rect 11000 29708 11020 29772
rect 11084 29708 11104 29772
rect 11000 29692 11104 29708
rect 11000 29628 11020 29692
rect 11084 29628 11104 29692
rect 11000 29612 11104 29628
rect 11000 29548 11020 29612
rect 11084 29548 11104 29612
rect 11000 29532 11104 29548
rect 11000 29468 11020 29532
rect 11084 29468 11104 29532
rect 11000 29452 11104 29468
rect 11000 29388 11020 29452
rect 11084 29388 11104 29452
rect 11000 29372 11104 29388
rect 11000 29308 11020 29372
rect 11084 29308 11104 29372
rect 11000 29292 11104 29308
rect 11000 29228 11020 29292
rect 11084 29228 11104 29292
rect 11000 29212 11104 29228
rect 11000 29148 11020 29212
rect 11084 29148 11104 29212
rect 11000 29132 11104 29148
rect 11000 29068 11020 29132
rect 11084 29068 11104 29132
rect 11000 29052 11104 29068
rect 11000 28988 11020 29052
rect 11084 28988 11104 29052
rect 11000 28972 11104 28988
rect 11000 28908 11020 28972
rect 11084 28908 11104 28972
rect 11000 28892 11104 28908
rect 11000 28828 11020 28892
rect 11084 28828 11104 28892
rect 11000 28812 11104 28828
rect 11000 28748 11020 28812
rect 11084 28748 11104 28812
rect 11000 28732 11104 28748
rect 11000 28668 11020 28732
rect 11084 28668 11104 28732
rect 11000 28652 11104 28668
rect 11000 28588 11020 28652
rect 11084 28588 11104 28652
rect 11000 28572 11104 28588
rect 11000 28508 11020 28572
rect 11084 28508 11104 28572
rect 11000 28492 11104 28508
rect 11000 28428 11020 28492
rect 11084 28428 11104 28492
rect 11000 28412 11104 28428
rect 11000 28348 11020 28412
rect 11084 28348 11104 28412
rect 11000 28332 11104 28348
rect 11000 28268 11020 28332
rect 11084 28268 11104 28332
rect 11000 28252 11104 28268
rect 11000 28188 11020 28252
rect 11084 28188 11104 28252
rect 11000 28172 11104 28188
rect 11000 28108 11020 28172
rect 11084 28108 11104 28172
rect 11000 28092 11104 28108
rect 11000 28028 11020 28092
rect 11084 28028 11104 28092
rect 11000 28012 11104 28028
rect 11000 27948 11020 28012
rect 11084 27948 11104 28012
rect 11000 27932 11104 27948
rect 11000 27868 11020 27932
rect 11084 27868 11104 27932
rect 11000 27852 11104 27868
rect 11000 27788 11020 27852
rect 11084 27788 11104 27852
rect 11000 27772 11104 27788
rect 11000 27708 11020 27772
rect 11084 27708 11104 27772
rect 11000 27692 11104 27708
rect 11000 27628 11020 27692
rect 11084 27628 11104 27692
rect 11000 27612 11104 27628
rect 11000 27548 11020 27612
rect 11084 27548 11104 27612
rect 11000 27532 11104 27548
rect 11000 27468 11020 27532
rect 11084 27468 11104 27532
rect 11000 27452 11104 27468
rect 11000 27388 11020 27452
rect 11084 27388 11104 27452
rect 11000 27372 11104 27388
rect 11000 27308 11020 27372
rect 11084 27308 11104 27372
rect 11000 27292 11104 27308
rect 11000 27228 11020 27292
rect 11084 27228 11104 27292
rect 11000 27212 11104 27228
rect 11000 27148 11020 27212
rect 11084 27148 11104 27212
rect 11000 27132 11104 27148
rect 11000 27068 11020 27132
rect 11084 27068 11104 27132
rect 11000 27052 11104 27068
rect 11000 26988 11020 27052
rect 11084 26988 11104 27052
rect 11000 26972 11104 26988
rect 11000 26908 11020 26972
rect 11084 26908 11104 26972
rect 11000 26892 11104 26908
rect 11000 26828 11020 26892
rect 11084 26828 11104 26892
rect 11000 26812 11104 26828
rect 5388 26452 5492 26748
rect -224 26372 -120 26388
rect -224 26308 -204 26372
rect -140 26308 -120 26372
rect -224 26292 -120 26308
rect -224 26228 -204 26292
rect -140 26228 -120 26292
rect -224 26212 -120 26228
rect -224 26148 -204 26212
rect -140 26148 -120 26212
rect -224 26132 -120 26148
rect -224 26068 -204 26132
rect -140 26068 -120 26132
rect -224 26052 -120 26068
rect -224 25988 -204 26052
rect -140 25988 -120 26052
rect -224 25972 -120 25988
rect -224 25908 -204 25972
rect -140 25908 -120 25972
rect -224 25892 -120 25908
rect -224 25828 -204 25892
rect -140 25828 -120 25892
rect -224 25812 -120 25828
rect -224 25748 -204 25812
rect -140 25748 -120 25812
rect -224 25732 -120 25748
rect -224 25668 -204 25732
rect -140 25668 -120 25732
rect -224 25652 -120 25668
rect -224 25588 -204 25652
rect -140 25588 -120 25652
rect -224 25572 -120 25588
rect -224 25508 -204 25572
rect -140 25508 -120 25572
rect -224 25492 -120 25508
rect -224 25428 -204 25492
rect -140 25428 -120 25492
rect -224 25412 -120 25428
rect -224 25348 -204 25412
rect -140 25348 -120 25412
rect -224 25332 -120 25348
rect -224 25268 -204 25332
rect -140 25268 -120 25332
rect -224 25252 -120 25268
rect -224 25188 -204 25252
rect -140 25188 -120 25252
rect -224 25172 -120 25188
rect -224 25108 -204 25172
rect -140 25108 -120 25172
rect -224 25092 -120 25108
rect -224 25028 -204 25092
rect -140 25028 -120 25092
rect -224 25012 -120 25028
rect -224 24948 -204 25012
rect -140 24948 -120 25012
rect -224 24932 -120 24948
rect -224 24868 -204 24932
rect -140 24868 -120 24932
rect -224 24852 -120 24868
rect -224 24788 -204 24852
rect -140 24788 -120 24852
rect -224 24772 -120 24788
rect -224 24708 -204 24772
rect -140 24708 -120 24772
rect -224 24692 -120 24708
rect -224 24628 -204 24692
rect -140 24628 -120 24692
rect -224 24612 -120 24628
rect -224 24548 -204 24612
rect -140 24548 -120 24612
rect -224 24532 -120 24548
rect -224 24468 -204 24532
rect -140 24468 -120 24532
rect -224 24452 -120 24468
rect -224 24388 -204 24452
rect -140 24388 -120 24452
rect -224 24372 -120 24388
rect -224 24308 -204 24372
rect -140 24308 -120 24372
rect -224 24292 -120 24308
rect -224 24228 -204 24292
rect -140 24228 -120 24292
rect -224 24212 -120 24228
rect -224 24148 -204 24212
rect -140 24148 -120 24212
rect -224 24132 -120 24148
rect -224 24068 -204 24132
rect -140 24068 -120 24132
rect -224 24052 -120 24068
rect -224 23988 -204 24052
rect -140 23988 -120 24052
rect -224 23972 -120 23988
rect -224 23908 -204 23972
rect -140 23908 -120 23972
rect -224 23892 -120 23908
rect -224 23828 -204 23892
rect -140 23828 -120 23892
rect -224 23812 -120 23828
rect -224 23748 -204 23812
rect -140 23748 -120 23812
rect -224 23732 -120 23748
rect -224 23668 -204 23732
rect -140 23668 -120 23732
rect -224 23652 -120 23668
rect -224 23588 -204 23652
rect -140 23588 -120 23652
rect -224 23572 -120 23588
rect -224 23508 -204 23572
rect -140 23508 -120 23572
rect -224 23492 -120 23508
rect -224 23428 -204 23492
rect -140 23428 -120 23492
rect -224 23412 -120 23428
rect -224 23348 -204 23412
rect -140 23348 -120 23412
rect -224 23332 -120 23348
rect -224 23268 -204 23332
rect -140 23268 -120 23332
rect -224 23252 -120 23268
rect -224 23188 -204 23252
rect -140 23188 -120 23252
rect -224 23172 -120 23188
rect -224 23108 -204 23172
rect -140 23108 -120 23172
rect -224 23092 -120 23108
rect -224 23028 -204 23092
rect -140 23028 -120 23092
rect -224 23012 -120 23028
rect -224 22948 -204 23012
rect -140 22948 -120 23012
rect -224 22932 -120 22948
rect -224 22868 -204 22932
rect -140 22868 -120 22932
rect -224 22852 -120 22868
rect -224 22788 -204 22852
rect -140 22788 -120 22852
rect -224 22772 -120 22788
rect -224 22708 -204 22772
rect -140 22708 -120 22772
rect -224 22692 -120 22708
rect -224 22628 -204 22692
rect -140 22628 -120 22692
rect -224 22612 -120 22628
rect -224 22548 -204 22612
rect -140 22548 -120 22612
rect -224 22532 -120 22548
rect -224 22468 -204 22532
rect -140 22468 -120 22532
rect -224 22452 -120 22468
rect -224 22388 -204 22452
rect -140 22388 -120 22452
rect -224 22372 -120 22388
rect -224 22308 -204 22372
rect -140 22308 -120 22372
rect -224 22292 -120 22308
rect -224 22228 -204 22292
rect -140 22228 -120 22292
rect -224 22212 -120 22228
rect -224 22148 -204 22212
rect -140 22148 -120 22212
rect -224 22132 -120 22148
rect -224 22068 -204 22132
rect -140 22068 -120 22132
rect -224 22052 -120 22068
rect -224 21988 -204 22052
rect -140 21988 -120 22052
rect -224 21972 -120 21988
rect -224 21908 -204 21972
rect -140 21908 -120 21972
rect -224 21892 -120 21908
rect -224 21828 -204 21892
rect -140 21828 -120 21892
rect -224 21812 -120 21828
rect -224 21748 -204 21812
rect -140 21748 -120 21812
rect -224 21732 -120 21748
rect -224 21668 -204 21732
rect -140 21668 -120 21732
rect -224 21652 -120 21668
rect -224 21588 -204 21652
rect -140 21588 -120 21652
rect -224 21572 -120 21588
rect -224 21508 -204 21572
rect -140 21508 -120 21572
rect -224 21492 -120 21508
rect -5836 21132 -5732 21428
rect -11448 21052 -11344 21068
rect -11448 20988 -11428 21052
rect -11364 20988 -11344 21052
rect -11448 20972 -11344 20988
rect -11448 20908 -11428 20972
rect -11364 20908 -11344 20972
rect -11448 20892 -11344 20908
rect -11448 20828 -11428 20892
rect -11364 20828 -11344 20892
rect -11448 20812 -11344 20828
rect -11448 20748 -11428 20812
rect -11364 20748 -11344 20812
rect -11448 20732 -11344 20748
rect -11448 20668 -11428 20732
rect -11364 20668 -11344 20732
rect -11448 20652 -11344 20668
rect -11448 20588 -11428 20652
rect -11364 20588 -11344 20652
rect -11448 20572 -11344 20588
rect -11448 20508 -11428 20572
rect -11364 20508 -11344 20572
rect -11448 20492 -11344 20508
rect -11448 20428 -11428 20492
rect -11364 20428 -11344 20492
rect -11448 20412 -11344 20428
rect -11448 20348 -11428 20412
rect -11364 20348 -11344 20412
rect -11448 20332 -11344 20348
rect -11448 20268 -11428 20332
rect -11364 20268 -11344 20332
rect -11448 20252 -11344 20268
rect -11448 20188 -11428 20252
rect -11364 20188 -11344 20252
rect -11448 20172 -11344 20188
rect -11448 20108 -11428 20172
rect -11364 20108 -11344 20172
rect -11448 20092 -11344 20108
rect -11448 20028 -11428 20092
rect -11364 20028 -11344 20092
rect -11448 20012 -11344 20028
rect -11448 19948 -11428 20012
rect -11364 19948 -11344 20012
rect -11448 19932 -11344 19948
rect -11448 19868 -11428 19932
rect -11364 19868 -11344 19932
rect -11448 19852 -11344 19868
rect -11448 19788 -11428 19852
rect -11364 19788 -11344 19852
rect -11448 19772 -11344 19788
rect -11448 19708 -11428 19772
rect -11364 19708 -11344 19772
rect -11448 19692 -11344 19708
rect -11448 19628 -11428 19692
rect -11364 19628 -11344 19692
rect -11448 19612 -11344 19628
rect -11448 19548 -11428 19612
rect -11364 19548 -11344 19612
rect -11448 19532 -11344 19548
rect -11448 19468 -11428 19532
rect -11364 19468 -11344 19532
rect -11448 19452 -11344 19468
rect -11448 19388 -11428 19452
rect -11364 19388 -11344 19452
rect -11448 19372 -11344 19388
rect -11448 19308 -11428 19372
rect -11364 19308 -11344 19372
rect -11448 19292 -11344 19308
rect -11448 19228 -11428 19292
rect -11364 19228 -11344 19292
rect -11448 19212 -11344 19228
rect -11448 19148 -11428 19212
rect -11364 19148 -11344 19212
rect -11448 19132 -11344 19148
rect -11448 19068 -11428 19132
rect -11364 19068 -11344 19132
rect -11448 19052 -11344 19068
rect -11448 18988 -11428 19052
rect -11364 18988 -11344 19052
rect -11448 18972 -11344 18988
rect -11448 18908 -11428 18972
rect -11364 18908 -11344 18972
rect -11448 18892 -11344 18908
rect -11448 18828 -11428 18892
rect -11364 18828 -11344 18892
rect -11448 18812 -11344 18828
rect -11448 18748 -11428 18812
rect -11364 18748 -11344 18812
rect -11448 18732 -11344 18748
rect -11448 18668 -11428 18732
rect -11364 18668 -11344 18732
rect -11448 18652 -11344 18668
rect -11448 18588 -11428 18652
rect -11364 18588 -11344 18652
rect -11448 18572 -11344 18588
rect -11448 18508 -11428 18572
rect -11364 18508 -11344 18572
rect -11448 18492 -11344 18508
rect -11448 18428 -11428 18492
rect -11364 18428 -11344 18492
rect -11448 18412 -11344 18428
rect -11448 18348 -11428 18412
rect -11364 18348 -11344 18412
rect -11448 18332 -11344 18348
rect -11448 18268 -11428 18332
rect -11364 18268 -11344 18332
rect -11448 18252 -11344 18268
rect -11448 18188 -11428 18252
rect -11364 18188 -11344 18252
rect -11448 18172 -11344 18188
rect -11448 18108 -11428 18172
rect -11364 18108 -11344 18172
rect -11448 18092 -11344 18108
rect -11448 18028 -11428 18092
rect -11364 18028 -11344 18092
rect -11448 18012 -11344 18028
rect -11448 17948 -11428 18012
rect -11364 17948 -11344 18012
rect -11448 17932 -11344 17948
rect -11448 17868 -11428 17932
rect -11364 17868 -11344 17932
rect -11448 17852 -11344 17868
rect -11448 17788 -11428 17852
rect -11364 17788 -11344 17852
rect -11448 17772 -11344 17788
rect -11448 17708 -11428 17772
rect -11364 17708 -11344 17772
rect -11448 17692 -11344 17708
rect -11448 17628 -11428 17692
rect -11364 17628 -11344 17692
rect -11448 17612 -11344 17628
rect -11448 17548 -11428 17612
rect -11364 17548 -11344 17612
rect -11448 17532 -11344 17548
rect -11448 17468 -11428 17532
rect -11364 17468 -11344 17532
rect -11448 17452 -11344 17468
rect -11448 17388 -11428 17452
rect -11364 17388 -11344 17452
rect -11448 17372 -11344 17388
rect -11448 17308 -11428 17372
rect -11364 17308 -11344 17372
rect -11448 17292 -11344 17308
rect -11448 17228 -11428 17292
rect -11364 17228 -11344 17292
rect -11448 17212 -11344 17228
rect -11448 17148 -11428 17212
rect -11364 17148 -11344 17212
rect -11448 17132 -11344 17148
rect -11448 17068 -11428 17132
rect -11364 17068 -11344 17132
rect -11448 17052 -11344 17068
rect -11448 16988 -11428 17052
rect -11364 16988 -11344 17052
rect -11448 16972 -11344 16988
rect -11448 16908 -11428 16972
rect -11364 16908 -11344 16972
rect -11448 16892 -11344 16908
rect -11448 16828 -11428 16892
rect -11364 16828 -11344 16892
rect -11448 16812 -11344 16828
rect -11448 16748 -11428 16812
rect -11364 16748 -11344 16812
rect -11448 16732 -11344 16748
rect -11448 16668 -11428 16732
rect -11364 16668 -11344 16732
rect -11448 16652 -11344 16668
rect -11448 16588 -11428 16652
rect -11364 16588 -11344 16652
rect -11448 16572 -11344 16588
rect -11448 16508 -11428 16572
rect -11364 16508 -11344 16572
rect -11448 16492 -11344 16508
rect -11448 16428 -11428 16492
rect -11364 16428 -11344 16492
rect -11448 16412 -11344 16428
rect -11448 16348 -11428 16412
rect -11364 16348 -11344 16412
rect -11448 16332 -11344 16348
rect -11448 16268 -11428 16332
rect -11364 16268 -11344 16332
rect -11448 16252 -11344 16268
rect -11448 16188 -11428 16252
rect -11364 16188 -11344 16252
rect -11448 16172 -11344 16188
rect -17060 15812 -16956 16108
rect -22672 15732 -22568 15748
rect -22672 15668 -22652 15732
rect -22588 15668 -22568 15732
rect -22672 15652 -22568 15668
rect -22672 15588 -22652 15652
rect -22588 15588 -22568 15652
rect -22672 15572 -22568 15588
rect -22672 15508 -22652 15572
rect -22588 15508 -22568 15572
rect -22672 15492 -22568 15508
rect -22672 15428 -22652 15492
rect -22588 15428 -22568 15492
rect -22672 15412 -22568 15428
rect -22672 15348 -22652 15412
rect -22588 15348 -22568 15412
rect -22672 15332 -22568 15348
rect -22672 15268 -22652 15332
rect -22588 15268 -22568 15332
rect -22672 15252 -22568 15268
rect -22672 15188 -22652 15252
rect -22588 15188 -22568 15252
rect -22672 15172 -22568 15188
rect -22672 15108 -22652 15172
rect -22588 15108 -22568 15172
rect -22672 15092 -22568 15108
rect -22672 15028 -22652 15092
rect -22588 15028 -22568 15092
rect -22672 15012 -22568 15028
rect -22672 14948 -22652 15012
rect -22588 14948 -22568 15012
rect -22672 14932 -22568 14948
rect -22672 14868 -22652 14932
rect -22588 14868 -22568 14932
rect -22672 14852 -22568 14868
rect -22672 14788 -22652 14852
rect -22588 14788 -22568 14852
rect -22672 14772 -22568 14788
rect -22672 14708 -22652 14772
rect -22588 14708 -22568 14772
rect -22672 14692 -22568 14708
rect -22672 14628 -22652 14692
rect -22588 14628 -22568 14692
rect -22672 14612 -22568 14628
rect -22672 14548 -22652 14612
rect -22588 14548 -22568 14612
rect -22672 14532 -22568 14548
rect -22672 14468 -22652 14532
rect -22588 14468 -22568 14532
rect -22672 14452 -22568 14468
rect -22672 14388 -22652 14452
rect -22588 14388 -22568 14452
rect -22672 14372 -22568 14388
rect -22672 14308 -22652 14372
rect -22588 14308 -22568 14372
rect -22672 14292 -22568 14308
rect -22672 14228 -22652 14292
rect -22588 14228 -22568 14292
rect -22672 14212 -22568 14228
rect -22672 14148 -22652 14212
rect -22588 14148 -22568 14212
rect -22672 14132 -22568 14148
rect -22672 14068 -22652 14132
rect -22588 14068 -22568 14132
rect -22672 14052 -22568 14068
rect -22672 13988 -22652 14052
rect -22588 13988 -22568 14052
rect -22672 13972 -22568 13988
rect -22672 13908 -22652 13972
rect -22588 13908 -22568 13972
rect -22672 13892 -22568 13908
rect -22672 13828 -22652 13892
rect -22588 13828 -22568 13892
rect -22672 13812 -22568 13828
rect -22672 13748 -22652 13812
rect -22588 13748 -22568 13812
rect -22672 13732 -22568 13748
rect -22672 13668 -22652 13732
rect -22588 13668 -22568 13732
rect -22672 13652 -22568 13668
rect -22672 13588 -22652 13652
rect -22588 13588 -22568 13652
rect -22672 13572 -22568 13588
rect -22672 13508 -22652 13572
rect -22588 13508 -22568 13572
rect -22672 13492 -22568 13508
rect -22672 13428 -22652 13492
rect -22588 13428 -22568 13492
rect -22672 13412 -22568 13428
rect -22672 13348 -22652 13412
rect -22588 13348 -22568 13412
rect -22672 13332 -22568 13348
rect -22672 13268 -22652 13332
rect -22588 13268 -22568 13332
rect -22672 13252 -22568 13268
rect -22672 13188 -22652 13252
rect -22588 13188 -22568 13252
rect -22672 13172 -22568 13188
rect -22672 13108 -22652 13172
rect -22588 13108 -22568 13172
rect -22672 13092 -22568 13108
rect -22672 13028 -22652 13092
rect -22588 13028 -22568 13092
rect -22672 13012 -22568 13028
rect -22672 12948 -22652 13012
rect -22588 12948 -22568 13012
rect -22672 12932 -22568 12948
rect -22672 12868 -22652 12932
rect -22588 12868 -22568 12932
rect -22672 12852 -22568 12868
rect -22672 12788 -22652 12852
rect -22588 12788 -22568 12852
rect -22672 12772 -22568 12788
rect -22672 12708 -22652 12772
rect -22588 12708 -22568 12772
rect -22672 12692 -22568 12708
rect -22672 12628 -22652 12692
rect -22588 12628 -22568 12692
rect -22672 12612 -22568 12628
rect -22672 12548 -22652 12612
rect -22588 12548 -22568 12612
rect -22672 12532 -22568 12548
rect -22672 12468 -22652 12532
rect -22588 12468 -22568 12532
rect -22672 12452 -22568 12468
rect -22672 12388 -22652 12452
rect -22588 12388 -22568 12452
rect -22672 12372 -22568 12388
rect -22672 12308 -22652 12372
rect -22588 12308 -22568 12372
rect -22672 12292 -22568 12308
rect -22672 12228 -22652 12292
rect -22588 12228 -22568 12292
rect -22672 12212 -22568 12228
rect -22672 12148 -22652 12212
rect -22588 12148 -22568 12212
rect -22672 12132 -22568 12148
rect -22672 12068 -22652 12132
rect -22588 12068 -22568 12132
rect -22672 12052 -22568 12068
rect -22672 11988 -22652 12052
rect -22588 11988 -22568 12052
rect -22672 11972 -22568 11988
rect -22672 11908 -22652 11972
rect -22588 11908 -22568 11972
rect -22672 11892 -22568 11908
rect -22672 11828 -22652 11892
rect -22588 11828 -22568 11892
rect -22672 11812 -22568 11828
rect -22672 11748 -22652 11812
rect -22588 11748 -22568 11812
rect -22672 11732 -22568 11748
rect -22672 11668 -22652 11732
rect -22588 11668 -22568 11732
rect -22672 11652 -22568 11668
rect -22672 11588 -22652 11652
rect -22588 11588 -22568 11652
rect -22672 11572 -22568 11588
rect -22672 11508 -22652 11572
rect -22588 11508 -22568 11572
rect -22672 11492 -22568 11508
rect -22672 11428 -22652 11492
rect -22588 11428 -22568 11492
rect -22672 11412 -22568 11428
rect -22672 11348 -22652 11412
rect -22588 11348 -22568 11412
rect -22672 11332 -22568 11348
rect -22672 11268 -22652 11332
rect -22588 11268 -22568 11332
rect -22672 11252 -22568 11268
rect -22672 11188 -22652 11252
rect -22588 11188 -22568 11252
rect -22672 11172 -22568 11188
rect -22672 11108 -22652 11172
rect -22588 11108 -22568 11172
rect -22672 11092 -22568 11108
rect -22672 11028 -22652 11092
rect -22588 11028 -22568 11092
rect -22672 11012 -22568 11028
rect -22672 10948 -22652 11012
rect -22588 10948 -22568 11012
rect -22672 10932 -22568 10948
rect -22672 10868 -22652 10932
rect -22588 10868 -22568 10932
rect -22672 10852 -22568 10868
rect -28284 10492 -28180 10788
rect -33896 10412 -33792 10428
rect -33896 10348 -33876 10412
rect -33812 10348 -33792 10412
rect -33896 10332 -33792 10348
rect -33896 10268 -33876 10332
rect -33812 10268 -33792 10332
rect -33896 10252 -33792 10268
rect -33896 10188 -33876 10252
rect -33812 10188 -33792 10252
rect -33896 10172 -33792 10188
rect -33896 10108 -33876 10172
rect -33812 10108 -33792 10172
rect -33896 10092 -33792 10108
rect -33896 10028 -33876 10092
rect -33812 10028 -33792 10092
rect -33896 10012 -33792 10028
rect -33896 9948 -33876 10012
rect -33812 9948 -33792 10012
rect -33896 9932 -33792 9948
rect -33896 9868 -33876 9932
rect -33812 9868 -33792 9932
rect -33896 9852 -33792 9868
rect -33896 9788 -33876 9852
rect -33812 9788 -33792 9852
rect -33896 9772 -33792 9788
rect -33896 9708 -33876 9772
rect -33812 9708 -33792 9772
rect -33896 9692 -33792 9708
rect -33896 9628 -33876 9692
rect -33812 9628 -33792 9692
rect -33896 9612 -33792 9628
rect -33896 9548 -33876 9612
rect -33812 9548 -33792 9612
rect -33896 9532 -33792 9548
rect -33896 9468 -33876 9532
rect -33812 9468 -33792 9532
rect -33896 9452 -33792 9468
rect -33896 9388 -33876 9452
rect -33812 9388 -33792 9452
rect -33896 9372 -33792 9388
rect -33896 9308 -33876 9372
rect -33812 9308 -33792 9372
rect -33896 9292 -33792 9308
rect -33896 9228 -33876 9292
rect -33812 9228 -33792 9292
rect -33896 9212 -33792 9228
rect -33896 9148 -33876 9212
rect -33812 9148 -33792 9212
rect -33896 9132 -33792 9148
rect -33896 9068 -33876 9132
rect -33812 9068 -33792 9132
rect -33896 9052 -33792 9068
rect -33896 8988 -33876 9052
rect -33812 8988 -33792 9052
rect -33896 8972 -33792 8988
rect -33896 8908 -33876 8972
rect -33812 8908 -33792 8972
rect -33896 8892 -33792 8908
rect -33896 8828 -33876 8892
rect -33812 8828 -33792 8892
rect -33896 8812 -33792 8828
rect -33896 8748 -33876 8812
rect -33812 8748 -33792 8812
rect -33896 8732 -33792 8748
rect -33896 8668 -33876 8732
rect -33812 8668 -33792 8732
rect -33896 8652 -33792 8668
rect -33896 8588 -33876 8652
rect -33812 8588 -33792 8652
rect -33896 8572 -33792 8588
rect -33896 8508 -33876 8572
rect -33812 8508 -33792 8572
rect -33896 8492 -33792 8508
rect -33896 8428 -33876 8492
rect -33812 8428 -33792 8492
rect -33896 8412 -33792 8428
rect -33896 8348 -33876 8412
rect -33812 8348 -33792 8412
rect -33896 8332 -33792 8348
rect -33896 8268 -33876 8332
rect -33812 8268 -33792 8332
rect -33896 8252 -33792 8268
rect -33896 8188 -33876 8252
rect -33812 8188 -33792 8252
rect -33896 8172 -33792 8188
rect -33896 8108 -33876 8172
rect -33812 8108 -33792 8172
rect -33896 8092 -33792 8108
rect -33896 8028 -33876 8092
rect -33812 8028 -33792 8092
rect -33896 8012 -33792 8028
rect -33896 7948 -33876 8012
rect -33812 7948 -33792 8012
rect -33896 7932 -33792 7948
rect -33896 7868 -33876 7932
rect -33812 7868 -33792 7932
rect -33896 7852 -33792 7868
rect -33896 7788 -33876 7852
rect -33812 7788 -33792 7852
rect -33896 7772 -33792 7788
rect -33896 7708 -33876 7772
rect -33812 7708 -33792 7772
rect -33896 7692 -33792 7708
rect -33896 7628 -33876 7692
rect -33812 7628 -33792 7692
rect -33896 7612 -33792 7628
rect -33896 7548 -33876 7612
rect -33812 7548 -33792 7612
rect -33896 7532 -33792 7548
rect -33896 7468 -33876 7532
rect -33812 7468 -33792 7532
rect -33896 7452 -33792 7468
rect -33896 7388 -33876 7452
rect -33812 7388 -33792 7452
rect -33896 7372 -33792 7388
rect -33896 7308 -33876 7372
rect -33812 7308 -33792 7372
rect -33896 7292 -33792 7308
rect -33896 7228 -33876 7292
rect -33812 7228 -33792 7292
rect -33896 7212 -33792 7228
rect -33896 7148 -33876 7212
rect -33812 7148 -33792 7212
rect -33896 7132 -33792 7148
rect -33896 7068 -33876 7132
rect -33812 7068 -33792 7132
rect -33896 7052 -33792 7068
rect -33896 6988 -33876 7052
rect -33812 6988 -33792 7052
rect -33896 6972 -33792 6988
rect -33896 6908 -33876 6972
rect -33812 6908 -33792 6972
rect -33896 6892 -33792 6908
rect -33896 6828 -33876 6892
rect -33812 6828 -33792 6892
rect -33896 6812 -33792 6828
rect -33896 6748 -33876 6812
rect -33812 6748 -33792 6812
rect -33896 6732 -33792 6748
rect -33896 6668 -33876 6732
rect -33812 6668 -33792 6732
rect -33896 6652 -33792 6668
rect -33896 6588 -33876 6652
rect -33812 6588 -33792 6652
rect -33896 6572 -33792 6588
rect -33896 6508 -33876 6572
rect -33812 6508 -33792 6572
rect -33896 6492 -33792 6508
rect -33896 6428 -33876 6492
rect -33812 6428 -33792 6492
rect -33896 6412 -33792 6428
rect -33896 6348 -33876 6412
rect -33812 6348 -33792 6412
rect -33896 6332 -33792 6348
rect -33896 6268 -33876 6332
rect -33812 6268 -33792 6332
rect -33896 6252 -33792 6268
rect -33896 6188 -33876 6252
rect -33812 6188 -33792 6252
rect -33896 6172 -33792 6188
rect -33896 6108 -33876 6172
rect -33812 6108 -33792 6172
rect -33896 6092 -33792 6108
rect -33896 6028 -33876 6092
rect -33812 6028 -33792 6092
rect -33896 6012 -33792 6028
rect -33896 5948 -33876 6012
rect -33812 5948 -33792 6012
rect -33896 5932 -33792 5948
rect -33896 5868 -33876 5932
rect -33812 5868 -33792 5932
rect -33896 5852 -33792 5868
rect -33896 5788 -33876 5852
rect -33812 5788 -33792 5852
rect -33896 5772 -33792 5788
rect -33896 5708 -33876 5772
rect -33812 5708 -33792 5772
rect -33896 5692 -33792 5708
rect -33896 5628 -33876 5692
rect -33812 5628 -33792 5692
rect -33896 5612 -33792 5628
rect -33896 5548 -33876 5612
rect -33812 5548 -33792 5612
rect -33896 5532 -33792 5548
rect -36676 5121 -36572 5519
rect -33896 5468 -33876 5532
rect -33812 5468 -33792 5532
rect -33473 10412 -28551 10441
rect -33473 5548 -33444 10412
rect -28580 5548 -28551 10412
rect -33473 5519 -28551 5548
rect -28284 10428 -28264 10492
rect -28200 10428 -28180 10492
rect -25452 10441 -25348 10839
rect -22672 10788 -22652 10852
rect -22588 10788 -22568 10852
rect -22249 15732 -17327 15761
rect -22249 10868 -22220 15732
rect -17356 10868 -17327 15732
rect -22249 10839 -17327 10868
rect -17060 15748 -17040 15812
rect -16976 15748 -16956 15812
rect -14228 15761 -14124 16159
rect -11448 16108 -11428 16172
rect -11364 16108 -11344 16172
rect -11025 21052 -6103 21081
rect -11025 16188 -10996 21052
rect -6132 16188 -6103 21052
rect -11025 16159 -6103 16188
rect -5836 21068 -5816 21132
rect -5752 21068 -5732 21132
rect -3004 21081 -2900 21479
rect -224 21428 -204 21492
rect -140 21428 -120 21492
rect 199 26372 5121 26401
rect 199 21508 228 26372
rect 5092 21508 5121 26372
rect 199 21479 5121 21508
rect 5388 26388 5408 26452
rect 5472 26388 5492 26452
rect 8220 26401 8324 26799
rect 11000 26748 11020 26812
rect 11084 26748 11104 26812
rect 11423 31692 16345 31721
rect 11423 26828 11452 31692
rect 16316 26828 16345 31692
rect 11423 26799 16345 26828
rect 16612 31708 16632 31772
rect 16696 31708 16716 31772
rect 19444 31721 19548 32119
rect 22224 32068 22244 32132
rect 22308 32068 22328 32132
rect 22647 37012 27569 37041
rect 22647 32148 22676 37012
rect 27540 32148 27569 37012
rect 22647 32119 27569 32148
rect 27836 37028 27856 37092
rect 27920 37028 27940 37092
rect 30668 37041 30772 37240
rect 33448 37092 33552 37240
rect 27836 37012 27940 37028
rect 27836 36948 27856 37012
rect 27920 36948 27940 37012
rect 27836 36932 27940 36948
rect 27836 36868 27856 36932
rect 27920 36868 27940 36932
rect 27836 36852 27940 36868
rect 27836 36788 27856 36852
rect 27920 36788 27940 36852
rect 27836 36772 27940 36788
rect 27836 36708 27856 36772
rect 27920 36708 27940 36772
rect 27836 36692 27940 36708
rect 27836 36628 27856 36692
rect 27920 36628 27940 36692
rect 27836 36612 27940 36628
rect 27836 36548 27856 36612
rect 27920 36548 27940 36612
rect 27836 36532 27940 36548
rect 27836 36468 27856 36532
rect 27920 36468 27940 36532
rect 27836 36452 27940 36468
rect 27836 36388 27856 36452
rect 27920 36388 27940 36452
rect 27836 36372 27940 36388
rect 27836 36308 27856 36372
rect 27920 36308 27940 36372
rect 27836 36292 27940 36308
rect 27836 36228 27856 36292
rect 27920 36228 27940 36292
rect 27836 36212 27940 36228
rect 27836 36148 27856 36212
rect 27920 36148 27940 36212
rect 27836 36132 27940 36148
rect 27836 36068 27856 36132
rect 27920 36068 27940 36132
rect 27836 36052 27940 36068
rect 27836 35988 27856 36052
rect 27920 35988 27940 36052
rect 27836 35972 27940 35988
rect 27836 35908 27856 35972
rect 27920 35908 27940 35972
rect 27836 35892 27940 35908
rect 27836 35828 27856 35892
rect 27920 35828 27940 35892
rect 27836 35812 27940 35828
rect 27836 35748 27856 35812
rect 27920 35748 27940 35812
rect 27836 35732 27940 35748
rect 27836 35668 27856 35732
rect 27920 35668 27940 35732
rect 27836 35652 27940 35668
rect 27836 35588 27856 35652
rect 27920 35588 27940 35652
rect 27836 35572 27940 35588
rect 27836 35508 27856 35572
rect 27920 35508 27940 35572
rect 27836 35492 27940 35508
rect 27836 35428 27856 35492
rect 27920 35428 27940 35492
rect 27836 35412 27940 35428
rect 27836 35348 27856 35412
rect 27920 35348 27940 35412
rect 27836 35332 27940 35348
rect 27836 35268 27856 35332
rect 27920 35268 27940 35332
rect 27836 35252 27940 35268
rect 27836 35188 27856 35252
rect 27920 35188 27940 35252
rect 27836 35172 27940 35188
rect 27836 35108 27856 35172
rect 27920 35108 27940 35172
rect 27836 35092 27940 35108
rect 27836 35028 27856 35092
rect 27920 35028 27940 35092
rect 27836 35012 27940 35028
rect 27836 34948 27856 35012
rect 27920 34948 27940 35012
rect 27836 34932 27940 34948
rect 27836 34868 27856 34932
rect 27920 34868 27940 34932
rect 27836 34852 27940 34868
rect 27836 34788 27856 34852
rect 27920 34788 27940 34852
rect 27836 34772 27940 34788
rect 27836 34708 27856 34772
rect 27920 34708 27940 34772
rect 27836 34692 27940 34708
rect 27836 34628 27856 34692
rect 27920 34628 27940 34692
rect 27836 34612 27940 34628
rect 27836 34548 27856 34612
rect 27920 34548 27940 34612
rect 27836 34532 27940 34548
rect 27836 34468 27856 34532
rect 27920 34468 27940 34532
rect 27836 34452 27940 34468
rect 27836 34388 27856 34452
rect 27920 34388 27940 34452
rect 27836 34372 27940 34388
rect 27836 34308 27856 34372
rect 27920 34308 27940 34372
rect 27836 34292 27940 34308
rect 27836 34228 27856 34292
rect 27920 34228 27940 34292
rect 27836 34212 27940 34228
rect 27836 34148 27856 34212
rect 27920 34148 27940 34212
rect 27836 34132 27940 34148
rect 27836 34068 27856 34132
rect 27920 34068 27940 34132
rect 27836 34052 27940 34068
rect 27836 33988 27856 34052
rect 27920 33988 27940 34052
rect 27836 33972 27940 33988
rect 27836 33908 27856 33972
rect 27920 33908 27940 33972
rect 27836 33892 27940 33908
rect 27836 33828 27856 33892
rect 27920 33828 27940 33892
rect 27836 33812 27940 33828
rect 27836 33748 27856 33812
rect 27920 33748 27940 33812
rect 27836 33732 27940 33748
rect 27836 33668 27856 33732
rect 27920 33668 27940 33732
rect 27836 33652 27940 33668
rect 27836 33588 27856 33652
rect 27920 33588 27940 33652
rect 27836 33572 27940 33588
rect 27836 33508 27856 33572
rect 27920 33508 27940 33572
rect 27836 33492 27940 33508
rect 27836 33428 27856 33492
rect 27920 33428 27940 33492
rect 27836 33412 27940 33428
rect 27836 33348 27856 33412
rect 27920 33348 27940 33412
rect 27836 33332 27940 33348
rect 27836 33268 27856 33332
rect 27920 33268 27940 33332
rect 27836 33252 27940 33268
rect 27836 33188 27856 33252
rect 27920 33188 27940 33252
rect 27836 33172 27940 33188
rect 27836 33108 27856 33172
rect 27920 33108 27940 33172
rect 27836 33092 27940 33108
rect 27836 33028 27856 33092
rect 27920 33028 27940 33092
rect 27836 33012 27940 33028
rect 27836 32948 27856 33012
rect 27920 32948 27940 33012
rect 27836 32932 27940 32948
rect 27836 32868 27856 32932
rect 27920 32868 27940 32932
rect 27836 32852 27940 32868
rect 27836 32788 27856 32852
rect 27920 32788 27940 32852
rect 27836 32772 27940 32788
rect 27836 32708 27856 32772
rect 27920 32708 27940 32772
rect 27836 32692 27940 32708
rect 27836 32628 27856 32692
rect 27920 32628 27940 32692
rect 27836 32612 27940 32628
rect 27836 32548 27856 32612
rect 27920 32548 27940 32612
rect 27836 32532 27940 32548
rect 27836 32468 27856 32532
rect 27920 32468 27940 32532
rect 27836 32452 27940 32468
rect 27836 32388 27856 32452
rect 27920 32388 27940 32452
rect 27836 32372 27940 32388
rect 27836 32308 27856 32372
rect 27920 32308 27940 32372
rect 27836 32292 27940 32308
rect 27836 32228 27856 32292
rect 27920 32228 27940 32292
rect 27836 32212 27940 32228
rect 27836 32148 27856 32212
rect 27920 32148 27940 32212
rect 27836 32132 27940 32148
rect 22224 31772 22328 32068
rect 16612 31692 16716 31708
rect 16612 31628 16632 31692
rect 16696 31628 16716 31692
rect 16612 31612 16716 31628
rect 16612 31548 16632 31612
rect 16696 31548 16716 31612
rect 16612 31532 16716 31548
rect 16612 31468 16632 31532
rect 16696 31468 16716 31532
rect 16612 31452 16716 31468
rect 16612 31388 16632 31452
rect 16696 31388 16716 31452
rect 16612 31372 16716 31388
rect 16612 31308 16632 31372
rect 16696 31308 16716 31372
rect 16612 31292 16716 31308
rect 16612 31228 16632 31292
rect 16696 31228 16716 31292
rect 16612 31212 16716 31228
rect 16612 31148 16632 31212
rect 16696 31148 16716 31212
rect 16612 31132 16716 31148
rect 16612 31068 16632 31132
rect 16696 31068 16716 31132
rect 16612 31052 16716 31068
rect 16612 30988 16632 31052
rect 16696 30988 16716 31052
rect 16612 30972 16716 30988
rect 16612 30908 16632 30972
rect 16696 30908 16716 30972
rect 16612 30892 16716 30908
rect 16612 30828 16632 30892
rect 16696 30828 16716 30892
rect 16612 30812 16716 30828
rect 16612 30748 16632 30812
rect 16696 30748 16716 30812
rect 16612 30732 16716 30748
rect 16612 30668 16632 30732
rect 16696 30668 16716 30732
rect 16612 30652 16716 30668
rect 16612 30588 16632 30652
rect 16696 30588 16716 30652
rect 16612 30572 16716 30588
rect 16612 30508 16632 30572
rect 16696 30508 16716 30572
rect 16612 30492 16716 30508
rect 16612 30428 16632 30492
rect 16696 30428 16716 30492
rect 16612 30412 16716 30428
rect 16612 30348 16632 30412
rect 16696 30348 16716 30412
rect 16612 30332 16716 30348
rect 16612 30268 16632 30332
rect 16696 30268 16716 30332
rect 16612 30252 16716 30268
rect 16612 30188 16632 30252
rect 16696 30188 16716 30252
rect 16612 30172 16716 30188
rect 16612 30108 16632 30172
rect 16696 30108 16716 30172
rect 16612 30092 16716 30108
rect 16612 30028 16632 30092
rect 16696 30028 16716 30092
rect 16612 30012 16716 30028
rect 16612 29948 16632 30012
rect 16696 29948 16716 30012
rect 16612 29932 16716 29948
rect 16612 29868 16632 29932
rect 16696 29868 16716 29932
rect 16612 29852 16716 29868
rect 16612 29788 16632 29852
rect 16696 29788 16716 29852
rect 16612 29772 16716 29788
rect 16612 29708 16632 29772
rect 16696 29708 16716 29772
rect 16612 29692 16716 29708
rect 16612 29628 16632 29692
rect 16696 29628 16716 29692
rect 16612 29612 16716 29628
rect 16612 29548 16632 29612
rect 16696 29548 16716 29612
rect 16612 29532 16716 29548
rect 16612 29468 16632 29532
rect 16696 29468 16716 29532
rect 16612 29452 16716 29468
rect 16612 29388 16632 29452
rect 16696 29388 16716 29452
rect 16612 29372 16716 29388
rect 16612 29308 16632 29372
rect 16696 29308 16716 29372
rect 16612 29292 16716 29308
rect 16612 29228 16632 29292
rect 16696 29228 16716 29292
rect 16612 29212 16716 29228
rect 16612 29148 16632 29212
rect 16696 29148 16716 29212
rect 16612 29132 16716 29148
rect 16612 29068 16632 29132
rect 16696 29068 16716 29132
rect 16612 29052 16716 29068
rect 16612 28988 16632 29052
rect 16696 28988 16716 29052
rect 16612 28972 16716 28988
rect 16612 28908 16632 28972
rect 16696 28908 16716 28972
rect 16612 28892 16716 28908
rect 16612 28828 16632 28892
rect 16696 28828 16716 28892
rect 16612 28812 16716 28828
rect 16612 28748 16632 28812
rect 16696 28748 16716 28812
rect 16612 28732 16716 28748
rect 16612 28668 16632 28732
rect 16696 28668 16716 28732
rect 16612 28652 16716 28668
rect 16612 28588 16632 28652
rect 16696 28588 16716 28652
rect 16612 28572 16716 28588
rect 16612 28508 16632 28572
rect 16696 28508 16716 28572
rect 16612 28492 16716 28508
rect 16612 28428 16632 28492
rect 16696 28428 16716 28492
rect 16612 28412 16716 28428
rect 16612 28348 16632 28412
rect 16696 28348 16716 28412
rect 16612 28332 16716 28348
rect 16612 28268 16632 28332
rect 16696 28268 16716 28332
rect 16612 28252 16716 28268
rect 16612 28188 16632 28252
rect 16696 28188 16716 28252
rect 16612 28172 16716 28188
rect 16612 28108 16632 28172
rect 16696 28108 16716 28172
rect 16612 28092 16716 28108
rect 16612 28028 16632 28092
rect 16696 28028 16716 28092
rect 16612 28012 16716 28028
rect 16612 27948 16632 28012
rect 16696 27948 16716 28012
rect 16612 27932 16716 27948
rect 16612 27868 16632 27932
rect 16696 27868 16716 27932
rect 16612 27852 16716 27868
rect 16612 27788 16632 27852
rect 16696 27788 16716 27852
rect 16612 27772 16716 27788
rect 16612 27708 16632 27772
rect 16696 27708 16716 27772
rect 16612 27692 16716 27708
rect 16612 27628 16632 27692
rect 16696 27628 16716 27692
rect 16612 27612 16716 27628
rect 16612 27548 16632 27612
rect 16696 27548 16716 27612
rect 16612 27532 16716 27548
rect 16612 27468 16632 27532
rect 16696 27468 16716 27532
rect 16612 27452 16716 27468
rect 16612 27388 16632 27452
rect 16696 27388 16716 27452
rect 16612 27372 16716 27388
rect 16612 27308 16632 27372
rect 16696 27308 16716 27372
rect 16612 27292 16716 27308
rect 16612 27228 16632 27292
rect 16696 27228 16716 27292
rect 16612 27212 16716 27228
rect 16612 27148 16632 27212
rect 16696 27148 16716 27212
rect 16612 27132 16716 27148
rect 16612 27068 16632 27132
rect 16696 27068 16716 27132
rect 16612 27052 16716 27068
rect 16612 26988 16632 27052
rect 16696 26988 16716 27052
rect 16612 26972 16716 26988
rect 16612 26908 16632 26972
rect 16696 26908 16716 26972
rect 16612 26892 16716 26908
rect 16612 26828 16632 26892
rect 16696 26828 16716 26892
rect 16612 26812 16716 26828
rect 11000 26452 11104 26748
rect 5388 26372 5492 26388
rect 5388 26308 5408 26372
rect 5472 26308 5492 26372
rect 5388 26292 5492 26308
rect 5388 26228 5408 26292
rect 5472 26228 5492 26292
rect 5388 26212 5492 26228
rect 5388 26148 5408 26212
rect 5472 26148 5492 26212
rect 5388 26132 5492 26148
rect 5388 26068 5408 26132
rect 5472 26068 5492 26132
rect 5388 26052 5492 26068
rect 5388 25988 5408 26052
rect 5472 25988 5492 26052
rect 5388 25972 5492 25988
rect 5388 25908 5408 25972
rect 5472 25908 5492 25972
rect 5388 25892 5492 25908
rect 5388 25828 5408 25892
rect 5472 25828 5492 25892
rect 5388 25812 5492 25828
rect 5388 25748 5408 25812
rect 5472 25748 5492 25812
rect 5388 25732 5492 25748
rect 5388 25668 5408 25732
rect 5472 25668 5492 25732
rect 5388 25652 5492 25668
rect 5388 25588 5408 25652
rect 5472 25588 5492 25652
rect 5388 25572 5492 25588
rect 5388 25508 5408 25572
rect 5472 25508 5492 25572
rect 5388 25492 5492 25508
rect 5388 25428 5408 25492
rect 5472 25428 5492 25492
rect 5388 25412 5492 25428
rect 5388 25348 5408 25412
rect 5472 25348 5492 25412
rect 5388 25332 5492 25348
rect 5388 25268 5408 25332
rect 5472 25268 5492 25332
rect 5388 25252 5492 25268
rect 5388 25188 5408 25252
rect 5472 25188 5492 25252
rect 5388 25172 5492 25188
rect 5388 25108 5408 25172
rect 5472 25108 5492 25172
rect 5388 25092 5492 25108
rect 5388 25028 5408 25092
rect 5472 25028 5492 25092
rect 5388 25012 5492 25028
rect 5388 24948 5408 25012
rect 5472 24948 5492 25012
rect 5388 24932 5492 24948
rect 5388 24868 5408 24932
rect 5472 24868 5492 24932
rect 5388 24852 5492 24868
rect 5388 24788 5408 24852
rect 5472 24788 5492 24852
rect 5388 24772 5492 24788
rect 5388 24708 5408 24772
rect 5472 24708 5492 24772
rect 5388 24692 5492 24708
rect 5388 24628 5408 24692
rect 5472 24628 5492 24692
rect 5388 24612 5492 24628
rect 5388 24548 5408 24612
rect 5472 24548 5492 24612
rect 5388 24532 5492 24548
rect 5388 24468 5408 24532
rect 5472 24468 5492 24532
rect 5388 24452 5492 24468
rect 5388 24388 5408 24452
rect 5472 24388 5492 24452
rect 5388 24372 5492 24388
rect 5388 24308 5408 24372
rect 5472 24308 5492 24372
rect 5388 24292 5492 24308
rect 5388 24228 5408 24292
rect 5472 24228 5492 24292
rect 5388 24212 5492 24228
rect 5388 24148 5408 24212
rect 5472 24148 5492 24212
rect 5388 24132 5492 24148
rect 5388 24068 5408 24132
rect 5472 24068 5492 24132
rect 5388 24052 5492 24068
rect 5388 23988 5408 24052
rect 5472 23988 5492 24052
rect 5388 23972 5492 23988
rect 5388 23908 5408 23972
rect 5472 23908 5492 23972
rect 5388 23892 5492 23908
rect 5388 23828 5408 23892
rect 5472 23828 5492 23892
rect 5388 23812 5492 23828
rect 5388 23748 5408 23812
rect 5472 23748 5492 23812
rect 5388 23732 5492 23748
rect 5388 23668 5408 23732
rect 5472 23668 5492 23732
rect 5388 23652 5492 23668
rect 5388 23588 5408 23652
rect 5472 23588 5492 23652
rect 5388 23572 5492 23588
rect 5388 23508 5408 23572
rect 5472 23508 5492 23572
rect 5388 23492 5492 23508
rect 5388 23428 5408 23492
rect 5472 23428 5492 23492
rect 5388 23412 5492 23428
rect 5388 23348 5408 23412
rect 5472 23348 5492 23412
rect 5388 23332 5492 23348
rect 5388 23268 5408 23332
rect 5472 23268 5492 23332
rect 5388 23252 5492 23268
rect 5388 23188 5408 23252
rect 5472 23188 5492 23252
rect 5388 23172 5492 23188
rect 5388 23108 5408 23172
rect 5472 23108 5492 23172
rect 5388 23092 5492 23108
rect 5388 23028 5408 23092
rect 5472 23028 5492 23092
rect 5388 23012 5492 23028
rect 5388 22948 5408 23012
rect 5472 22948 5492 23012
rect 5388 22932 5492 22948
rect 5388 22868 5408 22932
rect 5472 22868 5492 22932
rect 5388 22852 5492 22868
rect 5388 22788 5408 22852
rect 5472 22788 5492 22852
rect 5388 22772 5492 22788
rect 5388 22708 5408 22772
rect 5472 22708 5492 22772
rect 5388 22692 5492 22708
rect 5388 22628 5408 22692
rect 5472 22628 5492 22692
rect 5388 22612 5492 22628
rect 5388 22548 5408 22612
rect 5472 22548 5492 22612
rect 5388 22532 5492 22548
rect 5388 22468 5408 22532
rect 5472 22468 5492 22532
rect 5388 22452 5492 22468
rect 5388 22388 5408 22452
rect 5472 22388 5492 22452
rect 5388 22372 5492 22388
rect 5388 22308 5408 22372
rect 5472 22308 5492 22372
rect 5388 22292 5492 22308
rect 5388 22228 5408 22292
rect 5472 22228 5492 22292
rect 5388 22212 5492 22228
rect 5388 22148 5408 22212
rect 5472 22148 5492 22212
rect 5388 22132 5492 22148
rect 5388 22068 5408 22132
rect 5472 22068 5492 22132
rect 5388 22052 5492 22068
rect 5388 21988 5408 22052
rect 5472 21988 5492 22052
rect 5388 21972 5492 21988
rect 5388 21908 5408 21972
rect 5472 21908 5492 21972
rect 5388 21892 5492 21908
rect 5388 21828 5408 21892
rect 5472 21828 5492 21892
rect 5388 21812 5492 21828
rect 5388 21748 5408 21812
rect 5472 21748 5492 21812
rect 5388 21732 5492 21748
rect 5388 21668 5408 21732
rect 5472 21668 5492 21732
rect 5388 21652 5492 21668
rect 5388 21588 5408 21652
rect 5472 21588 5492 21652
rect 5388 21572 5492 21588
rect 5388 21508 5408 21572
rect 5472 21508 5492 21572
rect 5388 21492 5492 21508
rect -224 21132 -120 21428
rect -5836 21052 -5732 21068
rect -5836 20988 -5816 21052
rect -5752 20988 -5732 21052
rect -5836 20972 -5732 20988
rect -5836 20908 -5816 20972
rect -5752 20908 -5732 20972
rect -5836 20892 -5732 20908
rect -5836 20828 -5816 20892
rect -5752 20828 -5732 20892
rect -5836 20812 -5732 20828
rect -5836 20748 -5816 20812
rect -5752 20748 -5732 20812
rect -5836 20732 -5732 20748
rect -5836 20668 -5816 20732
rect -5752 20668 -5732 20732
rect -5836 20652 -5732 20668
rect -5836 20588 -5816 20652
rect -5752 20588 -5732 20652
rect -5836 20572 -5732 20588
rect -5836 20508 -5816 20572
rect -5752 20508 -5732 20572
rect -5836 20492 -5732 20508
rect -5836 20428 -5816 20492
rect -5752 20428 -5732 20492
rect -5836 20412 -5732 20428
rect -5836 20348 -5816 20412
rect -5752 20348 -5732 20412
rect -5836 20332 -5732 20348
rect -5836 20268 -5816 20332
rect -5752 20268 -5732 20332
rect -5836 20252 -5732 20268
rect -5836 20188 -5816 20252
rect -5752 20188 -5732 20252
rect -5836 20172 -5732 20188
rect -5836 20108 -5816 20172
rect -5752 20108 -5732 20172
rect -5836 20092 -5732 20108
rect -5836 20028 -5816 20092
rect -5752 20028 -5732 20092
rect -5836 20012 -5732 20028
rect -5836 19948 -5816 20012
rect -5752 19948 -5732 20012
rect -5836 19932 -5732 19948
rect -5836 19868 -5816 19932
rect -5752 19868 -5732 19932
rect -5836 19852 -5732 19868
rect -5836 19788 -5816 19852
rect -5752 19788 -5732 19852
rect -5836 19772 -5732 19788
rect -5836 19708 -5816 19772
rect -5752 19708 -5732 19772
rect -5836 19692 -5732 19708
rect -5836 19628 -5816 19692
rect -5752 19628 -5732 19692
rect -5836 19612 -5732 19628
rect -5836 19548 -5816 19612
rect -5752 19548 -5732 19612
rect -5836 19532 -5732 19548
rect -5836 19468 -5816 19532
rect -5752 19468 -5732 19532
rect -5836 19452 -5732 19468
rect -5836 19388 -5816 19452
rect -5752 19388 -5732 19452
rect -5836 19372 -5732 19388
rect -5836 19308 -5816 19372
rect -5752 19308 -5732 19372
rect -5836 19292 -5732 19308
rect -5836 19228 -5816 19292
rect -5752 19228 -5732 19292
rect -5836 19212 -5732 19228
rect -5836 19148 -5816 19212
rect -5752 19148 -5732 19212
rect -5836 19132 -5732 19148
rect -5836 19068 -5816 19132
rect -5752 19068 -5732 19132
rect -5836 19052 -5732 19068
rect -5836 18988 -5816 19052
rect -5752 18988 -5732 19052
rect -5836 18972 -5732 18988
rect -5836 18908 -5816 18972
rect -5752 18908 -5732 18972
rect -5836 18892 -5732 18908
rect -5836 18828 -5816 18892
rect -5752 18828 -5732 18892
rect -5836 18812 -5732 18828
rect -5836 18748 -5816 18812
rect -5752 18748 -5732 18812
rect -5836 18732 -5732 18748
rect -5836 18668 -5816 18732
rect -5752 18668 -5732 18732
rect -5836 18652 -5732 18668
rect -5836 18588 -5816 18652
rect -5752 18588 -5732 18652
rect -5836 18572 -5732 18588
rect -5836 18508 -5816 18572
rect -5752 18508 -5732 18572
rect -5836 18492 -5732 18508
rect -5836 18428 -5816 18492
rect -5752 18428 -5732 18492
rect -5836 18412 -5732 18428
rect -5836 18348 -5816 18412
rect -5752 18348 -5732 18412
rect -5836 18332 -5732 18348
rect -5836 18268 -5816 18332
rect -5752 18268 -5732 18332
rect -5836 18252 -5732 18268
rect -5836 18188 -5816 18252
rect -5752 18188 -5732 18252
rect -5836 18172 -5732 18188
rect -5836 18108 -5816 18172
rect -5752 18108 -5732 18172
rect -5836 18092 -5732 18108
rect -5836 18028 -5816 18092
rect -5752 18028 -5732 18092
rect -5836 18012 -5732 18028
rect -5836 17948 -5816 18012
rect -5752 17948 -5732 18012
rect -5836 17932 -5732 17948
rect -5836 17868 -5816 17932
rect -5752 17868 -5732 17932
rect -5836 17852 -5732 17868
rect -5836 17788 -5816 17852
rect -5752 17788 -5732 17852
rect -5836 17772 -5732 17788
rect -5836 17708 -5816 17772
rect -5752 17708 -5732 17772
rect -5836 17692 -5732 17708
rect -5836 17628 -5816 17692
rect -5752 17628 -5732 17692
rect -5836 17612 -5732 17628
rect -5836 17548 -5816 17612
rect -5752 17548 -5732 17612
rect -5836 17532 -5732 17548
rect -5836 17468 -5816 17532
rect -5752 17468 -5732 17532
rect -5836 17452 -5732 17468
rect -5836 17388 -5816 17452
rect -5752 17388 -5732 17452
rect -5836 17372 -5732 17388
rect -5836 17308 -5816 17372
rect -5752 17308 -5732 17372
rect -5836 17292 -5732 17308
rect -5836 17228 -5816 17292
rect -5752 17228 -5732 17292
rect -5836 17212 -5732 17228
rect -5836 17148 -5816 17212
rect -5752 17148 -5732 17212
rect -5836 17132 -5732 17148
rect -5836 17068 -5816 17132
rect -5752 17068 -5732 17132
rect -5836 17052 -5732 17068
rect -5836 16988 -5816 17052
rect -5752 16988 -5732 17052
rect -5836 16972 -5732 16988
rect -5836 16908 -5816 16972
rect -5752 16908 -5732 16972
rect -5836 16892 -5732 16908
rect -5836 16828 -5816 16892
rect -5752 16828 -5732 16892
rect -5836 16812 -5732 16828
rect -5836 16748 -5816 16812
rect -5752 16748 -5732 16812
rect -5836 16732 -5732 16748
rect -5836 16668 -5816 16732
rect -5752 16668 -5732 16732
rect -5836 16652 -5732 16668
rect -5836 16588 -5816 16652
rect -5752 16588 -5732 16652
rect -5836 16572 -5732 16588
rect -5836 16508 -5816 16572
rect -5752 16508 -5732 16572
rect -5836 16492 -5732 16508
rect -5836 16428 -5816 16492
rect -5752 16428 -5732 16492
rect -5836 16412 -5732 16428
rect -5836 16348 -5816 16412
rect -5752 16348 -5732 16412
rect -5836 16332 -5732 16348
rect -5836 16268 -5816 16332
rect -5752 16268 -5732 16332
rect -5836 16252 -5732 16268
rect -5836 16188 -5816 16252
rect -5752 16188 -5732 16252
rect -5836 16172 -5732 16188
rect -11448 15812 -11344 16108
rect -17060 15732 -16956 15748
rect -17060 15668 -17040 15732
rect -16976 15668 -16956 15732
rect -17060 15652 -16956 15668
rect -17060 15588 -17040 15652
rect -16976 15588 -16956 15652
rect -17060 15572 -16956 15588
rect -17060 15508 -17040 15572
rect -16976 15508 -16956 15572
rect -17060 15492 -16956 15508
rect -17060 15428 -17040 15492
rect -16976 15428 -16956 15492
rect -17060 15412 -16956 15428
rect -17060 15348 -17040 15412
rect -16976 15348 -16956 15412
rect -17060 15332 -16956 15348
rect -17060 15268 -17040 15332
rect -16976 15268 -16956 15332
rect -17060 15252 -16956 15268
rect -17060 15188 -17040 15252
rect -16976 15188 -16956 15252
rect -17060 15172 -16956 15188
rect -17060 15108 -17040 15172
rect -16976 15108 -16956 15172
rect -17060 15092 -16956 15108
rect -17060 15028 -17040 15092
rect -16976 15028 -16956 15092
rect -17060 15012 -16956 15028
rect -17060 14948 -17040 15012
rect -16976 14948 -16956 15012
rect -17060 14932 -16956 14948
rect -17060 14868 -17040 14932
rect -16976 14868 -16956 14932
rect -17060 14852 -16956 14868
rect -17060 14788 -17040 14852
rect -16976 14788 -16956 14852
rect -17060 14772 -16956 14788
rect -17060 14708 -17040 14772
rect -16976 14708 -16956 14772
rect -17060 14692 -16956 14708
rect -17060 14628 -17040 14692
rect -16976 14628 -16956 14692
rect -17060 14612 -16956 14628
rect -17060 14548 -17040 14612
rect -16976 14548 -16956 14612
rect -17060 14532 -16956 14548
rect -17060 14468 -17040 14532
rect -16976 14468 -16956 14532
rect -17060 14452 -16956 14468
rect -17060 14388 -17040 14452
rect -16976 14388 -16956 14452
rect -17060 14372 -16956 14388
rect -17060 14308 -17040 14372
rect -16976 14308 -16956 14372
rect -17060 14292 -16956 14308
rect -17060 14228 -17040 14292
rect -16976 14228 -16956 14292
rect -17060 14212 -16956 14228
rect -17060 14148 -17040 14212
rect -16976 14148 -16956 14212
rect -17060 14132 -16956 14148
rect -17060 14068 -17040 14132
rect -16976 14068 -16956 14132
rect -17060 14052 -16956 14068
rect -17060 13988 -17040 14052
rect -16976 13988 -16956 14052
rect -17060 13972 -16956 13988
rect -17060 13908 -17040 13972
rect -16976 13908 -16956 13972
rect -17060 13892 -16956 13908
rect -17060 13828 -17040 13892
rect -16976 13828 -16956 13892
rect -17060 13812 -16956 13828
rect -17060 13748 -17040 13812
rect -16976 13748 -16956 13812
rect -17060 13732 -16956 13748
rect -17060 13668 -17040 13732
rect -16976 13668 -16956 13732
rect -17060 13652 -16956 13668
rect -17060 13588 -17040 13652
rect -16976 13588 -16956 13652
rect -17060 13572 -16956 13588
rect -17060 13508 -17040 13572
rect -16976 13508 -16956 13572
rect -17060 13492 -16956 13508
rect -17060 13428 -17040 13492
rect -16976 13428 -16956 13492
rect -17060 13412 -16956 13428
rect -17060 13348 -17040 13412
rect -16976 13348 -16956 13412
rect -17060 13332 -16956 13348
rect -17060 13268 -17040 13332
rect -16976 13268 -16956 13332
rect -17060 13252 -16956 13268
rect -17060 13188 -17040 13252
rect -16976 13188 -16956 13252
rect -17060 13172 -16956 13188
rect -17060 13108 -17040 13172
rect -16976 13108 -16956 13172
rect -17060 13092 -16956 13108
rect -17060 13028 -17040 13092
rect -16976 13028 -16956 13092
rect -17060 13012 -16956 13028
rect -17060 12948 -17040 13012
rect -16976 12948 -16956 13012
rect -17060 12932 -16956 12948
rect -17060 12868 -17040 12932
rect -16976 12868 -16956 12932
rect -17060 12852 -16956 12868
rect -17060 12788 -17040 12852
rect -16976 12788 -16956 12852
rect -17060 12772 -16956 12788
rect -17060 12708 -17040 12772
rect -16976 12708 -16956 12772
rect -17060 12692 -16956 12708
rect -17060 12628 -17040 12692
rect -16976 12628 -16956 12692
rect -17060 12612 -16956 12628
rect -17060 12548 -17040 12612
rect -16976 12548 -16956 12612
rect -17060 12532 -16956 12548
rect -17060 12468 -17040 12532
rect -16976 12468 -16956 12532
rect -17060 12452 -16956 12468
rect -17060 12388 -17040 12452
rect -16976 12388 -16956 12452
rect -17060 12372 -16956 12388
rect -17060 12308 -17040 12372
rect -16976 12308 -16956 12372
rect -17060 12292 -16956 12308
rect -17060 12228 -17040 12292
rect -16976 12228 -16956 12292
rect -17060 12212 -16956 12228
rect -17060 12148 -17040 12212
rect -16976 12148 -16956 12212
rect -17060 12132 -16956 12148
rect -17060 12068 -17040 12132
rect -16976 12068 -16956 12132
rect -17060 12052 -16956 12068
rect -17060 11988 -17040 12052
rect -16976 11988 -16956 12052
rect -17060 11972 -16956 11988
rect -17060 11908 -17040 11972
rect -16976 11908 -16956 11972
rect -17060 11892 -16956 11908
rect -17060 11828 -17040 11892
rect -16976 11828 -16956 11892
rect -17060 11812 -16956 11828
rect -17060 11748 -17040 11812
rect -16976 11748 -16956 11812
rect -17060 11732 -16956 11748
rect -17060 11668 -17040 11732
rect -16976 11668 -16956 11732
rect -17060 11652 -16956 11668
rect -17060 11588 -17040 11652
rect -16976 11588 -16956 11652
rect -17060 11572 -16956 11588
rect -17060 11508 -17040 11572
rect -16976 11508 -16956 11572
rect -17060 11492 -16956 11508
rect -17060 11428 -17040 11492
rect -16976 11428 -16956 11492
rect -17060 11412 -16956 11428
rect -17060 11348 -17040 11412
rect -16976 11348 -16956 11412
rect -17060 11332 -16956 11348
rect -17060 11268 -17040 11332
rect -16976 11268 -16956 11332
rect -17060 11252 -16956 11268
rect -17060 11188 -17040 11252
rect -16976 11188 -16956 11252
rect -17060 11172 -16956 11188
rect -17060 11108 -17040 11172
rect -16976 11108 -16956 11172
rect -17060 11092 -16956 11108
rect -17060 11028 -17040 11092
rect -16976 11028 -16956 11092
rect -17060 11012 -16956 11028
rect -17060 10948 -17040 11012
rect -16976 10948 -16956 11012
rect -17060 10932 -16956 10948
rect -17060 10868 -17040 10932
rect -16976 10868 -16956 10932
rect -17060 10852 -16956 10868
rect -22672 10492 -22568 10788
rect -28284 10412 -28180 10428
rect -28284 10348 -28264 10412
rect -28200 10348 -28180 10412
rect -28284 10332 -28180 10348
rect -28284 10268 -28264 10332
rect -28200 10268 -28180 10332
rect -28284 10252 -28180 10268
rect -28284 10188 -28264 10252
rect -28200 10188 -28180 10252
rect -28284 10172 -28180 10188
rect -28284 10108 -28264 10172
rect -28200 10108 -28180 10172
rect -28284 10092 -28180 10108
rect -28284 10028 -28264 10092
rect -28200 10028 -28180 10092
rect -28284 10012 -28180 10028
rect -28284 9948 -28264 10012
rect -28200 9948 -28180 10012
rect -28284 9932 -28180 9948
rect -28284 9868 -28264 9932
rect -28200 9868 -28180 9932
rect -28284 9852 -28180 9868
rect -28284 9788 -28264 9852
rect -28200 9788 -28180 9852
rect -28284 9772 -28180 9788
rect -28284 9708 -28264 9772
rect -28200 9708 -28180 9772
rect -28284 9692 -28180 9708
rect -28284 9628 -28264 9692
rect -28200 9628 -28180 9692
rect -28284 9612 -28180 9628
rect -28284 9548 -28264 9612
rect -28200 9548 -28180 9612
rect -28284 9532 -28180 9548
rect -28284 9468 -28264 9532
rect -28200 9468 -28180 9532
rect -28284 9452 -28180 9468
rect -28284 9388 -28264 9452
rect -28200 9388 -28180 9452
rect -28284 9372 -28180 9388
rect -28284 9308 -28264 9372
rect -28200 9308 -28180 9372
rect -28284 9292 -28180 9308
rect -28284 9228 -28264 9292
rect -28200 9228 -28180 9292
rect -28284 9212 -28180 9228
rect -28284 9148 -28264 9212
rect -28200 9148 -28180 9212
rect -28284 9132 -28180 9148
rect -28284 9068 -28264 9132
rect -28200 9068 -28180 9132
rect -28284 9052 -28180 9068
rect -28284 8988 -28264 9052
rect -28200 8988 -28180 9052
rect -28284 8972 -28180 8988
rect -28284 8908 -28264 8972
rect -28200 8908 -28180 8972
rect -28284 8892 -28180 8908
rect -28284 8828 -28264 8892
rect -28200 8828 -28180 8892
rect -28284 8812 -28180 8828
rect -28284 8748 -28264 8812
rect -28200 8748 -28180 8812
rect -28284 8732 -28180 8748
rect -28284 8668 -28264 8732
rect -28200 8668 -28180 8732
rect -28284 8652 -28180 8668
rect -28284 8588 -28264 8652
rect -28200 8588 -28180 8652
rect -28284 8572 -28180 8588
rect -28284 8508 -28264 8572
rect -28200 8508 -28180 8572
rect -28284 8492 -28180 8508
rect -28284 8428 -28264 8492
rect -28200 8428 -28180 8492
rect -28284 8412 -28180 8428
rect -28284 8348 -28264 8412
rect -28200 8348 -28180 8412
rect -28284 8332 -28180 8348
rect -28284 8268 -28264 8332
rect -28200 8268 -28180 8332
rect -28284 8252 -28180 8268
rect -28284 8188 -28264 8252
rect -28200 8188 -28180 8252
rect -28284 8172 -28180 8188
rect -28284 8108 -28264 8172
rect -28200 8108 -28180 8172
rect -28284 8092 -28180 8108
rect -28284 8028 -28264 8092
rect -28200 8028 -28180 8092
rect -28284 8012 -28180 8028
rect -28284 7948 -28264 8012
rect -28200 7948 -28180 8012
rect -28284 7932 -28180 7948
rect -28284 7868 -28264 7932
rect -28200 7868 -28180 7932
rect -28284 7852 -28180 7868
rect -28284 7788 -28264 7852
rect -28200 7788 -28180 7852
rect -28284 7772 -28180 7788
rect -28284 7708 -28264 7772
rect -28200 7708 -28180 7772
rect -28284 7692 -28180 7708
rect -28284 7628 -28264 7692
rect -28200 7628 -28180 7692
rect -28284 7612 -28180 7628
rect -28284 7548 -28264 7612
rect -28200 7548 -28180 7612
rect -28284 7532 -28180 7548
rect -28284 7468 -28264 7532
rect -28200 7468 -28180 7532
rect -28284 7452 -28180 7468
rect -28284 7388 -28264 7452
rect -28200 7388 -28180 7452
rect -28284 7372 -28180 7388
rect -28284 7308 -28264 7372
rect -28200 7308 -28180 7372
rect -28284 7292 -28180 7308
rect -28284 7228 -28264 7292
rect -28200 7228 -28180 7292
rect -28284 7212 -28180 7228
rect -28284 7148 -28264 7212
rect -28200 7148 -28180 7212
rect -28284 7132 -28180 7148
rect -28284 7068 -28264 7132
rect -28200 7068 -28180 7132
rect -28284 7052 -28180 7068
rect -28284 6988 -28264 7052
rect -28200 6988 -28180 7052
rect -28284 6972 -28180 6988
rect -28284 6908 -28264 6972
rect -28200 6908 -28180 6972
rect -28284 6892 -28180 6908
rect -28284 6828 -28264 6892
rect -28200 6828 -28180 6892
rect -28284 6812 -28180 6828
rect -28284 6748 -28264 6812
rect -28200 6748 -28180 6812
rect -28284 6732 -28180 6748
rect -28284 6668 -28264 6732
rect -28200 6668 -28180 6732
rect -28284 6652 -28180 6668
rect -28284 6588 -28264 6652
rect -28200 6588 -28180 6652
rect -28284 6572 -28180 6588
rect -28284 6508 -28264 6572
rect -28200 6508 -28180 6572
rect -28284 6492 -28180 6508
rect -28284 6428 -28264 6492
rect -28200 6428 -28180 6492
rect -28284 6412 -28180 6428
rect -28284 6348 -28264 6412
rect -28200 6348 -28180 6412
rect -28284 6332 -28180 6348
rect -28284 6268 -28264 6332
rect -28200 6268 -28180 6332
rect -28284 6252 -28180 6268
rect -28284 6188 -28264 6252
rect -28200 6188 -28180 6252
rect -28284 6172 -28180 6188
rect -28284 6108 -28264 6172
rect -28200 6108 -28180 6172
rect -28284 6092 -28180 6108
rect -28284 6028 -28264 6092
rect -28200 6028 -28180 6092
rect -28284 6012 -28180 6028
rect -28284 5948 -28264 6012
rect -28200 5948 -28180 6012
rect -28284 5932 -28180 5948
rect -28284 5868 -28264 5932
rect -28200 5868 -28180 5932
rect -28284 5852 -28180 5868
rect -28284 5788 -28264 5852
rect -28200 5788 -28180 5852
rect -28284 5772 -28180 5788
rect -28284 5708 -28264 5772
rect -28200 5708 -28180 5772
rect -28284 5692 -28180 5708
rect -28284 5628 -28264 5692
rect -28200 5628 -28180 5692
rect -28284 5612 -28180 5628
rect -28284 5548 -28264 5612
rect -28200 5548 -28180 5612
rect -28284 5532 -28180 5548
rect -33896 5172 -33792 5468
rect -39085 5092 -34163 5121
rect -39085 228 -39056 5092
rect -34192 228 -34163 5092
rect -39085 199 -34163 228
rect -33896 5108 -33876 5172
rect -33812 5108 -33792 5172
rect -31064 5121 -30960 5519
rect -28284 5468 -28264 5532
rect -28200 5468 -28180 5532
rect -27861 10412 -22939 10441
rect -27861 5548 -27832 10412
rect -22968 5548 -22939 10412
rect -27861 5519 -22939 5548
rect -22672 10428 -22652 10492
rect -22588 10428 -22568 10492
rect -19840 10441 -19736 10839
rect -17060 10788 -17040 10852
rect -16976 10788 -16956 10852
rect -16637 15732 -11715 15761
rect -16637 10868 -16608 15732
rect -11744 10868 -11715 15732
rect -16637 10839 -11715 10868
rect -11448 15748 -11428 15812
rect -11364 15748 -11344 15812
rect -8616 15761 -8512 16159
rect -5836 16108 -5816 16172
rect -5752 16108 -5732 16172
rect -5413 21052 -491 21081
rect -5413 16188 -5384 21052
rect -520 16188 -491 21052
rect -5413 16159 -491 16188
rect -224 21068 -204 21132
rect -140 21068 -120 21132
rect 2608 21081 2712 21479
rect 5388 21428 5408 21492
rect 5472 21428 5492 21492
rect 5811 26372 10733 26401
rect 5811 21508 5840 26372
rect 10704 21508 10733 26372
rect 5811 21479 10733 21508
rect 11000 26388 11020 26452
rect 11084 26388 11104 26452
rect 13832 26401 13936 26799
rect 16612 26748 16632 26812
rect 16696 26748 16716 26812
rect 17035 31692 21957 31721
rect 17035 26828 17064 31692
rect 21928 26828 21957 31692
rect 17035 26799 21957 26828
rect 22224 31708 22244 31772
rect 22308 31708 22328 31772
rect 25056 31721 25160 32119
rect 27836 32068 27856 32132
rect 27920 32068 27940 32132
rect 28259 37012 33181 37041
rect 28259 32148 28288 37012
rect 33152 32148 33181 37012
rect 28259 32119 33181 32148
rect 33448 37028 33468 37092
rect 33532 37028 33552 37092
rect 36280 37041 36384 37240
rect 39060 37092 39164 37240
rect 33448 37012 33552 37028
rect 33448 36948 33468 37012
rect 33532 36948 33552 37012
rect 33448 36932 33552 36948
rect 33448 36868 33468 36932
rect 33532 36868 33552 36932
rect 33448 36852 33552 36868
rect 33448 36788 33468 36852
rect 33532 36788 33552 36852
rect 33448 36772 33552 36788
rect 33448 36708 33468 36772
rect 33532 36708 33552 36772
rect 33448 36692 33552 36708
rect 33448 36628 33468 36692
rect 33532 36628 33552 36692
rect 33448 36612 33552 36628
rect 33448 36548 33468 36612
rect 33532 36548 33552 36612
rect 33448 36532 33552 36548
rect 33448 36468 33468 36532
rect 33532 36468 33552 36532
rect 33448 36452 33552 36468
rect 33448 36388 33468 36452
rect 33532 36388 33552 36452
rect 33448 36372 33552 36388
rect 33448 36308 33468 36372
rect 33532 36308 33552 36372
rect 33448 36292 33552 36308
rect 33448 36228 33468 36292
rect 33532 36228 33552 36292
rect 33448 36212 33552 36228
rect 33448 36148 33468 36212
rect 33532 36148 33552 36212
rect 33448 36132 33552 36148
rect 33448 36068 33468 36132
rect 33532 36068 33552 36132
rect 33448 36052 33552 36068
rect 33448 35988 33468 36052
rect 33532 35988 33552 36052
rect 33448 35972 33552 35988
rect 33448 35908 33468 35972
rect 33532 35908 33552 35972
rect 33448 35892 33552 35908
rect 33448 35828 33468 35892
rect 33532 35828 33552 35892
rect 33448 35812 33552 35828
rect 33448 35748 33468 35812
rect 33532 35748 33552 35812
rect 33448 35732 33552 35748
rect 33448 35668 33468 35732
rect 33532 35668 33552 35732
rect 33448 35652 33552 35668
rect 33448 35588 33468 35652
rect 33532 35588 33552 35652
rect 33448 35572 33552 35588
rect 33448 35508 33468 35572
rect 33532 35508 33552 35572
rect 33448 35492 33552 35508
rect 33448 35428 33468 35492
rect 33532 35428 33552 35492
rect 33448 35412 33552 35428
rect 33448 35348 33468 35412
rect 33532 35348 33552 35412
rect 33448 35332 33552 35348
rect 33448 35268 33468 35332
rect 33532 35268 33552 35332
rect 33448 35252 33552 35268
rect 33448 35188 33468 35252
rect 33532 35188 33552 35252
rect 33448 35172 33552 35188
rect 33448 35108 33468 35172
rect 33532 35108 33552 35172
rect 33448 35092 33552 35108
rect 33448 35028 33468 35092
rect 33532 35028 33552 35092
rect 33448 35012 33552 35028
rect 33448 34948 33468 35012
rect 33532 34948 33552 35012
rect 33448 34932 33552 34948
rect 33448 34868 33468 34932
rect 33532 34868 33552 34932
rect 33448 34852 33552 34868
rect 33448 34788 33468 34852
rect 33532 34788 33552 34852
rect 33448 34772 33552 34788
rect 33448 34708 33468 34772
rect 33532 34708 33552 34772
rect 33448 34692 33552 34708
rect 33448 34628 33468 34692
rect 33532 34628 33552 34692
rect 33448 34612 33552 34628
rect 33448 34548 33468 34612
rect 33532 34548 33552 34612
rect 33448 34532 33552 34548
rect 33448 34468 33468 34532
rect 33532 34468 33552 34532
rect 33448 34452 33552 34468
rect 33448 34388 33468 34452
rect 33532 34388 33552 34452
rect 33448 34372 33552 34388
rect 33448 34308 33468 34372
rect 33532 34308 33552 34372
rect 33448 34292 33552 34308
rect 33448 34228 33468 34292
rect 33532 34228 33552 34292
rect 33448 34212 33552 34228
rect 33448 34148 33468 34212
rect 33532 34148 33552 34212
rect 33448 34132 33552 34148
rect 33448 34068 33468 34132
rect 33532 34068 33552 34132
rect 33448 34052 33552 34068
rect 33448 33988 33468 34052
rect 33532 33988 33552 34052
rect 33448 33972 33552 33988
rect 33448 33908 33468 33972
rect 33532 33908 33552 33972
rect 33448 33892 33552 33908
rect 33448 33828 33468 33892
rect 33532 33828 33552 33892
rect 33448 33812 33552 33828
rect 33448 33748 33468 33812
rect 33532 33748 33552 33812
rect 33448 33732 33552 33748
rect 33448 33668 33468 33732
rect 33532 33668 33552 33732
rect 33448 33652 33552 33668
rect 33448 33588 33468 33652
rect 33532 33588 33552 33652
rect 33448 33572 33552 33588
rect 33448 33508 33468 33572
rect 33532 33508 33552 33572
rect 33448 33492 33552 33508
rect 33448 33428 33468 33492
rect 33532 33428 33552 33492
rect 33448 33412 33552 33428
rect 33448 33348 33468 33412
rect 33532 33348 33552 33412
rect 33448 33332 33552 33348
rect 33448 33268 33468 33332
rect 33532 33268 33552 33332
rect 33448 33252 33552 33268
rect 33448 33188 33468 33252
rect 33532 33188 33552 33252
rect 33448 33172 33552 33188
rect 33448 33108 33468 33172
rect 33532 33108 33552 33172
rect 33448 33092 33552 33108
rect 33448 33028 33468 33092
rect 33532 33028 33552 33092
rect 33448 33012 33552 33028
rect 33448 32948 33468 33012
rect 33532 32948 33552 33012
rect 33448 32932 33552 32948
rect 33448 32868 33468 32932
rect 33532 32868 33552 32932
rect 33448 32852 33552 32868
rect 33448 32788 33468 32852
rect 33532 32788 33552 32852
rect 33448 32772 33552 32788
rect 33448 32708 33468 32772
rect 33532 32708 33552 32772
rect 33448 32692 33552 32708
rect 33448 32628 33468 32692
rect 33532 32628 33552 32692
rect 33448 32612 33552 32628
rect 33448 32548 33468 32612
rect 33532 32548 33552 32612
rect 33448 32532 33552 32548
rect 33448 32468 33468 32532
rect 33532 32468 33552 32532
rect 33448 32452 33552 32468
rect 33448 32388 33468 32452
rect 33532 32388 33552 32452
rect 33448 32372 33552 32388
rect 33448 32308 33468 32372
rect 33532 32308 33552 32372
rect 33448 32292 33552 32308
rect 33448 32228 33468 32292
rect 33532 32228 33552 32292
rect 33448 32212 33552 32228
rect 33448 32148 33468 32212
rect 33532 32148 33552 32212
rect 33448 32132 33552 32148
rect 27836 31772 27940 32068
rect 22224 31692 22328 31708
rect 22224 31628 22244 31692
rect 22308 31628 22328 31692
rect 22224 31612 22328 31628
rect 22224 31548 22244 31612
rect 22308 31548 22328 31612
rect 22224 31532 22328 31548
rect 22224 31468 22244 31532
rect 22308 31468 22328 31532
rect 22224 31452 22328 31468
rect 22224 31388 22244 31452
rect 22308 31388 22328 31452
rect 22224 31372 22328 31388
rect 22224 31308 22244 31372
rect 22308 31308 22328 31372
rect 22224 31292 22328 31308
rect 22224 31228 22244 31292
rect 22308 31228 22328 31292
rect 22224 31212 22328 31228
rect 22224 31148 22244 31212
rect 22308 31148 22328 31212
rect 22224 31132 22328 31148
rect 22224 31068 22244 31132
rect 22308 31068 22328 31132
rect 22224 31052 22328 31068
rect 22224 30988 22244 31052
rect 22308 30988 22328 31052
rect 22224 30972 22328 30988
rect 22224 30908 22244 30972
rect 22308 30908 22328 30972
rect 22224 30892 22328 30908
rect 22224 30828 22244 30892
rect 22308 30828 22328 30892
rect 22224 30812 22328 30828
rect 22224 30748 22244 30812
rect 22308 30748 22328 30812
rect 22224 30732 22328 30748
rect 22224 30668 22244 30732
rect 22308 30668 22328 30732
rect 22224 30652 22328 30668
rect 22224 30588 22244 30652
rect 22308 30588 22328 30652
rect 22224 30572 22328 30588
rect 22224 30508 22244 30572
rect 22308 30508 22328 30572
rect 22224 30492 22328 30508
rect 22224 30428 22244 30492
rect 22308 30428 22328 30492
rect 22224 30412 22328 30428
rect 22224 30348 22244 30412
rect 22308 30348 22328 30412
rect 22224 30332 22328 30348
rect 22224 30268 22244 30332
rect 22308 30268 22328 30332
rect 22224 30252 22328 30268
rect 22224 30188 22244 30252
rect 22308 30188 22328 30252
rect 22224 30172 22328 30188
rect 22224 30108 22244 30172
rect 22308 30108 22328 30172
rect 22224 30092 22328 30108
rect 22224 30028 22244 30092
rect 22308 30028 22328 30092
rect 22224 30012 22328 30028
rect 22224 29948 22244 30012
rect 22308 29948 22328 30012
rect 22224 29932 22328 29948
rect 22224 29868 22244 29932
rect 22308 29868 22328 29932
rect 22224 29852 22328 29868
rect 22224 29788 22244 29852
rect 22308 29788 22328 29852
rect 22224 29772 22328 29788
rect 22224 29708 22244 29772
rect 22308 29708 22328 29772
rect 22224 29692 22328 29708
rect 22224 29628 22244 29692
rect 22308 29628 22328 29692
rect 22224 29612 22328 29628
rect 22224 29548 22244 29612
rect 22308 29548 22328 29612
rect 22224 29532 22328 29548
rect 22224 29468 22244 29532
rect 22308 29468 22328 29532
rect 22224 29452 22328 29468
rect 22224 29388 22244 29452
rect 22308 29388 22328 29452
rect 22224 29372 22328 29388
rect 22224 29308 22244 29372
rect 22308 29308 22328 29372
rect 22224 29292 22328 29308
rect 22224 29228 22244 29292
rect 22308 29228 22328 29292
rect 22224 29212 22328 29228
rect 22224 29148 22244 29212
rect 22308 29148 22328 29212
rect 22224 29132 22328 29148
rect 22224 29068 22244 29132
rect 22308 29068 22328 29132
rect 22224 29052 22328 29068
rect 22224 28988 22244 29052
rect 22308 28988 22328 29052
rect 22224 28972 22328 28988
rect 22224 28908 22244 28972
rect 22308 28908 22328 28972
rect 22224 28892 22328 28908
rect 22224 28828 22244 28892
rect 22308 28828 22328 28892
rect 22224 28812 22328 28828
rect 22224 28748 22244 28812
rect 22308 28748 22328 28812
rect 22224 28732 22328 28748
rect 22224 28668 22244 28732
rect 22308 28668 22328 28732
rect 22224 28652 22328 28668
rect 22224 28588 22244 28652
rect 22308 28588 22328 28652
rect 22224 28572 22328 28588
rect 22224 28508 22244 28572
rect 22308 28508 22328 28572
rect 22224 28492 22328 28508
rect 22224 28428 22244 28492
rect 22308 28428 22328 28492
rect 22224 28412 22328 28428
rect 22224 28348 22244 28412
rect 22308 28348 22328 28412
rect 22224 28332 22328 28348
rect 22224 28268 22244 28332
rect 22308 28268 22328 28332
rect 22224 28252 22328 28268
rect 22224 28188 22244 28252
rect 22308 28188 22328 28252
rect 22224 28172 22328 28188
rect 22224 28108 22244 28172
rect 22308 28108 22328 28172
rect 22224 28092 22328 28108
rect 22224 28028 22244 28092
rect 22308 28028 22328 28092
rect 22224 28012 22328 28028
rect 22224 27948 22244 28012
rect 22308 27948 22328 28012
rect 22224 27932 22328 27948
rect 22224 27868 22244 27932
rect 22308 27868 22328 27932
rect 22224 27852 22328 27868
rect 22224 27788 22244 27852
rect 22308 27788 22328 27852
rect 22224 27772 22328 27788
rect 22224 27708 22244 27772
rect 22308 27708 22328 27772
rect 22224 27692 22328 27708
rect 22224 27628 22244 27692
rect 22308 27628 22328 27692
rect 22224 27612 22328 27628
rect 22224 27548 22244 27612
rect 22308 27548 22328 27612
rect 22224 27532 22328 27548
rect 22224 27468 22244 27532
rect 22308 27468 22328 27532
rect 22224 27452 22328 27468
rect 22224 27388 22244 27452
rect 22308 27388 22328 27452
rect 22224 27372 22328 27388
rect 22224 27308 22244 27372
rect 22308 27308 22328 27372
rect 22224 27292 22328 27308
rect 22224 27228 22244 27292
rect 22308 27228 22328 27292
rect 22224 27212 22328 27228
rect 22224 27148 22244 27212
rect 22308 27148 22328 27212
rect 22224 27132 22328 27148
rect 22224 27068 22244 27132
rect 22308 27068 22328 27132
rect 22224 27052 22328 27068
rect 22224 26988 22244 27052
rect 22308 26988 22328 27052
rect 22224 26972 22328 26988
rect 22224 26908 22244 26972
rect 22308 26908 22328 26972
rect 22224 26892 22328 26908
rect 22224 26828 22244 26892
rect 22308 26828 22328 26892
rect 22224 26812 22328 26828
rect 16612 26452 16716 26748
rect 11000 26372 11104 26388
rect 11000 26308 11020 26372
rect 11084 26308 11104 26372
rect 11000 26292 11104 26308
rect 11000 26228 11020 26292
rect 11084 26228 11104 26292
rect 11000 26212 11104 26228
rect 11000 26148 11020 26212
rect 11084 26148 11104 26212
rect 11000 26132 11104 26148
rect 11000 26068 11020 26132
rect 11084 26068 11104 26132
rect 11000 26052 11104 26068
rect 11000 25988 11020 26052
rect 11084 25988 11104 26052
rect 11000 25972 11104 25988
rect 11000 25908 11020 25972
rect 11084 25908 11104 25972
rect 11000 25892 11104 25908
rect 11000 25828 11020 25892
rect 11084 25828 11104 25892
rect 11000 25812 11104 25828
rect 11000 25748 11020 25812
rect 11084 25748 11104 25812
rect 11000 25732 11104 25748
rect 11000 25668 11020 25732
rect 11084 25668 11104 25732
rect 11000 25652 11104 25668
rect 11000 25588 11020 25652
rect 11084 25588 11104 25652
rect 11000 25572 11104 25588
rect 11000 25508 11020 25572
rect 11084 25508 11104 25572
rect 11000 25492 11104 25508
rect 11000 25428 11020 25492
rect 11084 25428 11104 25492
rect 11000 25412 11104 25428
rect 11000 25348 11020 25412
rect 11084 25348 11104 25412
rect 11000 25332 11104 25348
rect 11000 25268 11020 25332
rect 11084 25268 11104 25332
rect 11000 25252 11104 25268
rect 11000 25188 11020 25252
rect 11084 25188 11104 25252
rect 11000 25172 11104 25188
rect 11000 25108 11020 25172
rect 11084 25108 11104 25172
rect 11000 25092 11104 25108
rect 11000 25028 11020 25092
rect 11084 25028 11104 25092
rect 11000 25012 11104 25028
rect 11000 24948 11020 25012
rect 11084 24948 11104 25012
rect 11000 24932 11104 24948
rect 11000 24868 11020 24932
rect 11084 24868 11104 24932
rect 11000 24852 11104 24868
rect 11000 24788 11020 24852
rect 11084 24788 11104 24852
rect 11000 24772 11104 24788
rect 11000 24708 11020 24772
rect 11084 24708 11104 24772
rect 11000 24692 11104 24708
rect 11000 24628 11020 24692
rect 11084 24628 11104 24692
rect 11000 24612 11104 24628
rect 11000 24548 11020 24612
rect 11084 24548 11104 24612
rect 11000 24532 11104 24548
rect 11000 24468 11020 24532
rect 11084 24468 11104 24532
rect 11000 24452 11104 24468
rect 11000 24388 11020 24452
rect 11084 24388 11104 24452
rect 11000 24372 11104 24388
rect 11000 24308 11020 24372
rect 11084 24308 11104 24372
rect 11000 24292 11104 24308
rect 11000 24228 11020 24292
rect 11084 24228 11104 24292
rect 11000 24212 11104 24228
rect 11000 24148 11020 24212
rect 11084 24148 11104 24212
rect 11000 24132 11104 24148
rect 11000 24068 11020 24132
rect 11084 24068 11104 24132
rect 11000 24052 11104 24068
rect 11000 23988 11020 24052
rect 11084 23988 11104 24052
rect 11000 23972 11104 23988
rect 11000 23908 11020 23972
rect 11084 23908 11104 23972
rect 11000 23892 11104 23908
rect 11000 23828 11020 23892
rect 11084 23828 11104 23892
rect 11000 23812 11104 23828
rect 11000 23748 11020 23812
rect 11084 23748 11104 23812
rect 11000 23732 11104 23748
rect 11000 23668 11020 23732
rect 11084 23668 11104 23732
rect 11000 23652 11104 23668
rect 11000 23588 11020 23652
rect 11084 23588 11104 23652
rect 11000 23572 11104 23588
rect 11000 23508 11020 23572
rect 11084 23508 11104 23572
rect 11000 23492 11104 23508
rect 11000 23428 11020 23492
rect 11084 23428 11104 23492
rect 11000 23412 11104 23428
rect 11000 23348 11020 23412
rect 11084 23348 11104 23412
rect 11000 23332 11104 23348
rect 11000 23268 11020 23332
rect 11084 23268 11104 23332
rect 11000 23252 11104 23268
rect 11000 23188 11020 23252
rect 11084 23188 11104 23252
rect 11000 23172 11104 23188
rect 11000 23108 11020 23172
rect 11084 23108 11104 23172
rect 11000 23092 11104 23108
rect 11000 23028 11020 23092
rect 11084 23028 11104 23092
rect 11000 23012 11104 23028
rect 11000 22948 11020 23012
rect 11084 22948 11104 23012
rect 11000 22932 11104 22948
rect 11000 22868 11020 22932
rect 11084 22868 11104 22932
rect 11000 22852 11104 22868
rect 11000 22788 11020 22852
rect 11084 22788 11104 22852
rect 11000 22772 11104 22788
rect 11000 22708 11020 22772
rect 11084 22708 11104 22772
rect 11000 22692 11104 22708
rect 11000 22628 11020 22692
rect 11084 22628 11104 22692
rect 11000 22612 11104 22628
rect 11000 22548 11020 22612
rect 11084 22548 11104 22612
rect 11000 22532 11104 22548
rect 11000 22468 11020 22532
rect 11084 22468 11104 22532
rect 11000 22452 11104 22468
rect 11000 22388 11020 22452
rect 11084 22388 11104 22452
rect 11000 22372 11104 22388
rect 11000 22308 11020 22372
rect 11084 22308 11104 22372
rect 11000 22292 11104 22308
rect 11000 22228 11020 22292
rect 11084 22228 11104 22292
rect 11000 22212 11104 22228
rect 11000 22148 11020 22212
rect 11084 22148 11104 22212
rect 11000 22132 11104 22148
rect 11000 22068 11020 22132
rect 11084 22068 11104 22132
rect 11000 22052 11104 22068
rect 11000 21988 11020 22052
rect 11084 21988 11104 22052
rect 11000 21972 11104 21988
rect 11000 21908 11020 21972
rect 11084 21908 11104 21972
rect 11000 21892 11104 21908
rect 11000 21828 11020 21892
rect 11084 21828 11104 21892
rect 11000 21812 11104 21828
rect 11000 21748 11020 21812
rect 11084 21748 11104 21812
rect 11000 21732 11104 21748
rect 11000 21668 11020 21732
rect 11084 21668 11104 21732
rect 11000 21652 11104 21668
rect 11000 21588 11020 21652
rect 11084 21588 11104 21652
rect 11000 21572 11104 21588
rect 11000 21508 11020 21572
rect 11084 21508 11104 21572
rect 11000 21492 11104 21508
rect 5388 21132 5492 21428
rect -224 21052 -120 21068
rect -224 20988 -204 21052
rect -140 20988 -120 21052
rect -224 20972 -120 20988
rect -224 20908 -204 20972
rect -140 20908 -120 20972
rect -224 20892 -120 20908
rect -224 20828 -204 20892
rect -140 20828 -120 20892
rect -224 20812 -120 20828
rect -224 20748 -204 20812
rect -140 20748 -120 20812
rect -224 20732 -120 20748
rect -224 20668 -204 20732
rect -140 20668 -120 20732
rect -224 20652 -120 20668
rect -224 20588 -204 20652
rect -140 20588 -120 20652
rect -224 20572 -120 20588
rect -224 20508 -204 20572
rect -140 20508 -120 20572
rect -224 20492 -120 20508
rect -224 20428 -204 20492
rect -140 20428 -120 20492
rect -224 20412 -120 20428
rect -224 20348 -204 20412
rect -140 20348 -120 20412
rect -224 20332 -120 20348
rect -224 20268 -204 20332
rect -140 20268 -120 20332
rect -224 20252 -120 20268
rect -224 20188 -204 20252
rect -140 20188 -120 20252
rect -224 20172 -120 20188
rect -224 20108 -204 20172
rect -140 20108 -120 20172
rect -224 20092 -120 20108
rect -224 20028 -204 20092
rect -140 20028 -120 20092
rect -224 20012 -120 20028
rect -224 19948 -204 20012
rect -140 19948 -120 20012
rect -224 19932 -120 19948
rect -224 19868 -204 19932
rect -140 19868 -120 19932
rect -224 19852 -120 19868
rect -224 19788 -204 19852
rect -140 19788 -120 19852
rect -224 19772 -120 19788
rect -224 19708 -204 19772
rect -140 19708 -120 19772
rect -224 19692 -120 19708
rect -224 19628 -204 19692
rect -140 19628 -120 19692
rect -224 19612 -120 19628
rect -224 19548 -204 19612
rect -140 19548 -120 19612
rect -224 19532 -120 19548
rect -224 19468 -204 19532
rect -140 19468 -120 19532
rect -224 19452 -120 19468
rect -224 19388 -204 19452
rect -140 19388 -120 19452
rect -224 19372 -120 19388
rect -224 19308 -204 19372
rect -140 19308 -120 19372
rect -224 19292 -120 19308
rect -224 19228 -204 19292
rect -140 19228 -120 19292
rect -224 19212 -120 19228
rect -224 19148 -204 19212
rect -140 19148 -120 19212
rect -224 19132 -120 19148
rect -224 19068 -204 19132
rect -140 19068 -120 19132
rect -224 19052 -120 19068
rect -224 18988 -204 19052
rect -140 18988 -120 19052
rect -224 18972 -120 18988
rect -224 18908 -204 18972
rect -140 18908 -120 18972
rect -224 18892 -120 18908
rect -224 18828 -204 18892
rect -140 18828 -120 18892
rect -224 18812 -120 18828
rect -224 18748 -204 18812
rect -140 18748 -120 18812
rect -224 18732 -120 18748
rect -224 18668 -204 18732
rect -140 18668 -120 18732
rect -224 18652 -120 18668
rect -224 18588 -204 18652
rect -140 18588 -120 18652
rect -224 18572 -120 18588
rect -224 18508 -204 18572
rect -140 18508 -120 18572
rect -224 18492 -120 18508
rect -224 18428 -204 18492
rect -140 18428 -120 18492
rect -224 18412 -120 18428
rect -224 18348 -204 18412
rect -140 18348 -120 18412
rect -224 18332 -120 18348
rect -224 18268 -204 18332
rect -140 18268 -120 18332
rect -224 18252 -120 18268
rect -224 18188 -204 18252
rect -140 18188 -120 18252
rect -224 18172 -120 18188
rect -224 18108 -204 18172
rect -140 18108 -120 18172
rect -224 18092 -120 18108
rect -224 18028 -204 18092
rect -140 18028 -120 18092
rect -224 18012 -120 18028
rect -224 17948 -204 18012
rect -140 17948 -120 18012
rect -224 17932 -120 17948
rect -224 17868 -204 17932
rect -140 17868 -120 17932
rect -224 17852 -120 17868
rect -224 17788 -204 17852
rect -140 17788 -120 17852
rect -224 17772 -120 17788
rect -224 17708 -204 17772
rect -140 17708 -120 17772
rect -224 17692 -120 17708
rect -224 17628 -204 17692
rect -140 17628 -120 17692
rect -224 17612 -120 17628
rect -224 17548 -204 17612
rect -140 17548 -120 17612
rect -224 17532 -120 17548
rect -224 17468 -204 17532
rect -140 17468 -120 17532
rect -224 17452 -120 17468
rect -224 17388 -204 17452
rect -140 17388 -120 17452
rect -224 17372 -120 17388
rect -224 17308 -204 17372
rect -140 17308 -120 17372
rect -224 17292 -120 17308
rect -224 17228 -204 17292
rect -140 17228 -120 17292
rect -224 17212 -120 17228
rect -224 17148 -204 17212
rect -140 17148 -120 17212
rect -224 17132 -120 17148
rect -224 17068 -204 17132
rect -140 17068 -120 17132
rect -224 17052 -120 17068
rect -224 16988 -204 17052
rect -140 16988 -120 17052
rect -224 16972 -120 16988
rect -224 16908 -204 16972
rect -140 16908 -120 16972
rect -224 16892 -120 16908
rect -224 16828 -204 16892
rect -140 16828 -120 16892
rect -224 16812 -120 16828
rect -224 16748 -204 16812
rect -140 16748 -120 16812
rect -224 16732 -120 16748
rect -224 16668 -204 16732
rect -140 16668 -120 16732
rect -224 16652 -120 16668
rect -224 16588 -204 16652
rect -140 16588 -120 16652
rect -224 16572 -120 16588
rect -224 16508 -204 16572
rect -140 16508 -120 16572
rect -224 16492 -120 16508
rect -224 16428 -204 16492
rect -140 16428 -120 16492
rect -224 16412 -120 16428
rect -224 16348 -204 16412
rect -140 16348 -120 16412
rect -224 16332 -120 16348
rect -224 16268 -204 16332
rect -140 16268 -120 16332
rect -224 16252 -120 16268
rect -224 16188 -204 16252
rect -140 16188 -120 16252
rect -224 16172 -120 16188
rect -5836 15812 -5732 16108
rect -11448 15732 -11344 15748
rect -11448 15668 -11428 15732
rect -11364 15668 -11344 15732
rect -11448 15652 -11344 15668
rect -11448 15588 -11428 15652
rect -11364 15588 -11344 15652
rect -11448 15572 -11344 15588
rect -11448 15508 -11428 15572
rect -11364 15508 -11344 15572
rect -11448 15492 -11344 15508
rect -11448 15428 -11428 15492
rect -11364 15428 -11344 15492
rect -11448 15412 -11344 15428
rect -11448 15348 -11428 15412
rect -11364 15348 -11344 15412
rect -11448 15332 -11344 15348
rect -11448 15268 -11428 15332
rect -11364 15268 -11344 15332
rect -11448 15252 -11344 15268
rect -11448 15188 -11428 15252
rect -11364 15188 -11344 15252
rect -11448 15172 -11344 15188
rect -11448 15108 -11428 15172
rect -11364 15108 -11344 15172
rect -11448 15092 -11344 15108
rect -11448 15028 -11428 15092
rect -11364 15028 -11344 15092
rect -11448 15012 -11344 15028
rect -11448 14948 -11428 15012
rect -11364 14948 -11344 15012
rect -11448 14932 -11344 14948
rect -11448 14868 -11428 14932
rect -11364 14868 -11344 14932
rect -11448 14852 -11344 14868
rect -11448 14788 -11428 14852
rect -11364 14788 -11344 14852
rect -11448 14772 -11344 14788
rect -11448 14708 -11428 14772
rect -11364 14708 -11344 14772
rect -11448 14692 -11344 14708
rect -11448 14628 -11428 14692
rect -11364 14628 -11344 14692
rect -11448 14612 -11344 14628
rect -11448 14548 -11428 14612
rect -11364 14548 -11344 14612
rect -11448 14532 -11344 14548
rect -11448 14468 -11428 14532
rect -11364 14468 -11344 14532
rect -11448 14452 -11344 14468
rect -11448 14388 -11428 14452
rect -11364 14388 -11344 14452
rect -11448 14372 -11344 14388
rect -11448 14308 -11428 14372
rect -11364 14308 -11344 14372
rect -11448 14292 -11344 14308
rect -11448 14228 -11428 14292
rect -11364 14228 -11344 14292
rect -11448 14212 -11344 14228
rect -11448 14148 -11428 14212
rect -11364 14148 -11344 14212
rect -11448 14132 -11344 14148
rect -11448 14068 -11428 14132
rect -11364 14068 -11344 14132
rect -11448 14052 -11344 14068
rect -11448 13988 -11428 14052
rect -11364 13988 -11344 14052
rect -11448 13972 -11344 13988
rect -11448 13908 -11428 13972
rect -11364 13908 -11344 13972
rect -11448 13892 -11344 13908
rect -11448 13828 -11428 13892
rect -11364 13828 -11344 13892
rect -11448 13812 -11344 13828
rect -11448 13748 -11428 13812
rect -11364 13748 -11344 13812
rect -11448 13732 -11344 13748
rect -11448 13668 -11428 13732
rect -11364 13668 -11344 13732
rect -11448 13652 -11344 13668
rect -11448 13588 -11428 13652
rect -11364 13588 -11344 13652
rect -11448 13572 -11344 13588
rect -11448 13508 -11428 13572
rect -11364 13508 -11344 13572
rect -11448 13492 -11344 13508
rect -11448 13428 -11428 13492
rect -11364 13428 -11344 13492
rect -11448 13412 -11344 13428
rect -11448 13348 -11428 13412
rect -11364 13348 -11344 13412
rect -11448 13332 -11344 13348
rect -11448 13268 -11428 13332
rect -11364 13268 -11344 13332
rect -11448 13252 -11344 13268
rect -11448 13188 -11428 13252
rect -11364 13188 -11344 13252
rect -11448 13172 -11344 13188
rect -11448 13108 -11428 13172
rect -11364 13108 -11344 13172
rect -11448 13092 -11344 13108
rect -11448 13028 -11428 13092
rect -11364 13028 -11344 13092
rect -11448 13012 -11344 13028
rect -11448 12948 -11428 13012
rect -11364 12948 -11344 13012
rect -11448 12932 -11344 12948
rect -11448 12868 -11428 12932
rect -11364 12868 -11344 12932
rect -11448 12852 -11344 12868
rect -11448 12788 -11428 12852
rect -11364 12788 -11344 12852
rect -11448 12772 -11344 12788
rect -11448 12708 -11428 12772
rect -11364 12708 -11344 12772
rect -11448 12692 -11344 12708
rect -11448 12628 -11428 12692
rect -11364 12628 -11344 12692
rect -11448 12612 -11344 12628
rect -11448 12548 -11428 12612
rect -11364 12548 -11344 12612
rect -11448 12532 -11344 12548
rect -11448 12468 -11428 12532
rect -11364 12468 -11344 12532
rect -11448 12452 -11344 12468
rect -11448 12388 -11428 12452
rect -11364 12388 -11344 12452
rect -11448 12372 -11344 12388
rect -11448 12308 -11428 12372
rect -11364 12308 -11344 12372
rect -11448 12292 -11344 12308
rect -11448 12228 -11428 12292
rect -11364 12228 -11344 12292
rect -11448 12212 -11344 12228
rect -11448 12148 -11428 12212
rect -11364 12148 -11344 12212
rect -11448 12132 -11344 12148
rect -11448 12068 -11428 12132
rect -11364 12068 -11344 12132
rect -11448 12052 -11344 12068
rect -11448 11988 -11428 12052
rect -11364 11988 -11344 12052
rect -11448 11972 -11344 11988
rect -11448 11908 -11428 11972
rect -11364 11908 -11344 11972
rect -11448 11892 -11344 11908
rect -11448 11828 -11428 11892
rect -11364 11828 -11344 11892
rect -11448 11812 -11344 11828
rect -11448 11748 -11428 11812
rect -11364 11748 -11344 11812
rect -11448 11732 -11344 11748
rect -11448 11668 -11428 11732
rect -11364 11668 -11344 11732
rect -11448 11652 -11344 11668
rect -11448 11588 -11428 11652
rect -11364 11588 -11344 11652
rect -11448 11572 -11344 11588
rect -11448 11508 -11428 11572
rect -11364 11508 -11344 11572
rect -11448 11492 -11344 11508
rect -11448 11428 -11428 11492
rect -11364 11428 -11344 11492
rect -11448 11412 -11344 11428
rect -11448 11348 -11428 11412
rect -11364 11348 -11344 11412
rect -11448 11332 -11344 11348
rect -11448 11268 -11428 11332
rect -11364 11268 -11344 11332
rect -11448 11252 -11344 11268
rect -11448 11188 -11428 11252
rect -11364 11188 -11344 11252
rect -11448 11172 -11344 11188
rect -11448 11108 -11428 11172
rect -11364 11108 -11344 11172
rect -11448 11092 -11344 11108
rect -11448 11028 -11428 11092
rect -11364 11028 -11344 11092
rect -11448 11012 -11344 11028
rect -11448 10948 -11428 11012
rect -11364 10948 -11344 11012
rect -11448 10932 -11344 10948
rect -11448 10868 -11428 10932
rect -11364 10868 -11344 10932
rect -11448 10852 -11344 10868
rect -17060 10492 -16956 10788
rect -22672 10412 -22568 10428
rect -22672 10348 -22652 10412
rect -22588 10348 -22568 10412
rect -22672 10332 -22568 10348
rect -22672 10268 -22652 10332
rect -22588 10268 -22568 10332
rect -22672 10252 -22568 10268
rect -22672 10188 -22652 10252
rect -22588 10188 -22568 10252
rect -22672 10172 -22568 10188
rect -22672 10108 -22652 10172
rect -22588 10108 -22568 10172
rect -22672 10092 -22568 10108
rect -22672 10028 -22652 10092
rect -22588 10028 -22568 10092
rect -22672 10012 -22568 10028
rect -22672 9948 -22652 10012
rect -22588 9948 -22568 10012
rect -22672 9932 -22568 9948
rect -22672 9868 -22652 9932
rect -22588 9868 -22568 9932
rect -22672 9852 -22568 9868
rect -22672 9788 -22652 9852
rect -22588 9788 -22568 9852
rect -22672 9772 -22568 9788
rect -22672 9708 -22652 9772
rect -22588 9708 -22568 9772
rect -22672 9692 -22568 9708
rect -22672 9628 -22652 9692
rect -22588 9628 -22568 9692
rect -22672 9612 -22568 9628
rect -22672 9548 -22652 9612
rect -22588 9548 -22568 9612
rect -22672 9532 -22568 9548
rect -22672 9468 -22652 9532
rect -22588 9468 -22568 9532
rect -22672 9452 -22568 9468
rect -22672 9388 -22652 9452
rect -22588 9388 -22568 9452
rect -22672 9372 -22568 9388
rect -22672 9308 -22652 9372
rect -22588 9308 -22568 9372
rect -22672 9292 -22568 9308
rect -22672 9228 -22652 9292
rect -22588 9228 -22568 9292
rect -22672 9212 -22568 9228
rect -22672 9148 -22652 9212
rect -22588 9148 -22568 9212
rect -22672 9132 -22568 9148
rect -22672 9068 -22652 9132
rect -22588 9068 -22568 9132
rect -22672 9052 -22568 9068
rect -22672 8988 -22652 9052
rect -22588 8988 -22568 9052
rect -22672 8972 -22568 8988
rect -22672 8908 -22652 8972
rect -22588 8908 -22568 8972
rect -22672 8892 -22568 8908
rect -22672 8828 -22652 8892
rect -22588 8828 -22568 8892
rect -22672 8812 -22568 8828
rect -22672 8748 -22652 8812
rect -22588 8748 -22568 8812
rect -22672 8732 -22568 8748
rect -22672 8668 -22652 8732
rect -22588 8668 -22568 8732
rect -22672 8652 -22568 8668
rect -22672 8588 -22652 8652
rect -22588 8588 -22568 8652
rect -22672 8572 -22568 8588
rect -22672 8508 -22652 8572
rect -22588 8508 -22568 8572
rect -22672 8492 -22568 8508
rect -22672 8428 -22652 8492
rect -22588 8428 -22568 8492
rect -22672 8412 -22568 8428
rect -22672 8348 -22652 8412
rect -22588 8348 -22568 8412
rect -22672 8332 -22568 8348
rect -22672 8268 -22652 8332
rect -22588 8268 -22568 8332
rect -22672 8252 -22568 8268
rect -22672 8188 -22652 8252
rect -22588 8188 -22568 8252
rect -22672 8172 -22568 8188
rect -22672 8108 -22652 8172
rect -22588 8108 -22568 8172
rect -22672 8092 -22568 8108
rect -22672 8028 -22652 8092
rect -22588 8028 -22568 8092
rect -22672 8012 -22568 8028
rect -22672 7948 -22652 8012
rect -22588 7948 -22568 8012
rect -22672 7932 -22568 7948
rect -22672 7868 -22652 7932
rect -22588 7868 -22568 7932
rect -22672 7852 -22568 7868
rect -22672 7788 -22652 7852
rect -22588 7788 -22568 7852
rect -22672 7772 -22568 7788
rect -22672 7708 -22652 7772
rect -22588 7708 -22568 7772
rect -22672 7692 -22568 7708
rect -22672 7628 -22652 7692
rect -22588 7628 -22568 7692
rect -22672 7612 -22568 7628
rect -22672 7548 -22652 7612
rect -22588 7548 -22568 7612
rect -22672 7532 -22568 7548
rect -22672 7468 -22652 7532
rect -22588 7468 -22568 7532
rect -22672 7452 -22568 7468
rect -22672 7388 -22652 7452
rect -22588 7388 -22568 7452
rect -22672 7372 -22568 7388
rect -22672 7308 -22652 7372
rect -22588 7308 -22568 7372
rect -22672 7292 -22568 7308
rect -22672 7228 -22652 7292
rect -22588 7228 -22568 7292
rect -22672 7212 -22568 7228
rect -22672 7148 -22652 7212
rect -22588 7148 -22568 7212
rect -22672 7132 -22568 7148
rect -22672 7068 -22652 7132
rect -22588 7068 -22568 7132
rect -22672 7052 -22568 7068
rect -22672 6988 -22652 7052
rect -22588 6988 -22568 7052
rect -22672 6972 -22568 6988
rect -22672 6908 -22652 6972
rect -22588 6908 -22568 6972
rect -22672 6892 -22568 6908
rect -22672 6828 -22652 6892
rect -22588 6828 -22568 6892
rect -22672 6812 -22568 6828
rect -22672 6748 -22652 6812
rect -22588 6748 -22568 6812
rect -22672 6732 -22568 6748
rect -22672 6668 -22652 6732
rect -22588 6668 -22568 6732
rect -22672 6652 -22568 6668
rect -22672 6588 -22652 6652
rect -22588 6588 -22568 6652
rect -22672 6572 -22568 6588
rect -22672 6508 -22652 6572
rect -22588 6508 -22568 6572
rect -22672 6492 -22568 6508
rect -22672 6428 -22652 6492
rect -22588 6428 -22568 6492
rect -22672 6412 -22568 6428
rect -22672 6348 -22652 6412
rect -22588 6348 -22568 6412
rect -22672 6332 -22568 6348
rect -22672 6268 -22652 6332
rect -22588 6268 -22568 6332
rect -22672 6252 -22568 6268
rect -22672 6188 -22652 6252
rect -22588 6188 -22568 6252
rect -22672 6172 -22568 6188
rect -22672 6108 -22652 6172
rect -22588 6108 -22568 6172
rect -22672 6092 -22568 6108
rect -22672 6028 -22652 6092
rect -22588 6028 -22568 6092
rect -22672 6012 -22568 6028
rect -22672 5948 -22652 6012
rect -22588 5948 -22568 6012
rect -22672 5932 -22568 5948
rect -22672 5868 -22652 5932
rect -22588 5868 -22568 5932
rect -22672 5852 -22568 5868
rect -22672 5788 -22652 5852
rect -22588 5788 -22568 5852
rect -22672 5772 -22568 5788
rect -22672 5708 -22652 5772
rect -22588 5708 -22568 5772
rect -22672 5692 -22568 5708
rect -22672 5628 -22652 5692
rect -22588 5628 -22568 5692
rect -22672 5612 -22568 5628
rect -22672 5548 -22652 5612
rect -22588 5548 -22568 5612
rect -22672 5532 -22568 5548
rect -28284 5172 -28180 5468
rect -33896 5092 -33792 5108
rect -33896 5028 -33876 5092
rect -33812 5028 -33792 5092
rect -33896 5012 -33792 5028
rect -33896 4948 -33876 5012
rect -33812 4948 -33792 5012
rect -33896 4932 -33792 4948
rect -33896 4868 -33876 4932
rect -33812 4868 -33792 4932
rect -33896 4852 -33792 4868
rect -33896 4788 -33876 4852
rect -33812 4788 -33792 4852
rect -33896 4772 -33792 4788
rect -33896 4708 -33876 4772
rect -33812 4708 -33792 4772
rect -33896 4692 -33792 4708
rect -33896 4628 -33876 4692
rect -33812 4628 -33792 4692
rect -33896 4612 -33792 4628
rect -33896 4548 -33876 4612
rect -33812 4548 -33792 4612
rect -33896 4532 -33792 4548
rect -33896 4468 -33876 4532
rect -33812 4468 -33792 4532
rect -33896 4452 -33792 4468
rect -33896 4388 -33876 4452
rect -33812 4388 -33792 4452
rect -33896 4372 -33792 4388
rect -33896 4308 -33876 4372
rect -33812 4308 -33792 4372
rect -33896 4292 -33792 4308
rect -33896 4228 -33876 4292
rect -33812 4228 -33792 4292
rect -33896 4212 -33792 4228
rect -33896 4148 -33876 4212
rect -33812 4148 -33792 4212
rect -33896 4132 -33792 4148
rect -33896 4068 -33876 4132
rect -33812 4068 -33792 4132
rect -33896 4052 -33792 4068
rect -33896 3988 -33876 4052
rect -33812 3988 -33792 4052
rect -33896 3972 -33792 3988
rect -33896 3908 -33876 3972
rect -33812 3908 -33792 3972
rect -33896 3892 -33792 3908
rect -33896 3828 -33876 3892
rect -33812 3828 -33792 3892
rect -33896 3812 -33792 3828
rect -33896 3748 -33876 3812
rect -33812 3748 -33792 3812
rect -33896 3732 -33792 3748
rect -33896 3668 -33876 3732
rect -33812 3668 -33792 3732
rect -33896 3652 -33792 3668
rect -33896 3588 -33876 3652
rect -33812 3588 -33792 3652
rect -33896 3572 -33792 3588
rect -33896 3508 -33876 3572
rect -33812 3508 -33792 3572
rect -33896 3492 -33792 3508
rect -33896 3428 -33876 3492
rect -33812 3428 -33792 3492
rect -33896 3412 -33792 3428
rect -33896 3348 -33876 3412
rect -33812 3348 -33792 3412
rect -33896 3332 -33792 3348
rect -33896 3268 -33876 3332
rect -33812 3268 -33792 3332
rect -33896 3252 -33792 3268
rect -33896 3188 -33876 3252
rect -33812 3188 -33792 3252
rect -33896 3172 -33792 3188
rect -33896 3108 -33876 3172
rect -33812 3108 -33792 3172
rect -33896 3092 -33792 3108
rect -33896 3028 -33876 3092
rect -33812 3028 -33792 3092
rect -33896 3012 -33792 3028
rect -33896 2948 -33876 3012
rect -33812 2948 -33792 3012
rect -33896 2932 -33792 2948
rect -33896 2868 -33876 2932
rect -33812 2868 -33792 2932
rect -33896 2852 -33792 2868
rect -33896 2788 -33876 2852
rect -33812 2788 -33792 2852
rect -33896 2772 -33792 2788
rect -33896 2708 -33876 2772
rect -33812 2708 -33792 2772
rect -33896 2692 -33792 2708
rect -33896 2628 -33876 2692
rect -33812 2628 -33792 2692
rect -33896 2612 -33792 2628
rect -33896 2548 -33876 2612
rect -33812 2548 -33792 2612
rect -33896 2532 -33792 2548
rect -33896 2468 -33876 2532
rect -33812 2468 -33792 2532
rect -33896 2452 -33792 2468
rect -33896 2388 -33876 2452
rect -33812 2388 -33792 2452
rect -33896 2372 -33792 2388
rect -33896 2308 -33876 2372
rect -33812 2308 -33792 2372
rect -33896 2292 -33792 2308
rect -33896 2228 -33876 2292
rect -33812 2228 -33792 2292
rect -33896 2212 -33792 2228
rect -33896 2148 -33876 2212
rect -33812 2148 -33792 2212
rect -33896 2132 -33792 2148
rect -33896 2068 -33876 2132
rect -33812 2068 -33792 2132
rect -33896 2052 -33792 2068
rect -33896 1988 -33876 2052
rect -33812 1988 -33792 2052
rect -33896 1972 -33792 1988
rect -33896 1908 -33876 1972
rect -33812 1908 -33792 1972
rect -33896 1892 -33792 1908
rect -33896 1828 -33876 1892
rect -33812 1828 -33792 1892
rect -33896 1812 -33792 1828
rect -33896 1748 -33876 1812
rect -33812 1748 -33792 1812
rect -33896 1732 -33792 1748
rect -33896 1668 -33876 1732
rect -33812 1668 -33792 1732
rect -33896 1652 -33792 1668
rect -33896 1588 -33876 1652
rect -33812 1588 -33792 1652
rect -33896 1572 -33792 1588
rect -33896 1508 -33876 1572
rect -33812 1508 -33792 1572
rect -33896 1492 -33792 1508
rect -33896 1428 -33876 1492
rect -33812 1428 -33792 1492
rect -33896 1412 -33792 1428
rect -33896 1348 -33876 1412
rect -33812 1348 -33792 1412
rect -33896 1332 -33792 1348
rect -33896 1268 -33876 1332
rect -33812 1268 -33792 1332
rect -33896 1252 -33792 1268
rect -33896 1188 -33876 1252
rect -33812 1188 -33792 1252
rect -33896 1172 -33792 1188
rect -33896 1108 -33876 1172
rect -33812 1108 -33792 1172
rect -33896 1092 -33792 1108
rect -33896 1028 -33876 1092
rect -33812 1028 -33792 1092
rect -33896 1012 -33792 1028
rect -33896 948 -33876 1012
rect -33812 948 -33792 1012
rect -33896 932 -33792 948
rect -33896 868 -33876 932
rect -33812 868 -33792 932
rect -33896 852 -33792 868
rect -33896 788 -33876 852
rect -33812 788 -33792 852
rect -33896 772 -33792 788
rect -33896 708 -33876 772
rect -33812 708 -33792 772
rect -33896 692 -33792 708
rect -33896 628 -33876 692
rect -33812 628 -33792 692
rect -33896 612 -33792 628
rect -33896 548 -33876 612
rect -33812 548 -33792 612
rect -33896 532 -33792 548
rect -33896 468 -33876 532
rect -33812 468 -33792 532
rect -33896 452 -33792 468
rect -33896 388 -33876 452
rect -33812 388 -33792 452
rect -33896 372 -33792 388
rect -33896 308 -33876 372
rect -33812 308 -33792 372
rect -33896 292 -33792 308
rect -33896 228 -33876 292
rect -33812 228 -33792 292
rect -33896 212 -33792 228
rect -36676 -199 -36572 199
rect -33896 148 -33876 212
rect -33812 148 -33792 212
rect -33473 5092 -28551 5121
rect -33473 228 -33444 5092
rect -28580 228 -28551 5092
rect -33473 199 -28551 228
rect -28284 5108 -28264 5172
rect -28200 5108 -28180 5172
rect -25452 5121 -25348 5519
rect -22672 5468 -22652 5532
rect -22588 5468 -22568 5532
rect -22249 10412 -17327 10441
rect -22249 5548 -22220 10412
rect -17356 5548 -17327 10412
rect -22249 5519 -17327 5548
rect -17060 10428 -17040 10492
rect -16976 10428 -16956 10492
rect -14228 10441 -14124 10839
rect -11448 10788 -11428 10852
rect -11364 10788 -11344 10852
rect -11025 15732 -6103 15761
rect -11025 10868 -10996 15732
rect -6132 10868 -6103 15732
rect -11025 10839 -6103 10868
rect -5836 15748 -5816 15812
rect -5752 15748 -5732 15812
rect -3004 15761 -2900 16159
rect -224 16108 -204 16172
rect -140 16108 -120 16172
rect 199 21052 5121 21081
rect 199 16188 228 21052
rect 5092 16188 5121 21052
rect 199 16159 5121 16188
rect 5388 21068 5408 21132
rect 5472 21068 5492 21132
rect 8220 21081 8324 21479
rect 11000 21428 11020 21492
rect 11084 21428 11104 21492
rect 11423 26372 16345 26401
rect 11423 21508 11452 26372
rect 16316 21508 16345 26372
rect 11423 21479 16345 21508
rect 16612 26388 16632 26452
rect 16696 26388 16716 26452
rect 19444 26401 19548 26799
rect 22224 26748 22244 26812
rect 22308 26748 22328 26812
rect 22647 31692 27569 31721
rect 22647 26828 22676 31692
rect 27540 26828 27569 31692
rect 22647 26799 27569 26828
rect 27836 31708 27856 31772
rect 27920 31708 27940 31772
rect 30668 31721 30772 32119
rect 33448 32068 33468 32132
rect 33532 32068 33552 32132
rect 33871 37012 38793 37041
rect 33871 32148 33900 37012
rect 38764 32148 38793 37012
rect 33871 32119 38793 32148
rect 39060 37028 39080 37092
rect 39144 37028 39164 37092
rect 39060 37012 39164 37028
rect 39060 36948 39080 37012
rect 39144 36948 39164 37012
rect 39060 36932 39164 36948
rect 39060 36868 39080 36932
rect 39144 36868 39164 36932
rect 39060 36852 39164 36868
rect 39060 36788 39080 36852
rect 39144 36788 39164 36852
rect 39060 36772 39164 36788
rect 39060 36708 39080 36772
rect 39144 36708 39164 36772
rect 39060 36692 39164 36708
rect 39060 36628 39080 36692
rect 39144 36628 39164 36692
rect 39060 36612 39164 36628
rect 39060 36548 39080 36612
rect 39144 36548 39164 36612
rect 39060 36532 39164 36548
rect 39060 36468 39080 36532
rect 39144 36468 39164 36532
rect 39060 36452 39164 36468
rect 39060 36388 39080 36452
rect 39144 36388 39164 36452
rect 39060 36372 39164 36388
rect 39060 36308 39080 36372
rect 39144 36308 39164 36372
rect 39060 36292 39164 36308
rect 39060 36228 39080 36292
rect 39144 36228 39164 36292
rect 39060 36212 39164 36228
rect 39060 36148 39080 36212
rect 39144 36148 39164 36212
rect 39060 36132 39164 36148
rect 39060 36068 39080 36132
rect 39144 36068 39164 36132
rect 39060 36052 39164 36068
rect 39060 35988 39080 36052
rect 39144 35988 39164 36052
rect 39060 35972 39164 35988
rect 39060 35908 39080 35972
rect 39144 35908 39164 35972
rect 39060 35892 39164 35908
rect 39060 35828 39080 35892
rect 39144 35828 39164 35892
rect 39060 35812 39164 35828
rect 39060 35748 39080 35812
rect 39144 35748 39164 35812
rect 39060 35732 39164 35748
rect 39060 35668 39080 35732
rect 39144 35668 39164 35732
rect 39060 35652 39164 35668
rect 39060 35588 39080 35652
rect 39144 35588 39164 35652
rect 39060 35572 39164 35588
rect 39060 35508 39080 35572
rect 39144 35508 39164 35572
rect 39060 35492 39164 35508
rect 39060 35428 39080 35492
rect 39144 35428 39164 35492
rect 39060 35412 39164 35428
rect 39060 35348 39080 35412
rect 39144 35348 39164 35412
rect 39060 35332 39164 35348
rect 39060 35268 39080 35332
rect 39144 35268 39164 35332
rect 39060 35252 39164 35268
rect 39060 35188 39080 35252
rect 39144 35188 39164 35252
rect 39060 35172 39164 35188
rect 39060 35108 39080 35172
rect 39144 35108 39164 35172
rect 39060 35092 39164 35108
rect 39060 35028 39080 35092
rect 39144 35028 39164 35092
rect 39060 35012 39164 35028
rect 39060 34948 39080 35012
rect 39144 34948 39164 35012
rect 39060 34932 39164 34948
rect 39060 34868 39080 34932
rect 39144 34868 39164 34932
rect 39060 34852 39164 34868
rect 39060 34788 39080 34852
rect 39144 34788 39164 34852
rect 39060 34772 39164 34788
rect 39060 34708 39080 34772
rect 39144 34708 39164 34772
rect 39060 34692 39164 34708
rect 39060 34628 39080 34692
rect 39144 34628 39164 34692
rect 39060 34612 39164 34628
rect 39060 34548 39080 34612
rect 39144 34548 39164 34612
rect 39060 34532 39164 34548
rect 39060 34468 39080 34532
rect 39144 34468 39164 34532
rect 39060 34452 39164 34468
rect 39060 34388 39080 34452
rect 39144 34388 39164 34452
rect 39060 34372 39164 34388
rect 39060 34308 39080 34372
rect 39144 34308 39164 34372
rect 39060 34292 39164 34308
rect 39060 34228 39080 34292
rect 39144 34228 39164 34292
rect 39060 34212 39164 34228
rect 39060 34148 39080 34212
rect 39144 34148 39164 34212
rect 39060 34132 39164 34148
rect 39060 34068 39080 34132
rect 39144 34068 39164 34132
rect 39060 34052 39164 34068
rect 39060 33988 39080 34052
rect 39144 33988 39164 34052
rect 39060 33972 39164 33988
rect 39060 33908 39080 33972
rect 39144 33908 39164 33972
rect 39060 33892 39164 33908
rect 39060 33828 39080 33892
rect 39144 33828 39164 33892
rect 39060 33812 39164 33828
rect 39060 33748 39080 33812
rect 39144 33748 39164 33812
rect 39060 33732 39164 33748
rect 39060 33668 39080 33732
rect 39144 33668 39164 33732
rect 39060 33652 39164 33668
rect 39060 33588 39080 33652
rect 39144 33588 39164 33652
rect 39060 33572 39164 33588
rect 39060 33508 39080 33572
rect 39144 33508 39164 33572
rect 39060 33492 39164 33508
rect 39060 33428 39080 33492
rect 39144 33428 39164 33492
rect 39060 33412 39164 33428
rect 39060 33348 39080 33412
rect 39144 33348 39164 33412
rect 39060 33332 39164 33348
rect 39060 33268 39080 33332
rect 39144 33268 39164 33332
rect 39060 33252 39164 33268
rect 39060 33188 39080 33252
rect 39144 33188 39164 33252
rect 39060 33172 39164 33188
rect 39060 33108 39080 33172
rect 39144 33108 39164 33172
rect 39060 33092 39164 33108
rect 39060 33028 39080 33092
rect 39144 33028 39164 33092
rect 39060 33012 39164 33028
rect 39060 32948 39080 33012
rect 39144 32948 39164 33012
rect 39060 32932 39164 32948
rect 39060 32868 39080 32932
rect 39144 32868 39164 32932
rect 39060 32852 39164 32868
rect 39060 32788 39080 32852
rect 39144 32788 39164 32852
rect 39060 32772 39164 32788
rect 39060 32708 39080 32772
rect 39144 32708 39164 32772
rect 39060 32692 39164 32708
rect 39060 32628 39080 32692
rect 39144 32628 39164 32692
rect 39060 32612 39164 32628
rect 39060 32548 39080 32612
rect 39144 32548 39164 32612
rect 39060 32532 39164 32548
rect 39060 32468 39080 32532
rect 39144 32468 39164 32532
rect 39060 32452 39164 32468
rect 39060 32388 39080 32452
rect 39144 32388 39164 32452
rect 39060 32372 39164 32388
rect 39060 32308 39080 32372
rect 39144 32308 39164 32372
rect 39060 32292 39164 32308
rect 39060 32228 39080 32292
rect 39144 32228 39164 32292
rect 39060 32212 39164 32228
rect 39060 32148 39080 32212
rect 39144 32148 39164 32212
rect 39060 32132 39164 32148
rect 33448 31772 33552 32068
rect 27836 31692 27940 31708
rect 27836 31628 27856 31692
rect 27920 31628 27940 31692
rect 27836 31612 27940 31628
rect 27836 31548 27856 31612
rect 27920 31548 27940 31612
rect 27836 31532 27940 31548
rect 27836 31468 27856 31532
rect 27920 31468 27940 31532
rect 27836 31452 27940 31468
rect 27836 31388 27856 31452
rect 27920 31388 27940 31452
rect 27836 31372 27940 31388
rect 27836 31308 27856 31372
rect 27920 31308 27940 31372
rect 27836 31292 27940 31308
rect 27836 31228 27856 31292
rect 27920 31228 27940 31292
rect 27836 31212 27940 31228
rect 27836 31148 27856 31212
rect 27920 31148 27940 31212
rect 27836 31132 27940 31148
rect 27836 31068 27856 31132
rect 27920 31068 27940 31132
rect 27836 31052 27940 31068
rect 27836 30988 27856 31052
rect 27920 30988 27940 31052
rect 27836 30972 27940 30988
rect 27836 30908 27856 30972
rect 27920 30908 27940 30972
rect 27836 30892 27940 30908
rect 27836 30828 27856 30892
rect 27920 30828 27940 30892
rect 27836 30812 27940 30828
rect 27836 30748 27856 30812
rect 27920 30748 27940 30812
rect 27836 30732 27940 30748
rect 27836 30668 27856 30732
rect 27920 30668 27940 30732
rect 27836 30652 27940 30668
rect 27836 30588 27856 30652
rect 27920 30588 27940 30652
rect 27836 30572 27940 30588
rect 27836 30508 27856 30572
rect 27920 30508 27940 30572
rect 27836 30492 27940 30508
rect 27836 30428 27856 30492
rect 27920 30428 27940 30492
rect 27836 30412 27940 30428
rect 27836 30348 27856 30412
rect 27920 30348 27940 30412
rect 27836 30332 27940 30348
rect 27836 30268 27856 30332
rect 27920 30268 27940 30332
rect 27836 30252 27940 30268
rect 27836 30188 27856 30252
rect 27920 30188 27940 30252
rect 27836 30172 27940 30188
rect 27836 30108 27856 30172
rect 27920 30108 27940 30172
rect 27836 30092 27940 30108
rect 27836 30028 27856 30092
rect 27920 30028 27940 30092
rect 27836 30012 27940 30028
rect 27836 29948 27856 30012
rect 27920 29948 27940 30012
rect 27836 29932 27940 29948
rect 27836 29868 27856 29932
rect 27920 29868 27940 29932
rect 27836 29852 27940 29868
rect 27836 29788 27856 29852
rect 27920 29788 27940 29852
rect 27836 29772 27940 29788
rect 27836 29708 27856 29772
rect 27920 29708 27940 29772
rect 27836 29692 27940 29708
rect 27836 29628 27856 29692
rect 27920 29628 27940 29692
rect 27836 29612 27940 29628
rect 27836 29548 27856 29612
rect 27920 29548 27940 29612
rect 27836 29532 27940 29548
rect 27836 29468 27856 29532
rect 27920 29468 27940 29532
rect 27836 29452 27940 29468
rect 27836 29388 27856 29452
rect 27920 29388 27940 29452
rect 27836 29372 27940 29388
rect 27836 29308 27856 29372
rect 27920 29308 27940 29372
rect 27836 29292 27940 29308
rect 27836 29228 27856 29292
rect 27920 29228 27940 29292
rect 27836 29212 27940 29228
rect 27836 29148 27856 29212
rect 27920 29148 27940 29212
rect 27836 29132 27940 29148
rect 27836 29068 27856 29132
rect 27920 29068 27940 29132
rect 27836 29052 27940 29068
rect 27836 28988 27856 29052
rect 27920 28988 27940 29052
rect 27836 28972 27940 28988
rect 27836 28908 27856 28972
rect 27920 28908 27940 28972
rect 27836 28892 27940 28908
rect 27836 28828 27856 28892
rect 27920 28828 27940 28892
rect 27836 28812 27940 28828
rect 27836 28748 27856 28812
rect 27920 28748 27940 28812
rect 27836 28732 27940 28748
rect 27836 28668 27856 28732
rect 27920 28668 27940 28732
rect 27836 28652 27940 28668
rect 27836 28588 27856 28652
rect 27920 28588 27940 28652
rect 27836 28572 27940 28588
rect 27836 28508 27856 28572
rect 27920 28508 27940 28572
rect 27836 28492 27940 28508
rect 27836 28428 27856 28492
rect 27920 28428 27940 28492
rect 27836 28412 27940 28428
rect 27836 28348 27856 28412
rect 27920 28348 27940 28412
rect 27836 28332 27940 28348
rect 27836 28268 27856 28332
rect 27920 28268 27940 28332
rect 27836 28252 27940 28268
rect 27836 28188 27856 28252
rect 27920 28188 27940 28252
rect 27836 28172 27940 28188
rect 27836 28108 27856 28172
rect 27920 28108 27940 28172
rect 27836 28092 27940 28108
rect 27836 28028 27856 28092
rect 27920 28028 27940 28092
rect 27836 28012 27940 28028
rect 27836 27948 27856 28012
rect 27920 27948 27940 28012
rect 27836 27932 27940 27948
rect 27836 27868 27856 27932
rect 27920 27868 27940 27932
rect 27836 27852 27940 27868
rect 27836 27788 27856 27852
rect 27920 27788 27940 27852
rect 27836 27772 27940 27788
rect 27836 27708 27856 27772
rect 27920 27708 27940 27772
rect 27836 27692 27940 27708
rect 27836 27628 27856 27692
rect 27920 27628 27940 27692
rect 27836 27612 27940 27628
rect 27836 27548 27856 27612
rect 27920 27548 27940 27612
rect 27836 27532 27940 27548
rect 27836 27468 27856 27532
rect 27920 27468 27940 27532
rect 27836 27452 27940 27468
rect 27836 27388 27856 27452
rect 27920 27388 27940 27452
rect 27836 27372 27940 27388
rect 27836 27308 27856 27372
rect 27920 27308 27940 27372
rect 27836 27292 27940 27308
rect 27836 27228 27856 27292
rect 27920 27228 27940 27292
rect 27836 27212 27940 27228
rect 27836 27148 27856 27212
rect 27920 27148 27940 27212
rect 27836 27132 27940 27148
rect 27836 27068 27856 27132
rect 27920 27068 27940 27132
rect 27836 27052 27940 27068
rect 27836 26988 27856 27052
rect 27920 26988 27940 27052
rect 27836 26972 27940 26988
rect 27836 26908 27856 26972
rect 27920 26908 27940 26972
rect 27836 26892 27940 26908
rect 27836 26828 27856 26892
rect 27920 26828 27940 26892
rect 27836 26812 27940 26828
rect 22224 26452 22328 26748
rect 16612 26372 16716 26388
rect 16612 26308 16632 26372
rect 16696 26308 16716 26372
rect 16612 26292 16716 26308
rect 16612 26228 16632 26292
rect 16696 26228 16716 26292
rect 16612 26212 16716 26228
rect 16612 26148 16632 26212
rect 16696 26148 16716 26212
rect 16612 26132 16716 26148
rect 16612 26068 16632 26132
rect 16696 26068 16716 26132
rect 16612 26052 16716 26068
rect 16612 25988 16632 26052
rect 16696 25988 16716 26052
rect 16612 25972 16716 25988
rect 16612 25908 16632 25972
rect 16696 25908 16716 25972
rect 16612 25892 16716 25908
rect 16612 25828 16632 25892
rect 16696 25828 16716 25892
rect 16612 25812 16716 25828
rect 16612 25748 16632 25812
rect 16696 25748 16716 25812
rect 16612 25732 16716 25748
rect 16612 25668 16632 25732
rect 16696 25668 16716 25732
rect 16612 25652 16716 25668
rect 16612 25588 16632 25652
rect 16696 25588 16716 25652
rect 16612 25572 16716 25588
rect 16612 25508 16632 25572
rect 16696 25508 16716 25572
rect 16612 25492 16716 25508
rect 16612 25428 16632 25492
rect 16696 25428 16716 25492
rect 16612 25412 16716 25428
rect 16612 25348 16632 25412
rect 16696 25348 16716 25412
rect 16612 25332 16716 25348
rect 16612 25268 16632 25332
rect 16696 25268 16716 25332
rect 16612 25252 16716 25268
rect 16612 25188 16632 25252
rect 16696 25188 16716 25252
rect 16612 25172 16716 25188
rect 16612 25108 16632 25172
rect 16696 25108 16716 25172
rect 16612 25092 16716 25108
rect 16612 25028 16632 25092
rect 16696 25028 16716 25092
rect 16612 25012 16716 25028
rect 16612 24948 16632 25012
rect 16696 24948 16716 25012
rect 16612 24932 16716 24948
rect 16612 24868 16632 24932
rect 16696 24868 16716 24932
rect 16612 24852 16716 24868
rect 16612 24788 16632 24852
rect 16696 24788 16716 24852
rect 16612 24772 16716 24788
rect 16612 24708 16632 24772
rect 16696 24708 16716 24772
rect 16612 24692 16716 24708
rect 16612 24628 16632 24692
rect 16696 24628 16716 24692
rect 16612 24612 16716 24628
rect 16612 24548 16632 24612
rect 16696 24548 16716 24612
rect 16612 24532 16716 24548
rect 16612 24468 16632 24532
rect 16696 24468 16716 24532
rect 16612 24452 16716 24468
rect 16612 24388 16632 24452
rect 16696 24388 16716 24452
rect 16612 24372 16716 24388
rect 16612 24308 16632 24372
rect 16696 24308 16716 24372
rect 16612 24292 16716 24308
rect 16612 24228 16632 24292
rect 16696 24228 16716 24292
rect 16612 24212 16716 24228
rect 16612 24148 16632 24212
rect 16696 24148 16716 24212
rect 16612 24132 16716 24148
rect 16612 24068 16632 24132
rect 16696 24068 16716 24132
rect 16612 24052 16716 24068
rect 16612 23988 16632 24052
rect 16696 23988 16716 24052
rect 16612 23972 16716 23988
rect 16612 23908 16632 23972
rect 16696 23908 16716 23972
rect 16612 23892 16716 23908
rect 16612 23828 16632 23892
rect 16696 23828 16716 23892
rect 16612 23812 16716 23828
rect 16612 23748 16632 23812
rect 16696 23748 16716 23812
rect 16612 23732 16716 23748
rect 16612 23668 16632 23732
rect 16696 23668 16716 23732
rect 16612 23652 16716 23668
rect 16612 23588 16632 23652
rect 16696 23588 16716 23652
rect 16612 23572 16716 23588
rect 16612 23508 16632 23572
rect 16696 23508 16716 23572
rect 16612 23492 16716 23508
rect 16612 23428 16632 23492
rect 16696 23428 16716 23492
rect 16612 23412 16716 23428
rect 16612 23348 16632 23412
rect 16696 23348 16716 23412
rect 16612 23332 16716 23348
rect 16612 23268 16632 23332
rect 16696 23268 16716 23332
rect 16612 23252 16716 23268
rect 16612 23188 16632 23252
rect 16696 23188 16716 23252
rect 16612 23172 16716 23188
rect 16612 23108 16632 23172
rect 16696 23108 16716 23172
rect 16612 23092 16716 23108
rect 16612 23028 16632 23092
rect 16696 23028 16716 23092
rect 16612 23012 16716 23028
rect 16612 22948 16632 23012
rect 16696 22948 16716 23012
rect 16612 22932 16716 22948
rect 16612 22868 16632 22932
rect 16696 22868 16716 22932
rect 16612 22852 16716 22868
rect 16612 22788 16632 22852
rect 16696 22788 16716 22852
rect 16612 22772 16716 22788
rect 16612 22708 16632 22772
rect 16696 22708 16716 22772
rect 16612 22692 16716 22708
rect 16612 22628 16632 22692
rect 16696 22628 16716 22692
rect 16612 22612 16716 22628
rect 16612 22548 16632 22612
rect 16696 22548 16716 22612
rect 16612 22532 16716 22548
rect 16612 22468 16632 22532
rect 16696 22468 16716 22532
rect 16612 22452 16716 22468
rect 16612 22388 16632 22452
rect 16696 22388 16716 22452
rect 16612 22372 16716 22388
rect 16612 22308 16632 22372
rect 16696 22308 16716 22372
rect 16612 22292 16716 22308
rect 16612 22228 16632 22292
rect 16696 22228 16716 22292
rect 16612 22212 16716 22228
rect 16612 22148 16632 22212
rect 16696 22148 16716 22212
rect 16612 22132 16716 22148
rect 16612 22068 16632 22132
rect 16696 22068 16716 22132
rect 16612 22052 16716 22068
rect 16612 21988 16632 22052
rect 16696 21988 16716 22052
rect 16612 21972 16716 21988
rect 16612 21908 16632 21972
rect 16696 21908 16716 21972
rect 16612 21892 16716 21908
rect 16612 21828 16632 21892
rect 16696 21828 16716 21892
rect 16612 21812 16716 21828
rect 16612 21748 16632 21812
rect 16696 21748 16716 21812
rect 16612 21732 16716 21748
rect 16612 21668 16632 21732
rect 16696 21668 16716 21732
rect 16612 21652 16716 21668
rect 16612 21588 16632 21652
rect 16696 21588 16716 21652
rect 16612 21572 16716 21588
rect 16612 21508 16632 21572
rect 16696 21508 16716 21572
rect 16612 21492 16716 21508
rect 11000 21132 11104 21428
rect 5388 21052 5492 21068
rect 5388 20988 5408 21052
rect 5472 20988 5492 21052
rect 5388 20972 5492 20988
rect 5388 20908 5408 20972
rect 5472 20908 5492 20972
rect 5388 20892 5492 20908
rect 5388 20828 5408 20892
rect 5472 20828 5492 20892
rect 5388 20812 5492 20828
rect 5388 20748 5408 20812
rect 5472 20748 5492 20812
rect 5388 20732 5492 20748
rect 5388 20668 5408 20732
rect 5472 20668 5492 20732
rect 5388 20652 5492 20668
rect 5388 20588 5408 20652
rect 5472 20588 5492 20652
rect 5388 20572 5492 20588
rect 5388 20508 5408 20572
rect 5472 20508 5492 20572
rect 5388 20492 5492 20508
rect 5388 20428 5408 20492
rect 5472 20428 5492 20492
rect 5388 20412 5492 20428
rect 5388 20348 5408 20412
rect 5472 20348 5492 20412
rect 5388 20332 5492 20348
rect 5388 20268 5408 20332
rect 5472 20268 5492 20332
rect 5388 20252 5492 20268
rect 5388 20188 5408 20252
rect 5472 20188 5492 20252
rect 5388 20172 5492 20188
rect 5388 20108 5408 20172
rect 5472 20108 5492 20172
rect 5388 20092 5492 20108
rect 5388 20028 5408 20092
rect 5472 20028 5492 20092
rect 5388 20012 5492 20028
rect 5388 19948 5408 20012
rect 5472 19948 5492 20012
rect 5388 19932 5492 19948
rect 5388 19868 5408 19932
rect 5472 19868 5492 19932
rect 5388 19852 5492 19868
rect 5388 19788 5408 19852
rect 5472 19788 5492 19852
rect 5388 19772 5492 19788
rect 5388 19708 5408 19772
rect 5472 19708 5492 19772
rect 5388 19692 5492 19708
rect 5388 19628 5408 19692
rect 5472 19628 5492 19692
rect 5388 19612 5492 19628
rect 5388 19548 5408 19612
rect 5472 19548 5492 19612
rect 5388 19532 5492 19548
rect 5388 19468 5408 19532
rect 5472 19468 5492 19532
rect 5388 19452 5492 19468
rect 5388 19388 5408 19452
rect 5472 19388 5492 19452
rect 5388 19372 5492 19388
rect 5388 19308 5408 19372
rect 5472 19308 5492 19372
rect 5388 19292 5492 19308
rect 5388 19228 5408 19292
rect 5472 19228 5492 19292
rect 5388 19212 5492 19228
rect 5388 19148 5408 19212
rect 5472 19148 5492 19212
rect 5388 19132 5492 19148
rect 5388 19068 5408 19132
rect 5472 19068 5492 19132
rect 5388 19052 5492 19068
rect 5388 18988 5408 19052
rect 5472 18988 5492 19052
rect 5388 18972 5492 18988
rect 5388 18908 5408 18972
rect 5472 18908 5492 18972
rect 5388 18892 5492 18908
rect 5388 18828 5408 18892
rect 5472 18828 5492 18892
rect 5388 18812 5492 18828
rect 5388 18748 5408 18812
rect 5472 18748 5492 18812
rect 5388 18732 5492 18748
rect 5388 18668 5408 18732
rect 5472 18668 5492 18732
rect 5388 18652 5492 18668
rect 5388 18588 5408 18652
rect 5472 18588 5492 18652
rect 5388 18572 5492 18588
rect 5388 18508 5408 18572
rect 5472 18508 5492 18572
rect 5388 18492 5492 18508
rect 5388 18428 5408 18492
rect 5472 18428 5492 18492
rect 5388 18412 5492 18428
rect 5388 18348 5408 18412
rect 5472 18348 5492 18412
rect 5388 18332 5492 18348
rect 5388 18268 5408 18332
rect 5472 18268 5492 18332
rect 5388 18252 5492 18268
rect 5388 18188 5408 18252
rect 5472 18188 5492 18252
rect 5388 18172 5492 18188
rect 5388 18108 5408 18172
rect 5472 18108 5492 18172
rect 5388 18092 5492 18108
rect 5388 18028 5408 18092
rect 5472 18028 5492 18092
rect 5388 18012 5492 18028
rect 5388 17948 5408 18012
rect 5472 17948 5492 18012
rect 5388 17932 5492 17948
rect 5388 17868 5408 17932
rect 5472 17868 5492 17932
rect 5388 17852 5492 17868
rect 5388 17788 5408 17852
rect 5472 17788 5492 17852
rect 5388 17772 5492 17788
rect 5388 17708 5408 17772
rect 5472 17708 5492 17772
rect 5388 17692 5492 17708
rect 5388 17628 5408 17692
rect 5472 17628 5492 17692
rect 5388 17612 5492 17628
rect 5388 17548 5408 17612
rect 5472 17548 5492 17612
rect 5388 17532 5492 17548
rect 5388 17468 5408 17532
rect 5472 17468 5492 17532
rect 5388 17452 5492 17468
rect 5388 17388 5408 17452
rect 5472 17388 5492 17452
rect 5388 17372 5492 17388
rect 5388 17308 5408 17372
rect 5472 17308 5492 17372
rect 5388 17292 5492 17308
rect 5388 17228 5408 17292
rect 5472 17228 5492 17292
rect 5388 17212 5492 17228
rect 5388 17148 5408 17212
rect 5472 17148 5492 17212
rect 5388 17132 5492 17148
rect 5388 17068 5408 17132
rect 5472 17068 5492 17132
rect 5388 17052 5492 17068
rect 5388 16988 5408 17052
rect 5472 16988 5492 17052
rect 5388 16972 5492 16988
rect 5388 16908 5408 16972
rect 5472 16908 5492 16972
rect 5388 16892 5492 16908
rect 5388 16828 5408 16892
rect 5472 16828 5492 16892
rect 5388 16812 5492 16828
rect 5388 16748 5408 16812
rect 5472 16748 5492 16812
rect 5388 16732 5492 16748
rect 5388 16668 5408 16732
rect 5472 16668 5492 16732
rect 5388 16652 5492 16668
rect 5388 16588 5408 16652
rect 5472 16588 5492 16652
rect 5388 16572 5492 16588
rect 5388 16508 5408 16572
rect 5472 16508 5492 16572
rect 5388 16492 5492 16508
rect 5388 16428 5408 16492
rect 5472 16428 5492 16492
rect 5388 16412 5492 16428
rect 5388 16348 5408 16412
rect 5472 16348 5492 16412
rect 5388 16332 5492 16348
rect 5388 16268 5408 16332
rect 5472 16268 5492 16332
rect 5388 16252 5492 16268
rect 5388 16188 5408 16252
rect 5472 16188 5492 16252
rect 5388 16172 5492 16188
rect -224 15812 -120 16108
rect -5836 15732 -5732 15748
rect -5836 15668 -5816 15732
rect -5752 15668 -5732 15732
rect -5836 15652 -5732 15668
rect -5836 15588 -5816 15652
rect -5752 15588 -5732 15652
rect -5836 15572 -5732 15588
rect -5836 15508 -5816 15572
rect -5752 15508 -5732 15572
rect -5836 15492 -5732 15508
rect -5836 15428 -5816 15492
rect -5752 15428 -5732 15492
rect -5836 15412 -5732 15428
rect -5836 15348 -5816 15412
rect -5752 15348 -5732 15412
rect -5836 15332 -5732 15348
rect -5836 15268 -5816 15332
rect -5752 15268 -5732 15332
rect -5836 15252 -5732 15268
rect -5836 15188 -5816 15252
rect -5752 15188 -5732 15252
rect -5836 15172 -5732 15188
rect -5836 15108 -5816 15172
rect -5752 15108 -5732 15172
rect -5836 15092 -5732 15108
rect -5836 15028 -5816 15092
rect -5752 15028 -5732 15092
rect -5836 15012 -5732 15028
rect -5836 14948 -5816 15012
rect -5752 14948 -5732 15012
rect -5836 14932 -5732 14948
rect -5836 14868 -5816 14932
rect -5752 14868 -5732 14932
rect -5836 14852 -5732 14868
rect -5836 14788 -5816 14852
rect -5752 14788 -5732 14852
rect -5836 14772 -5732 14788
rect -5836 14708 -5816 14772
rect -5752 14708 -5732 14772
rect -5836 14692 -5732 14708
rect -5836 14628 -5816 14692
rect -5752 14628 -5732 14692
rect -5836 14612 -5732 14628
rect -5836 14548 -5816 14612
rect -5752 14548 -5732 14612
rect -5836 14532 -5732 14548
rect -5836 14468 -5816 14532
rect -5752 14468 -5732 14532
rect -5836 14452 -5732 14468
rect -5836 14388 -5816 14452
rect -5752 14388 -5732 14452
rect -5836 14372 -5732 14388
rect -5836 14308 -5816 14372
rect -5752 14308 -5732 14372
rect -5836 14292 -5732 14308
rect -5836 14228 -5816 14292
rect -5752 14228 -5732 14292
rect -5836 14212 -5732 14228
rect -5836 14148 -5816 14212
rect -5752 14148 -5732 14212
rect -5836 14132 -5732 14148
rect -5836 14068 -5816 14132
rect -5752 14068 -5732 14132
rect -5836 14052 -5732 14068
rect -5836 13988 -5816 14052
rect -5752 13988 -5732 14052
rect -5836 13972 -5732 13988
rect -5836 13908 -5816 13972
rect -5752 13908 -5732 13972
rect -5836 13892 -5732 13908
rect -5836 13828 -5816 13892
rect -5752 13828 -5732 13892
rect -5836 13812 -5732 13828
rect -5836 13748 -5816 13812
rect -5752 13748 -5732 13812
rect -5836 13732 -5732 13748
rect -5836 13668 -5816 13732
rect -5752 13668 -5732 13732
rect -5836 13652 -5732 13668
rect -5836 13588 -5816 13652
rect -5752 13588 -5732 13652
rect -5836 13572 -5732 13588
rect -5836 13508 -5816 13572
rect -5752 13508 -5732 13572
rect -5836 13492 -5732 13508
rect -5836 13428 -5816 13492
rect -5752 13428 -5732 13492
rect -5836 13412 -5732 13428
rect -5836 13348 -5816 13412
rect -5752 13348 -5732 13412
rect -5836 13332 -5732 13348
rect -5836 13268 -5816 13332
rect -5752 13268 -5732 13332
rect -5836 13252 -5732 13268
rect -5836 13188 -5816 13252
rect -5752 13188 -5732 13252
rect -5836 13172 -5732 13188
rect -5836 13108 -5816 13172
rect -5752 13108 -5732 13172
rect -5836 13092 -5732 13108
rect -5836 13028 -5816 13092
rect -5752 13028 -5732 13092
rect -5836 13012 -5732 13028
rect -5836 12948 -5816 13012
rect -5752 12948 -5732 13012
rect -5836 12932 -5732 12948
rect -5836 12868 -5816 12932
rect -5752 12868 -5732 12932
rect -5836 12852 -5732 12868
rect -5836 12788 -5816 12852
rect -5752 12788 -5732 12852
rect -5836 12772 -5732 12788
rect -5836 12708 -5816 12772
rect -5752 12708 -5732 12772
rect -5836 12692 -5732 12708
rect -5836 12628 -5816 12692
rect -5752 12628 -5732 12692
rect -5836 12612 -5732 12628
rect -5836 12548 -5816 12612
rect -5752 12548 -5732 12612
rect -5836 12532 -5732 12548
rect -5836 12468 -5816 12532
rect -5752 12468 -5732 12532
rect -5836 12452 -5732 12468
rect -5836 12388 -5816 12452
rect -5752 12388 -5732 12452
rect -5836 12372 -5732 12388
rect -5836 12308 -5816 12372
rect -5752 12308 -5732 12372
rect -5836 12292 -5732 12308
rect -5836 12228 -5816 12292
rect -5752 12228 -5732 12292
rect -5836 12212 -5732 12228
rect -5836 12148 -5816 12212
rect -5752 12148 -5732 12212
rect -5836 12132 -5732 12148
rect -5836 12068 -5816 12132
rect -5752 12068 -5732 12132
rect -5836 12052 -5732 12068
rect -5836 11988 -5816 12052
rect -5752 11988 -5732 12052
rect -5836 11972 -5732 11988
rect -5836 11908 -5816 11972
rect -5752 11908 -5732 11972
rect -5836 11892 -5732 11908
rect -5836 11828 -5816 11892
rect -5752 11828 -5732 11892
rect -5836 11812 -5732 11828
rect -5836 11748 -5816 11812
rect -5752 11748 -5732 11812
rect -5836 11732 -5732 11748
rect -5836 11668 -5816 11732
rect -5752 11668 -5732 11732
rect -5836 11652 -5732 11668
rect -5836 11588 -5816 11652
rect -5752 11588 -5732 11652
rect -5836 11572 -5732 11588
rect -5836 11508 -5816 11572
rect -5752 11508 -5732 11572
rect -5836 11492 -5732 11508
rect -5836 11428 -5816 11492
rect -5752 11428 -5732 11492
rect -5836 11412 -5732 11428
rect -5836 11348 -5816 11412
rect -5752 11348 -5732 11412
rect -5836 11332 -5732 11348
rect -5836 11268 -5816 11332
rect -5752 11268 -5732 11332
rect -5836 11252 -5732 11268
rect -5836 11188 -5816 11252
rect -5752 11188 -5732 11252
rect -5836 11172 -5732 11188
rect -5836 11108 -5816 11172
rect -5752 11108 -5732 11172
rect -5836 11092 -5732 11108
rect -5836 11028 -5816 11092
rect -5752 11028 -5732 11092
rect -5836 11012 -5732 11028
rect -5836 10948 -5816 11012
rect -5752 10948 -5732 11012
rect -5836 10932 -5732 10948
rect -5836 10868 -5816 10932
rect -5752 10868 -5732 10932
rect -5836 10852 -5732 10868
rect -11448 10492 -11344 10788
rect -17060 10412 -16956 10428
rect -17060 10348 -17040 10412
rect -16976 10348 -16956 10412
rect -17060 10332 -16956 10348
rect -17060 10268 -17040 10332
rect -16976 10268 -16956 10332
rect -17060 10252 -16956 10268
rect -17060 10188 -17040 10252
rect -16976 10188 -16956 10252
rect -17060 10172 -16956 10188
rect -17060 10108 -17040 10172
rect -16976 10108 -16956 10172
rect -17060 10092 -16956 10108
rect -17060 10028 -17040 10092
rect -16976 10028 -16956 10092
rect -17060 10012 -16956 10028
rect -17060 9948 -17040 10012
rect -16976 9948 -16956 10012
rect -17060 9932 -16956 9948
rect -17060 9868 -17040 9932
rect -16976 9868 -16956 9932
rect -17060 9852 -16956 9868
rect -17060 9788 -17040 9852
rect -16976 9788 -16956 9852
rect -17060 9772 -16956 9788
rect -17060 9708 -17040 9772
rect -16976 9708 -16956 9772
rect -17060 9692 -16956 9708
rect -17060 9628 -17040 9692
rect -16976 9628 -16956 9692
rect -17060 9612 -16956 9628
rect -17060 9548 -17040 9612
rect -16976 9548 -16956 9612
rect -17060 9532 -16956 9548
rect -17060 9468 -17040 9532
rect -16976 9468 -16956 9532
rect -17060 9452 -16956 9468
rect -17060 9388 -17040 9452
rect -16976 9388 -16956 9452
rect -17060 9372 -16956 9388
rect -17060 9308 -17040 9372
rect -16976 9308 -16956 9372
rect -17060 9292 -16956 9308
rect -17060 9228 -17040 9292
rect -16976 9228 -16956 9292
rect -17060 9212 -16956 9228
rect -17060 9148 -17040 9212
rect -16976 9148 -16956 9212
rect -17060 9132 -16956 9148
rect -17060 9068 -17040 9132
rect -16976 9068 -16956 9132
rect -17060 9052 -16956 9068
rect -17060 8988 -17040 9052
rect -16976 8988 -16956 9052
rect -17060 8972 -16956 8988
rect -17060 8908 -17040 8972
rect -16976 8908 -16956 8972
rect -17060 8892 -16956 8908
rect -17060 8828 -17040 8892
rect -16976 8828 -16956 8892
rect -17060 8812 -16956 8828
rect -17060 8748 -17040 8812
rect -16976 8748 -16956 8812
rect -17060 8732 -16956 8748
rect -17060 8668 -17040 8732
rect -16976 8668 -16956 8732
rect -17060 8652 -16956 8668
rect -17060 8588 -17040 8652
rect -16976 8588 -16956 8652
rect -17060 8572 -16956 8588
rect -17060 8508 -17040 8572
rect -16976 8508 -16956 8572
rect -17060 8492 -16956 8508
rect -17060 8428 -17040 8492
rect -16976 8428 -16956 8492
rect -17060 8412 -16956 8428
rect -17060 8348 -17040 8412
rect -16976 8348 -16956 8412
rect -17060 8332 -16956 8348
rect -17060 8268 -17040 8332
rect -16976 8268 -16956 8332
rect -17060 8252 -16956 8268
rect -17060 8188 -17040 8252
rect -16976 8188 -16956 8252
rect -17060 8172 -16956 8188
rect -17060 8108 -17040 8172
rect -16976 8108 -16956 8172
rect -17060 8092 -16956 8108
rect -17060 8028 -17040 8092
rect -16976 8028 -16956 8092
rect -17060 8012 -16956 8028
rect -17060 7948 -17040 8012
rect -16976 7948 -16956 8012
rect -17060 7932 -16956 7948
rect -17060 7868 -17040 7932
rect -16976 7868 -16956 7932
rect -17060 7852 -16956 7868
rect -17060 7788 -17040 7852
rect -16976 7788 -16956 7852
rect -17060 7772 -16956 7788
rect -17060 7708 -17040 7772
rect -16976 7708 -16956 7772
rect -17060 7692 -16956 7708
rect -17060 7628 -17040 7692
rect -16976 7628 -16956 7692
rect -17060 7612 -16956 7628
rect -17060 7548 -17040 7612
rect -16976 7548 -16956 7612
rect -17060 7532 -16956 7548
rect -17060 7468 -17040 7532
rect -16976 7468 -16956 7532
rect -17060 7452 -16956 7468
rect -17060 7388 -17040 7452
rect -16976 7388 -16956 7452
rect -17060 7372 -16956 7388
rect -17060 7308 -17040 7372
rect -16976 7308 -16956 7372
rect -17060 7292 -16956 7308
rect -17060 7228 -17040 7292
rect -16976 7228 -16956 7292
rect -17060 7212 -16956 7228
rect -17060 7148 -17040 7212
rect -16976 7148 -16956 7212
rect -17060 7132 -16956 7148
rect -17060 7068 -17040 7132
rect -16976 7068 -16956 7132
rect -17060 7052 -16956 7068
rect -17060 6988 -17040 7052
rect -16976 6988 -16956 7052
rect -17060 6972 -16956 6988
rect -17060 6908 -17040 6972
rect -16976 6908 -16956 6972
rect -17060 6892 -16956 6908
rect -17060 6828 -17040 6892
rect -16976 6828 -16956 6892
rect -17060 6812 -16956 6828
rect -17060 6748 -17040 6812
rect -16976 6748 -16956 6812
rect -17060 6732 -16956 6748
rect -17060 6668 -17040 6732
rect -16976 6668 -16956 6732
rect -17060 6652 -16956 6668
rect -17060 6588 -17040 6652
rect -16976 6588 -16956 6652
rect -17060 6572 -16956 6588
rect -17060 6508 -17040 6572
rect -16976 6508 -16956 6572
rect -17060 6492 -16956 6508
rect -17060 6428 -17040 6492
rect -16976 6428 -16956 6492
rect -17060 6412 -16956 6428
rect -17060 6348 -17040 6412
rect -16976 6348 -16956 6412
rect -17060 6332 -16956 6348
rect -17060 6268 -17040 6332
rect -16976 6268 -16956 6332
rect -17060 6252 -16956 6268
rect -17060 6188 -17040 6252
rect -16976 6188 -16956 6252
rect -17060 6172 -16956 6188
rect -17060 6108 -17040 6172
rect -16976 6108 -16956 6172
rect -17060 6092 -16956 6108
rect -17060 6028 -17040 6092
rect -16976 6028 -16956 6092
rect -17060 6012 -16956 6028
rect -17060 5948 -17040 6012
rect -16976 5948 -16956 6012
rect -17060 5932 -16956 5948
rect -17060 5868 -17040 5932
rect -16976 5868 -16956 5932
rect -17060 5852 -16956 5868
rect -17060 5788 -17040 5852
rect -16976 5788 -16956 5852
rect -17060 5772 -16956 5788
rect -17060 5708 -17040 5772
rect -16976 5708 -16956 5772
rect -17060 5692 -16956 5708
rect -17060 5628 -17040 5692
rect -16976 5628 -16956 5692
rect -17060 5612 -16956 5628
rect -17060 5548 -17040 5612
rect -16976 5548 -16956 5612
rect -17060 5532 -16956 5548
rect -22672 5172 -22568 5468
rect -28284 5092 -28180 5108
rect -28284 5028 -28264 5092
rect -28200 5028 -28180 5092
rect -28284 5012 -28180 5028
rect -28284 4948 -28264 5012
rect -28200 4948 -28180 5012
rect -28284 4932 -28180 4948
rect -28284 4868 -28264 4932
rect -28200 4868 -28180 4932
rect -28284 4852 -28180 4868
rect -28284 4788 -28264 4852
rect -28200 4788 -28180 4852
rect -28284 4772 -28180 4788
rect -28284 4708 -28264 4772
rect -28200 4708 -28180 4772
rect -28284 4692 -28180 4708
rect -28284 4628 -28264 4692
rect -28200 4628 -28180 4692
rect -28284 4612 -28180 4628
rect -28284 4548 -28264 4612
rect -28200 4548 -28180 4612
rect -28284 4532 -28180 4548
rect -28284 4468 -28264 4532
rect -28200 4468 -28180 4532
rect -28284 4452 -28180 4468
rect -28284 4388 -28264 4452
rect -28200 4388 -28180 4452
rect -28284 4372 -28180 4388
rect -28284 4308 -28264 4372
rect -28200 4308 -28180 4372
rect -28284 4292 -28180 4308
rect -28284 4228 -28264 4292
rect -28200 4228 -28180 4292
rect -28284 4212 -28180 4228
rect -28284 4148 -28264 4212
rect -28200 4148 -28180 4212
rect -28284 4132 -28180 4148
rect -28284 4068 -28264 4132
rect -28200 4068 -28180 4132
rect -28284 4052 -28180 4068
rect -28284 3988 -28264 4052
rect -28200 3988 -28180 4052
rect -28284 3972 -28180 3988
rect -28284 3908 -28264 3972
rect -28200 3908 -28180 3972
rect -28284 3892 -28180 3908
rect -28284 3828 -28264 3892
rect -28200 3828 -28180 3892
rect -28284 3812 -28180 3828
rect -28284 3748 -28264 3812
rect -28200 3748 -28180 3812
rect -28284 3732 -28180 3748
rect -28284 3668 -28264 3732
rect -28200 3668 -28180 3732
rect -28284 3652 -28180 3668
rect -28284 3588 -28264 3652
rect -28200 3588 -28180 3652
rect -28284 3572 -28180 3588
rect -28284 3508 -28264 3572
rect -28200 3508 -28180 3572
rect -28284 3492 -28180 3508
rect -28284 3428 -28264 3492
rect -28200 3428 -28180 3492
rect -28284 3412 -28180 3428
rect -28284 3348 -28264 3412
rect -28200 3348 -28180 3412
rect -28284 3332 -28180 3348
rect -28284 3268 -28264 3332
rect -28200 3268 -28180 3332
rect -28284 3252 -28180 3268
rect -28284 3188 -28264 3252
rect -28200 3188 -28180 3252
rect -28284 3172 -28180 3188
rect -28284 3108 -28264 3172
rect -28200 3108 -28180 3172
rect -28284 3092 -28180 3108
rect -28284 3028 -28264 3092
rect -28200 3028 -28180 3092
rect -28284 3012 -28180 3028
rect -28284 2948 -28264 3012
rect -28200 2948 -28180 3012
rect -28284 2932 -28180 2948
rect -28284 2868 -28264 2932
rect -28200 2868 -28180 2932
rect -28284 2852 -28180 2868
rect -28284 2788 -28264 2852
rect -28200 2788 -28180 2852
rect -28284 2772 -28180 2788
rect -28284 2708 -28264 2772
rect -28200 2708 -28180 2772
rect -28284 2692 -28180 2708
rect -28284 2628 -28264 2692
rect -28200 2628 -28180 2692
rect -28284 2612 -28180 2628
rect -28284 2548 -28264 2612
rect -28200 2548 -28180 2612
rect -28284 2532 -28180 2548
rect -28284 2468 -28264 2532
rect -28200 2468 -28180 2532
rect -28284 2452 -28180 2468
rect -28284 2388 -28264 2452
rect -28200 2388 -28180 2452
rect -28284 2372 -28180 2388
rect -28284 2308 -28264 2372
rect -28200 2308 -28180 2372
rect -28284 2292 -28180 2308
rect -28284 2228 -28264 2292
rect -28200 2228 -28180 2292
rect -28284 2212 -28180 2228
rect -28284 2148 -28264 2212
rect -28200 2148 -28180 2212
rect -28284 2132 -28180 2148
rect -28284 2068 -28264 2132
rect -28200 2068 -28180 2132
rect -28284 2052 -28180 2068
rect -28284 1988 -28264 2052
rect -28200 1988 -28180 2052
rect -28284 1972 -28180 1988
rect -28284 1908 -28264 1972
rect -28200 1908 -28180 1972
rect -28284 1892 -28180 1908
rect -28284 1828 -28264 1892
rect -28200 1828 -28180 1892
rect -28284 1812 -28180 1828
rect -28284 1748 -28264 1812
rect -28200 1748 -28180 1812
rect -28284 1732 -28180 1748
rect -28284 1668 -28264 1732
rect -28200 1668 -28180 1732
rect -28284 1652 -28180 1668
rect -28284 1588 -28264 1652
rect -28200 1588 -28180 1652
rect -28284 1572 -28180 1588
rect -28284 1508 -28264 1572
rect -28200 1508 -28180 1572
rect -28284 1492 -28180 1508
rect -28284 1428 -28264 1492
rect -28200 1428 -28180 1492
rect -28284 1412 -28180 1428
rect -28284 1348 -28264 1412
rect -28200 1348 -28180 1412
rect -28284 1332 -28180 1348
rect -28284 1268 -28264 1332
rect -28200 1268 -28180 1332
rect -28284 1252 -28180 1268
rect -28284 1188 -28264 1252
rect -28200 1188 -28180 1252
rect -28284 1172 -28180 1188
rect -28284 1108 -28264 1172
rect -28200 1108 -28180 1172
rect -28284 1092 -28180 1108
rect -28284 1028 -28264 1092
rect -28200 1028 -28180 1092
rect -28284 1012 -28180 1028
rect -28284 948 -28264 1012
rect -28200 948 -28180 1012
rect -28284 932 -28180 948
rect -28284 868 -28264 932
rect -28200 868 -28180 932
rect -28284 852 -28180 868
rect -28284 788 -28264 852
rect -28200 788 -28180 852
rect -28284 772 -28180 788
rect -28284 708 -28264 772
rect -28200 708 -28180 772
rect -28284 692 -28180 708
rect -28284 628 -28264 692
rect -28200 628 -28180 692
rect -28284 612 -28180 628
rect -28284 548 -28264 612
rect -28200 548 -28180 612
rect -28284 532 -28180 548
rect -28284 468 -28264 532
rect -28200 468 -28180 532
rect -28284 452 -28180 468
rect -28284 388 -28264 452
rect -28200 388 -28180 452
rect -28284 372 -28180 388
rect -28284 308 -28264 372
rect -28200 308 -28180 372
rect -28284 292 -28180 308
rect -28284 228 -28264 292
rect -28200 228 -28180 292
rect -28284 212 -28180 228
rect -33896 -148 -33792 148
rect -39085 -228 -34163 -199
rect -39085 -5092 -39056 -228
rect -34192 -5092 -34163 -228
rect -39085 -5121 -34163 -5092
rect -33896 -212 -33876 -148
rect -33812 -212 -33792 -148
rect -31064 -199 -30960 199
rect -28284 148 -28264 212
rect -28200 148 -28180 212
rect -27861 5092 -22939 5121
rect -27861 228 -27832 5092
rect -22968 228 -22939 5092
rect -27861 199 -22939 228
rect -22672 5108 -22652 5172
rect -22588 5108 -22568 5172
rect -19840 5121 -19736 5519
rect -17060 5468 -17040 5532
rect -16976 5468 -16956 5532
rect -16637 10412 -11715 10441
rect -16637 5548 -16608 10412
rect -11744 5548 -11715 10412
rect -16637 5519 -11715 5548
rect -11448 10428 -11428 10492
rect -11364 10428 -11344 10492
rect -8616 10441 -8512 10839
rect -5836 10788 -5816 10852
rect -5752 10788 -5732 10852
rect -5413 15732 -491 15761
rect -5413 10868 -5384 15732
rect -520 10868 -491 15732
rect -5413 10839 -491 10868
rect -224 15748 -204 15812
rect -140 15748 -120 15812
rect 2608 15761 2712 16159
rect 5388 16108 5408 16172
rect 5472 16108 5492 16172
rect 5811 21052 10733 21081
rect 5811 16188 5840 21052
rect 10704 16188 10733 21052
rect 5811 16159 10733 16188
rect 11000 21068 11020 21132
rect 11084 21068 11104 21132
rect 13832 21081 13936 21479
rect 16612 21428 16632 21492
rect 16696 21428 16716 21492
rect 17035 26372 21957 26401
rect 17035 21508 17064 26372
rect 21928 21508 21957 26372
rect 17035 21479 21957 21508
rect 22224 26388 22244 26452
rect 22308 26388 22328 26452
rect 25056 26401 25160 26799
rect 27836 26748 27856 26812
rect 27920 26748 27940 26812
rect 28259 31692 33181 31721
rect 28259 26828 28288 31692
rect 33152 26828 33181 31692
rect 28259 26799 33181 26828
rect 33448 31708 33468 31772
rect 33532 31708 33552 31772
rect 36280 31721 36384 32119
rect 39060 32068 39080 32132
rect 39144 32068 39164 32132
rect 39060 31772 39164 32068
rect 33448 31692 33552 31708
rect 33448 31628 33468 31692
rect 33532 31628 33552 31692
rect 33448 31612 33552 31628
rect 33448 31548 33468 31612
rect 33532 31548 33552 31612
rect 33448 31532 33552 31548
rect 33448 31468 33468 31532
rect 33532 31468 33552 31532
rect 33448 31452 33552 31468
rect 33448 31388 33468 31452
rect 33532 31388 33552 31452
rect 33448 31372 33552 31388
rect 33448 31308 33468 31372
rect 33532 31308 33552 31372
rect 33448 31292 33552 31308
rect 33448 31228 33468 31292
rect 33532 31228 33552 31292
rect 33448 31212 33552 31228
rect 33448 31148 33468 31212
rect 33532 31148 33552 31212
rect 33448 31132 33552 31148
rect 33448 31068 33468 31132
rect 33532 31068 33552 31132
rect 33448 31052 33552 31068
rect 33448 30988 33468 31052
rect 33532 30988 33552 31052
rect 33448 30972 33552 30988
rect 33448 30908 33468 30972
rect 33532 30908 33552 30972
rect 33448 30892 33552 30908
rect 33448 30828 33468 30892
rect 33532 30828 33552 30892
rect 33448 30812 33552 30828
rect 33448 30748 33468 30812
rect 33532 30748 33552 30812
rect 33448 30732 33552 30748
rect 33448 30668 33468 30732
rect 33532 30668 33552 30732
rect 33448 30652 33552 30668
rect 33448 30588 33468 30652
rect 33532 30588 33552 30652
rect 33448 30572 33552 30588
rect 33448 30508 33468 30572
rect 33532 30508 33552 30572
rect 33448 30492 33552 30508
rect 33448 30428 33468 30492
rect 33532 30428 33552 30492
rect 33448 30412 33552 30428
rect 33448 30348 33468 30412
rect 33532 30348 33552 30412
rect 33448 30332 33552 30348
rect 33448 30268 33468 30332
rect 33532 30268 33552 30332
rect 33448 30252 33552 30268
rect 33448 30188 33468 30252
rect 33532 30188 33552 30252
rect 33448 30172 33552 30188
rect 33448 30108 33468 30172
rect 33532 30108 33552 30172
rect 33448 30092 33552 30108
rect 33448 30028 33468 30092
rect 33532 30028 33552 30092
rect 33448 30012 33552 30028
rect 33448 29948 33468 30012
rect 33532 29948 33552 30012
rect 33448 29932 33552 29948
rect 33448 29868 33468 29932
rect 33532 29868 33552 29932
rect 33448 29852 33552 29868
rect 33448 29788 33468 29852
rect 33532 29788 33552 29852
rect 33448 29772 33552 29788
rect 33448 29708 33468 29772
rect 33532 29708 33552 29772
rect 33448 29692 33552 29708
rect 33448 29628 33468 29692
rect 33532 29628 33552 29692
rect 33448 29612 33552 29628
rect 33448 29548 33468 29612
rect 33532 29548 33552 29612
rect 33448 29532 33552 29548
rect 33448 29468 33468 29532
rect 33532 29468 33552 29532
rect 33448 29452 33552 29468
rect 33448 29388 33468 29452
rect 33532 29388 33552 29452
rect 33448 29372 33552 29388
rect 33448 29308 33468 29372
rect 33532 29308 33552 29372
rect 33448 29292 33552 29308
rect 33448 29228 33468 29292
rect 33532 29228 33552 29292
rect 33448 29212 33552 29228
rect 33448 29148 33468 29212
rect 33532 29148 33552 29212
rect 33448 29132 33552 29148
rect 33448 29068 33468 29132
rect 33532 29068 33552 29132
rect 33448 29052 33552 29068
rect 33448 28988 33468 29052
rect 33532 28988 33552 29052
rect 33448 28972 33552 28988
rect 33448 28908 33468 28972
rect 33532 28908 33552 28972
rect 33448 28892 33552 28908
rect 33448 28828 33468 28892
rect 33532 28828 33552 28892
rect 33448 28812 33552 28828
rect 33448 28748 33468 28812
rect 33532 28748 33552 28812
rect 33448 28732 33552 28748
rect 33448 28668 33468 28732
rect 33532 28668 33552 28732
rect 33448 28652 33552 28668
rect 33448 28588 33468 28652
rect 33532 28588 33552 28652
rect 33448 28572 33552 28588
rect 33448 28508 33468 28572
rect 33532 28508 33552 28572
rect 33448 28492 33552 28508
rect 33448 28428 33468 28492
rect 33532 28428 33552 28492
rect 33448 28412 33552 28428
rect 33448 28348 33468 28412
rect 33532 28348 33552 28412
rect 33448 28332 33552 28348
rect 33448 28268 33468 28332
rect 33532 28268 33552 28332
rect 33448 28252 33552 28268
rect 33448 28188 33468 28252
rect 33532 28188 33552 28252
rect 33448 28172 33552 28188
rect 33448 28108 33468 28172
rect 33532 28108 33552 28172
rect 33448 28092 33552 28108
rect 33448 28028 33468 28092
rect 33532 28028 33552 28092
rect 33448 28012 33552 28028
rect 33448 27948 33468 28012
rect 33532 27948 33552 28012
rect 33448 27932 33552 27948
rect 33448 27868 33468 27932
rect 33532 27868 33552 27932
rect 33448 27852 33552 27868
rect 33448 27788 33468 27852
rect 33532 27788 33552 27852
rect 33448 27772 33552 27788
rect 33448 27708 33468 27772
rect 33532 27708 33552 27772
rect 33448 27692 33552 27708
rect 33448 27628 33468 27692
rect 33532 27628 33552 27692
rect 33448 27612 33552 27628
rect 33448 27548 33468 27612
rect 33532 27548 33552 27612
rect 33448 27532 33552 27548
rect 33448 27468 33468 27532
rect 33532 27468 33552 27532
rect 33448 27452 33552 27468
rect 33448 27388 33468 27452
rect 33532 27388 33552 27452
rect 33448 27372 33552 27388
rect 33448 27308 33468 27372
rect 33532 27308 33552 27372
rect 33448 27292 33552 27308
rect 33448 27228 33468 27292
rect 33532 27228 33552 27292
rect 33448 27212 33552 27228
rect 33448 27148 33468 27212
rect 33532 27148 33552 27212
rect 33448 27132 33552 27148
rect 33448 27068 33468 27132
rect 33532 27068 33552 27132
rect 33448 27052 33552 27068
rect 33448 26988 33468 27052
rect 33532 26988 33552 27052
rect 33448 26972 33552 26988
rect 33448 26908 33468 26972
rect 33532 26908 33552 26972
rect 33448 26892 33552 26908
rect 33448 26828 33468 26892
rect 33532 26828 33552 26892
rect 33448 26812 33552 26828
rect 27836 26452 27940 26748
rect 22224 26372 22328 26388
rect 22224 26308 22244 26372
rect 22308 26308 22328 26372
rect 22224 26292 22328 26308
rect 22224 26228 22244 26292
rect 22308 26228 22328 26292
rect 22224 26212 22328 26228
rect 22224 26148 22244 26212
rect 22308 26148 22328 26212
rect 22224 26132 22328 26148
rect 22224 26068 22244 26132
rect 22308 26068 22328 26132
rect 22224 26052 22328 26068
rect 22224 25988 22244 26052
rect 22308 25988 22328 26052
rect 22224 25972 22328 25988
rect 22224 25908 22244 25972
rect 22308 25908 22328 25972
rect 22224 25892 22328 25908
rect 22224 25828 22244 25892
rect 22308 25828 22328 25892
rect 22224 25812 22328 25828
rect 22224 25748 22244 25812
rect 22308 25748 22328 25812
rect 22224 25732 22328 25748
rect 22224 25668 22244 25732
rect 22308 25668 22328 25732
rect 22224 25652 22328 25668
rect 22224 25588 22244 25652
rect 22308 25588 22328 25652
rect 22224 25572 22328 25588
rect 22224 25508 22244 25572
rect 22308 25508 22328 25572
rect 22224 25492 22328 25508
rect 22224 25428 22244 25492
rect 22308 25428 22328 25492
rect 22224 25412 22328 25428
rect 22224 25348 22244 25412
rect 22308 25348 22328 25412
rect 22224 25332 22328 25348
rect 22224 25268 22244 25332
rect 22308 25268 22328 25332
rect 22224 25252 22328 25268
rect 22224 25188 22244 25252
rect 22308 25188 22328 25252
rect 22224 25172 22328 25188
rect 22224 25108 22244 25172
rect 22308 25108 22328 25172
rect 22224 25092 22328 25108
rect 22224 25028 22244 25092
rect 22308 25028 22328 25092
rect 22224 25012 22328 25028
rect 22224 24948 22244 25012
rect 22308 24948 22328 25012
rect 22224 24932 22328 24948
rect 22224 24868 22244 24932
rect 22308 24868 22328 24932
rect 22224 24852 22328 24868
rect 22224 24788 22244 24852
rect 22308 24788 22328 24852
rect 22224 24772 22328 24788
rect 22224 24708 22244 24772
rect 22308 24708 22328 24772
rect 22224 24692 22328 24708
rect 22224 24628 22244 24692
rect 22308 24628 22328 24692
rect 22224 24612 22328 24628
rect 22224 24548 22244 24612
rect 22308 24548 22328 24612
rect 22224 24532 22328 24548
rect 22224 24468 22244 24532
rect 22308 24468 22328 24532
rect 22224 24452 22328 24468
rect 22224 24388 22244 24452
rect 22308 24388 22328 24452
rect 22224 24372 22328 24388
rect 22224 24308 22244 24372
rect 22308 24308 22328 24372
rect 22224 24292 22328 24308
rect 22224 24228 22244 24292
rect 22308 24228 22328 24292
rect 22224 24212 22328 24228
rect 22224 24148 22244 24212
rect 22308 24148 22328 24212
rect 22224 24132 22328 24148
rect 22224 24068 22244 24132
rect 22308 24068 22328 24132
rect 22224 24052 22328 24068
rect 22224 23988 22244 24052
rect 22308 23988 22328 24052
rect 22224 23972 22328 23988
rect 22224 23908 22244 23972
rect 22308 23908 22328 23972
rect 22224 23892 22328 23908
rect 22224 23828 22244 23892
rect 22308 23828 22328 23892
rect 22224 23812 22328 23828
rect 22224 23748 22244 23812
rect 22308 23748 22328 23812
rect 22224 23732 22328 23748
rect 22224 23668 22244 23732
rect 22308 23668 22328 23732
rect 22224 23652 22328 23668
rect 22224 23588 22244 23652
rect 22308 23588 22328 23652
rect 22224 23572 22328 23588
rect 22224 23508 22244 23572
rect 22308 23508 22328 23572
rect 22224 23492 22328 23508
rect 22224 23428 22244 23492
rect 22308 23428 22328 23492
rect 22224 23412 22328 23428
rect 22224 23348 22244 23412
rect 22308 23348 22328 23412
rect 22224 23332 22328 23348
rect 22224 23268 22244 23332
rect 22308 23268 22328 23332
rect 22224 23252 22328 23268
rect 22224 23188 22244 23252
rect 22308 23188 22328 23252
rect 22224 23172 22328 23188
rect 22224 23108 22244 23172
rect 22308 23108 22328 23172
rect 22224 23092 22328 23108
rect 22224 23028 22244 23092
rect 22308 23028 22328 23092
rect 22224 23012 22328 23028
rect 22224 22948 22244 23012
rect 22308 22948 22328 23012
rect 22224 22932 22328 22948
rect 22224 22868 22244 22932
rect 22308 22868 22328 22932
rect 22224 22852 22328 22868
rect 22224 22788 22244 22852
rect 22308 22788 22328 22852
rect 22224 22772 22328 22788
rect 22224 22708 22244 22772
rect 22308 22708 22328 22772
rect 22224 22692 22328 22708
rect 22224 22628 22244 22692
rect 22308 22628 22328 22692
rect 22224 22612 22328 22628
rect 22224 22548 22244 22612
rect 22308 22548 22328 22612
rect 22224 22532 22328 22548
rect 22224 22468 22244 22532
rect 22308 22468 22328 22532
rect 22224 22452 22328 22468
rect 22224 22388 22244 22452
rect 22308 22388 22328 22452
rect 22224 22372 22328 22388
rect 22224 22308 22244 22372
rect 22308 22308 22328 22372
rect 22224 22292 22328 22308
rect 22224 22228 22244 22292
rect 22308 22228 22328 22292
rect 22224 22212 22328 22228
rect 22224 22148 22244 22212
rect 22308 22148 22328 22212
rect 22224 22132 22328 22148
rect 22224 22068 22244 22132
rect 22308 22068 22328 22132
rect 22224 22052 22328 22068
rect 22224 21988 22244 22052
rect 22308 21988 22328 22052
rect 22224 21972 22328 21988
rect 22224 21908 22244 21972
rect 22308 21908 22328 21972
rect 22224 21892 22328 21908
rect 22224 21828 22244 21892
rect 22308 21828 22328 21892
rect 22224 21812 22328 21828
rect 22224 21748 22244 21812
rect 22308 21748 22328 21812
rect 22224 21732 22328 21748
rect 22224 21668 22244 21732
rect 22308 21668 22328 21732
rect 22224 21652 22328 21668
rect 22224 21588 22244 21652
rect 22308 21588 22328 21652
rect 22224 21572 22328 21588
rect 22224 21508 22244 21572
rect 22308 21508 22328 21572
rect 22224 21492 22328 21508
rect 16612 21132 16716 21428
rect 11000 21052 11104 21068
rect 11000 20988 11020 21052
rect 11084 20988 11104 21052
rect 11000 20972 11104 20988
rect 11000 20908 11020 20972
rect 11084 20908 11104 20972
rect 11000 20892 11104 20908
rect 11000 20828 11020 20892
rect 11084 20828 11104 20892
rect 11000 20812 11104 20828
rect 11000 20748 11020 20812
rect 11084 20748 11104 20812
rect 11000 20732 11104 20748
rect 11000 20668 11020 20732
rect 11084 20668 11104 20732
rect 11000 20652 11104 20668
rect 11000 20588 11020 20652
rect 11084 20588 11104 20652
rect 11000 20572 11104 20588
rect 11000 20508 11020 20572
rect 11084 20508 11104 20572
rect 11000 20492 11104 20508
rect 11000 20428 11020 20492
rect 11084 20428 11104 20492
rect 11000 20412 11104 20428
rect 11000 20348 11020 20412
rect 11084 20348 11104 20412
rect 11000 20332 11104 20348
rect 11000 20268 11020 20332
rect 11084 20268 11104 20332
rect 11000 20252 11104 20268
rect 11000 20188 11020 20252
rect 11084 20188 11104 20252
rect 11000 20172 11104 20188
rect 11000 20108 11020 20172
rect 11084 20108 11104 20172
rect 11000 20092 11104 20108
rect 11000 20028 11020 20092
rect 11084 20028 11104 20092
rect 11000 20012 11104 20028
rect 11000 19948 11020 20012
rect 11084 19948 11104 20012
rect 11000 19932 11104 19948
rect 11000 19868 11020 19932
rect 11084 19868 11104 19932
rect 11000 19852 11104 19868
rect 11000 19788 11020 19852
rect 11084 19788 11104 19852
rect 11000 19772 11104 19788
rect 11000 19708 11020 19772
rect 11084 19708 11104 19772
rect 11000 19692 11104 19708
rect 11000 19628 11020 19692
rect 11084 19628 11104 19692
rect 11000 19612 11104 19628
rect 11000 19548 11020 19612
rect 11084 19548 11104 19612
rect 11000 19532 11104 19548
rect 11000 19468 11020 19532
rect 11084 19468 11104 19532
rect 11000 19452 11104 19468
rect 11000 19388 11020 19452
rect 11084 19388 11104 19452
rect 11000 19372 11104 19388
rect 11000 19308 11020 19372
rect 11084 19308 11104 19372
rect 11000 19292 11104 19308
rect 11000 19228 11020 19292
rect 11084 19228 11104 19292
rect 11000 19212 11104 19228
rect 11000 19148 11020 19212
rect 11084 19148 11104 19212
rect 11000 19132 11104 19148
rect 11000 19068 11020 19132
rect 11084 19068 11104 19132
rect 11000 19052 11104 19068
rect 11000 18988 11020 19052
rect 11084 18988 11104 19052
rect 11000 18972 11104 18988
rect 11000 18908 11020 18972
rect 11084 18908 11104 18972
rect 11000 18892 11104 18908
rect 11000 18828 11020 18892
rect 11084 18828 11104 18892
rect 11000 18812 11104 18828
rect 11000 18748 11020 18812
rect 11084 18748 11104 18812
rect 11000 18732 11104 18748
rect 11000 18668 11020 18732
rect 11084 18668 11104 18732
rect 11000 18652 11104 18668
rect 11000 18588 11020 18652
rect 11084 18588 11104 18652
rect 11000 18572 11104 18588
rect 11000 18508 11020 18572
rect 11084 18508 11104 18572
rect 11000 18492 11104 18508
rect 11000 18428 11020 18492
rect 11084 18428 11104 18492
rect 11000 18412 11104 18428
rect 11000 18348 11020 18412
rect 11084 18348 11104 18412
rect 11000 18332 11104 18348
rect 11000 18268 11020 18332
rect 11084 18268 11104 18332
rect 11000 18252 11104 18268
rect 11000 18188 11020 18252
rect 11084 18188 11104 18252
rect 11000 18172 11104 18188
rect 11000 18108 11020 18172
rect 11084 18108 11104 18172
rect 11000 18092 11104 18108
rect 11000 18028 11020 18092
rect 11084 18028 11104 18092
rect 11000 18012 11104 18028
rect 11000 17948 11020 18012
rect 11084 17948 11104 18012
rect 11000 17932 11104 17948
rect 11000 17868 11020 17932
rect 11084 17868 11104 17932
rect 11000 17852 11104 17868
rect 11000 17788 11020 17852
rect 11084 17788 11104 17852
rect 11000 17772 11104 17788
rect 11000 17708 11020 17772
rect 11084 17708 11104 17772
rect 11000 17692 11104 17708
rect 11000 17628 11020 17692
rect 11084 17628 11104 17692
rect 11000 17612 11104 17628
rect 11000 17548 11020 17612
rect 11084 17548 11104 17612
rect 11000 17532 11104 17548
rect 11000 17468 11020 17532
rect 11084 17468 11104 17532
rect 11000 17452 11104 17468
rect 11000 17388 11020 17452
rect 11084 17388 11104 17452
rect 11000 17372 11104 17388
rect 11000 17308 11020 17372
rect 11084 17308 11104 17372
rect 11000 17292 11104 17308
rect 11000 17228 11020 17292
rect 11084 17228 11104 17292
rect 11000 17212 11104 17228
rect 11000 17148 11020 17212
rect 11084 17148 11104 17212
rect 11000 17132 11104 17148
rect 11000 17068 11020 17132
rect 11084 17068 11104 17132
rect 11000 17052 11104 17068
rect 11000 16988 11020 17052
rect 11084 16988 11104 17052
rect 11000 16972 11104 16988
rect 11000 16908 11020 16972
rect 11084 16908 11104 16972
rect 11000 16892 11104 16908
rect 11000 16828 11020 16892
rect 11084 16828 11104 16892
rect 11000 16812 11104 16828
rect 11000 16748 11020 16812
rect 11084 16748 11104 16812
rect 11000 16732 11104 16748
rect 11000 16668 11020 16732
rect 11084 16668 11104 16732
rect 11000 16652 11104 16668
rect 11000 16588 11020 16652
rect 11084 16588 11104 16652
rect 11000 16572 11104 16588
rect 11000 16508 11020 16572
rect 11084 16508 11104 16572
rect 11000 16492 11104 16508
rect 11000 16428 11020 16492
rect 11084 16428 11104 16492
rect 11000 16412 11104 16428
rect 11000 16348 11020 16412
rect 11084 16348 11104 16412
rect 11000 16332 11104 16348
rect 11000 16268 11020 16332
rect 11084 16268 11104 16332
rect 11000 16252 11104 16268
rect 11000 16188 11020 16252
rect 11084 16188 11104 16252
rect 11000 16172 11104 16188
rect 5388 15812 5492 16108
rect -224 15732 -120 15748
rect -224 15668 -204 15732
rect -140 15668 -120 15732
rect -224 15652 -120 15668
rect -224 15588 -204 15652
rect -140 15588 -120 15652
rect -224 15572 -120 15588
rect -224 15508 -204 15572
rect -140 15508 -120 15572
rect -224 15492 -120 15508
rect -224 15428 -204 15492
rect -140 15428 -120 15492
rect -224 15412 -120 15428
rect -224 15348 -204 15412
rect -140 15348 -120 15412
rect -224 15332 -120 15348
rect -224 15268 -204 15332
rect -140 15268 -120 15332
rect -224 15252 -120 15268
rect -224 15188 -204 15252
rect -140 15188 -120 15252
rect -224 15172 -120 15188
rect -224 15108 -204 15172
rect -140 15108 -120 15172
rect -224 15092 -120 15108
rect -224 15028 -204 15092
rect -140 15028 -120 15092
rect -224 15012 -120 15028
rect -224 14948 -204 15012
rect -140 14948 -120 15012
rect -224 14932 -120 14948
rect -224 14868 -204 14932
rect -140 14868 -120 14932
rect -224 14852 -120 14868
rect -224 14788 -204 14852
rect -140 14788 -120 14852
rect -224 14772 -120 14788
rect -224 14708 -204 14772
rect -140 14708 -120 14772
rect -224 14692 -120 14708
rect -224 14628 -204 14692
rect -140 14628 -120 14692
rect -224 14612 -120 14628
rect -224 14548 -204 14612
rect -140 14548 -120 14612
rect -224 14532 -120 14548
rect -224 14468 -204 14532
rect -140 14468 -120 14532
rect -224 14452 -120 14468
rect -224 14388 -204 14452
rect -140 14388 -120 14452
rect -224 14372 -120 14388
rect -224 14308 -204 14372
rect -140 14308 -120 14372
rect -224 14292 -120 14308
rect -224 14228 -204 14292
rect -140 14228 -120 14292
rect -224 14212 -120 14228
rect -224 14148 -204 14212
rect -140 14148 -120 14212
rect -224 14132 -120 14148
rect -224 14068 -204 14132
rect -140 14068 -120 14132
rect -224 14052 -120 14068
rect -224 13988 -204 14052
rect -140 13988 -120 14052
rect -224 13972 -120 13988
rect -224 13908 -204 13972
rect -140 13908 -120 13972
rect -224 13892 -120 13908
rect -224 13828 -204 13892
rect -140 13828 -120 13892
rect -224 13812 -120 13828
rect -224 13748 -204 13812
rect -140 13748 -120 13812
rect -224 13732 -120 13748
rect -224 13668 -204 13732
rect -140 13668 -120 13732
rect -224 13652 -120 13668
rect -224 13588 -204 13652
rect -140 13588 -120 13652
rect -224 13572 -120 13588
rect -224 13508 -204 13572
rect -140 13508 -120 13572
rect -224 13492 -120 13508
rect -224 13428 -204 13492
rect -140 13428 -120 13492
rect -224 13412 -120 13428
rect -224 13348 -204 13412
rect -140 13348 -120 13412
rect -224 13332 -120 13348
rect -224 13268 -204 13332
rect -140 13268 -120 13332
rect -224 13252 -120 13268
rect -224 13188 -204 13252
rect -140 13188 -120 13252
rect -224 13172 -120 13188
rect -224 13108 -204 13172
rect -140 13108 -120 13172
rect -224 13092 -120 13108
rect -224 13028 -204 13092
rect -140 13028 -120 13092
rect -224 13012 -120 13028
rect -224 12948 -204 13012
rect -140 12948 -120 13012
rect -224 12932 -120 12948
rect -224 12868 -204 12932
rect -140 12868 -120 12932
rect -224 12852 -120 12868
rect -224 12788 -204 12852
rect -140 12788 -120 12852
rect -224 12772 -120 12788
rect -224 12708 -204 12772
rect -140 12708 -120 12772
rect -224 12692 -120 12708
rect -224 12628 -204 12692
rect -140 12628 -120 12692
rect -224 12612 -120 12628
rect -224 12548 -204 12612
rect -140 12548 -120 12612
rect -224 12532 -120 12548
rect -224 12468 -204 12532
rect -140 12468 -120 12532
rect -224 12452 -120 12468
rect -224 12388 -204 12452
rect -140 12388 -120 12452
rect -224 12372 -120 12388
rect -224 12308 -204 12372
rect -140 12308 -120 12372
rect -224 12292 -120 12308
rect -224 12228 -204 12292
rect -140 12228 -120 12292
rect -224 12212 -120 12228
rect -224 12148 -204 12212
rect -140 12148 -120 12212
rect -224 12132 -120 12148
rect -224 12068 -204 12132
rect -140 12068 -120 12132
rect -224 12052 -120 12068
rect -224 11988 -204 12052
rect -140 11988 -120 12052
rect -224 11972 -120 11988
rect -224 11908 -204 11972
rect -140 11908 -120 11972
rect -224 11892 -120 11908
rect -224 11828 -204 11892
rect -140 11828 -120 11892
rect -224 11812 -120 11828
rect -224 11748 -204 11812
rect -140 11748 -120 11812
rect -224 11732 -120 11748
rect -224 11668 -204 11732
rect -140 11668 -120 11732
rect -224 11652 -120 11668
rect -224 11588 -204 11652
rect -140 11588 -120 11652
rect -224 11572 -120 11588
rect -224 11508 -204 11572
rect -140 11508 -120 11572
rect -224 11492 -120 11508
rect -224 11428 -204 11492
rect -140 11428 -120 11492
rect -224 11412 -120 11428
rect -224 11348 -204 11412
rect -140 11348 -120 11412
rect -224 11332 -120 11348
rect -224 11268 -204 11332
rect -140 11268 -120 11332
rect -224 11252 -120 11268
rect -224 11188 -204 11252
rect -140 11188 -120 11252
rect -224 11172 -120 11188
rect -224 11108 -204 11172
rect -140 11108 -120 11172
rect -224 11092 -120 11108
rect -224 11028 -204 11092
rect -140 11028 -120 11092
rect -224 11012 -120 11028
rect -224 10948 -204 11012
rect -140 10948 -120 11012
rect -224 10932 -120 10948
rect -224 10868 -204 10932
rect -140 10868 -120 10932
rect -224 10852 -120 10868
rect -5836 10492 -5732 10788
rect -11448 10412 -11344 10428
rect -11448 10348 -11428 10412
rect -11364 10348 -11344 10412
rect -11448 10332 -11344 10348
rect -11448 10268 -11428 10332
rect -11364 10268 -11344 10332
rect -11448 10252 -11344 10268
rect -11448 10188 -11428 10252
rect -11364 10188 -11344 10252
rect -11448 10172 -11344 10188
rect -11448 10108 -11428 10172
rect -11364 10108 -11344 10172
rect -11448 10092 -11344 10108
rect -11448 10028 -11428 10092
rect -11364 10028 -11344 10092
rect -11448 10012 -11344 10028
rect -11448 9948 -11428 10012
rect -11364 9948 -11344 10012
rect -11448 9932 -11344 9948
rect -11448 9868 -11428 9932
rect -11364 9868 -11344 9932
rect -11448 9852 -11344 9868
rect -11448 9788 -11428 9852
rect -11364 9788 -11344 9852
rect -11448 9772 -11344 9788
rect -11448 9708 -11428 9772
rect -11364 9708 -11344 9772
rect -11448 9692 -11344 9708
rect -11448 9628 -11428 9692
rect -11364 9628 -11344 9692
rect -11448 9612 -11344 9628
rect -11448 9548 -11428 9612
rect -11364 9548 -11344 9612
rect -11448 9532 -11344 9548
rect -11448 9468 -11428 9532
rect -11364 9468 -11344 9532
rect -11448 9452 -11344 9468
rect -11448 9388 -11428 9452
rect -11364 9388 -11344 9452
rect -11448 9372 -11344 9388
rect -11448 9308 -11428 9372
rect -11364 9308 -11344 9372
rect -11448 9292 -11344 9308
rect -11448 9228 -11428 9292
rect -11364 9228 -11344 9292
rect -11448 9212 -11344 9228
rect -11448 9148 -11428 9212
rect -11364 9148 -11344 9212
rect -11448 9132 -11344 9148
rect -11448 9068 -11428 9132
rect -11364 9068 -11344 9132
rect -11448 9052 -11344 9068
rect -11448 8988 -11428 9052
rect -11364 8988 -11344 9052
rect -11448 8972 -11344 8988
rect -11448 8908 -11428 8972
rect -11364 8908 -11344 8972
rect -11448 8892 -11344 8908
rect -11448 8828 -11428 8892
rect -11364 8828 -11344 8892
rect -11448 8812 -11344 8828
rect -11448 8748 -11428 8812
rect -11364 8748 -11344 8812
rect -11448 8732 -11344 8748
rect -11448 8668 -11428 8732
rect -11364 8668 -11344 8732
rect -11448 8652 -11344 8668
rect -11448 8588 -11428 8652
rect -11364 8588 -11344 8652
rect -11448 8572 -11344 8588
rect -11448 8508 -11428 8572
rect -11364 8508 -11344 8572
rect -11448 8492 -11344 8508
rect -11448 8428 -11428 8492
rect -11364 8428 -11344 8492
rect -11448 8412 -11344 8428
rect -11448 8348 -11428 8412
rect -11364 8348 -11344 8412
rect -11448 8332 -11344 8348
rect -11448 8268 -11428 8332
rect -11364 8268 -11344 8332
rect -11448 8252 -11344 8268
rect -11448 8188 -11428 8252
rect -11364 8188 -11344 8252
rect -11448 8172 -11344 8188
rect -11448 8108 -11428 8172
rect -11364 8108 -11344 8172
rect -11448 8092 -11344 8108
rect -11448 8028 -11428 8092
rect -11364 8028 -11344 8092
rect -11448 8012 -11344 8028
rect -11448 7948 -11428 8012
rect -11364 7948 -11344 8012
rect -11448 7932 -11344 7948
rect -11448 7868 -11428 7932
rect -11364 7868 -11344 7932
rect -11448 7852 -11344 7868
rect -11448 7788 -11428 7852
rect -11364 7788 -11344 7852
rect -11448 7772 -11344 7788
rect -11448 7708 -11428 7772
rect -11364 7708 -11344 7772
rect -11448 7692 -11344 7708
rect -11448 7628 -11428 7692
rect -11364 7628 -11344 7692
rect -11448 7612 -11344 7628
rect -11448 7548 -11428 7612
rect -11364 7548 -11344 7612
rect -11448 7532 -11344 7548
rect -11448 7468 -11428 7532
rect -11364 7468 -11344 7532
rect -11448 7452 -11344 7468
rect -11448 7388 -11428 7452
rect -11364 7388 -11344 7452
rect -11448 7372 -11344 7388
rect -11448 7308 -11428 7372
rect -11364 7308 -11344 7372
rect -11448 7292 -11344 7308
rect -11448 7228 -11428 7292
rect -11364 7228 -11344 7292
rect -11448 7212 -11344 7228
rect -11448 7148 -11428 7212
rect -11364 7148 -11344 7212
rect -11448 7132 -11344 7148
rect -11448 7068 -11428 7132
rect -11364 7068 -11344 7132
rect -11448 7052 -11344 7068
rect -11448 6988 -11428 7052
rect -11364 6988 -11344 7052
rect -11448 6972 -11344 6988
rect -11448 6908 -11428 6972
rect -11364 6908 -11344 6972
rect -11448 6892 -11344 6908
rect -11448 6828 -11428 6892
rect -11364 6828 -11344 6892
rect -11448 6812 -11344 6828
rect -11448 6748 -11428 6812
rect -11364 6748 -11344 6812
rect -11448 6732 -11344 6748
rect -11448 6668 -11428 6732
rect -11364 6668 -11344 6732
rect -11448 6652 -11344 6668
rect -11448 6588 -11428 6652
rect -11364 6588 -11344 6652
rect -11448 6572 -11344 6588
rect -11448 6508 -11428 6572
rect -11364 6508 -11344 6572
rect -11448 6492 -11344 6508
rect -11448 6428 -11428 6492
rect -11364 6428 -11344 6492
rect -11448 6412 -11344 6428
rect -11448 6348 -11428 6412
rect -11364 6348 -11344 6412
rect -11448 6332 -11344 6348
rect -11448 6268 -11428 6332
rect -11364 6268 -11344 6332
rect -11448 6252 -11344 6268
rect -11448 6188 -11428 6252
rect -11364 6188 -11344 6252
rect -11448 6172 -11344 6188
rect -11448 6108 -11428 6172
rect -11364 6108 -11344 6172
rect -11448 6092 -11344 6108
rect -11448 6028 -11428 6092
rect -11364 6028 -11344 6092
rect -11448 6012 -11344 6028
rect -11448 5948 -11428 6012
rect -11364 5948 -11344 6012
rect -11448 5932 -11344 5948
rect -11448 5868 -11428 5932
rect -11364 5868 -11344 5932
rect -11448 5852 -11344 5868
rect -11448 5788 -11428 5852
rect -11364 5788 -11344 5852
rect -11448 5772 -11344 5788
rect -11448 5708 -11428 5772
rect -11364 5708 -11344 5772
rect -11448 5692 -11344 5708
rect -11448 5628 -11428 5692
rect -11364 5628 -11344 5692
rect -11448 5612 -11344 5628
rect -11448 5548 -11428 5612
rect -11364 5548 -11344 5612
rect -11448 5532 -11344 5548
rect -17060 5172 -16956 5468
rect -22672 5092 -22568 5108
rect -22672 5028 -22652 5092
rect -22588 5028 -22568 5092
rect -22672 5012 -22568 5028
rect -22672 4948 -22652 5012
rect -22588 4948 -22568 5012
rect -22672 4932 -22568 4948
rect -22672 4868 -22652 4932
rect -22588 4868 -22568 4932
rect -22672 4852 -22568 4868
rect -22672 4788 -22652 4852
rect -22588 4788 -22568 4852
rect -22672 4772 -22568 4788
rect -22672 4708 -22652 4772
rect -22588 4708 -22568 4772
rect -22672 4692 -22568 4708
rect -22672 4628 -22652 4692
rect -22588 4628 -22568 4692
rect -22672 4612 -22568 4628
rect -22672 4548 -22652 4612
rect -22588 4548 -22568 4612
rect -22672 4532 -22568 4548
rect -22672 4468 -22652 4532
rect -22588 4468 -22568 4532
rect -22672 4452 -22568 4468
rect -22672 4388 -22652 4452
rect -22588 4388 -22568 4452
rect -22672 4372 -22568 4388
rect -22672 4308 -22652 4372
rect -22588 4308 -22568 4372
rect -22672 4292 -22568 4308
rect -22672 4228 -22652 4292
rect -22588 4228 -22568 4292
rect -22672 4212 -22568 4228
rect -22672 4148 -22652 4212
rect -22588 4148 -22568 4212
rect -22672 4132 -22568 4148
rect -22672 4068 -22652 4132
rect -22588 4068 -22568 4132
rect -22672 4052 -22568 4068
rect -22672 3988 -22652 4052
rect -22588 3988 -22568 4052
rect -22672 3972 -22568 3988
rect -22672 3908 -22652 3972
rect -22588 3908 -22568 3972
rect -22672 3892 -22568 3908
rect -22672 3828 -22652 3892
rect -22588 3828 -22568 3892
rect -22672 3812 -22568 3828
rect -22672 3748 -22652 3812
rect -22588 3748 -22568 3812
rect -22672 3732 -22568 3748
rect -22672 3668 -22652 3732
rect -22588 3668 -22568 3732
rect -22672 3652 -22568 3668
rect -22672 3588 -22652 3652
rect -22588 3588 -22568 3652
rect -22672 3572 -22568 3588
rect -22672 3508 -22652 3572
rect -22588 3508 -22568 3572
rect -22672 3492 -22568 3508
rect -22672 3428 -22652 3492
rect -22588 3428 -22568 3492
rect -22672 3412 -22568 3428
rect -22672 3348 -22652 3412
rect -22588 3348 -22568 3412
rect -22672 3332 -22568 3348
rect -22672 3268 -22652 3332
rect -22588 3268 -22568 3332
rect -22672 3252 -22568 3268
rect -22672 3188 -22652 3252
rect -22588 3188 -22568 3252
rect -22672 3172 -22568 3188
rect -22672 3108 -22652 3172
rect -22588 3108 -22568 3172
rect -22672 3092 -22568 3108
rect -22672 3028 -22652 3092
rect -22588 3028 -22568 3092
rect -22672 3012 -22568 3028
rect -22672 2948 -22652 3012
rect -22588 2948 -22568 3012
rect -22672 2932 -22568 2948
rect -22672 2868 -22652 2932
rect -22588 2868 -22568 2932
rect -22672 2852 -22568 2868
rect -22672 2788 -22652 2852
rect -22588 2788 -22568 2852
rect -22672 2772 -22568 2788
rect -22672 2708 -22652 2772
rect -22588 2708 -22568 2772
rect -22672 2692 -22568 2708
rect -22672 2628 -22652 2692
rect -22588 2628 -22568 2692
rect -22672 2612 -22568 2628
rect -22672 2548 -22652 2612
rect -22588 2548 -22568 2612
rect -22672 2532 -22568 2548
rect -22672 2468 -22652 2532
rect -22588 2468 -22568 2532
rect -22672 2452 -22568 2468
rect -22672 2388 -22652 2452
rect -22588 2388 -22568 2452
rect -22672 2372 -22568 2388
rect -22672 2308 -22652 2372
rect -22588 2308 -22568 2372
rect -22672 2292 -22568 2308
rect -22672 2228 -22652 2292
rect -22588 2228 -22568 2292
rect -22672 2212 -22568 2228
rect -22672 2148 -22652 2212
rect -22588 2148 -22568 2212
rect -22672 2132 -22568 2148
rect -22672 2068 -22652 2132
rect -22588 2068 -22568 2132
rect -22672 2052 -22568 2068
rect -22672 1988 -22652 2052
rect -22588 1988 -22568 2052
rect -22672 1972 -22568 1988
rect -22672 1908 -22652 1972
rect -22588 1908 -22568 1972
rect -22672 1892 -22568 1908
rect -22672 1828 -22652 1892
rect -22588 1828 -22568 1892
rect -22672 1812 -22568 1828
rect -22672 1748 -22652 1812
rect -22588 1748 -22568 1812
rect -22672 1732 -22568 1748
rect -22672 1668 -22652 1732
rect -22588 1668 -22568 1732
rect -22672 1652 -22568 1668
rect -22672 1588 -22652 1652
rect -22588 1588 -22568 1652
rect -22672 1572 -22568 1588
rect -22672 1508 -22652 1572
rect -22588 1508 -22568 1572
rect -22672 1492 -22568 1508
rect -22672 1428 -22652 1492
rect -22588 1428 -22568 1492
rect -22672 1412 -22568 1428
rect -22672 1348 -22652 1412
rect -22588 1348 -22568 1412
rect -22672 1332 -22568 1348
rect -22672 1268 -22652 1332
rect -22588 1268 -22568 1332
rect -22672 1252 -22568 1268
rect -22672 1188 -22652 1252
rect -22588 1188 -22568 1252
rect -22672 1172 -22568 1188
rect -22672 1108 -22652 1172
rect -22588 1108 -22568 1172
rect -22672 1092 -22568 1108
rect -22672 1028 -22652 1092
rect -22588 1028 -22568 1092
rect -22672 1012 -22568 1028
rect -22672 948 -22652 1012
rect -22588 948 -22568 1012
rect -22672 932 -22568 948
rect -22672 868 -22652 932
rect -22588 868 -22568 932
rect -22672 852 -22568 868
rect -22672 788 -22652 852
rect -22588 788 -22568 852
rect -22672 772 -22568 788
rect -22672 708 -22652 772
rect -22588 708 -22568 772
rect -22672 692 -22568 708
rect -22672 628 -22652 692
rect -22588 628 -22568 692
rect -22672 612 -22568 628
rect -22672 548 -22652 612
rect -22588 548 -22568 612
rect -22672 532 -22568 548
rect -22672 468 -22652 532
rect -22588 468 -22568 532
rect -22672 452 -22568 468
rect -22672 388 -22652 452
rect -22588 388 -22568 452
rect -22672 372 -22568 388
rect -22672 308 -22652 372
rect -22588 308 -22568 372
rect -22672 292 -22568 308
rect -22672 228 -22652 292
rect -22588 228 -22568 292
rect -22672 212 -22568 228
rect -28284 -148 -28180 148
rect -33896 -228 -33792 -212
rect -33896 -292 -33876 -228
rect -33812 -292 -33792 -228
rect -33896 -308 -33792 -292
rect -33896 -372 -33876 -308
rect -33812 -372 -33792 -308
rect -33896 -388 -33792 -372
rect -33896 -452 -33876 -388
rect -33812 -452 -33792 -388
rect -33896 -468 -33792 -452
rect -33896 -532 -33876 -468
rect -33812 -532 -33792 -468
rect -33896 -548 -33792 -532
rect -33896 -612 -33876 -548
rect -33812 -612 -33792 -548
rect -33896 -628 -33792 -612
rect -33896 -692 -33876 -628
rect -33812 -692 -33792 -628
rect -33896 -708 -33792 -692
rect -33896 -772 -33876 -708
rect -33812 -772 -33792 -708
rect -33896 -788 -33792 -772
rect -33896 -852 -33876 -788
rect -33812 -852 -33792 -788
rect -33896 -868 -33792 -852
rect -33896 -932 -33876 -868
rect -33812 -932 -33792 -868
rect -33896 -948 -33792 -932
rect -33896 -1012 -33876 -948
rect -33812 -1012 -33792 -948
rect -33896 -1028 -33792 -1012
rect -33896 -1092 -33876 -1028
rect -33812 -1092 -33792 -1028
rect -33896 -1108 -33792 -1092
rect -33896 -1172 -33876 -1108
rect -33812 -1172 -33792 -1108
rect -33896 -1188 -33792 -1172
rect -33896 -1252 -33876 -1188
rect -33812 -1252 -33792 -1188
rect -33896 -1268 -33792 -1252
rect -33896 -1332 -33876 -1268
rect -33812 -1332 -33792 -1268
rect -33896 -1348 -33792 -1332
rect -33896 -1412 -33876 -1348
rect -33812 -1412 -33792 -1348
rect -33896 -1428 -33792 -1412
rect -33896 -1492 -33876 -1428
rect -33812 -1492 -33792 -1428
rect -33896 -1508 -33792 -1492
rect -33896 -1572 -33876 -1508
rect -33812 -1572 -33792 -1508
rect -33896 -1588 -33792 -1572
rect -33896 -1652 -33876 -1588
rect -33812 -1652 -33792 -1588
rect -33896 -1668 -33792 -1652
rect -33896 -1732 -33876 -1668
rect -33812 -1732 -33792 -1668
rect -33896 -1748 -33792 -1732
rect -33896 -1812 -33876 -1748
rect -33812 -1812 -33792 -1748
rect -33896 -1828 -33792 -1812
rect -33896 -1892 -33876 -1828
rect -33812 -1892 -33792 -1828
rect -33896 -1908 -33792 -1892
rect -33896 -1972 -33876 -1908
rect -33812 -1972 -33792 -1908
rect -33896 -1988 -33792 -1972
rect -33896 -2052 -33876 -1988
rect -33812 -2052 -33792 -1988
rect -33896 -2068 -33792 -2052
rect -33896 -2132 -33876 -2068
rect -33812 -2132 -33792 -2068
rect -33896 -2148 -33792 -2132
rect -33896 -2212 -33876 -2148
rect -33812 -2212 -33792 -2148
rect -33896 -2228 -33792 -2212
rect -33896 -2292 -33876 -2228
rect -33812 -2292 -33792 -2228
rect -33896 -2308 -33792 -2292
rect -33896 -2372 -33876 -2308
rect -33812 -2372 -33792 -2308
rect -33896 -2388 -33792 -2372
rect -33896 -2452 -33876 -2388
rect -33812 -2452 -33792 -2388
rect -33896 -2468 -33792 -2452
rect -33896 -2532 -33876 -2468
rect -33812 -2532 -33792 -2468
rect -33896 -2548 -33792 -2532
rect -33896 -2612 -33876 -2548
rect -33812 -2612 -33792 -2548
rect -33896 -2628 -33792 -2612
rect -33896 -2692 -33876 -2628
rect -33812 -2692 -33792 -2628
rect -33896 -2708 -33792 -2692
rect -33896 -2772 -33876 -2708
rect -33812 -2772 -33792 -2708
rect -33896 -2788 -33792 -2772
rect -33896 -2852 -33876 -2788
rect -33812 -2852 -33792 -2788
rect -33896 -2868 -33792 -2852
rect -33896 -2932 -33876 -2868
rect -33812 -2932 -33792 -2868
rect -33896 -2948 -33792 -2932
rect -33896 -3012 -33876 -2948
rect -33812 -3012 -33792 -2948
rect -33896 -3028 -33792 -3012
rect -33896 -3092 -33876 -3028
rect -33812 -3092 -33792 -3028
rect -33896 -3108 -33792 -3092
rect -33896 -3172 -33876 -3108
rect -33812 -3172 -33792 -3108
rect -33896 -3188 -33792 -3172
rect -33896 -3252 -33876 -3188
rect -33812 -3252 -33792 -3188
rect -33896 -3268 -33792 -3252
rect -33896 -3332 -33876 -3268
rect -33812 -3332 -33792 -3268
rect -33896 -3348 -33792 -3332
rect -33896 -3412 -33876 -3348
rect -33812 -3412 -33792 -3348
rect -33896 -3428 -33792 -3412
rect -33896 -3492 -33876 -3428
rect -33812 -3492 -33792 -3428
rect -33896 -3508 -33792 -3492
rect -33896 -3572 -33876 -3508
rect -33812 -3572 -33792 -3508
rect -33896 -3588 -33792 -3572
rect -33896 -3652 -33876 -3588
rect -33812 -3652 -33792 -3588
rect -33896 -3668 -33792 -3652
rect -33896 -3732 -33876 -3668
rect -33812 -3732 -33792 -3668
rect -33896 -3748 -33792 -3732
rect -33896 -3812 -33876 -3748
rect -33812 -3812 -33792 -3748
rect -33896 -3828 -33792 -3812
rect -33896 -3892 -33876 -3828
rect -33812 -3892 -33792 -3828
rect -33896 -3908 -33792 -3892
rect -33896 -3972 -33876 -3908
rect -33812 -3972 -33792 -3908
rect -33896 -3988 -33792 -3972
rect -33896 -4052 -33876 -3988
rect -33812 -4052 -33792 -3988
rect -33896 -4068 -33792 -4052
rect -33896 -4132 -33876 -4068
rect -33812 -4132 -33792 -4068
rect -33896 -4148 -33792 -4132
rect -33896 -4212 -33876 -4148
rect -33812 -4212 -33792 -4148
rect -33896 -4228 -33792 -4212
rect -33896 -4292 -33876 -4228
rect -33812 -4292 -33792 -4228
rect -33896 -4308 -33792 -4292
rect -33896 -4372 -33876 -4308
rect -33812 -4372 -33792 -4308
rect -33896 -4388 -33792 -4372
rect -33896 -4452 -33876 -4388
rect -33812 -4452 -33792 -4388
rect -33896 -4468 -33792 -4452
rect -33896 -4532 -33876 -4468
rect -33812 -4532 -33792 -4468
rect -33896 -4548 -33792 -4532
rect -33896 -4612 -33876 -4548
rect -33812 -4612 -33792 -4548
rect -33896 -4628 -33792 -4612
rect -33896 -4692 -33876 -4628
rect -33812 -4692 -33792 -4628
rect -33896 -4708 -33792 -4692
rect -33896 -4772 -33876 -4708
rect -33812 -4772 -33792 -4708
rect -33896 -4788 -33792 -4772
rect -33896 -4852 -33876 -4788
rect -33812 -4852 -33792 -4788
rect -33896 -4868 -33792 -4852
rect -33896 -4932 -33876 -4868
rect -33812 -4932 -33792 -4868
rect -33896 -4948 -33792 -4932
rect -33896 -5012 -33876 -4948
rect -33812 -5012 -33792 -4948
rect -33896 -5028 -33792 -5012
rect -33896 -5092 -33876 -5028
rect -33812 -5092 -33792 -5028
rect -33896 -5108 -33792 -5092
rect -36676 -5519 -36572 -5121
rect -33896 -5172 -33876 -5108
rect -33812 -5172 -33792 -5108
rect -33473 -228 -28551 -199
rect -33473 -5092 -33444 -228
rect -28580 -5092 -28551 -228
rect -33473 -5121 -28551 -5092
rect -28284 -212 -28264 -148
rect -28200 -212 -28180 -148
rect -25452 -199 -25348 199
rect -22672 148 -22652 212
rect -22588 148 -22568 212
rect -22249 5092 -17327 5121
rect -22249 228 -22220 5092
rect -17356 228 -17327 5092
rect -22249 199 -17327 228
rect -17060 5108 -17040 5172
rect -16976 5108 -16956 5172
rect -14228 5121 -14124 5519
rect -11448 5468 -11428 5532
rect -11364 5468 -11344 5532
rect -11025 10412 -6103 10441
rect -11025 5548 -10996 10412
rect -6132 5548 -6103 10412
rect -11025 5519 -6103 5548
rect -5836 10428 -5816 10492
rect -5752 10428 -5732 10492
rect -3004 10441 -2900 10839
rect -224 10788 -204 10852
rect -140 10788 -120 10852
rect 199 15732 5121 15761
rect 199 10868 228 15732
rect 5092 10868 5121 15732
rect 199 10839 5121 10868
rect 5388 15748 5408 15812
rect 5472 15748 5492 15812
rect 8220 15761 8324 16159
rect 11000 16108 11020 16172
rect 11084 16108 11104 16172
rect 11423 21052 16345 21081
rect 11423 16188 11452 21052
rect 16316 16188 16345 21052
rect 11423 16159 16345 16188
rect 16612 21068 16632 21132
rect 16696 21068 16716 21132
rect 19444 21081 19548 21479
rect 22224 21428 22244 21492
rect 22308 21428 22328 21492
rect 22647 26372 27569 26401
rect 22647 21508 22676 26372
rect 27540 21508 27569 26372
rect 22647 21479 27569 21508
rect 27836 26388 27856 26452
rect 27920 26388 27940 26452
rect 30668 26401 30772 26799
rect 33448 26748 33468 26812
rect 33532 26748 33552 26812
rect 33871 31692 38793 31721
rect 33871 26828 33900 31692
rect 38764 26828 38793 31692
rect 33871 26799 38793 26828
rect 39060 31708 39080 31772
rect 39144 31708 39164 31772
rect 39060 31692 39164 31708
rect 39060 31628 39080 31692
rect 39144 31628 39164 31692
rect 39060 31612 39164 31628
rect 39060 31548 39080 31612
rect 39144 31548 39164 31612
rect 39060 31532 39164 31548
rect 39060 31468 39080 31532
rect 39144 31468 39164 31532
rect 39060 31452 39164 31468
rect 39060 31388 39080 31452
rect 39144 31388 39164 31452
rect 39060 31372 39164 31388
rect 39060 31308 39080 31372
rect 39144 31308 39164 31372
rect 39060 31292 39164 31308
rect 39060 31228 39080 31292
rect 39144 31228 39164 31292
rect 39060 31212 39164 31228
rect 39060 31148 39080 31212
rect 39144 31148 39164 31212
rect 39060 31132 39164 31148
rect 39060 31068 39080 31132
rect 39144 31068 39164 31132
rect 39060 31052 39164 31068
rect 39060 30988 39080 31052
rect 39144 30988 39164 31052
rect 39060 30972 39164 30988
rect 39060 30908 39080 30972
rect 39144 30908 39164 30972
rect 39060 30892 39164 30908
rect 39060 30828 39080 30892
rect 39144 30828 39164 30892
rect 39060 30812 39164 30828
rect 39060 30748 39080 30812
rect 39144 30748 39164 30812
rect 39060 30732 39164 30748
rect 39060 30668 39080 30732
rect 39144 30668 39164 30732
rect 39060 30652 39164 30668
rect 39060 30588 39080 30652
rect 39144 30588 39164 30652
rect 39060 30572 39164 30588
rect 39060 30508 39080 30572
rect 39144 30508 39164 30572
rect 39060 30492 39164 30508
rect 39060 30428 39080 30492
rect 39144 30428 39164 30492
rect 39060 30412 39164 30428
rect 39060 30348 39080 30412
rect 39144 30348 39164 30412
rect 39060 30332 39164 30348
rect 39060 30268 39080 30332
rect 39144 30268 39164 30332
rect 39060 30252 39164 30268
rect 39060 30188 39080 30252
rect 39144 30188 39164 30252
rect 39060 30172 39164 30188
rect 39060 30108 39080 30172
rect 39144 30108 39164 30172
rect 39060 30092 39164 30108
rect 39060 30028 39080 30092
rect 39144 30028 39164 30092
rect 39060 30012 39164 30028
rect 39060 29948 39080 30012
rect 39144 29948 39164 30012
rect 39060 29932 39164 29948
rect 39060 29868 39080 29932
rect 39144 29868 39164 29932
rect 39060 29852 39164 29868
rect 39060 29788 39080 29852
rect 39144 29788 39164 29852
rect 39060 29772 39164 29788
rect 39060 29708 39080 29772
rect 39144 29708 39164 29772
rect 39060 29692 39164 29708
rect 39060 29628 39080 29692
rect 39144 29628 39164 29692
rect 39060 29612 39164 29628
rect 39060 29548 39080 29612
rect 39144 29548 39164 29612
rect 39060 29532 39164 29548
rect 39060 29468 39080 29532
rect 39144 29468 39164 29532
rect 39060 29452 39164 29468
rect 39060 29388 39080 29452
rect 39144 29388 39164 29452
rect 39060 29372 39164 29388
rect 39060 29308 39080 29372
rect 39144 29308 39164 29372
rect 39060 29292 39164 29308
rect 39060 29228 39080 29292
rect 39144 29228 39164 29292
rect 39060 29212 39164 29228
rect 39060 29148 39080 29212
rect 39144 29148 39164 29212
rect 39060 29132 39164 29148
rect 39060 29068 39080 29132
rect 39144 29068 39164 29132
rect 39060 29052 39164 29068
rect 39060 28988 39080 29052
rect 39144 28988 39164 29052
rect 39060 28972 39164 28988
rect 39060 28908 39080 28972
rect 39144 28908 39164 28972
rect 39060 28892 39164 28908
rect 39060 28828 39080 28892
rect 39144 28828 39164 28892
rect 39060 28812 39164 28828
rect 39060 28748 39080 28812
rect 39144 28748 39164 28812
rect 39060 28732 39164 28748
rect 39060 28668 39080 28732
rect 39144 28668 39164 28732
rect 39060 28652 39164 28668
rect 39060 28588 39080 28652
rect 39144 28588 39164 28652
rect 39060 28572 39164 28588
rect 39060 28508 39080 28572
rect 39144 28508 39164 28572
rect 39060 28492 39164 28508
rect 39060 28428 39080 28492
rect 39144 28428 39164 28492
rect 39060 28412 39164 28428
rect 39060 28348 39080 28412
rect 39144 28348 39164 28412
rect 39060 28332 39164 28348
rect 39060 28268 39080 28332
rect 39144 28268 39164 28332
rect 39060 28252 39164 28268
rect 39060 28188 39080 28252
rect 39144 28188 39164 28252
rect 39060 28172 39164 28188
rect 39060 28108 39080 28172
rect 39144 28108 39164 28172
rect 39060 28092 39164 28108
rect 39060 28028 39080 28092
rect 39144 28028 39164 28092
rect 39060 28012 39164 28028
rect 39060 27948 39080 28012
rect 39144 27948 39164 28012
rect 39060 27932 39164 27948
rect 39060 27868 39080 27932
rect 39144 27868 39164 27932
rect 39060 27852 39164 27868
rect 39060 27788 39080 27852
rect 39144 27788 39164 27852
rect 39060 27772 39164 27788
rect 39060 27708 39080 27772
rect 39144 27708 39164 27772
rect 39060 27692 39164 27708
rect 39060 27628 39080 27692
rect 39144 27628 39164 27692
rect 39060 27612 39164 27628
rect 39060 27548 39080 27612
rect 39144 27548 39164 27612
rect 39060 27532 39164 27548
rect 39060 27468 39080 27532
rect 39144 27468 39164 27532
rect 39060 27452 39164 27468
rect 39060 27388 39080 27452
rect 39144 27388 39164 27452
rect 39060 27372 39164 27388
rect 39060 27308 39080 27372
rect 39144 27308 39164 27372
rect 39060 27292 39164 27308
rect 39060 27228 39080 27292
rect 39144 27228 39164 27292
rect 39060 27212 39164 27228
rect 39060 27148 39080 27212
rect 39144 27148 39164 27212
rect 39060 27132 39164 27148
rect 39060 27068 39080 27132
rect 39144 27068 39164 27132
rect 39060 27052 39164 27068
rect 39060 26988 39080 27052
rect 39144 26988 39164 27052
rect 39060 26972 39164 26988
rect 39060 26908 39080 26972
rect 39144 26908 39164 26972
rect 39060 26892 39164 26908
rect 39060 26828 39080 26892
rect 39144 26828 39164 26892
rect 39060 26812 39164 26828
rect 33448 26452 33552 26748
rect 27836 26372 27940 26388
rect 27836 26308 27856 26372
rect 27920 26308 27940 26372
rect 27836 26292 27940 26308
rect 27836 26228 27856 26292
rect 27920 26228 27940 26292
rect 27836 26212 27940 26228
rect 27836 26148 27856 26212
rect 27920 26148 27940 26212
rect 27836 26132 27940 26148
rect 27836 26068 27856 26132
rect 27920 26068 27940 26132
rect 27836 26052 27940 26068
rect 27836 25988 27856 26052
rect 27920 25988 27940 26052
rect 27836 25972 27940 25988
rect 27836 25908 27856 25972
rect 27920 25908 27940 25972
rect 27836 25892 27940 25908
rect 27836 25828 27856 25892
rect 27920 25828 27940 25892
rect 27836 25812 27940 25828
rect 27836 25748 27856 25812
rect 27920 25748 27940 25812
rect 27836 25732 27940 25748
rect 27836 25668 27856 25732
rect 27920 25668 27940 25732
rect 27836 25652 27940 25668
rect 27836 25588 27856 25652
rect 27920 25588 27940 25652
rect 27836 25572 27940 25588
rect 27836 25508 27856 25572
rect 27920 25508 27940 25572
rect 27836 25492 27940 25508
rect 27836 25428 27856 25492
rect 27920 25428 27940 25492
rect 27836 25412 27940 25428
rect 27836 25348 27856 25412
rect 27920 25348 27940 25412
rect 27836 25332 27940 25348
rect 27836 25268 27856 25332
rect 27920 25268 27940 25332
rect 27836 25252 27940 25268
rect 27836 25188 27856 25252
rect 27920 25188 27940 25252
rect 27836 25172 27940 25188
rect 27836 25108 27856 25172
rect 27920 25108 27940 25172
rect 27836 25092 27940 25108
rect 27836 25028 27856 25092
rect 27920 25028 27940 25092
rect 27836 25012 27940 25028
rect 27836 24948 27856 25012
rect 27920 24948 27940 25012
rect 27836 24932 27940 24948
rect 27836 24868 27856 24932
rect 27920 24868 27940 24932
rect 27836 24852 27940 24868
rect 27836 24788 27856 24852
rect 27920 24788 27940 24852
rect 27836 24772 27940 24788
rect 27836 24708 27856 24772
rect 27920 24708 27940 24772
rect 27836 24692 27940 24708
rect 27836 24628 27856 24692
rect 27920 24628 27940 24692
rect 27836 24612 27940 24628
rect 27836 24548 27856 24612
rect 27920 24548 27940 24612
rect 27836 24532 27940 24548
rect 27836 24468 27856 24532
rect 27920 24468 27940 24532
rect 27836 24452 27940 24468
rect 27836 24388 27856 24452
rect 27920 24388 27940 24452
rect 27836 24372 27940 24388
rect 27836 24308 27856 24372
rect 27920 24308 27940 24372
rect 27836 24292 27940 24308
rect 27836 24228 27856 24292
rect 27920 24228 27940 24292
rect 27836 24212 27940 24228
rect 27836 24148 27856 24212
rect 27920 24148 27940 24212
rect 27836 24132 27940 24148
rect 27836 24068 27856 24132
rect 27920 24068 27940 24132
rect 27836 24052 27940 24068
rect 27836 23988 27856 24052
rect 27920 23988 27940 24052
rect 27836 23972 27940 23988
rect 27836 23908 27856 23972
rect 27920 23908 27940 23972
rect 27836 23892 27940 23908
rect 27836 23828 27856 23892
rect 27920 23828 27940 23892
rect 27836 23812 27940 23828
rect 27836 23748 27856 23812
rect 27920 23748 27940 23812
rect 27836 23732 27940 23748
rect 27836 23668 27856 23732
rect 27920 23668 27940 23732
rect 27836 23652 27940 23668
rect 27836 23588 27856 23652
rect 27920 23588 27940 23652
rect 27836 23572 27940 23588
rect 27836 23508 27856 23572
rect 27920 23508 27940 23572
rect 27836 23492 27940 23508
rect 27836 23428 27856 23492
rect 27920 23428 27940 23492
rect 27836 23412 27940 23428
rect 27836 23348 27856 23412
rect 27920 23348 27940 23412
rect 27836 23332 27940 23348
rect 27836 23268 27856 23332
rect 27920 23268 27940 23332
rect 27836 23252 27940 23268
rect 27836 23188 27856 23252
rect 27920 23188 27940 23252
rect 27836 23172 27940 23188
rect 27836 23108 27856 23172
rect 27920 23108 27940 23172
rect 27836 23092 27940 23108
rect 27836 23028 27856 23092
rect 27920 23028 27940 23092
rect 27836 23012 27940 23028
rect 27836 22948 27856 23012
rect 27920 22948 27940 23012
rect 27836 22932 27940 22948
rect 27836 22868 27856 22932
rect 27920 22868 27940 22932
rect 27836 22852 27940 22868
rect 27836 22788 27856 22852
rect 27920 22788 27940 22852
rect 27836 22772 27940 22788
rect 27836 22708 27856 22772
rect 27920 22708 27940 22772
rect 27836 22692 27940 22708
rect 27836 22628 27856 22692
rect 27920 22628 27940 22692
rect 27836 22612 27940 22628
rect 27836 22548 27856 22612
rect 27920 22548 27940 22612
rect 27836 22532 27940 22548
rect 27836 22468 27856 22532
rect 27920 22468 27940 22532
rect 27836 22452 27940 22468
rect 27836 22388 27856 22452
rect 27920 22388 27940 22452
rect 27836 22372 27940 22388
rect 27836 22308 27856 22372
rect 27920 22308 27940 22372
rect 27836 22292 27940 22308
rect 27836 22228 27856 22292
rect 27920 22228 27940 22292
rect 27836 22212 27940 22228
rect 27836 22148 27856 22212
rect 27920 22148 27940 22212
rect 27836 22132 27940 22148
rect 27836 22068 27856 22132
rect 27920 22068 27940 22132
rect 27836 22052 27940 22068
rect 27836 21988 27856 22052
rect 27920 21988 27940 22052
rect 27836 21972 27940 21988
rect 27836 21908 27856 21972
rect 27920 21908 27940 21972
rect 27836 21892 27940 21908
rect 27836 21828 27856 21892
rect 27920 21828 27940 21892
rect 27836 21812 27940 21828
rect 27836 21748 27856 21812
rect 27920 21748 27940 21812
rect 27836 21732 27940 21748
rect 27836 21668 27856 21732
rect 27920 21668 27940 21732
rect 27836 21652 27940 21668
rect 27836 21588 27856 21652
rect 27920 21588 27940 21652
rect 27836 21572 27940 21588
rect 27836 21508 27856 21572
rect 27920 21508 27940 21572
rect 27836 21492 27940 21508
rect 22224 21132 22328 21428
rect 16612 21052 16716 21068
rect 16612 20988 16632 21052
rect 16696 20988 16716 21052
rect 16612 20972 16716 20988
rect 16612 20908 16632 20972
rect 16696 20908 16716 20972
rect 16612 20892 16716 20908
rect 16612 20828 16632 20892
rect 16696 20828 16716 20892
rect 16612 20812 16716 20828
rect 16612 20748 16632 20812
rect 16696 20748 16716 20812
rect 16612 20732 16716 20748
rect 16612 20668 16632 20732
rect 16696 20668 16716 20732
rect 16612 20652 16716 20668
rect 16612 20588 16632 20652
rect 16696 20588 16716 20652
rect 16612 20572 16716 20588
rect 16612 20508 16632 20572
rect 16696 20508 16716 20572
rect 16612 20492 16716 20508
rect 16612 20428 16632 20492
rect 16696 20428 16716 20492
rect 16612 20412 16716 20428
rect 16612 20348 16632 20412
rect 16696 20348 16716 20412
rect 16612 20332 16716 20348
rect 16612 20268 16632 20332
rect 16696 20268 16716 20332
rect 16612 20252 16716 20268
rect 16612 20188 16632 20252
rect 16696 20188 16716 20252
rect 16612 20172 16716 20188
rect 16612 20108 16632 20172
rect 16696 20108 16716 20172
rect 16612 20092 16716 20108
rect 16612 20028 16632 20092
rect 16696 20028 16716 20092
rect 16612 20012 16716 20028
rect 16612 19948 16632 20012
rect 16696 19948 16716 20012
rect 16612 19932 16716 19948
rect 16612 19868 16632 19932
rect 16696 19868 16716 19932
rect 16612 19852 16716 19868
rect 16612 19788 16632 19852
rect 16696 19788 16716 19852
rect 16612 19772 16716 19788
rect 16612 19708 16632 19772
rect 16696 19708 16716 19772
rect 16612 19692 16716 19708
rect 16612 19628 16632 19692
rect 16696 19628 16716 19692
rect 16612 19612 16716 19628
rect 16612 19548 16632 19612
rect 16696 19548 16716 19612
rect 16612 19532 16716 19548
rect 16612 19468 16632 19532
rect 16696 19468 16716 19532
rect 16612 19452 16716 19468
rect 16612 19388 16632 19452
rect 16696 19388 16716 19452
rect 16612 19372 16716 19388
rect 16612 19308 16632 19372
rect 16696 19308 16716 19372
rect 16612 19292 16716 19308
rect 16612 19228 16632 19292
rect 16696 19228 16716 19292
rect 16612 19212 16716 19228
rect 16612 19148 16632 19212
rect 16696 19148 16716 19212
rect 16612 19132 16716 19148
rect 16612 19068 16632 19132
rect 16696 19068 16716 19132
rect 16612 19052 16716 19068
rect 16612 18988 16632 19052
rect 16696 18988 16716 19052
rect 16612 18972 16716 18988
rect 16612 18908 16632 18972
rect 16696 18908 16716 18972
rect 16612 18892 16716 18908
rect 16612 18828 16632 18892
rect 16696 18828 16716 18892
rect 16612 18812 16716 18828
rect 16612 18748 16632 18812
rect 16696 18748 16716 18812
rect 16612 18732 16716 18748
rect 16612 18668 16632 18732
rect 16696 18668 16716 18732
rect 16612 18652 16716 18668
rect 16612 18588 16632 18652
rect 16696 18588 16716 18652
rect 16612 18572 16716 18588
rect 16612 18508 16632 18572
rect 16696 18508 16716 18572
rect 16612 18492 16716 18508
rect 16612 18428 16632 18492
rect 16696 18428 16716 18492
rect 16612 18412 16716 18428
rect 16612 18348 16632 18412
rect 16696 18348 16716 18412
rect 16612 18332 16716 18348
rect 16612 18268 16632 18332
rect 16696 18268 16716 18332
rect 16612 18252 16716 18268
rect 16612 18188 16632 18252
rect 16696 18188 16716 18252
rect 16612 18172 16716 18188
rect 16612 18108 16632 18172
rect 16696 18108 16716 18172
rect 16612 18092 16716 18108
rect 16612 18028 16632 18092
rect 16696 18028 16716 18092
rect 16612 18012 16716 18028
rect 16612 17948 16632 18012
rect 16696 17948 16716 18012
rect 16612 17932 16716 17948
rect 16612 17868 16632 17932
rect 16696 17868 16716 17932
rect 16612 17852 16716 17868
rect 16612 17788 16632 17852
rect 16696 17788 16716 17852
rect 16612 17772 16716 17788
rect 16612 17708 16632 17772
rect 16696 17708 16716 17772
rect 16612 17692 16716 17708
rect 16612 17628 16632 17692
rect 16696 17628 16716 17692
rect 16612 17612 16716 17628
rect 16612 17548 16632 17612
rect 16696 17548 16716 17612
rect 16612 17532 16716 17548
rect 16612 17468 16632 17532
rect 16696 17468 16716 17532
rect 16612 17452 16716 17468
rect 16612 17388 16632 17452
rect 16696 17388 16716 17452
rect 16612 17372 16716 17388
rect 16612 17308 16632 17372
rect 16696 17308 16716 17372
rect 16612 17292 16716 17308
rect 16612 17228 16632 17292
rect 16696 17228 16716 17292
rect 16612 17212 16716 17228
rect 16612 17148 16632 17212
rect 16696 17148 16716 17212
rect 16612 17132 16716 17148
rect 16612 17068 16632 17132
rect 16696 17068 16716 17132
rect 16612 17052 16716 17068
rect 16612 16988 16632 17052
rect 16696 16988 16716 17052
rect 16612 16972 16716 16988
rect 16612 16908 16632 16972
rect 16696 16908 16716 16972
rect 16612 16892 16716 16908
rect 16612 16828 16632 16892
rect 16696 16828 16716 16892
rect 16612 16812 16716 16828
rect 16612 16748 16632 16812
rect 16696 16748 16716 16812
rect 16612 16732 16716 16748
rect 16612 16668 16632 16732
rect 16696 16668 16716 16732
rect 16612 16652 16716 16668
rect 16612 16588 16632 16652
rect 16696 16588 16716 16652
rect 16612 16572 16716 16588
rect 16612 16508 16632 16572
rect 16696 16508 16716 16572
rect 16612 16492 16716 16508
rect 16612 16428 16632 16492
rect 16696 16428 16716 16492
rect 16612 16412 16716 16428
rect 16612 16348 16632 16412
rect 16696 16348 16716 16412
rect 16612 16332 16716 16348
rect 16612 16268 16632 16332
rect 16696 16268 16716 16332
rect 16612 16252 16716 16268
rect 16612 16188 16632 16252
rect 16696 16188 16716 16252
rect 16612 16172 16716 16188
rect 11000 15812 11104 16108
rect 5388 15732 5492 15748
rect 5388 15668 5408 15732
rect 5472 15668 5492 15732
rect 5388 15652 5492 15668
rect 5388 15588 5408 15652
rect 5472 15588 5492 15652
rect 5388 15572 5492 15588
rect 5388 15508 5408 15572
rect 5472 15508 5492 15572
rect 5388 15492 5492 15508
rect 5388 15428 5408 15492
rect 5472 15428 5492 15492
rect 5388 15412 5492 15428
rect 5388 15348 5408 15412
rect 5472 15348 5492 15412
rect 5388 15332 5492 15348
rect 5388 15268 5408 15332
rect 5472 15268 5492 15332
rect 5388 15252 5492 15268
rect 5388 15188 5408 15252
rect 5472 15188 5492 15252
rect 5388 15172 5492 15188
rect 5388 15108 5408 15172
rect 5472 15108 5492 15172
rect 5388 15092 5492 15108
rect 5388 15028 5408 15092
rect 5472 15028 5492 15092
rect 5388 15012 5492 15028
rect 5388 14948 5408 15012
rect 5472 14948 5492 15012
rect 5388 14932 5492 14948
rect 5388 14868 5408 14932
rect 5472 14868 5492 14932
rect 5388 14852 5492 14868
rect 5388 14788 5408 14852
rect 5472 14788 5492 14852
rect 5388 14772 5492 14788
rect 5388 14708 5408 14772
rect 5472 14708 5492 14772
rect 5388 14692 5492 14708
rect 5388 14628 5408 14692
rect 5472 14628 5492 14692
rect 5388 14612 5492 14628
rect 5388 14548 5408 14612
rect 5472 14548 5492 14612
rect 5388 14532 5492 14548
rect 5388 14468 5408 14532
rect 5472 14468 5492 14532
rect 5388 14452 5492 14468
rect 5388 14388 5408 14452
rect 5472 14388 5492 14452
rect 5388 14372 5492 14388
rect 5388 14308 5408 14372
rect 5472 14308 5492 14372
rect 5388 14292 5492 14308
rect 5388 14228 5408 14292
rect 5472 14228 5492 14292
rect 5388 14212 5492 14228
rect 5388 14148 5408 14212
rect 5472 14148 5492 14212
rect 5388 14132 5492 14148
rect 5388 14068 5408 14132
rect 5472 14068 5492 14132
rect 5388 14052 5492 14068
rect 5388 13988 5408 14052
rect 5472 13988 5492 14052
rect 5388 13972 5492 13988
rect 5388 13908 5408 13972
rect 5472 13908 5492 13972
rect 5388 13892 5492 13908
rect 5388 13828 5408 13892
rect 5472 13828 5492 13892
rect 5388 13812 5492 13828
rect 5388 13748 5408 13812
rect 5472 13748 5492 13812
rect 5388 13732 5492 13748
rect 5388 13668 5408 13732
rect 5472 13668 5492 13732
rect 5388 13652 5492 13668
rect 5388 13588 5408 13652
rect 5472 13588 5492 13652
rect 5388 13572 5492 13588
rect 5388 13508 5408 13572
rect 5472 13508 5492 13572
rect 5388 13492 5492 13508
rect 5388 13428 5408 13492
rect 5472 13428 5492 13492
rect 5388 13412 5492 13428
rect 5388 13348 5408 13412
rect 5472 13348 5492 13412
rect 5388 13332 5492 13348
rect 5388 13268 5408 13332
rect 5472 13268 5492 13332
rect 5388 13252 5492 13268
rect 5388 13188 5408 13252
rect 5472 13188 5492 13252
rect 5388 13172 5492 13188
rect 5388 13108 5408 13172
rect 5472 13108 5492 13172
rect 5388 13092 5492 13108
rect 5388 13028 5408 13092
rect 5472 13028 5492 13092
rect 5388 13012 5492 13028
rect 5388 12948 5408 13012
rect 5472 12948 5492 13012
rect 5388 12932 5492 12948
rect 5388 12868 5408 12932
rect 5472 12868 5492 12932
rect 5388 12852 5492 12868
rect 5388 12788 5408 12852
rect 5472 12788 5492 12852
rect 5388 12772 5492 12788
rect 5388 12708 5408 12772
rect 5472 12708 5492 12772
rect 5388 12692 5492 12708
rect 5388 12628 5408 12692
rect 5472 12628 5492 12692
rect 5388 12612 5492 12628
rect 5388 12548 5408 12612
rect 5472 12548 5492 12612
rect 5388 12532 5492 12548
rect 5388 12468 5408 12532
rect 5472 12468 5492 12532
rect 5388 12452 5492 12468
rect 5388 12388 5408 12452
rect 5472 12388 5492 12452
rect 5388 12372 5492 12388
rect 5388 12308 5408 12372
rect 5472 12308 5492 12372
rect 5388 12292 5492 12308
rect 5388 12228 5408 12292
rect 5472 12228 5492 12292
rect 5388 12212 5492 12228
rect 5388 12148 5408 12212
rect 5472 12148 5492 12212
rect 5388 12132 5492 12148
rect 5388 12068 5408 12132
rect 5472 12068 5492 12132
rect 5388 12052 5492 12068
rect 5388 11988 5408 12052
rect 5472 11988 5492 12052
rect 5388 11972 5492 11988
rect 5388 11908 5408 11972
rect 5472 11908 5492 11972
rect 5388 11892 5492 11908
rect 5388 11828 5408 11892
rect 5472 11828 5492 11892
rect 5388 11812 5492 11828
rect 5388 11748 5408 11812
rect 5472 11748 5492 11812
rect 5388 11732 5492 11748
rect 5388 11668 5408 11732
rect 5472 11668 5492 11732
rect 5388 11652 5492 11668
rect 5388 11588 5408 11652
rect 5472 11588 5492 11652
rect 5388 11572 5492 11588
rect 5388 11508 5408 11572
rect 5472 11508 5492 11572
rect 5388 11492 5492 11508
rect 5388 11428 5408 11492
rect 5472 11428 5492 11492
rect 5388 11412 5492 11428
rect 5388 11348 5408 11412
rect 5472 11348 5492 11412
rect 5388 11332 5492 11348
rect 5388 11268 5408 11332
rect 5472 11268 5492 11332
rect 5388 11252 5492 11268
rect 5388 11188 5408 11252
rect 5472 11188 5492 11252
rect 5388 11172 5492 11188
rect 5388 11108 5408 11172
rect 5472 11108 5492 11172
rect 5388 11092 5492 11108
rect 5388 11028 5408 11092
rect 5472 11028 5492 11092
rect 5388 11012 5492 11028
rect 5388 10948 5408 11012
rect 5472 10948 5492 11012
rect 5388 10932 5492 10948
rect 5388 10868 5408 10932
rect 5472 10868 5492 10932
rect 5388 10852 5492 10868
rect -224 10492 -120 10788
rect -5836 10412 -5732 10428
rect -5836 10348 -5816 10412
rect -5752 10348 -5732 10412
rect -5836 10332 -5732 10348
rect -5836 10268 -5816 10332
rect -5752 10268 -5732 10332
rect -5836 10252 -5732 10268
rect -5836 10188 -5816 10252
rect -5752 10188 -5732 10252
rect -5836 10172 -5732 10188
rect -5836 10108 -5816 10172
rect -5752 10108 -5732 10172
rect -5836 10092 -5732 10108
rect -5836 10028 -5816 10092
rect -5752 10028 -5732 10092
rect -5836 10012 -5732 10028
rect -5836 9948 -5816 10012
rect -5752 9948 -5732 10012
rect -5836 9932 -5732 9948
rect -5836 9868 -5816 9932
rect -5752 9868 -5732 9932
rect -5836 9852 -5732 9868
rect -5836 9788 -5816 9852
rect -5752 9788 -5732 9852
rect -5836 9772 -5732 9788
rect -5836 9708 -5816 9772
rect -5752 9708 -5732 9772
rect -5836 9692 -5732 9708
rect -5836 9628 -5816 9692
rect -5752 9628 -5732 9692
rect -5836 9612 -5732 9628
rect -5836 9548 -5816 9612
rect -5752 9548 -5732 9612
rect -5836 9532 -5732 9548
rect -5836 9468 -5816 9532
rect -5752 9468 -5732 9532
rect -5836 9452 -5732 9468
rect -5836 9388 -5816 9452
rect -5752 9388 -5732 9452
rect -5836 9372 -5732 9388
rect -5836 9308 -5816 9372
rect -5752 9308 -5732 9372
rect -5836 9292 -5732 9308
rect -5836 9228 -5816 9292
rect -5752 9228 -5732 9292
rect -5836 9212 -5732 9228
rect -5836 9148 -5816 9212
rect -5752 9148 -5732 9212
rect -5836 9132 -5732 9148
rect -5836 9068 -5816 9132
rect -5752 9068 -5732 9132
rect -5836 9052 -5732 9068
rect -5836 8988 -5816 9052
rect -5752 8988 -5732 9052
rect -5836 8972 -5732 8988
rect -5836 8908 -5816 8972
rect -5752 8908 -5732 8972
rect -5836 8892 -5732 8908
rect -5836 8828 -5816 8892
rect -5752 8828 -5732 8892
rect -5836 8812 -5732 8828
rect -5836 8748 -5816 8812
rect -5752 8748 -5732 8812
rect -5836 8732 -5732 8748
rect -5836 8668 -5816 8732
rect -5752 8668 -5732 8732
rect -5836 8652 -5732 8668
rect -5836 8588 -5816 8652
rect -5752 8588 -5732 8652
rect -5836 8572 -5732 8588
rect -5836 8508 -5816 8572
rect -5752 8508 -5732 8572
rect -5836 8492 -5732 8508
rect -5836 8428 -5816 8492
rect -5752 8428 -5732 8492
rect -5836 8412 -5732 8428
rect -5836 8348 -5816 8412
rect -5752 8348 -5732 8412
rect -5836 8332 -5732 8348
rect -5836 8268 -5816 8332
rect -5752 8268 -5732 8332
rect -5836 8252 -5732 8268
rect -5836 8188 -5816 8252
rect -5752 8188 -5732 8252
rect -5836 8172 -5732 8188
rect -5836 8108 -5816 8172
rect -5752 8108 -5732 8172
rect -5836 8092 -5732 8108
rect -5836 8028 -5816 8092
rect -5752 8028 -5732 8092
rect -5836 8012 -5732 8028
rect -5836 7948 -5816 8012
rect -5752 7948 -5732 8012
rect -5836 7932 -5732 7948
rect -5836 7868 -5816 7932
rect -5752 7868 -5732 7932
rect -5836 7852 -5732 7868
rect -5836 7788 -5816 7852
rect -5752 7788 -5732 7852
rect -5836 7772 -5732 7788
rect -5836 7708 -5816 7772
rect -5752 7708 -5732 7772
rect -5836 7692 -5732 7708
rect -5836 7628 -5816 7692
rect -5752 7628 -5732 7692
rect -5836 7612 -5732 7628
rect -5836 7548 -5816 7612
rect -5752 7548 -5732 7612
rect -5836 7532 -5732 7548
rect -5836 7468 -5816 7532
rect -5752 7468 -5732 7532
rect -5836 7452 -5732 7468
rect -5836 7388 -5816 7452
rect -5752 7388 -5732 7452
rect -5836 7372 -5732 7388
rect -5836 7308 -5816 7372
rect -5752 7308 -5732 7372
rect -5836 7292 -5732 7308
rect -5836 7228 -5816 7292
rect -5752 7228 -5732 7292
rect -5836 7212 -5732 7228
rect -5836 7148 -5816 7212
rect -5752 7148 -5732 7212
rect -5836 7132 -5732 7148
rect -5836 7068 -5816 7132
rect -5752 7068 -5732 7132
rect -5836 7052 -5732 7068
rect -5836 6988 -5816 7052
rect -5752 6988 -5732 7052
rect -5836 6972 -5732 6988
rect -5836 6908 -5816 6972
rect -5752 6908 -5732 6972
rect -5836 6892 -5732 6908
rect -5836 6828 -5816 6892
rect -5752 6828 -5732 6892
rect -5836 6812 -5732 6828
rect -5836 6748 -5816 6812
rect -5752 6748 -5732 6812
rect -5836 6732 -5732 6748
rect -5836 6668 -5816 6732
rect -5752 6668 -5732 6732
rect -5836 6652 -5732 6668
rect -5836 6588 -5816 6652
rect -5752 6588 -5732 6652
rect -5836 6572 -5732 6588
rect -5836 6508 -5816 6572
rect -5752 6508 -5732 6572
rect -5836 6492 -5732 6508
rect -5836 6428 -5816 6492
rect -5752 6428 -5732 6492
rect -5836 6412 -5732 6428
rect -5836 6348 -5816 6412
rect -5752 6348 -5732 6412
rect -5836 6332 -5732 6348
rect -5836 6268 -5816 6332
rect -5752 6268 -5732 6332
rect -5836 6252 -5732 6268
rect -5836 6188 -5816 6252
rect -5752 6188 -5732 6252
rect -5836 6172 -5732 6188
rect -5836 6108 -5816 6172
rect -5752 6108 -5732 6172
rect -5836 6092 -5732 6108
rect -5836 6028 -5816 6092
rect -5752 6028 -5732 6092
rect -5836 6012 -5732 6028
rect -5836 5948 -5816 6012
rect -5752 5948 -5732 6012
rect -5836 5932 -5732 5948
rect -5836 5868 -5816 5932
rect -5752 5868 -5732 5932
rect -5836 5852 -5732 5868
rect -5836 5788 -5816 5852
rect -5752 5788 -5732 5852
rect -5836 5772 -5732 5788
rect -5836 5708 -5816 5772
rect -5752 5708 -5732 5772
rect -5836 5692 -5732 5708
rect -5836 5628 -5816 5692
rect -5752 5628 -5732 5692
rect -5836 5612 -5732 5628
rect -5836 5548 -5816 5612
rect -5752 5548 -5732 5612
rect -5836 5532 -5732 5548
rect -11448 5172 -11344 5468
rect -17060 5092 -16956 5108
rect -17060 5028 -17040 5092
rect -16976 5028 -16956 5092
rect -17060 5012 -16956 5028
rect -17060 4948 -17040 5012
rect -16976 4948 -16956 5012
rect -17060 4932 -16956 4948
rect -17060 4868 -17040 4932
rect -16976 4868 -16956 4932
rect -17060 4852 -16956 4868
rect -17060 4788 -17040 4852
rect -16976 4788 -16956 4852
rect -17060 4772 -16956 4788
rect -17060 4708 -17040 4772
rect -16976 4708 -16956 4772
rect -17060 4692 -16956 4708
rect -17060 4628 -17040 4692
rect -16976 4628 -16956 4692
rect -17060 4612 -16956 4628
rect -17060 4548 -17040 4612
rect -16976 4548 -16956 4612
rect -17060 4532 -16956 4548
rect -17060 4468 -17040 4532
rect -16976 4468 -16956 4532
rect -17060 4452 -16956 4468
rect -17060 4388 -17040 4452
rect -16976 4388 -16956 4452
rect -17060 4372 -16956 4388
rect -17060 4308 -17040 4372
rect -16976 4308 -16956 4372
rect -17060 4292 -16956 4308
rect -17060 4228 -17040 4292
rect -16976 4228 -16956 4292
rect -17060 4212 -16956 4228
rect -17060 4148 -17040 4212
rect -16976 4148 -16956 4212
rect -17060 4132 -16956 4148
rect -17060 4068 -17040 4132
rect -16976 4068 -16956 4132
rect -17060 4052 -16956 4068
rect -17060 3988 -17040 4052
rect -16976 3988 -16956 4052
rect -17060 3972 -16956 3988
rect -17060 3908 -17040 3972
rect -16976 3908 -16956 3972
rect -17060 3892 -16956 3908
rect -17060 3828 -17040 3892
rect -16976 3828 -16956 3892
rect -17060 3812 -16956 3828
rect -17060 3748 -17040 3812
rect -16976 3748 -16956 3812
rect -17060 3732 -16956 3748
rect -17060 3668 -17040 3732
rect -16976 3668 -16956 3732
rect -17060 3652 -16956 3668
rect -17060 3588 -17040 3652
rect -16976 3588 -16956 3652
rect -17060 3572 -16956 3588
rect -17060 3508 -17040 3572
rect -16976 3508 -16956 3572
rect -17060 3492 -16956 3508
rect -17060 3428 -17040 3492
rect -16976 3428 -16956 3492
rect -17060 3412 -16956 3428
rect -17060 3348 -17040 3412
rect -16976 3348 -16956 3412
rect -17060 3332 -16956 3348
rect -17060 3268 -17040 3332
rect -16976 3268 -16956 3332
rect -17060 3252 -16956 3268
rect -17060 3188 -17040 3252
rect -16976 3188 -16956 3252
rect -17060 3172 -16956 3188
rect -17060 3108 -17040 3172
rect -16976 3108 -16956 3172
rect -17060 3092 -16956 3108
rect -17060 3028 -17040 3092
rect -16976 3028 -16956 3092
rect -17060 3012 -16956 3028
rect -17060 2948 -17040 3012
rect -16976 2948 -16956 3012
rect -17060 2932 -16956 2948
rect -17060 2868 -17040 2932
rect -16976 2868 -16956 2932
rect -17060 2852 -16956 2868
rect -17060 2788 -17040 2852
rect -16976 2788 -16956 2852
rect -17060 2772 -16956 2788
rect -17060 2708 -17040 2772
rect -16976 2708 -16956 2772
rect -17060 2692 -16956 2708
rect -17060 2628 -17040 2692
rect -16976 2628 -16956 2692
rect -17060 2612 -16956 2628
rect -17060 2548 -17040 2612
rect -16976 2548 -16956 2612
rect -17060 2532 -16956 2548
rect -17060 2468 -17040 2532
rect -16976 2468 -16956 2532
rect -17060 2452 -16956 2468
rect -17060 2388 -17040 2452
rect -16976 2388 -16956 2452
rect -17060 2372 -16956 2388
rect -17060 2308 -17040 2372
rect -16976 2308 -16956 2372
rect -17060 2292 -16956 2308
rect -17060 2228 -17040 2292
rect -16976 2228 -16956 2292
rect -17060 2212 -16956 2228
rect -17060 2148 -17040 2212
rect -16976 2148 -16956 2212
rect -17060 2132 -16956 2148
rect -17060 2068 -17040 2132
rect -16976 2068 -16956 2132
rect -17060 2052 -16956 2068
rect -17060 1988 -17040 2052
rect -16976 1988 -16956 2052
rect -17060 1972 -16956 1988
rect -17060 1908 -17040 1972
rect -16976 1908 -16956 1972
rect -17060 1892 -16956 1908
rect -17060 1828 -17040 1892
rect -16976 1828 -16956 1892
rect -17060 1812 -16956 1828
rect -17060 1748 -17040 1812
rect -16976 1748 -16956 1812
rect -17060 1732 -16956 1748
rect -17060 1668 -17040 1732
rect -16976 1668 -16956 1732
rect -17060 1652 -16956 1668
rect -17060 1588 -17040 1652
rect -16976 1588 -16956 1652
rect -17060 1572 -16956 1588
rect -17060 1508 -17040 1572
rect -16976 1508 -16956 1572
rect -17060 1492 -16956 1508
rect -17060 1428 -17040 1492
rect -16976 1428 -16956 1492
rect -17060 1412 -16956 1428
rect -17060 1348 -17040 1412
rect -16976 1348 -16956 1412
rect -17060 1332 -16956 1348
rect -17060 1268 -17040 1332
rect -16976 1268 -16956 1332
rect -17060 1252 -16956 1268
rect -17060 1188 -17040 1252
rect -16976 1188 -16956 1252
rect -17060 1172 -16956 1188
rect -17060 1108 -17040 1172
rect -16976 1108 -16956 1172
rect -17060 1092 -16956 1108
rect -17060 1028 -17040 1092
rect -16976 1028 -16956 1092
rect -17060 1012 -16956 1028
rect -17060 948 -17040 1012
rect -16976 948 -16956 1012
rect -17060 932 -16956 948
rect -17060 868 -17040 932
rect -16976 868 -16956 932
rect -17060 852 -16956 868
rect -17060 788 -17040 852
rect -16976 788 -16956 852
rect -17060 772 -16956 788
rect -17060 708 -17040 772
rect -16976 708 -16956 772
rect -17060 692 -16956 708
rect -17060 628 -17040 692
rect -16976 628 -16956 692
rect -17060 612 -16956 628
rect -17060 548 -17040 612
rect -16976 548 -16956 612
rect -17060 532 -16956 548
rect -17060 468 -17040 532
rect -16976 468 -16956 532
rect -17060 452 -16956 468
rect -17060 388 -17040 452
rect -16976 388 -16956 452
rect -17060 372 -16956 388
rect -17060 308 -17040 372
rect -16976 308 -16956 372
rect -17060 292 -16956 308
rect -17060 228 -17040 292
rect -16976 228 -16956 292
rect -17060 212 -16956 228
rect -22672 -148 -22568 148
rect -28284 -228 -28180 -212
rect -28284 -292 -28264 -228
rect -28200 -292 -28180 -228
rect -28284 -308 -28180 -292
rect -28284 -372 -28264 -308
rect -28200 -372 -28180 -308
rect -28284 -388 -28180 -372
rect -28284 -452 -28264 -388
rect -28200 -452 -28180 -388
rect -28284 -468 -28180 -452
rect -28284 -532 -28264 -468
rect -28200 -532 -28180 -468
rect -28284 -548 -28180 -532
rect -28284 -612 -28264 -548
rect -28200 -612 -28180 -548
rect -28284 -628 -28180 -612
rect -28284 -692 -28264 -628
rect -28200 -692 -28180 -628
rect -28284 -708 -28180 -692
rect -28284 -772 -28264 -708
rect -28200 -772 -28180 -708
rect -28284 -788 -28180 -772
rect -28284 -852 -28264 -788
rect -28200 -852 -28180 -788
rect -28284 -868 -28180 -852
rect -28284 -932 -28264 -868
rect -28200 -932 -28180 -868
rect -28284 -948 -28180 -932
rect -28284 -1012 -28264 -948
rect -28200 -1012 -28180 -948
rect -28284 -1028 -28180 -1012
rect -28284 -1092 -28264 -1028
rect -28200 -1092 -28180 -1028
rect -28284 -1108 -28180 -1092
rect -28284 -1172 -28264 -1108
rect -28200 -1172 -28180 -1108
rect -28284 -1188 -28180 -1172
rect -28284 -1252 -28264 -1188
rect -28200 -1252 -28180 -1188
rect -28284 -1268 -28180 -1252
rect -28284 -1332 -28264 -1268
rect -28200 -1332 -28180 -1268
rect -28284 -1348 -28180 -1332
rect -28284 -1412 -28264 -1348
rect -28200 -1412 -28180 -1348
rect -28284 -1428 -28180 -1412
rect -28284 -1492 -28264 -1428
rect -28200 -1492 -28180 -1428
rect -28284 -1508 -28180 -1492
rect -28284 -1572 -28264 -1508
rect -28200 -1572 -28180 -1508
rect -28284 -1588 -28180 -1572
rect -28284 -1652 -28264 -1588
rect -28200 -1652 -28180 -1588
rect -28284 -1668 -28180 -1652
rect -28284 -1732 -28264 -1668
rect -28200 -1732 -28180 -1668
rect -28284 -1748 -28180 -1732
rect -28284 -1812 -28264 -1748
rect -28200 -1812 -28180 -1748
rect -28284 -1828 -28180 -1812
rect -28284 -1892 -28264 -1828
rect -28200 -1892 -28180 -1828
rect -28284 -1908 -28180 -1892
rect -28284 -1972 -28264 -1908
rect -28200 -1972 -28180 -1908
rect -28284 -1988 -28180 -1972
rect -28284 -2052 -28264 -1988
rect -28200 -2052 -28180 -1988
rect -28284 -2068 -28180 -2052
rect -28284 -2132 -28264 -2068
rect -28200 -2132 -28180 -2068
rect -28284 -2148 -28180 -2132
rect -28284 -2212 -28264 -2148
rect -28200 -2212 -28180 -2148
rect -28284 -2228 -28180 -2212
rect -28284 -2292 -28264 -2228
rect -28200 -2292 -28180 -2228
rect -28284 -2308 -28180 -2292
rect -28284 -2372 -28264 -2308
rect -28200 -2372 -28180 -2308
rect -28284 -2388 -28180 -2372
rect -28284 -2452 -28264 -2388
rect -28200 -2452 -28180 -2388
rect -28284 -2468 -28180 -2452
rect -28284 -2532 -28264 -2468
rect -28200 -2532 -28180 -2468
rect -28284 -2548 -28180 -2532
rect -28284 -2612 -28264 -2548
rect -28200 -2612 -28180 -2548
rect -28284 -2628 -28180 -2612
rect -28284 -2692 -28264 -2628
rect -28200 -2692 -28180 -2628
rect -28284 -2708 -28180 -2692
rect -28284 -2772 -28264 -2708
rect -28200 -2772 -28180 -2708
rect -28284 -2788 -28180 -2772
rect -28284 -2852 -28264 -2788
rect -28200 -2852 -28180 -2788
rect -28284 -2868 -28180 -2852
rect -28284 -2932 -28264 -2868
rect -28200 -2932 -28180 -2868
rect -28284 -2948 -28180 -2932
rect -28284 -3012 -28264 -2948
rect -28200 -3012 -28180 -2948
rect -28284 -3028 -28180 -3012
rect -28284 -3092 -28264 -3028
rect -28200 -3092 -28180 -3028
rect -28284 -3108 -28180 -3092
rect -28284 -3172 -28264 -3108
rect -28200 -3172 -28180 -3108
rect -28284 -3188 -28180 -3172
rect -28284 -3252 -28264 -3188
rect -28200 -3252 -28180 -3188
rect -28284 -3268 -28180 -3252
rect -28284 -3332 -28264 -3268
rect -28200 -3332 -28180 -3268
rect -28284 -3348 -28180 -3332
rect -28284 -3412 -28264 -3348
rect -28200 -3412 -28180 -3348
rect -28284 -3428 -28180 -3412
rect -28284 -3492 -28264 -3428
rect -28200 -3492 -28180 -3428
rect -28284 -3508 -28180 -3492
rect -28284 -3572 -28264 -3508
rect -28200 -3572 -28180 -3508
rect -28284 -3588 -28180 -3572
rect -28284 -3652 -28264 -3588
rect -28200 -3652 -28180 -3588
rect -28284 -3668 -28180 -3652
rect -28284 -3732 -28264 -3668
rect -28200 -3732 -28180 -3668
rect -28284 -3748 -28180 -3732
rect -28284 -3812 -28264 -3748
rect -28200 -3812 -28180 -3748
rect -28284 -3828 -28180 -3812
rect -28284 -3892 -28264 -3828
rect -28200 -3892 -28180 -3828
rect -28284 -3908 -28180 -3892
rect -28284 -3972 -28264 -3908
rect -28200 -3972 -28180 -3908
rect -28284 -3988 -28180 -3972
rect -28284 -4052 -28264 -3988
rect -28200 -4052 -28180 -3988
rect -28284 -4068 -28180 -4052
rect -28284 -4132 -28264 -4068
rect -28200 -4132 -28180 -4068
rect -28284 -4148 -28180 -4132
rect -28284 -4212 -28264 -4148
rect -28200 -4212 -28180 -4148
rect -28284 -4228 -28180 -4212
rect -28284 -4292 -28264 -4228
rect -28200 -4292 -28180 -4228
rect -28284 -4308 -28180 -4292
rect -28284 -4372 -28264 -4308
rect -28200 -4372 -28180 -4308
rect -28284 -4388 -28180 -4372
rect -28284 -4452 -28264 -4388
rect -28200 -4452 -28180 -4388
rect -28284 -4468 -28180 -4452
rect -28284 -4532 -28264 -4468
rect -28200 -4532 -28180 -4468
rect -28284 -4548 -28180 -4532
rect -28284 -4612 -28264 -4548
rect -28200 -4612 -28180 -4548
rect -28284 -4628 -28180 -4612
rect -28284 -4692 -28264 -4628
rect -28200 -4692 -28180 -4628
rect -28284 -4708 -28180 -4692
rect -28284 -4772 -28264 -4708
rect -28200 -4772 -28180 -4708
rect -28284 -4788 -28180 -4772
rect -28284 -4852 -28264 -4788
rect -28200 -4852 -28180 -4788
rect -28284 -4868 -28180 -4852
rect -28284 -4932 -28264 -4868
rect -28200 -4932 -28180 -4868
rect -28284 -4948 -28180 -4932
rect -28284 -5012 -28264 -4948
rect -28200 -5012 -28180 -4948
rect -28284 -5028 -28180 -5012
rect -28284 -5092 -28264 -5028
rect -28200 -5092 -28180 -5028
rect -28284 -5108 -28180 -5092
rect -33896 -5468 -33792 -5172
rect -39085 -5548 -34163 -5519
rect -39085 -10412 -39056 -5548
rect -34192 -10412 -34163 -5548
rect -39085 -10441 -34163 -10412
rect -33896 -5532 -33876 -5468
rect -33812 -5532 -33792 -5468
rect -31064 -5519 -30960 -5121
rect -28284 -5172 -28264 -5108
rect -28200 -5172 -28180 -5108
rect -27861 -228 -22939 -199
rect -27861 -5092 -27832 -228
rect -22968 -5092 -22939 -228
rect -27861 -5121 -22939 -5092
rect -22672 -212 -22652 -148
rect -22588 -212 -22568 -148
rect -19840 -199 -19736 199
rect -17060 148 -17040 212
rect -16976 148 -16956 212
rect -16637 5092 -11715 5121
rect -16637 228 -16608 5092
rect -11744 228 -11715 5092
rect -16637 199 -11715 228
rect -11448 5108 -11428 5172
rect -11364 5108 -11344 5172
rect -8616 5121 -8512 5519
rect -5836 5468 -5816 5532
rect -5752 5468 -5732 5532
rect -5413 10412 -491 10441
rect -5413 5548 -5384 10412
rect -520 5548 -491 10412
rect -5413 5519 -491 5548
rect -224 10428 -204 10492
rect -140 10428 -120 10492
rect 2608 10441 2712 10839
rect 5388 10788 5408 10852
rect 5472 10788 5492 10852
rect 5811 15732 10733 15761
rect 5811 10868 5840 15732
rect 10704 10868 10733 15732
rect 5811 10839 10733 10868
rect 11000 15748 11020 15812
rect 11084 15748 11104 15812
rect 13832 15761 13936 16159
rect 16612 16108 16632 16172
rect 16696 16108 16716 16172
rect 17035 21052 21957 21081
rect 17035 16188 17064 21052
rect 21928 16188 21957 21052
rect 17035 16159 21957 16188
rect 22224 21068 22244 21132
rect 22308 21068 22328 21132
rect 25056 21081 25160 21479
rect 27836 21428 27856 21492
rect 27920 21428 27940 21492
rect 28259 26372 33181 26401
rect 28259 21508 28288 26372
rect 33152 21508 33181 26372
rect 28259 21479 33181 21508
rect 33448 26388 33468 26452
rect 33532 26388 33552 26452
rect 36280 26401 36384 26799
rect 39060 26748 39080 26812
rect 39144 26748 39164 26812
rect 39060 26452 39164 26748
rect 33448 26372 33552 26388
rect 33448 26308 33468 26372
rect 33532 26308 33552 26372
rect 33448 26292 33552 26308
rect 33448 26228 33468 26292
rect 33532 26228 33552 26292
rect 33448 26212 33552 26228
rect 33448 26148 33468 26212
rect 33532 26148 33552 26212
rect 33448 26132 33552 26148
rect 33448 26068 33468 26132
rect 33532 26068 33552 26132
rect 33448 26052 33552 26068
rect 33448 25988 33468 26052
rect 33532 25988 33552 26052
rect 33448 25972 33552 25988
rect 33448 25908 33468 25972
rect 33532 25908 33552 25972
rect 33448 25892 33552 25908
rect 33448 25828 33468 25892
rect 33532 25828 33552 25892
rect 33448 25812 33552 25828
rect 33448 25748 33468 25812
rect 33532 25748 33552 25812
rect 33448 25732 33552 25748
rect 33448 25668 33468 25732
rect 33532 25668 33552 25732
rect 33448 25652 33552 25668
rect 33448 25588 33468 25652
rect 33532 25588 33552 25652
rect 33448 25572 33552 25588
rect 33448 25508 33468 25572
rect 33532 25508 33552 25572
rect 33448 25492 33552 25508
rect 33448 25428 33468 25492
rect 33532 25428 33552 25492
rect 33448 25412 33552 25428
rect 33448 25348 33468 25412
rect 33532 25348 33552 25412
rect 33448 25332 33552 25348
rect 33448 25268 33468 25332
rect 33532 25268 33552 25332
rect 33448 25252 33552 25268
rect 33448 25188 33468 25252
rect 33532 25188 33552 25252
rect 33448 25172 33552 25188
rect 33448 25108 33468 25172
rect 33532 25108 33552 25172
rect 33448 25092 33552 25108
rect 33448 25028 33468 25092
rect 33532 25028 33552 25092
rect 33448 25012 33552 25028
rect 33448 24948 33468 25012
rect 33532 24948 33552 25012
rect 33448 24932 33552 24948
rect 33448 24868 33468 24932
rect 33532 24868 33552 24932
rect 33448 24852 33552 24868
rect 33448 24788 33468 24852
rect 33532 24788 33552 24852
rect 33448 24772 33552 24788
rect 33448 24708 33468 24772
rect 33532 24708 33552 24772
rect 33448 24692 33552 24708
rect 33448 24628 33468 24692
rect 33532 24628 33552 24692
rect 33448 24612 33552 24628
rect 33448 24548 33468 24612
rect 33532 24548 33552 24612
rect 33448 24532 33552 24548
rect 33448 24468 33468 24532
rect 33532 24468 33552 24532
rect 33448 24452 33552 24468
rect 33448 24388 33468 24452
rect 33532 24388 33552 24452
rect 33448 24372 33552 24388
rect 33448 24308 33468 24372
rect 33532 24308 33552 24372
rect 33448 24292 33552 24308
rect 33448 24228 33468 24292
rect 33532 24228 33552 24292
rect 33448 24212 33552 24228
rect 33448 24148 33468 24212
rect 33532 24148 33552 24212
rect 33448 24132 33552 24148
rect 33448 24068 33468 24132
rect 33532 24068 33552 24132
rect 33448 24052 33552 24068
rect 33448 23988 33468 24052
rect 33532 23988 33552 24052
rect 33448 23972 33552 23988
rect 33448 23908 33468 23972
rect 33532 23908 33552 23972
rect 33448 23892 33552 23908
rect 33448 23828 33468 23892
rect 33532 23828 33552 23892
rect 33448 23812 33552 23828
rect 33448 23748 33468 23812
rect 33532 23748 33552 23812
rect 33448 23732 33552 23748
rect 33448 23668 33468 23732
rect 33532 23668 33552 23732
rect 33448 23652 33552 23668
rect 33448 23588 33468 23652
rect 33532 23588 33552 23652
rect 33448 23572 33552 23588
rect 33448 23508 33468 23572
rect 33532 23508 33552 23572
rect 33448 23492 33552 23508
rect 33448 23428 33468 23492
rect 33532 23428 33552 23492
rect 33448 23412 33552 23428
rect 33448 23348 33468 23412
rect 33532 23348 33552 23412
rect 33448 23332 33552 23348
rect 33448 23268 33468 23332
rect 33532 23268 33552 23332
rect 33448 23252 33552 23268
rect 33448 23188 33468 23252
rect 33532 23188 33552 23252
rect 33448 23172 33552 23188
rect 33448 23108 33468 23172
rect 33532 23108 33552 23172
rect 33448 23092 33552 23108
rect 33448 23028 33468 23092
rect 33532 23028 33552 23092
rect 33448 23012 33552 23028
rect 33448 22948 33468 23012
rect 33532 22948 33552 23012
rect 33448 22932 33552 22948
rect 33448 22868 33468 22932
rect 33532 22868 33552 22932
rect 33448 22852 33552 22868
rect 33448 22788 33468 22852
rect 33532 22788 33552 22852
rect 33448 22772 33552 22788
rect 33448 22708 33468 22772
rect 33532 22708 33552 22772
rect 33448 22692 33552 22708
rect 33448 22628 33468 22692
rect 33532 22628 33552 22692
rect 33448 22612 33552 22628
rect 33448 22548 33468 22612
rect 33532 22548 33552 22612
rect 33448 22532 33552 22548
rect 33448 22468 33468 22532
rect 33532 22468 33552 22532
rect 33448 22452 33552 22468
rect 33448 22388 33468 22452
rect 33532 22388 33552 22452
rect 33448 22372 33552 22388
rect 33448 22308 33468 22372
rect 33532 22308 33552 22372
rect 33448 22292 33552 22308
rect 33448 22228 33468 22292
rect 33532 22228 33552 22292
rect 33448 22212 33552 22228
rect 33448 22148 33468 22212
rect 33532 22148 33552 22212
rect 33448 22132 33552 22148
rect 33448 22068 33468 22132
rect 33532 22068 33552 22132
rect 33448 22052 33552 22068
rect 33448 21988 33468 22052
rect 33532 21988 33552 22052
rect 33448 21972 33552 21988
rect 33448 21908 33468 21972
rect 33532 21908 33552 21972
rect 33448 21892 33552 21908
rect 33448 21828 33468 21892
rect 33532 21828 33552 21892
rect 33448 21812 33552 21828
rect 33448 21748 33468 21812
rect 33532 21748 33552 21812
rect 33448 21732 33552 21748
rect 33448 21668 33468 21732
rect 33532 21668 33552 21732
rect 33448 21652 33552 21668
rect 33448 21588 33468 21652
rect 33532 21588 33552 21652
rect 33448 21572 33552 21588
rect 33448 21508 33468 21572
rect 33532 21508 33552 21572
rect 33448 21492 33552 21508
rect 27836 21132 27940 21428
rect 22224 21052 22328 21068
rect 22224 20988 22244 21052
rect 22308 20988 22328 21052
rect 22224 20972 22328 20988
rect 22224 20908 22244 20972
rect 22308 20908 22328 20972
rect 22224 20892 22328 20908
rect 22224 20828 22244 20892
rect 22308 20828 22328 20892
rect 22224 20812 22328 20828
rect 22224 20748 22244 20812
rect 22308 20748 22328 20812
rect 22224 20732 22328 20748
rect 22224 20668 22244 20732
rect 22308 20668 22328 20732
rect 22224 20652 22328 20668
rect 22224 20588 22244 20652
rect 22308 20588 22328 20652
rect 22224 20572 22328 20588
rect 22224 20508 22244 20572
rect 22308 20508 22328 20572
rect 22224 20492 22328 20508
rect 22224 20428 22244 20492
rect 22308 20428 22328 20492
rect 22224 20412 22328 20428
rect 22224 20348 22244 20412
rect 22308 20348 22328 20412
rect 22224 20332 22328 20348
rect 22224 20268 22244 20332
rect 22308 20268 22328 20332
rect 22224 20252 22328 20268
rect 22224 20188 22244 20252
rect 22308 20188 22328 20252
rect 22224 20172 22328 20188
rect 22224 20108 22244 20172
rect 22308 20108 22328 20172
rect 22224 20092 22328 20108
rect 22224 20028 22244 20092
rect 22308 20028 22328 20092
rect 22224 20012 22328 20028
rect 22224 19948 22244 20012
rect 22308 19948 22328 20012
rect 22224 19932 22328 19948
rect 22224 19868 22244 19932
rect 22308 19868 22328 19932
rect 22224 19852 22328 19868
rect 22224 19788 22244 19852
rect 22308 19788 22328 19852
rect 22224 19772 22328 19788
rect 22224 19708 22244 19772
rect 22308 19708 22328 19772
rect 22224 19692 22328 19708
rect 22224 19628 22244 19692
rect 22308 19628 22328 19692
rect 22224 19612 22328 19628
rect 22224 19548 22244 19612
rect 22308 19548 22328 19612
rect 22224 19532 22328 19548
rect 22224 19468 22244 19532
rect 22308 19468 22328 19532
rect 22224 19452 22328 19468
rect 22224 19388 22244 19452
rect 22308 19388 22328 19452
rect 22224 19372 22328 19388
rect 22224 19308 22244 19372
rect 22308 19308 22328 19372
rect 22224 19292 22328 19308
rect 22224 19228 22244 19292
rect 22308 19228 22328 19292
rect 22224 19212 22328 19228
rect 22224 19148 22244 19212
rect 22308 19148 22328 19212
rect 22224 19132 22328 19148
rect 22224 19068 22244 19132
rect 22308 19068 22328 19132
rect 22224 19052 22328 19068
rect 22224 18988 22244 19052
rect 22308 18988 22328 19052
rect 22224 18972 22328 18988
rect 22224 18908 22244 18972
rect 22308 18908 22328 18972
rect 22224 18892 22328 18908
rect 22224 18828 22244 18892
rect 22308 18828 22328 18892
rect 22224 18812 22328 18828
rect 22224 18748 22244 18812
rect 22308 18748 22328 18812
rect 22224 18732 22328 18748
rect 22224 18668 22244 18732
rect 22308 18668 22328 18732
rect 22224 18652 22328 18668
rect 22224 18588 22244 18652
rect 22308 18588 22328 18652
rect 22224 18572 22328 18588
rect 22224 18508 22244 18572
rect 22308 18508 22328 18572
rect 22224 18492 22328 18508
rect 22224 18428 22244 18492
rect 22308 18428 22328 18492
rect 22224 18412 22328 18428
rect 22224 18348 22244 18412
rect 22308 18348 22328 18412
rect 22224 18332 22328 18348
rect 22224 18268 22244 18332
rect 22308 18268 22328 18332
rect 22224 18252 22328 18268
rect 22224 18188 22244 18252
rect 22308 18188 22328 18252
rect 22224 18172 22328 18188
rect 22224 18108 22244 18172
rect 22308 18108 22328 18172
rect 22224 18092 22328 18108
rect 22224 18028 22244 18092
rect 22308 18028 22328 18092
rect 22224 18012 22328 18028
rect 22224 17948 22244 18012
rect 22308 17948 22328 18012
rect 22224 17932 22328 17948
rect 22224 17868 22244 17932
rect 22308 17868 22328 17932
rect 22224 17852 22328 17868
rect 22224 17788 22244 17852
rect 22308 17788 22328 17852
rect 22224 17772 22328 17788
rect 22224 17708 22244 17772
rect 22308 17708 22328 17772
rect 22224 17692 22328 17708
rect 22224 17628 22244 17692
rect 22308 17628 22328 17692
rect 22224 17612 22328 17628
rect 22224 17548 22244 17612
rect 22308 17548 22328 17612
rect 22224 17532 22328 17548
rect 22224 17468 22244 17532
rect 22308 17468 22328 17532
rect 22224 17452 22328 17468
rect 22224 17388 22244 17452
rect 22308 17388 22328 17452
rect 22224 17372 22328 17388
rect 22224 17308 22244 17372
rect 22308 17308 22328 17372
rect 22224 17292 22328 17308
rect 22224 17228 22244 17292
rect 22308 17228 22328 17292
rect 22224 17212 22328 17228
rect 22224 17148 22244 17212
rect 22308 17148 22328 17212
rect 22224 17132 22328 17148
rect 22224 17068 22244 17132
rect 22308 17068 22328 17132
rect 22224 17052 22328 17068
rect 22224 16988 22244 17052
rect 22308 16988 22328 17052
rect 22224 16972 22328 16988
rect 22224 16908 22244 16972
rect 22308 16908 22328 16972
rect 22224 16892 22328 16908
rect 22224 16828 22244 16892
rect 22308 16828 22328 16892
rect 22224 16812 22328 16828
rect 22224 16748 22244 16812
rect 22308 16748 22328 16812
rect 22224 16732 22328 16748
rect 22224 16668 22244 16732
rect 22308 16668 22328 16732
rect 22224 16652 22328 16668
rect 22224 16588 22244 16652
rect 22308 16588 22328 16652
rect 22224 16572 22328 16588
rect 22224 16508 22244 16572
rect 22308 16508 22328 16572
rect 22224 16492 22328 16508
rect 22224 16428 22244 16492
rect 22308 16428 22328 16492
rect 22224 16412 22328 16428
rect 22224 16348 22244 16412
rect 22308 16348 22328 16412
rect 22224 16332 22328 16348
rect 22224 16268 22244 16332
rect 22308 16268 22328 16332
rect 22224 16252 22328 16268
rect 22224 16188 22244 16252
rect 22308 16188 22328 16252
rect 22224 16172 22328 16188
rect 16612 15812 16716 16108
rect 11000 15732 11104 15748
rect 11000 15668 11020 15732
rect 11084 15668 11104 15732
rect 11000 15652 11104 15668
rect 11000 15588 11020 15652
rect 11084 15588 11104 15652
rect 11000 15572 11104 15588
rect 11000 15508 11020 15572
rect 11084 15508 11104 15572
rect 11000 15492 11104 15508
rect 11000 15428 11020 15492
rect 11084 15428 11104 15492
rect 11000 15412 11104 15428
rect 11000 15348 11020 15412
rect 11084 15348 11104 15412
rect 11000 15332 11104 15348
rect 11000 15268 11020 15332
rect 11084 15268 11104 15332
rect 11000 15252 11104 15268
rect 11000 15188 11020 15252
rect 11084 15188 11104 15252
rect 11000 15172 11104 15188
rect 11000 15108 11020 15172
rect 11084 15108 11104 15172
rect 11000 15092 11104 15108
rect 11000 15028 11020 15092
rect 11084 15028 11104 15092
rect 11000 15012 11104 15028
rect 11000 14948 11020 15012
rect 11084 14948 11104 15012
rect 11000 14932 11104 14948
rect 11000 14868 11020 14932
rect 11084 14868 11104 14932
rect 11000 14852 11104 14868
rect 11000 14788 11020 14852
rect 11084 14788 11104 14852
rect 11000 14772 11104 14788
rect 11000 14708 11020 14772
rect 11084 14708 11104 14772
rect 11000 14692 11104 14708
rect 11000 14628 11020 14692
rect 11084 14628 11104 14692
rect 11000 14612 11104 14628
rect 11000 14548 11020 14612
rect 11084 14548 11104 14612
rect 11000 14532 11104 14548
rect 11000 14468 11020 14532
rect 11084 14468 11104 14532
rect 11000 14452 11104 14468
rect 11000 14388 11020 14452
rect 11084 14388 11104 14452
rect 11000 14372 11104 14388
rect 11000 14308 11020 14372
rect 11084 14308 11104 14372
rect 11000 14292 11104 14308
rect 11000 14228 11020 14292
rect 11084 14228 11104 14292
rect 11000 14212 11104 14228
rect 11000 14148 11020 14212
rect 11084 14148 11104 14212
rect 11000 14132 11104 14148
rect 11000 14068 11020 14132
rect 11084 14068 11104 14132
rect 11000 14052 11104 14068
rect 11000 13988 11020 14052
rect 11084 13988 11104 14052
rect 11000 13972 11104 13988
rect 11000 13908 11020 13972
rect 11084 13908 11104 13972
rect 11000 13892 11104 13908
rect 11000 13828 11020 13892
rect 11084 13828 11104 13892
rect 11000 13812 11104 13828
rect 11000 13748 11020 13812
rect 11084 13748 11104 13812
rect 11000 13732 11104 13748
rect 11000 13668 11020 13732
rect 11084 13668 11104 13732
rect 11000 13652 11104 13668
rect 11000 13588 11020 13652
rect 11084 13588 11104 13652
rect 11000 13572 11104 13588
rect 11000 13508 11020 13572
rect 11084 13508 11104 13572
rect 11000 13492 11104 13508
rect 11000 13428 11020 13492
rect 11084 13428 11104 13492
rect 11000 13412 11104 13428
rect 11000 13348 11020 13412
rect 11084 13348 11104 13412
rect 11000 13332 11104 13348
rect 11000 13268 11020 13332
rect 11084 13268 11104 13332
rect 11000 13252 11104 13268
rect 11000 13188 11020 13252
rect 11084 13188 11104 13252
rect 11000 13172 11104 13188
rect 11000 13108 11020 13172
rect 11084 13108 11104 13172
rect 11000 13092 11104 13108
rect 11000 13028 11020 13092
rect 11084 13028 11104 13092
rect 11000 13012 11104 13028
rect 11000 12948 11020 13012
rect 11084 12948 11104 13012
rect 11000 12932 11104 12948
rect 11000 12868 11020 12932
rect 11084 12868 11104 12932
rect 11000 12852 11104 12868
rect 11000 12788 11020 12852
rect 11084 12788 11104 12852
rect 11000 12772 11104 12788
rect 11000 12708 11020 12772
rect 11084 12708 11104 12772
rect 11000 12692 11104 12708
rect 11000 12628 11020 12692
rect 11084 12628 11104 12692
rect 11000 12612 11104 12628
rect 11000 12548 11020 12612
rect 11084 12548 11104 12612
rect 11000 12532 11104 12548
rect 11000 12468 11020 12532
rect 11084 12468 11104 12532
rect 11000 12452 11104 12468
rect 11000 12388 11020 12452
rect 11084 12388 11104 12452
rect 11000 12372 11104 12388
rect 11000 12308 11020 12372
rect 11084 12308 11104 12372
rect 11000 12292 11104 12308
rect 11000 12228 11020 12292
rect 11084 12228 11104 12292
rect 11000 12212 11104 12228
rect 11000 12148 11020 12212
rect 11084 12148 11104 12212
rect 11000 12132 11104 12148
rect 11000 12068 11020 12132
rect 11084 12068 11104 12132
rect 11000 12052 11104 12068
rect 11000 11988 11020 12052
rect 11084 11988 11104 12052
rect 11000 11972 11104 11988
rect 11000 11908 11020 11972
rect 11084 11908 11104 11972
rect 11000 11892 11104 11908
rect 11000 11828 11020 11892
rect 11084 11828 11104 11892
rect 11000 11812 11104 11828
rect 11000 11748 11020 11812
rect 11084 11748 11104 11812
rect 11000 11732 11104 11748
rect 11000 11668 11020 11732
rect 11084 11668 11104 11732
rect 11000 11652 11104 11668
rect 11000 11588 11020 11652
rect 11084 11588 11104 11652
rect 11000 11572 11104 11588
rect 11000 11508 11020 11572
rect 11084 11508 11104 11572
rect 11000 11492 11104 11508
rect 11000 11428 11020 11492
rect 11084 11428 11104 11492
rect 11000 11412 11104 11428
rect 11000 11348 11020 11412
rect 11084 11348 11104 11412
rect 11000 11332 11104 11348
rect 11000 11268 11020 11332
rect 11084 11268 11104 11332
rect 11000 11252 11104 11268
rect 11000 11188 11020 11252
rect 11084 11188 11104 11252
rect 11000 11172 11104 11188
rect 11000 11108 11020 11172
rect 11084 11108 11104 11172
rect 11000 11092 11104 11108
rect 11000 11028 11020 11092
rect 11084 11028 11104 11092
rect 11000 11012 11104 11028
rect 11000 10948 11020 11012
rect 11084 10948 11104 11012
rect 11000 10932 11104 10948
rect 11000 10868 11020 10932
rect 11084 10868 11104 10932
rect 11000 10852 11104 10868
rect 5388 10492 5492 10788
rect -224 10412 -120 10428
rect -224 10348 -204 10412
rect -140 10348 -120 10412
rect -224 10332 -120 10348
rect -224 10268 -204 10332
rect -140 10268 -120 10332
rect -224 10252 -120 10268
rect -224 10188 -204 10252
rect -140 10188 -120 10252
rect -224 10172 -120 10188
rect -224 10108 -204 10172
rect -140 10108 -120 10172
rect -224 10092 -120 10108
rect -224 10028 -204 10092
rect -140 10028 -120 10092
rect -224 10012 -120 10028
rect -224 9948 -204 10012
rect -140 9948 -120 10012
rect -224 9932 -120 9948
rect -224 9868 -204 9932
rect -140 9868 -120 9932
rect -224 9852 -120 9868
rect -224 9788 -204 9852
rect -140 9788 -120 9852
rect -224 9772 -120 9788
rect -224 9708 -204 9772
rect -140 9708 -120 9772
rect -224 9692 -120 9708
rect -224 9628 -204 9692
rect -140 9628 -120 9692
rect -224 9612 -120 9628
rect -224 9548 -204 9612
rect -140 9548 -120 9612
rect -224 9532 -120 9548
rect -224 9468 -204 9532
rect -140 9468 -120 9532
rect -224 9452 -120 9468
rect -224 9388 -204 9452
rect -140 9388 -120 9452
rect -224 9372 -120 9388
rect -224 9308 -204 9372
rect -140 9308 -120 9372
rect -224 9292 -120 9308
rect -224 9228 -204 9292
rect -140 9228 -120 9292
rect -224 9212 -120 9228
rect -224 9148 -204 9212
rect -140 9148 -120 9212
rect -224 9132 -120 9148
rect -224 9068 -204 9132
rect -140 9068 -120 9132
rect -224 9052 -120 9068
rect -224 8988 -204 9052
rect -140 8988 -120 9052
rect -224 8972 -120 8988
rect -224 8908 -204 8972
rect -140 8908 -120 8972
rect -224 8892 -120 8908
rect -224 8828 -204 8892
rect -140 8828 -120 8892
rect -224 8812 -120 8828
rect -224 8748 -204 8812
rect -140 8748 -120 8812
rect -224 8732 -120 8748
rect -224 8668 -204 8732
rect -140 8668 -120 8732
rect -224 8652 -120 8668
rect -224 8588 -204 8652
rect -140 8588 -120 8652
rect -224 8572 -120 8588
rect -224 8508 -204 8572
rect -140 8508 -120 8572
rect -224 8492 -120 8508
rect -224 8428 -204 8492
rect -140 8428 -120 8492
rect -224 8412 -120 8428
rect -224 8348 -204 8412
rect -140 8348 -120 8412
rect -224 8332 -120 8348
rect -224 8268 -204 8332
rect -140 8268 -120 8332
rect -224 8252 -120 8268
rect -224 8188 -204 8252
rect -140 8188 -120 8252
rect -224 8172 -120 8188
rect -224 8108 -204 8172
rect -140 8108 -120 8172
rect -224 8092 -120 8108
rect -224 8028 -204 8092
rect -140 8028 -120 8092
rect -224 8012 -120 8028
rect -224 7948 -204 8012
rect -140 7948 -120 8012
rect -224 7932 -120 7948
rect -224 7868 -204 7932
rect -140 7868 -120 7932
rect -224 7852 -120 7868
rect -224 7788 -204 7852
rect -140 7788 -120 7852
rect -224 7772 -120 7788
rect -224 7708 -204 7772
rect -140 7708 -120 7772
rect -224 7692 -120 7708
rect -224 7628 -204 7692
rect -140 7628 -120 7692
rect -224 7612 -120 7628
rect -224 7548 -204 7612
rect -140 7548 -120 7612
rect -224 7532 -120 7548
rect -224 7468 -204 7532
rect -140 7468 -120 7532
rect -224 7452 -120 7468
rect -224 7388 -204 7452
rect -140 7388 -120 7452
rect -224 7372 -120 7388
rect -224 7308 -204 7372
rect -140 7308 -120 7372
rect -224 7292 -120 7308
rect -224 7228 -204 7292
rect -140 7228 -120 7292
rect -224 7212 -120 7228
rect -224 7148 -204 7212
rect -140 7148 -120 7212
rect -224 7132 -120 7148
rect -224 7068 -204 7132
rect -140 7068 -120 7132
rect -224 7052 -120 7068
rect -224 6988 -204 7052
rect -140 6988 -120 7052
rect -224 6972 -120 6988
rect -224 6908 -204 6972
rect -140 6908 -120 6972
rect -224 6892 -120 6908
rect -224 6828 -204 6892
rect -140 6828 -120 6892
rect -224 6812 -120 6828
rect -224 6748 -204 6812
rect -140 6748 -120 6812
rect -224 6732 -120 6748
rect -224 6668 -204 6732
rect -140 6668 -120 6732
rect -224 6652 -120 6668
rect -224 6588 -204 6652
rect -140 6588 -120 6652
rect -224 6572 -120 6588
rect -224 6508 -204 6572
rect -140 6508 -120 6572
rect -224 6492 -120 6508
rect -224 6428 -204 6492
rect -140 6428 -120 6492
rect -224 6412 -120 6428
rect -224 6348 -204 6412
rect -140 6348 -120 6412
rect -224 6332 -120 6348
rect -224 6268 -204 6332
rect -140 6268 -120 6332
rect -224 6252 -120 6268
rect -224 6188 -204 6252
rect -140 6188 -120 6252
rect -224 6172 -120 6188
rect -224 6108 -204 6172
rect -140 6108 -120 6172
rect -224 6092 -120 6108
rect -224 6028 -204 6092
rect -140 6028 -120 6092
rect -224 6012 -120 6028
rect -224 5948 -204 6012
rect -140 5948 -120 6012
rect -224 5932 -120 5948
rect -224 5868 -204 5932
rect -140 5868 -120 5932
rect -224 5852 -120 5868
rect -224 5788 -204 5852
rect -140 5788 -120 5852
rect -224 5772 -120 5788
rect -224 5708 -204 5772
rect -140 5708 -120 5772
rect -224 5692 -120 5708
rect -224 5628 -204 5692
rect -140 5628 -120 5692
rect -224 5612 -120 5628
rect -224 5548 -204 5612
rect -140 5548 -120 5612
rect -224 5532 -120 5548
rect -5836 5172 -5732 5468
rect -11448 5092 -11344 5108
rect -11448 5028 -11428 5092
rect -11364 5028 -11344 5092
rect -11448 5012 -11344 5028
rect -11448 4948 -11428 5012
rect -11364 4948 -11344 5012
rect -11448 4932 -11344 4948
rect -11448 4868 -11428 4932
rect -11364 4868 -11344 4932
rect -11448 4852 -11344 4868
rect -11448 4788 -11428 4852
rect -11364 4788 -11344 4852
rect -11448 4772 -11344 4788
rect -11448 4708 -11428 4772
rect -11364 4708 -11344 4772
rect -11448 4692 -11344 4708
rect -11448 4628 -11428 4692
rect -11364 4628 -11344 4692
rect -11448 4612 -11344 4628
rect -11448 4548 -11428 4612
rect -11364 4548 -11344 4612
rect -11448 4532 -11344 4548
rect -11448 4468 -11428 4532
rect -11364 4468 -11344 4532
rect -11448 4452 -11344 4468
rect -11448 4388 -11428 4452
rect -11364 4388 -11344 4452
rect -11448 4372 -11344 4388
rect -11448 4308 -11428 4372
rect -11364 4308 -11344 4372
rect -11448 4292 -11344 4308
rect -11448 4228 -11428 4292
rect -11364 4228 -11344 4292
rect -11448 4212 -11344 4228
rect -11448 4148 -11428 4212
rect -11364 4148 -11344 4212
rect -11448 4132 -11344 4148
rect -11448 4068 -11428 4132
rect -11364 4068 -11344 4132
rect -11448 4052 -11344 4068
rect -11448 3988 -11428 4052
rect -11364 3988 -11344 4052
rect -11448 3972 -11344 3988
rect -11448 3908 -11428 3972
rect -11364 3908 -11344 3972
rect -11448 3892 -11344 3908
rect -11448 3828 -11428 3892
rect -11364 3828 -11344 3892
rect -11448 3812 -11344 3828
rect -11448 3748 -11428 3812
rect -11364 3748 -11344 3812
rect -11448 3732 -11344 3748
rect -11448 3668 -11428 3732
rect -11364 3668 -11344 3732
rect -11448 3652 -11344 3668
rect -11448 3588 -11428 3652
rect -11364 3588 -11344 3652
rect -11448 3572 -11344 3588
rect -11448 3508 -11428 3572
rect -11364 3508 -11344 3572
rect -11448 3492 -11344 3508
rect -11448 3428 -11428 3492
rect -11364 3428 -11344 3492
rect -11448 3412 -11344 3428
rect -11448 3348 -11428 3412
rect -11364 3348 -11344 3412
rect -11448 3332 -11344 3348
rect -11448 3268 -11428 3332
rect -11364 3268 -11344 3332
rect -11448 3252 -11344 3268
rect -11448 3188 -11428 3252
rect -11364 3188 -11344 3252
rect -11448 3172 -11344 3188
rect -11448 3108 -11428 3172
rect -11364 3108 -11344 3172
rect -11448 3092 -11344 3108
rect -11448 3028 -11428 3092
rect -11364 3028 -11344 3092
rect -11448 3012 -11344 3028
rect -11448 2948 -11428 3012
rect -11364 2948 -11344 3012
rect -11448 2932 -11344 2948
rect -11448 2868 -11428 2932
rect -11364 2868 -11344 2932
rect -11448 2852 -11344 2868
rect -11448 2788 -11428 2852
rect -11364 2788 -11344 2852
rect -11448 2772 -11344 2788
rect -11448 2708 -11428 2772
rect -11364 2708 -11344 2772
rect -11448 2692 -11344 2708
rect -11448 2628 -11428 2692
rect -11364 2628 -11344 2692
rect -11448 2612 -11344 2628
rect -11448 2548 -11428 2612
rect -11364 2548 -11344 2612
rect -11448 2532 -11344 2548
rect -11448 2468 -11428 2532
rect -11364 2468 -11344 2532
rect -11448 2452 -11344 2468
rect -11448 2388 -11428 2452
rect -11364 2388 -11344 2452
rect -11448 2372 -11344 2388
rect -11448 2308 -11428 2372
rect -11364 2308 -11344 2372
rect -11448 2292 -11344 2308
rect -11448 2228 -11428 2292
rect -11364 2228 -11344 2292
rect -11448 2212 -11344 2228
rect -11448 2148 -11428 2212
rect -11364 2148 -11344 2212
rect -11448 2132 -11344 2148
rect -11448 2068 -11428 2132
rect -11364 2068 -11344 2132
rect -11448 2052 -11344 2068
rect -11448 1988 -11428 2052
rect -11364 1988 -11344 2052
rect -11448 1972 -11344 1988
rect -11448 1908 -11428 1972
rect -11364 1908 -11344 1972
rect -11448 1892 -11344 1908
rect -11448 1828 -11428 1892
rect -11364 1828 -11344 1892
rect -11448 1812 -11344 1828
rect -11448 1748 -11428 1812
rect -11364 1748 -11344 1812
rect -11448 1732 -11344 1748
rect -11448 1668 -11428 1732
rect -11364 1668 -11344 1732
rect -11448 1652 -11344 1668
rect -11448 1588 -11428 1652
rect -11364 1588 -11344 1652
rect -11448 1572 -11344 1588
rect -11448 1508 -11428 1572
rect -11364 1508 -11344 1572
rect -11448 1492 -11344 1508
rect -11448 1428 -11428 1492
rect -11364 1428 -11344 1492
rect -11448 1412 -11344 1428
rect -11448 1348 -11428 1412
rect -11364 1348 -11344 1412
rect -11448 1332 -11344 1348
rect -11448 1268 -11428 1332
rect -11364 1268 -11344 1332
rect -11448 1252 -11344 1268
rect -11448 1188 -11428 1252
rect -11364 1188 -11344 1252
rect -11448 1172 -11344 1188
rect -11448 1108 -11428 1172
rect -11364 1108 -11344 1172
rect -11448 1092 -11344 1108
rect -11448 1028 -11428 1092
rect -11364 1028 -11344 1092
rect -11448 1012 -11344 1028
rect -11448 948 -11428 1012
rect -11364 948 -11344 1012
rect -11448 932 -11344 948
rect -11448 868 -11428 932
rect -11364 868 -11344 932
rect -11448 852 -11344 868
rect -11448 788 -11428 852
rect -11364 788 -11344 852
rect -11448 772 -11344 788
rect -11448 708 -11428 772
rect -11364 708 -11344 772
rect -11448 692 -11344 708
rect -11448 628 -11428 692
rect -11364 628 -11344 692
rect -11448 612 -11344 628
rect -11448 548 -11428 612
rect -11364 548 -11344 612
rect -11448 532 -11344 548
rect -11448 468 -11428 532
rect -11364 468 -11344 532
rect -11448 452 -11344 468
rect -11448 388 -11428 452
rect -11364 388 -11344 452
rect -11448 372 -11344 388
rect -11448 308 -11428 372
rect -11364 308 -11344 372
rect -11448 292 -11344 308
rect -11448 228 -11428 292
rect -11364 228 -11344 292
rect -11448 212 -11344 228
rect -17060 -148 -16956 148
rect -22672 -228 -22568 -212
rect -22672 -292 -22652 -228
rect -22588 -292 -22568 -228
rect -22672 -308 -22568 -292
rect -22672 -372 -22652 -308
rect -22588 -372 -22568 -308
rect -22672 -388 -22568 -372
rect -22672 -452 -22652 -388
rect -22588 -452 -22568 -388
rect -22672 -468 -22568 -452
rect -22672 -532 -22652 -468
rect -22588 -532 -22568 -468
rect -22672 -548 -22568 -532
rect -22672 -612 -22652 -548
rect -22588 -612 -22568 -548
rect -22672 -628 -22568 -612
rect -22672 -692 -22652 -628
rect -22588 -692 -22568 -628
rect -22672 -708 -22568 -692
rect -22672 -772 -22652 -708
rect -22588 -772 -22568 -708
rect -22672 -788 -22568 -772
rect -22672 -852 -22652 -788
rect -22588 -852 -22568 -788
rect -22672 -868 -22568 -852
rect -22672 -932 -22652 -868
rect -22588 -932 -22568 -868
rect -22672 -948 -22568 -932
rect -22672 -1012 -22652 -948
rect -22588 -1012 -22568 -948
rect -22672 -1028 -22568 -1012
rect -22672 -1092 -22652 -1028
rect -22588 -1092 -22568 -1028
rect -22672 -1108 -22568 -1092
rect -22672 -1172 -22652 -1108
rect -22588 -1172 -22568 -1108
rect -22672 -1188 -22568 -1172
rect -22672 -1252 -22652 -1188
rect -22588 -1252 -22568 -1188
rect -22672 -1268 -22568 -1252
rect -22672 -1332 -22652 -1268
rect -22588 -1332 -22568 -1268
rect -22672 -1348 -22568 -1332
rect -22672 -1412 -22652 -1348
rect -22588 -1412 -22568 -1348
rect -22672 -1428 -22568 -1412
rect -22672 -1492 -22652 -1428
rect -22588 -1492 -22568 -1428
rect -22672 -1508 -22568 -1492
rect -22672 -1572 -22652 -1508
rect -22588 -1572 -22568 -1508
rect -22672 -1588 -22568 -1572
rect -22672 -1652 -22652 -1588
rect -22588 -1652 -22568 -1588
rect -22672 -1668 -22568 -1652
rect -22672 -1732 -22652 -1668
rect -22588 -1732 -22568 -1668
rect -22672 -1748 -22568 -1732
rect -22672 -1812 -22652 -1748
rect -22588 -1812 -22568 -1748
rect -22672 -1828 -22568 -1812
rect -22672 -1892 -22652 -1828
rect -22588 -1892 -22568 -1828
rect -22672 -1908 -22568 -1892
rect -22672 -1972 -22652 -1908
rect -22588 -1972 -22568 -1908
rect -22672 -1988 -22568 -1972
rect -22672 -2052 -22652 -1988
rect -22588 -2052 -22568 -1988
rect -22672 -2068 -22568 -2052
rect -22672 -2132 -22652 -2068
rect -22588 -2132 -22568 -2068
rect -22672 -2148 -22568 -2132
rect -22672 -2212 -22652 -2148
rect -22588 -2212 -22568 -2148
rect -22672 -2228 -22568 -2212
rect -22672 -2292 -22652 -2228
rect -22588 -2292 -22568 -2228
rect -22672 -2308 -22568 -2292
rect -22672 -2372 -22652 -2308
rect -22588 -2372 -22568 -2308
rect -22672 -2388 -22568 -2372
rect -22672 -2452 -22652 -2388
rect -22588 -2452 -22568 -2388
rect -22672 -2468 -22568 -2452
rect -22672 -2532 -22652 -2468
rect -22588 -2532 -22568 -2468
rect -22672 -2548 -22568 -2532
rect -22672 -2612 -22652 -2548
rect -22588 -2612 -22568 -2548
rect -22672 -2628 -22568 -2612
rect -22672 -2692 -22652 -2628
rect -22588 -2692 -22568 -2628
rect -22672 -2708 -22568 -2692
rect -22672 -2772 -22652 -2708
rect -22588 -2772 -22568 -2708
rect -22672 -2788 -22568 -2772
rect -22672 -2852 -22652 -2788
rect -22588 -2852 -22568 -2788
rect -22672 -2868 -22568 -2852
rect -22672 -2932 -22652 -2868
rect -22588 -2932 -22568 -2868
rect -22672 -2948 -22568 -2932
rect -22672 -3012 -22652 -2948
rect -22588 -3012 -22568 -2948
rect -22672 -3028 -22568 -3012
rect -22672 -3092 -22652 -3028
rect -22588 -3092 -22568 -3028
rect -22672 -3108 -22568 -3092
rect -22672 -3172 -22652 -3108
rect -22588 -3172 -22568 -3108
rect -22672 -3188 -22568 -3172
rect -22672 -3252 -22652 -3188
rect -22588 -3252 -22568 -3188
rect -22672 -3268 -22568 -3252
rect -22672 -3332 -22652 -3268
rect -22588 -3332 -22568 -3268
rect -22672 -3348 -22568 -3332
rect -22672 -3412 -22652 -3348
rect -22588 -3412 -22568 -3348
rect -22672 -3428 -22568 -3412
rect -22672 -3492 -22652 -3428
rect -22588 -3492 -22568 -3428
rect -22672 -3508 -22568 -3492
rect -22672 -3572 -22652 -3508
rect -22588 -3572 -22568 -3508
rect -22672 -3588 -22568 -3572
rect -22672 -3652 -22652 -3588
rect -22588 -3652 -22568 -3588
rect -22672 -3668 -22568 -3652
rect -22672 -3732 -22652 -3668
rect -22588 -3732 -22568 -3668
rect -22672 -3748 -22568 -3732
rect -22672 -3812 -22652 -3748
rect -22588 -3812 -22568 -3748
rect -22672 -3828 -22568 -3812
rect -22672 -3892 -22652 -3828
rect -22588 -3892 -22568 -3828
rect -22672 -3908 -22568 -3892
rect -22672 -3972 -22652 -3908
rect -22588 -3972 -22568 -3908
rect -22672 -3988 -22568 -3972
rect -22672 -4052 -22652 -3988
rect -22588 -4052 -22568 -3988
rect -22672 -4068 -22568 -4052
rect -22672 -4132 -22652 -4068
rect -22588 -4132 -22568 -4068
rect -22672 -4148 -22568 -4132
rect -22672 -4212 -22652 -4148
rect -22588 -4212 -22568 -4148
rect -22672 -4228 -22568 -4212
rect -22672 -4292 -22652 -4228
rect -22588 -4292 -22568 -4228
rect -22672 -4308 -22568 -4292
rect -22672 -4372 -22652 -4308
rect -22588 -4372 -22568 -4308
rect -22672 -4388 -22568 -4372
rect -22672 -4452 -22652 -4388
rect -22588 -4452 -22568 -4388
rect -22672 -4468 -22568 -4452
rect -22672 -4532 -22652 -4468
rect -22588 -4532 -22568 -4468
rect -22672 -4548 -22568 -4532
rect -22672 -4612 -22652 -4548
rect -22588 -4612 -22568 -4548
rect -22672 -4628 -22568 -4612
rect -22672 -4692 -22652 -4628
rect -22588 -4692 -22568 -4628
rect -22672 -4708 -22568 -4692
rect -22672 -4772 -22652 -4708
rect -22588 -4772 -22568 -4708
rect -22672 -4788 -22568 -4772
rect -22672 -4852 -22652 -4788
rect -22588 -4852 -22568 -4788
rect -22672 -4868 -22568 -4852
rect -22672 -4932 -22652 -4868
rect -22588 -4932 -22568 -4868
rect -22672 -4948 -22568 -4932
rect -22672 -5012 -22652 -4948
rect -22588 -5012 -22568 -4948
rect -22672 -5028 -22568 -5012
rect -22672 -5092 -22652 -5028
rect -22588 -5092 -22568 -5028
rect -22672 -5108 -22568 -5092
rect -28284 -5468 -28180 -5172
rect -33896 -5548 -33792 -5532
rect -33896 -5612 -33876 -5548
rect -33812 -5612 -33792 -5548
rect -33896 -5628 -33792 -5612
rect -33896 -5692 -33876 -5628
rect -33812 -5692 -33792 -5628
rect -33896 -5708 -33792 -5692
rect -33896 -5772 -33876 -5708
rect -33812 -5772 -33792 -5708
rect -33896 -5788 -33792 -5772
rect -33896 -5852 -33876 -5788
rect -33812 -5852 -33792 -5788
rect -33896 -5868 -33792 -5852
rect -33896 -5932 -33876 -5868
rect -33812 -5932 -33792 -5868
rect -33896 -5948 -33792 -5932
rect -33896 -6012 -33876 -5948
rect -33812 -6012 -33792 -5948
rect -33896 -6028 -33792 -6012
rect -33896 -6092 -33876 -6028
rect -33812 -6092 -33792 -6028
rect -33896 -6108 -33792 -6092
rect -33896 -6172 -33876 -6108
rect -33812 -6172 -33792 -6108
rect -33896 -6188 -33792 -6172
rect -33896 -6252 -33876 -6188
rect -33812 -6252 -33792 -6188
rect -33896 -6268 -33792 -6252
rect -33896 -6332 -33876 -6268
rect -33812 -6332 -33792 -6268
rect -33896 -6348 -33792 -6332
rect -33896 -6412 -33876 -6348
rect -33812 -6412 -33792 -6348
rect -33896 -6428 -33792 -6412
rect -33896 -6492 -33876 -6428
rect -33812 -6492 -33792 -6428
rect -33896 -6508 -33792 -6492
rect -33896 -6572 -33876 -6508
rect -33812 -6572 -33792 -6508
rect -33896 -6588 -33792 -6572
rect -33896 -6652 -33876 -6588
rect -33812 -6652 -33792 -6588
rect -33896 -6668 -33792 -6652
rect -33896 -6732 -33876 -6668
rect -33812 -6732 -33792 -6668
rect -33896 -6748 -33792 -6732
rect -33896 -6812 -33876 -6748
rect -33812 -6812 -33792 -6748
rect -33896 -6828 -33792 -6812
rect -33896 -6892 -33876 -6828
rect -33812 -6892 -33792 -6828
rect -33896 -6908 -33792 -6892
rect -33896 -6972 -33876 -6908
rect -33812 -6972 -33792 -6908
rect -33896 -6988 -33792 -6972
rect -33896 -7052 -33876 -6988
rect -33812 -7052 -33792 -6988
rect -33896 -7068 -33792 -7052
rect -33896 -7132 -33876 -7068
rect -33812 -7132 -33792 -7068
rect -33896 -7148 -33792 -7132
rect -33896 -7212 -33876 -7148
rect -33812 -7212 -33792 -7148
rect -33896 -7228 -33792 -7212
rect -33896 -7292 -33876 -7228
rect -33812 -7292 -33792 -7228
rect -33896 -7308 -33792 -7292
rect -33896 -7372 -33876 -7308
rect -33812 -7372 -33792 -7308
rect -33896 -7388 -33792 -7372
rect -33896 -7452 -33876 -7388
rect -33812 -7452 -33792 -7388
rect -33896 -7468 -33792 -7452
rect -33896 -7532 -33876 -7468
rect -33812 -7532 -33792 -7468
rect -33896 -7548 -33792 -7532
rect -33896 -7612 -33876 -7548
rect -33812 -7612 -33792 -7548
rect -33896 -7628 -33792 -7612
rect -33896 -7692 -33876 -7628
rect -33812 -7692 -33792 -7628
rect -33896 -7708 -33792 -7692
rect -33896 -7772 -33876 -7708
rect -33812 -7772 -33792 -7708
rect -33896 -7788 -33792 -7772
rect -33896 -7852 -33876 -7788
rect -33812 -7852 -33792 -7788
rect -33896 -7868 -33792 -7852
rect -33896 -7932 -33876 -7868
rect -33812 -7932 -33792 -7868
rect -33896 -7948 -33792 -7932
rect -33896 -8012 -33876 -7948
rect -33812 -8012 -33792 -7948
rect -33896 -8028 -33792 -8012
rect -33896 -8092 -33876 -8028
rect -33812 -8092 -33792 -8028
rect -33896 -8108 -33792 -8092
rect -33896 -8172 -33876 -8108
rect -33812 -8172 -33792 -8108
rect -33896 -8188 -33792 -8172
rect -33896 -8252 -33876 -8188
rect -33812 -8252 -33792 -8188
rect -33896 -8268 -33792 -8252
rect -33896 -8332 -33876 -8268
rect -33812 -8332 -33792 -8268
rect -33896 -8348 -33792 -8332
rect -33896 -8412 -33876 -8348
rect -33812 -8412 -33792 -8348
rect -33896 -8428 -33792 -8412
rect -33896 -8492 -33876 -8428
rect -33812 -8492 -33792 -8428
rect -33896 -8508 -33792 -8492
rect -33896 -8572 -33876 -8508
rect -33812 -8572 -33792 -8508
rect -33896 -8588 -33792 -8572
rect -33896 -8652 -33876 -8588
rect -33812 -8652 -33792 -8588
rect -33896 -8668 -33792 -8652
rect -33896 -8732 -33876 -8668
rect -33812 -8732 -33792 -8668
rect -33896 -8748 -33792 -8732
rect -33896 -8812 -33876 -8748
rect -33812 -8812 -33792 -8748
rect -33896 -8828 -33792 -8812
rect -33896 -8892 -33876 -8828
rect -33812 -8892 -33792 -8828
rect -33896 -8908 -33792 -8892
rect -33896 -8972 -33876 -8908
rect -33812 -8972 -33792 -8908
rect -33896 -8988 -33792 -8972
rect -33896 -9052 -33876 -8988
rect -33812 -9052 -33792 -8988
rect -33896 -9068 -33792 -9052
rect -33896 -9132 -33876 -9068
rect -33812 -9132 -33792 -9068
rect -33896 -9148 -33792 -9132
rect -33896 -9212 -33876 -9148
rect -33812 -9212 -33792 -9148
rect -33896 -9228 -33792 -9212
rect -33896 -9292 -33876 -9228
rect -33812 -9292 -33792 -9228
rect -33896 -9308 -33792 -9292
rect -33896 -9372 -33876 -9308
rect -33812 -9372 -33792 -9308
rect -33896 -9388 -33792 -9372
rect -33896 -9452 -33876 -9388
rect -33812 -9452 -33792 -9388
rect -33896 -9468 -33792 -9452
rect -33896 -9532 -33876 -9468
rect -33812 -9532 -33792 -9468
rect -33896 -9548 -33792 -9532
rect -33896 -9612 -33876 -9548
rect -33812 -9612 -33792 -9548
rect -33896 -9628 -33792 -9612
rect -33896 -9692 -33876 -9628
rect -33812 -9692 -33792 -9628
rect -33896 -9708 -33792 -9692
rect -33896 -9772 -33876 -9708
rect -33812 -9772 -33792 -9708
rect -33896 -9788 -33792 -9772
rect -33896 -9852 -33876 -9788
rect -33812 -9852 -33792 -9788
rect -33896 -9868 -33792 -9852
rect -33896 -9932 -33876 -9868
rect -33812 -9932 -33792 -9868
rect -33896 -9948 -33792 -9932
rect -33896 -10012 -33876 -9948
rect -33812 -10012 -33792 -9948
rect -33896 -10028 -33792 -10012
rect -33896 -10092 -33876 -10028
rect -33812 -10092 -33792 -10028
rect -33896 -10108 -33792 -10092
rect -33896 -10172 -33876 -10108
rect -33812 -10172 -33792 -10108
rect -33896 -10188 -33792 -10172
rect -33896 -10252 -33876 -10188
rect -33812 -10252 -33792 -10188
rect -33896 -10268 -33792 -10252
rect -33896 -10332 -33876 -10268
rect -33812 -10332 -33792 -10268
rect -33896 -10348 -33792 -10332
rect -33896 -10412 -33876 -10348
rect -33812 -10412 -33792 -10348
rect -33896 -10428 -33792 -10412
rect -36676 -10839 -36572 -10441
rect -33896 -10492 -33876 -10428
rect -33812 -10492 -33792 -10428
rect -33473 -5548 -28551 -5519
rect -33473 -10412 -33444 -5548
rect -28580 -10412 -28551 -5548
rect -33473 -10441 -28551 -10412
rect -28284 -5532 -28264 -5468
rect -28200 -5532 -28180 -5468
rect -25452 -5519 -25348 -5121
rect -22672 -5172 -22652 -5108
rect -22588 -5172 -22568 -5108
rect -22249 -228 -17327 -199
rect -22249 -5092 -22220 -228
rect -17356 -5092 -17327 -228
rect -22249 -5121 -17327 -5092
rect -17060 -212 -17040 -148
rect -16976 -212 -16956 -148
rect -14228 -199 -14124 199
rect -11448 148 -11428 212
rect -11364 148 -11344 212
rect -11025 5092 -6103 5121
rect -11025 228 -10996 5092
rect -6132 228 -6103 5092
rect -11025 199 -6103 228
rect -5836 5108 -5816 5172
rect -5752 5108 -5732 5172
rect -3004 5121 -2900 5519
rect -224 5468 -204 5532
rect -140 5468 -120 5532
rect 199 10412 5121 10441
rect 199 5548 228 10412
rect 5092 5548 5121 10412
rect 199 5519 5121 5548
rect 5388 10428 5408 10492
rect 5472 10428 5492 10492
rect 8220 10441 8324 10839
rect 11000 10788 11020 10852
rect 11084 10788 11104 10852
rect 11423 15732 16345 15761
rect 11423 10868 11452 15732
rect 16316 10868 16345 15732
rect 11423 10839 16345 10868
rect 16612 15748 16632 15812
rect 16696 15748 16716 15812
rect 19444 15761 19548 16159
rect 22224 16108 22244 16172
rect 22308 16108 22328 16172
rect 22647 21052 27569 21081
rect 22647 16188 22676 21052
rect 27540 16188 27569 21052
rect 22647 16159 27569 16188
rect 27836 21068 27856 21132
rect 27920 21068 27940 21132
rect 30668 21081 30772 21479
rect 33448 21428 33468 21492
rect 33532 21428 33552 21492
rect 33871 26372 38793 26401
rect 33871 21508 33900 26372
rect 38764 21508 38793 26372
rect 33871 21479 38793 21508
rect 39060 26388 39080 26452
rect 39144 26388 39164 26452
rect 39060 26372 39164 26388
rect 39060 26308 39080 26372
rect 39144 26308 39164 26372
rect 39060 26292 39164 26308
rect 39060 26228 39080 26292
rect 39144 26228 39164 26292
rect 39060 26212 39164 26228
rect 39060 26148 39080 26212
rect 39144 26148 39164 26212
rect 39060 26132 39164 26148
rect 39060 26068 39080 26132
rect 39144 26068 39164 26132
rect 39060 26052 39164 26068
rect 39060 25988 39080 26052
rect 39144 25988 39164 26052
rect 39060 25972 39164 25988
rect 39060 25908 39080 25972
rect 39144 25908 39164 25972
rect 39060 25892 39164 25908
rect 39060 25828 39080 25892
rect 39144 25828 39164 25892
rect 39060 25812 39164 25828
rect 39060 25748 39080 25812
rect 39144 25748 39164 25812
rect 39060 25732 39164 25748
rect 39060 25668 39080 25732
rect 39144 25668 39164 25732
rect 39060 25652 39164 25668
rect 39060 25588 39080 25652
rect 39144 25588 39164 25652
rect 39060 25572 39164 25588
rect 39060 25508 39080 25572
rect 39144 25508 39164 25572
rect 39060 25492 39164 25508
rect 39060 25428 39080 25492
rect 39144 25428 39164 25492
rect 39060 25412 39164 25428
rect 39060 25348 39080 25412
rect 39144 25348 39164 25412
rect 39060 25332 39164 25348
rect 39060 25268 39080 25332
rect 39144 25268 39164 25332
rect 39060 25252 39164 25268
rect 39060 25188 39080 25252
rect 39144 25188 39164 25252
rect 39060 25172 39164 25188
rect 39060 25108 39080 25172
rect 39144 25108 39164 25172
rect 39060 25092 39164 25108
rect 39060 25028 39080 25092
rect 39144 25028 39164 25092
rect 39060 25012 39164 25028
rect 39060 24948 39080 25012
rect 39144 24948 39164 25012
rect 39060 24932 39164 24948
rect 39060 24868 39080 24932
rect 39144 24868 39164 24932
rect 39060 24852 39164 24868
rect 39060 24788 39080 24852
rect 39144 24788 39164 24852
rect 39060 24772 39164 24788
rect 39060 24708 39080 24772
rect 39144 24708 39164 24772
rect 39060 24692 39164 24708
rect 39060 24628 39080 24692
rect 39144 24628 39164 24692
rect 39060 24612 39164 24628
rect 39060 24548 39080 24612
rect 39144 24548 39164 24612
rect 39060 24532 39164 24548
rect 39060 24468 39080 24532
rect 39144 24468 39164 24532
rect 39060 24452 39164 24468
rect 39060 24388 39080 24452
rect 39144 24388 39164 24452
rect 39060 24372 39164 24388
rect 39060 24308 39080 24372
rect 39144 24308 39164 24372
rect 39060 24292 39164 24308
rect 39060 24228 39080 24292
rect 39144 24228 39164 24292
rect 39060 24212 39164 24228
rect 39060 24148 39080 24212
rect 39144 24148 39164 24212
rect 39060 24132 39164 24148
rect 39060 24068 39080 24132
rect 39144 24068 39164 24132
rect 39060 24052 39164 24068
rect 39060 23988 39080 24052
rect 39144 23988 39164 24052
rect 39060 23972 39164 23988
rect 39060 23908 39080 23972
rect 39144 23908 39164 23972
rect 39060 23892 39164 23908
rect 39060 23828 39080 23892
rect 39144 23828 39164 23892
rect 39060 23812 39164 23828
rect 39060 23748 39080 23812
rect 39144 23748 39164 23812
rect 39060 23732 39164 23748
rect 39060 23668 39080 23732
rect 39144 23668 39164 23732
rect 39060 23652 39164 23668
rect 39060 23588 39080 23652
rect 39144 23588 39164 23652
rect 39060 23572 39164 23588
rect 39060 23508 39080 23572
rect 39144 23508 39164 23572
rect 39060 23492 39164 23508
rect 39060 23428 39080 23492
rect 39144 23428 39164 23492
rect 39060 23412 39164 23428
rect 39060 23348 39080 23412
rect 39144 23348 39164 23412
rect 39060 23332 39164 23348
rect 39060 23268 39080 23332
rect 39144 23268 39164 23332
rect 39060 23252 39164 23268
rect 39060 23188 39080 23252
rect 39144 23188 39164 23252
rect 39060 23172 39164 23188
rect 39060 23108 39080 23172
rect 39144 23108 39164 23172
rect 39060 23092 39164 23108
rect 39060 23028 39080 23092
rect 39144 23028 39164 23092
rect 39060 23012 39164 23028
rect 39060 22948 39080 23012
rect 39144 22948 39164 23012
rect 39060 22932 39164 22948
rect 39060 22868 39080 22932
rect 39144 22868 39164 22932
rect 39060 22852 39164 22868
rect 39060 22788 39080 22852
rect 39144 22788 39164 22852
rect 39060 22772 39164 22788
rect 39060 22708 39080 22772
rect 39144 22708 39164 22772
rect 39060 22692 39164 22708
rect 39060 22628 39080 22692
rect 39144 22628 39164 22692
rect 39060 22612 39164 22628
rect 39060 22548 39080 22612
rect 39144 22548 39164 22612
rect 39060 22532 39164 22548
rect 39060 22468 39080 22532
rect 39144 22468 39164 22532
rect 39060 22452 39164 22468
rect 39060 22388 39080 22452
rect 39144 22388 39164 22452
rect 39060 22372 39164 22388
rect 39060 22308 39080 22372
rect 39144 22308 39164 22372
rect 39060 22292 39164 22308
rect 39060 22228 39080 22292
rect 39144 22228 39164 22292
rect 39060 22212 39164 22228
rect 39060 22148 39080 22212
rect 39144 22148 39164 22212
rect 39060 22132 39164 22148
rect 39060 22068 39080 22132
rect 39144 22068 39164 22132
rect 39060 22052 39164 22068
rect 39060 21988 39080 22052
rect 39144 21988 39164 22052
rect 39060 21972 39164 21988
rect 39060 21908 39080 21972
rect 39144 21908 39164 21972
rect 39060 21892 39164 21908
rect 39060 21828 39080 21892
rect 39144 21828 39164 21892
rect 39060 21812 39164 21828
rect 39060 21748 39080 21812
rect 39144 21748 39164 21812
rect 39060 21732 39164 21748
rect 39060 21668 39080 21732
rect 39144 21668 39164 21732
rect 39060 21652 39164 21668
rect 39060 21588 39080 21652
rect 39144 21588 39164 21652
rect 39060 21572 39164 21588
rect 39060 21508 39080 21572
rect 39144 21508 39164 21572
rect 39060 21492 39164 21508
rect 33448 21132 33552 21428
rect 27836 21052 27940 21068
rect 27836 20988 27856 21052
rect 27920 20988 27940 21052
rect 27836 20972 27940 20988
rect 27836 20908 27856 20972
rect 27920 20908 27940 20972
rect 27836 20892 27940 20908
rect 27836 20828 27856 20892
rect 27920 20828 27940 20892
rect 27836 20812 27940 20828
rect 27836 20748 27856 20812
rect 27920 20748 27940 20812
rect 27836 20732 27940 20748
rect 27836 20668 27856 20732
rect 27920 20668 27940 20732
rect 27836 20652 27940 20668
rect 27836 20588 27856 20652
rect 27920 20588 27940 20652
rect 27836 20572 27940 20588
rect 27836 20508 27856 20572
rect 27920 20508 27940 20572
rect 27836 20492 27940 20508
rect 27836 20428 27856 20492
rect 27920 20428 27940 20492
rect 27836 20412 27940 20428
rect 27836 20348 27856 20412
rect 27920 20348 27940 20412
rect 27836 20332 27940 20348
rect 27836 20268 27856 20332
rect 27920 20268 27940 20332
rect 27836 20252 27940 20268
rect 27836 20188 27856 20252
rect 27920 20188 27940 20252
rect 27836 20172 27940 20188
rect 27836 20108 27856 20172
rect 27920 20108 27940 20172
rect 27836 20092 27940 20108
rect 27836 20028 27856 20092
rect 27920 20028 27940 20092
rect 27836 20012 27940 20028
rect 27836 19948 27856 20012
rect 27920 19948 27940 20012
rect 27836 19932 27940 19948
rect 27836 19868 27856 19932
rect 27920 19868 27940 19932
rect 27836 19852 27940 19868
rect 27836 19788 27856 19852
rect 27920 19788 27940 19852
rect 27836 19772 27940 19788
rect 27836 19708 27856 19772
rect 27920 19708 27940 19772
rect 27836 19692 27940 19708
rect 27836 19628 27856 19692
rect 27920 19628 27940 19692
rect 27836 19612 27940 19628
rect 27836 19548 27856 19612
rect 27920 19548 27940 19612
rect 27836 19532 27940 19548
rect 27836 19468 27856 19532
rect 27920 19468 27940 19532
rect 27836 19452 27940 19468
rect 27836 19388 27856 19452
rect 27920 19388 27940 19452
rect 27836 19372 27940 19388
rect 27836 19308 27856 19372
rect 27920 19308 27940 19372
rect 27836 19292 27940 19308
rect 27836 19228 27856 19292
rect 27920 19228 27940 19292
rect 27836 19212 27940 19228
rect 27836 19148 27856 19212
rect 27920 19148 27940 19212
rect 27836 19132 27940 19148
rect 27836 19068 27856 19132
rect 27920 19068 27940 19132
rect 27836 19052 27940 19068
rect 27836 18988 27856 19052
rect 27920 18988 27940 19052
rect 27836 18972 27940 18988
rect 27836 18908 27856 18972
rect 27920 18908 27940 18972
rect 27836 18892 27940 18908
rect 27836 18828 27856 18892
rect 27920 18828 27940 18892
rect 27836 18812 27940 18828
rect 27836 18748 27856 18812
rect 27920 18748 27940 18812
rect 27836 18732 27940 18748
rect 27836 18668 27856 18732
rect 27920 18668 27940 18732
rect 27836 18652 27940 18668
rect 27836 18588 27856 18652
rect 27920 18588 27940 18652
rect 27836 18572 27940 18588
rect 27836 18508 27856 18572
rect 27920 18508 27940 18572
rect 27836 18492 27940 18508
rect 27836 18428 27856 18492
rect 27920 18428 27940 18492
rect 27836 18412 27940 18428
rect 27836 18348 27856 18412
rect 27920 18348 27940 18412
rect 27836 18332 27940 18348
rect 27836 18268 27856 18332
rect 27920 18268 27940 18332
rect 27836 18252 27940 18268
rect 27836 18188 27856 18252
rect 27920 18188 27940 18252
rect 27836 18172 27940 18188
rect 27836 18108 27856 18172
rect 27920 18108 27940 18172
rect 27836 18092 27940 18108
rect 27836 18028 27856 18092
rect 27920 18028 27940 18092
rect 27836 18012 27940 18028
rect 27836 17948 27856 18012
rect 27920 17948 27940 18012
rect 27836 17932 27940 17948
rect 27836 17868 27856 17932
rect 27920 17868 27940 17932
rect 27836 17852 27940 17868
rect 27836 17788 27856 17852
rect 27920 17788 27940 17852
rect 27836 17772 27940 17788
rect 27836 17708 27856 17772
rect 27920 17708 27940 17772
rect 27836 17692 27940 17708
rect 27836 17628 27856 17692
rect 27920 17628 27940 17692
rect 27836 17612 27940 17628
rect 27836 17548 27856 17612
rect 27920 17548 27940 17612
rect 27836 17532 27940 17548
rect 27836 17468 27856 17532
rect 27920 17468 27940 17532
rect 27836 17452 27940 17468
rect 27836 17388 27856 17452
rect 27920 17388 27940 17452
rect 27836 17372 27940 17388
rect 27836 17308 27856 17372
rect 27920 17308 27940 17372
rect 27836 17292 27940 17308
rect 27836 17228 27856 17292
rect 27920 17228 27940 17292
rect 27836 17212 27940 17228
rect 27836 17148 27856 17212
rect 27920 17148 27940 17212
rect 27836 17132 27940 17148
rect 27836 17068 27856 17132
rect 27920 17068 27940 17132
rect 27836 17052 27940 17068
rect 27836 16988 27856 17052
rect 27920 16988 27940 17052
rect 27836 16972 27940 16988
rect 27836 16908 27856 16972
rect 27920 16908 27940 16972
rect 27836 16892 27940 16908
rect 27836 16828 27856 16892
rect 27920 16828 27940 16892
rect 27836 16812 27940 16828
rect 27836 16748 27856 16812
rect 27920 16748 27940 16812
rect 27836 16732 27940 16748
rect 27836 16668 27856 16732
rect 27920 16668 27940 16732
rect 27836 16652 27940 16668
rect 27836 16588 27856 16652
rect 27920 16588 27940 16652
rect 27836 16572 27940 16588
rect 27836 16508 27856 16572
rect 27920 16508 27940 16572
rect 27836 16492 27940 16508
rect 27836 16428 27856 16492
rect 27920 16428 27940 16492
rect 27836 16412 27940 16428
rect 27836 16348 27856 16412
rect 27920 16348 27940 16412
rect 27836 16332 27940 16348
rect 27836 16268 27856 16332
rect 27920 16268 27940 16332
rect 27836 16252 27940 16268
rect 27836 16188 27856 16252
rect 27920 16188 27940 16252
rect 27836 16172 27940 16188
rect 22224 15812 22328 16108
rect 16612 15732 16716 15748
rect 16612 15668 16632 15732
rect 16696 15668 16716 15732
rect 16612 15652 16716 15668
rect 16612 15588 16632 15652
rect 16696 15588 16716 15652
rect 16612 15572 16716 15588
rect 16612 15508 16632 15572
rect 16696 15508 16716 15572
rect 16612 15492 16716 15508
rect 16612 15428 16632 15492
rect 16696 15428 16716 15492
rect 16612 15412 16716 15428
rect 16612 15348 16632 15412
rect 16696 15348 16716 15412
rect 16612 15332 16716 15348
rect 16612 15268 16632 15332
rect 16696 15268 16716 15332
rect 16612 15252 16716 15268
rect 16612 15188 16632 15252
rect 16696 15188 16716 15252
rect 16612 15172 16716 15188
rect 16612 15108 16632 15172
rect 16696 15108 16716 15172
rect 16612 15092 16716 15108
rect 16612 15028 16632 15092
rect 16696 15028 16716 15092
rect 16612 15012 16716 15028
rect 16612 14948 16632 15012
rect 16696 14948 16716 15012
rect 16612 14932 16716 14948
rect 16612 14868 16632 14932
rect 16696 14868 16716 14932
rect 16612 14852 16716 14868
rect 16612 14788 16632 14852
rect 16696 14788 16716 14852
rect 16612 14772 16716 14788
rect 16612 14708 16632 14772
rect 16696 14708 16716 14772
rect 16612 14692 16716 14708
rect 16612 14628 16632 14692
rect 16696 14628 16716 14692
rect 16612 14612 16716 14628
rect 16612 14548 16632 14612
rect 16696 14548 16716 14612
rect 16612 14532 16716 14548
rect 16612 14468 16632 14532
rect 16696 14468 16716 14532
rect 16612 14452 16716 14468
rect 16612 14388 16632 14452
rect 16696 14388 16716 14452
rect 16612 14372 16716 14388
rect 16612 14308 16632 14372
rect 16696 14308 16716 14372
rect 16612 14292 16716 14308
rect 16612 14228 16632 14292
rect 16696 14228 16716 14292
rect 16612 14212 16716 14228
rect 16612 14148 16632 14212
rect 16696 14148 16716 14212
rect 16612 14132 16716 14148
rect 16612 14068 16632 14132
rect 16696 14068 16716 14132
rect 16612 14052 16716 14068
rect 16612 13988 16632 14052
rect 16696 13988 16716 14052
rect 16612 13972 16716 13988
rect 16612 13908 16632 13972
rect 16696 13908 16716 13972
rect 16612 13892 16716 13908
rect 16612 13828 16632 13892
rect 16696 13828 16716 13892
rect 16612 13812 16716 13828
rect 16612 13748 16632 13812
rect 16696 13748 16716 13812
rect 16612 13732 16716 13748
rect 16612 13668 16632 13732
rect 16696 13668 16716 13732
rect 16612 13652 16716 13668
rect 16612 13588 16632 13652
rect 16696 13588 16716 13652
rect 16612 13572 16716 13588
rect 16612 13508 16632 13572
rect 16696 13508 16716 13572
rect 16612 13492 16716 13508
rect 16612 13428 16632 13492
rect 16696 13428 16716 13492
rect 16612 13412 16716 13428
rect 16612 13348 16632 13412
rect 16696 13348 16716 13412
rect 16612 13332 16716 13348
rect 16612 13268 16632 13332
rect 16696 13268 16716 13332
rect 16612 13252 16716 13268
rect 16612 13188 16632 13252
rect 16696 13188 16716 13252
rect 16612 13172 16716 13188
rect 16612 13108 16632 13172
rect 16696 13108 16716 13172
rect 16612 13092 16716 13108
rect 16612 13028 16632 13092
rect 16696 13028 16716 13092
rect 16612 13012 16716 13028
rect 16612 12948 16632 13012
rect 16696 12948 16716 13012
rect 16612 12932 16716 12948
rect 16612 12868 16632 12932
rect 16696 12868 16716 12932
rect 16612 12852 16716 12868
rect 16612 12788 16632 12852
rect 16696 12788 16716 12852
rect 16612 12772 16716 12788
rect 16612 12708 16632 12772
rect 16696 12708 16716 12772
rect 16612 12692 16716 12708
rect 16612 12628 16632 12692
rect 16696 12628 16716 12692
rect 16612 12612 16716 12628
rect 16612 12548 16632 12612
rect 16696 12548 16716 12612
rect 16612 12532 16716 12548
rect 16612 12468 16632 12532
rect 16696 12468 16716 12532
rect 16612 12452 16716 12468
rect 16612 12388 16632 12452
rect 16696 12388 16716 12452
rect 16612 12372 16716 12388
rect 16612 12308 16632 12372
rect 16696 12308 16716 12372
rect 16612 12292 16716 12308
rect 16612 12228 16632 12292
rect 16696 12228 16716 12292
rect 16612 12212 16716 12228
rect 16612 12148 16632 12212
rect 16696 12148 16716 12212
rect 16612 12132 16716 12148
rect 16612 12068 16632 12132
rect 16696 12068 16716 12132
rect 16612 12052 16716 12068
rect 16612 11988 16632 12052
rect 16696 11988 16716 12052
rect 16612 11972 16716 11988
rect 16612 11908 16632 11972
rect 16696 11908 16716 11972
rect 16612 11892 16716 11908
rect 16612 11828 16632 11892
rect 16696 11828 16716 11892
rect 16612 11812 16716 11828
rect 16612 11748 16632 11812
rect 16696 11748 16716 11812
rect 16612 11732 16716 11748
rect 16612 11668 16632 11732
rect 16696 11668 16716 11732
rect 16612 11652 16716 11668
rect 16612 11588 16632 11652
rect 16696 11588 16716 11652
rect 16612 11572 16716 11588
rect 16612 11508 16632 11572
rect 16696 11508 16716 11572
rect 16612 11492 16716 11508
rect 16612 11428 16632 11492
rect 16696 11428 16716 11492
rect 16612 11412 16716 11428
rect 16612 11348 16632 11412
rect 16696 11348 16716 11412
rect 16612 11332 16716 11348
rect 16612 11268 16632 11332
rect 16696 11268 16716 11332
rect 16612 11252 16716 11268
rect 16612 11188 16632 11252
rect 16696 11188 16716 11252
rect 16612 11172 16716 11188
rect 16612 11108 16632 11172
rect 16696 11108 16716 11172
rect 16612 11092 16716 11108
rect 16612 11028 16632 11092
rect 16696 11028 16716 11092
rect 16612 11012 16716 11028
rect 16612 10948 16632 11012
rect 16696 10948 16716 11012
rect 16612 10932 16716 10948
rect 16612 10868 16632 10932
rect 16696 10868 16716 10932
rect 16612 10852 16716 10868
rect 11000 10492 11104 10788
rect 5388 10412 5492 10428
rect 5388 10348 5408 10412
rect 5472 10348 5492 10412
rect 5388 10332 5492 10348
rect 5388 10268 5408 10332
rect 5472 10268 5492 10332
rect 5388 10252 5492 10268
rect 5388 10188 5408 10252
rect 5472 10188 5492 10252
rect 5388 10172 5492 10188
rect 5388 10108 5408 10172
rect 5472 10108 5492 10172
rect 5388 10092 5492 10108
rect 5388 10028 5408 10092
rect 5472 10028 5492 10092
rect 5388 10012 5492 10028
rect 5388 9948 5408 10012
rect 5472 9948 5492 10012
rect 5388 9932 5492 9948
rect 5388 9868 5408 9932
rect 5472 9868 5492 9932
rect 5388 9852 5492 9868
rect 5388 9788 5408 9852
rect 5472 9788 5492 9852
rect 5388 9772 5492 9788
rect 5388 9708 5408 9772
rect 5472 9708 5492 9772
rect 5388 9692 5492 9708
rect 5388 9628 5408 9692
rect 5472 9628 5492 9692
rect 5388 9612 5492 9628
rect 5388 9548 5408 9612
rect 5472 9548 5492 9612
rect 5388 9532 5492 9548
rect 5388 9468 5408 9532
rect 5472 9468 5492 9532
rect 5388 9452 5492 9468
rect 5388 9388 5408 9452
rect 5472 9388 5492 9452
rect 5388 9372 5492 9388
rect 5388 9308 5408 9372
rect 5472 9308 5492 9372
rect 5388 9292 5492 9308
rect 5388 9228 5408 9292
rect 5472 9228 5492 9292
rect 5388 9212 5492 9228
rect 5388 9148 5408 9212
rect 5472 9148 5492 9212
rect 5388 9132 5492 9148
rect 5388 9068 5408 9132
rect 5472 9068 5492 9132
rect 5388 9052 5492 9068
rect 5388 8988 5408 9052
rect 5472 8988 5492 9052
rect 5388 8972 5492 8988
rect 5388 8908 5408 8972
rect 5472 8908 5492 8972
rect 5388 8892 5492 8908
rect 5388 8828 5408 8892
rect 5472 8828 5492 8892
rect 5388 8812 5492 8828
rect 5388 8748 5408 8812
rect 5472 8748 5492 8812
rect 5388 8732 5492 8748
rect 5388 8668 5408 8732
rect 5472 8668 5492 8732
rect 5388 8652 5492 8668
rect 5388 8588 5408 8652
rect 5472 8588 5492 8652
rect 5388 8572 5492 8588
rect 5388 8508 5408 8572
rect 5472 8508 5492 8572
rect 5388 8492 5492 8508
rect 5388 8428 5408 8492
rect 5472 8428 5492 8492
rect 5388 8412 5492 8428
rect 5388 8348 5408 8412
rect 5472 8348 5492 8412
rect 5388 8332 5492 8348
rect 5388 8268 5408 8332
rect 5472 8268 5492 8332
rect 5388 8252 5492 8268
rect 5388 8188 5408 8252
rect 5472 8188 5492 8252
rect 5388 8172 5492 8188
rect 5388 8108 5408 8172
rect 5472 8108 5492 8172
rect 5388 8092 5492 8108
rect 5388 8028 5408 8092
rect 5472 8028 5492 8092
rect 5388 8012 5492 8028
rect 5388 7948 5408 8012
rect 5472 7948 5492 8012
rect 5388 7932 5492 7948
rect 5388 7868 5408 7932
rect 5472 7868 5492 7932
rect 5388 7852 5492 7868
rect 5388 7788 5408 7852
rect 5472 7788 5492 7852
rect 5388 7772 5492 7788
rect 5388 7708 5408 7772
rect 5472 7708 5492 7772
rect 5388 7692 5492 7708
rect 5388 7628 5408 7692
rect 5472 7628 5492 7692
rect 5388 7612 5492 7628
rect 5388 7548 5408 7612
rect 5472 7548 5492 7612
rect 5388 7532 5492 7548
rect 5388 7468 5408 7532
rect 5472 7468 5492 7532
rect 5388 7452 5492 7468
rect 5388 7388 5408 7452
rect 5472 7388 5492 7452
rect 5388 7372 5492 7388
rect 5388 7308 5408 7372
rect 5472 7308 5492 7372
rect 5388 7292 5492 7308
rect 5388 7228 5408 7292
rect 5472 7228 5492 7292
rect 5388 7212 5492 7228
rect 5388 7148 5408 7212
rect 5472 7148 5492 7212
rect 5388 7132 5492 7148
rect 5388 7068 5408 7132
rect 5472 7068 5492 7132
rect 5388 7052 5492 7068
rect 5388 6988 5408 7052
rect 5472 6988 5492 7052
rect 5388 6972 5492 6988
rect 5388 6908 5408 6972
rect 5472 6908 5492 6972
rect 5388 6892 5492 6908
rect 5388 6828 5408 6892
rect 5472 6828 5492 6892
rect 5388 6812 5492 6828
rect 5388 6748 5408 6812
rect 5472 6748 5492 6812
rect 5388 6732 5492 6748
rect 5388 6668 5408 6732
rect 5472 6668 5492 6732
rect 5388 6652 5492 6668
rect 5388 6588 5408 6652
rect 5472 6588 5492 6652
rect 5388 6572 5492 6588
rect 5388 6508 5408 6572
rect 5472 6508 5492 6572
rect 5388 6492 5492 6508
rect 5388 6428 5408 6492
rect 5472 6428 5492 6492
rect 5388 6412 5492 6428
rect 5388 6348 5408 6412
rect 5472 6348 5492 6412
rect 5388 6332 5492 6348
rect 5388 6268 5408 6332
rect 5472 6268 5492 6332
rect 5388 6252 5492 6268
rect 5388 6188 5408 6252
rect 5472 6188 5492 6252
rect 5388 6172 5492 6188
rect 5388 6108 5408 6172
rect 5472 6108 5492 6172
rect 5388 6092 5492 6108
rect 5388 6028 5408 6092
rect 5472 6028 5492 6092
rect 5388 6012 5492 6028
rect 5388 5948 5408 6012
rect 5472 5948 5492 6012
rect 5388 5932 5492 5948
rect 5388 5868 5408 5932
rect 5472 5868 5492 5932
rect 5388 5852 5492 5868
rect 5388 5788 5408 5852
rect 5472 5788 5492 5852
rect 5388 5772 5492 5788
rect 5388 5708 5408 5772
rect 5472 5708 5492 5772
rect 5388 5692 5492 5708
rect 5388 5628 5408 5692
rect 5472 5628 5492 5692
rect 5388 5612 5492 5628
rect 5388 5548 5408 5612
rect 5472 5548 5492 5612
rect 5388 5532 5492 5548
rect -224 5172 -120 5468
rect -5836 5092 -5732 5108
rect -5836 5028 -5816 5092
rect -5752 5028 -5732 5092
rect -5836 5012 -5732 5028
rect -5836 4948 -5816 5012
rect -5752 4948 -5732 5012
rect -5836 4932 -5732 4948
rect -5836 4868 -5816 4932
rect -5752 4868 -5732 4932
rect -5836 4852 -5732 4868
rect -5836 4788 -5816 4852
rect -5752 4788 -5732 4852
rect -5836 4772 -5732 4788
rect -5836 4708 -5816 4772
rect -5752 4708 -5732 4772
rect -5836 4692 -5732 4708
rect -5836 4628 -5816 4692
rect -5752 4628 -5732 4692
rect -5836 4612 -5732 4628
rect -5836 4548 -5816 4612
rect -5752 4548 -5732 4612
rect -5836 4532 -5732 4548
rect -5836 4468 -5816 4532
rect -5752 4468 -5732 4532
rect -5836 4452 -5732 4468
rect -5836 4388 -5816 4452
rect -5752 4388 -5732 4452
rect -5836 4372 -5732 4388
rect -5836 4308 -5816 4372
rect -5752 4308 -5732 4372
rect -5836 4292 -5732 4308
rect -5836 4228 -5816 4292
rect -5752 4228 -5732 4292
rect -5836 4212 -5732 4228
rect -5836 4148 -5816 4212
rect -5752 4148 -5732 4212
rect -5836 4132 -5732 4148
rect -5836 4068 -5816 4132
rect -5752 4068 -5732 4132
rect -5836 4052 -5732 4068
rect -5836 3988 -5816 4052
rect -5752 3988 -5732 4052
rect -5836 3972 -5732 3988
rect -5836 3908 -5816 3972
rect -5752 3908 -5732 3972
rect -5836 3892 -5732 3908
rect -5836 3828 -5816 3892
rect -5752 3828 -5732 3892
rect -5836 3812 -5732 3828
rect -5836 3748 -5816 3812
rect -5752 3748 -5732 3812
rect -5836 3732 -5732 3748
rect -5836 3668 -5816 3732
rect -5752 3668 -5732 3732
rect -5836 3652 -5732 3668
rect -5836 3588 -5816 3652
rect -5752 3588 -5732 3652
rect -5836 3572 -5732 3588
rect -5836 3508 -5816 3572
rect -5752 3508 -5732 3572
rect -5836 3492 -5732 3508
rect -5836 3428 -5816 3492
rect -5752 3428 -5732 3492
rect -5836 3412 -5732 3428
rect -5836 3348 -5816 3412
rect -5752 3348 -5732 3412
rect -5836 3332 -5732 3348
rect -5836 3268 -5816 3332
rect -5752 3268 -5732 3332
rect -5836 3252 -5732 3268
rect -5836 3188 -5816 3252
rect -5752 3188 -5732 3252
rect -5836 3172 -5732 3188
rect -5836 3108 -5816 3172
rect -5752 3108 -5732 3172
rect -5836 3092 -5732 3108
rect -5836 3028 -5816 3092
rect -5752 3028 -5732 3092
rect -5836 3012 -5732 3028
rect -5836 2948 -5816 3012
rect -5752 2948 -5732 3012
rect -5836 2932 -5732 2948
rect -5836 2868 -5816 2932
rect -5752 2868 -5732 2932
rect -5836 2852 -5732 2868
rect -5836 2788 -5816 2852
rect -5752 2788 -5732 2852
rect -5836 2772 -5732 2788
rect -5836 2708 -5816 2772
rect -5752 2708 -5732 2772
rect -5836 2692 -5732 2708
rect -5836 2628 -5816 2692
rect -5752 2628 -5732 2692
rect -5836 2612 -5732 2628
rect -5836 2548 -5816 2612
rect -5752 2548 -5732 2612
rect -5836 2532 -5732 2548
rect -5836 2468 -5816 2532
rect -5752 2468 -5732 2532
rect -5836 2452 -5732 2468
rect -5836 2388 -5816 2452
rect -5752 2388 -5732 2452
rect -5836 2372 -5732 2388
rect -5836 2308 -5816 2372
rect -5752 2308 -5732 2372
rect -5836 2292 -5732 2308
rect -5836 2228 -5816 2292
rect -5752 2228 -5732 2292
rect -5836 2212 -5732 2228
rect -5836 2148 -5816 2212
rect -5752 2148 -5732 2212
rect -5836 2132 -5732 2148
rect -5836 2068 -5816 2132
rect -5752 2068 -5732 2132
rect -5836 2052 -5732 2068
rect -5836 1988 -5816 2052
rect -5752 1988 -5732 2052
rect -5836 1972 -5732 1988
rect -5836 1908 -5816 1972
rect -5752 1908 -5732 1972
rect -5836 1892 -5732 1908
rect -5836 1828 -5816 1892
rect -5752 1828 -5732 1892
rect -5836 1812 -5732 1828
rect -5836 1748 -5816 1812
rect -5752 1748 -5732 1812
rect -5836 1732 -5732 1748
rect -5836 1668 -5816 1732
rect -5752 1668 -5732 1732
rect -5836 1652 -5732 1668
rect -5836 1588 -5816 1652
rect -5752 1588 -5732 1652
rect -5836 1572 -5732 1588
rect -5836 1508 -5816 1572
rect -5752 1508 -5732 1572
rect -5836 1492 -5732 1508
rect -5836 1428 -5816 1492
rect -5752 1428 -5732 1492
rect -5836 1412 -5732 1428
rect -5836 1348 -5816 1412
rect -5752 1348 -5732 1412
rect -5836 1332 -5732 1348
rect -5836 1268 -5816 1332
rect -5752 1268 -5732 1332
rect -5836 1252 -5732 1268
rect -5836 1188 -5816 1252
rect -5752 1188 -5732 1252
rect -5836 1172 -5732 1188
rect -5836 1108 -5816 1172
rect -5752 1108 -5732 1172
rect -5836 1092 -5732 1108
rect -5836 1028 -5816 1092
rect -5752 1028 -5732 1092
rect -5836 1012 -5732 1028
rect -5836 948 -5816 1012
rect -5752 948 -5732 1012
rect -5836 932 -5732 948
rect -5836 868 -5816 932
rect -5752 868 -5732 932
rect -5836 852 -5732 868
rect -5836 788 -5816 852
rect -5752 788 -5732 852
rect -5836 772 -5732 788
rect -5836 708 -5816 772
rect -5752 708 -5732 772
rect -5836 692 -5732 708
rect -5836 628 -5816 692
rect -5752 628 -5732 692
rect -5836 612 -5732 628
rect -5836 548 -5816 612
rect -5752 548 -5732 612
rect -5836 532 -5732 548
rect -5836 468 -5816 532
rect -5752 468 -5732 532
rect -5836 452 -5732 468
rect -5836 388 -5816 452
rect -5752 388 -5732 452
rect -5836 372 -5732 388
rect -5836 308 -5816 372
rect -5752 308 -5732 372
rect -5836 292 -5732 308
rect -5836 228 -5816 292
rect -5752 228 -5732 292
rect -5836 212 -5732 228
rect -11448 -148 -11344 148
rect -17060 -228 -16956 -212
rect -17060 -292 -17040 -228
rect -16976 -292 -16956 -228
rect -17060 -308 -16956 -292
rect -17060 -372 -17040 -308
rect -16976 -372 -16956 -308
rect -17060 -388 -16956 -372
rect -17060 -452 -17040 -388
rect -16976 -452 -16956 -388
rect -17060 -468 -16956 -452
rect -17060 -532 -17040 -468
rect -16976 -532 -16956 -468
rect -17060 -548 -16956 -532
rect -17060 -612 -17040 -548
rect -16976 -612 -16956 -548
rect -17060 -628 -16956 -612
rect -17060 -692 -17040 -628
rect -16976 -692 -16956 -628
rect -17060 -708 -16956 -692
rect -17060 -772 -17040 -708
rect -16976 -772 -16956 -708
rect -17060 -788 -16956 -772
rect -17060 -852 -17040 -788
rect -16976 -852 -16956 -788
rect -17060 -868 -16956 -852
rect -17060 -932 -17040 -868
rect -16976 -932 -16956 -868
rect -17060 -948 -16956 -932
rect -17060 -1012 -17040 -948
rect -16976 -1012 -16956 -948
rect -17060 -1028 -16956 -1012
rect -17060 -1092 -17040 -1028
rect -16976 -1092 -16956 -1028
rect -17060 -1108 -16956 -1092
rect -17060 -1172 -17040 -1108
rect -16976 -1172 -16956 -1108
rect -17060 -1188 -16956 -1172
rect -17060 -1252 -17040 -1188
rect -16976 -1252 -16956 -1188
rect -17060 -1268 -16956 -1252
rect -17060 -1332 -17040 -1268
rect -16976 -1332 -16956 -1268
rect -17060 -1348 -16956 -1332
rect -17060 -1412 -17040 -1348
rect -16976 -1412 -16956 -1348
rect -17060 -1428 -16956 -1412
rect -17060 -1492 -17040 -1428
rect -16976 -1492 -16956 -1428
rect -17060 -1508 -16956 -1492
rect -17060 -1572 -17040 -1508
rect -16976 -1572 -16956 -1508
rect -17060 -1588 -16956 -1572
rect -17060 -1652 -17040 -1588
rect -16976 -1652 -16956 -1588
rect -17060 -1668 -16956 -1652
rect -17060 -1732 -17040 -1668
rect -16976 -1732 -16956 -1668
rect -17060 -1748 -16956 -1732
rect -17060 -1812 -17040 -1748
rect -16976 -1812 -16956 -1748
rect -17060 -1828 -16956 -1812
rect -17060 -1892 -17040 -1828
rect -16976 -1892 -16956 -1828
rect -17060 -1908 -16956 -1892
rect -17060 -1972 -17040 -1908
rect -16976 -1972 -16956 -1908
rect -17060 -1988 -16956 -1972
rect -17060 -2052 -17040 -1988
rect -16976 -2052 -16956 -1988
rect -17060 -2068 -16956 -2052
rect -17060 -2132 -17040 -2068
rect -16976 -2132 -16956 -2068
rect -17060 -2148 -16956 -2132
rect -17060 -2212 -17040 -2148
rect -16976 -2212 -16956 -2148
rect -17060 -2228 -16956 -2212
rect -17060 -2292 -17040 -2228
rect -16976 -2292 -16956 -2228
rect -17060 -2308 -16956 -2292
rect -17060 -2372 -17040 -2308
rect -16976 -2372 -16956 -2308
rect -17060 -2388 -16956 -2372
rect -17060 -2452 -17040 -2388
rect -16976 -2452 -16956 -2388
rect -17060 -2468 -16956 -2452
rect -17060 -2532 -17040 -2468
rect -16976 -2532 -16956 -2468
rect -17060 -2548 -16956 -2532
rect -17060 -2612 -17040 -2548
rect -16976 -2612 -16956 -2548
rect -17060 -2628 -16956 -2612
rect -17060 -2692 -17040 -2628
rect -16976 -2692 -16956 -2628
rect -17060 -2708 -16956 -2692
rect -17060 -2772 -17040 -2708
rect -16976 -2772 -16956 -2708
rect -17060 -2788 -16956 -2772
rect -17060 -2852 -17040 -2788
rect -16976 -2852 -16956 -2788
rect -17060 -2868 -16956 -2852
rect -17060 -2932 -17040 -2868
rect -16976 -2932 -16956 -2868
rect -17060 -2948 -16956 -2932
rect -17060 -3012 -17040 -2948
rect -16976 -3012 -16956 -2948
rect -17060 -3028 -16956 -3012
rect -17060 -3092 -17040 -3028
rect -16976 -3092 -16956 -3028
rect -17060 -3108 -16956 -3092
rect -17060 -3172 -17040 -3108
rect -16976 -3172 -16956 -3108
rect -17060 -3188 -16956 -3172
rect -17060 -3252 -17040 -3188
rect -16976 -3252 -16956 -3188
rect -17060 -3268 -16956 -3252
rect -17060 -3332 -17040 -3268
rect -16976 -3332 -16956 -3268
rect -17060 -3348 -16956 -3332
rect -17060 -3412 -17040 -3348
rect -16976 -3412 -16956 -3348
rect -17060 -3428 -16956 -3412
rect -17060 -3492 -17040 -3428
rect -16976 -3492 -16956 -3428
rect -17060 -3508 -16956 -3492
rect -17060 -3572 -17040 -3508
rect -16976 -3572 -16956 -3508
rect -17060 -3588 -16956 -3572
rect -17060 -3652 -17040 -3588
rect -16976 -3652 -16956 -3588
rect -17060 -3668 -16956 -3652
rect -17060 -3732 -17040 -3668
rect -16976 -3732 -16956 -3668
rect -17060 -3748 -16956 -3732
rect -17060 -3812 -17040 -3748
rect -16976 -3812 -16956 -3748
rect -17060 -3828 -16956 -3812
rect -17060 -3892 -17040 -3828
rect -16976 -3892 -16956 -3828
rect -17060 -3908 -16956 -3892
rect -17060 -3972 -17040 -3908
rect -16976 -3972 -16956 -3908
rect -17060 -3988 -16956 -3972
rect -17060 -4052 -17040 -3988
rect -16976 -4052 -16956 -3988
rect -17060 -4068 -16956 -4052
rect -17060 -4132 -17040 -4068
rect -16976 -4132 -16956 -4068
rect -17060 -4148 -16956 -4132
rect -17060 -4212 -17040 -4148
rect -16976 -4212 -16956 -4148
rect -17060 -4228 -16956 -4212
rect -17060 -4292 -17040 -4228
rect -16976 -4292 -16956 -4228
rect -17060 -4308 -16956 -4292
rect -17060 -4372 -17040 -4308
rect -16976 -4372 -16956 -4308
rect -17060 -4388 -16956 -4372
rect -17060 -4452 -17040 -4388
rect -16976 -4452 -16956 -4388
rect -17060 -4468 -16956 -4452
rect -17060 -4532 -17040 -4468
rect -16976 -4532 -16956 -4468
rect -17060 -4548 -16956 -4532
rect -17060 -4612 -17040 -4548
rect -16976 -4612 -16956 -4548
rect -17060 -4628 -16956 -4612
rect -17060 -4692 -17040 -4628
rect -16976 -4692 -16956 -4628
rect -17060 -4708 -16956 -4692
rect -17060 -4772 -17040 -4708
rect -16976 -4772 -16956 -4708
rect -17060 -4788 -16956 -4772
rect -17060 -4852 -17040 -4788
rect -16976 -4852 -16956 -4788
rect -17060 -4868 -16956 -4852
rect -17060 -4932 -17040 -4868
rect -16976 -4932 -16956 -4868
rect -17060 -4948 -16956 -4932
rect -17060 -5012 -17040 -4948
rect -16976 -5012 -16956 -4948
rect -17060 -5028 -16956 -5012
rect -17060 -5092 -17040 -5028
rect -16976 -5092 -16956 -5028
rect -17060 -5108 -16956 -5092
rect -22672 -5468 -22568 -5172
rect -28284 -5548 -28180 -5532
rect -28284 -5612 -28264 -5548
rect -28200 -5612 -28180 -5548
rect -28284 -5628 -28180 -5612
rect -28284 -5692 -28264 -5628
rect -28200 -5692 -28180 -5628
rect -28284 -5708 -28180 -5692
rect -28284 -5772 -28264 -5708
rect -28200 -5772 -28180 -5708
rect -28284 -5788 -28180 -5772
rect -28284 -5852 -28264 -5788
rect -28200 -5852 -28180 -5788
rect -28284 -5868 -28180 -5852
rect -28284 -5932 -28264 -5868
rect -28200 -5932 -28180 -5868
rect -28284 -5948 -28180 -5932
rect -28284 -6012 -28264 -5948
rect -28200 -6012 -28180 -5948
rect -28284 -6028 -28180 -6012
rect -28284 -6092 -28264 -6028
rect -28200 -6092 -28180 -6028
rect -28284 -6108 -28180 -6092
rect -28284 -6172 -28264 -6108
rect -28200 -6172 -28180 -6108
rect -28284 -6188 -28180 -6172
rect -28284 -6252 -28264 -6188
rect -28200 -6252 -28180 -6188
rect -28284 -6268 -28180 -6252
rect -28284 -6332 -28264 -6268
rect -28200 -6332 -28180 -6268
rect -28284 -6348 -28180 -6332
rect -28284 -6412 -28264 -6348
rect -28200 -6412 -28180 -6348
rect -28284 -6428 -28180 -6412
rect -28284 -6492 -28264 -6428
rect -28200 -6492 -28180 -6428
rect -28284 -6508 -28180 -6492
rect -28284 -6572 -28264 -6508
rect -28200 -6572 -28180 -6508
rect -28284 -6588 -28180 -6572
rect -28284 -6652 -28264 -6588
rect -28200 -6652 -28180 -6588
rect -28284 -6668 -28180 -6652
rect -28284 -6732 -28264 -6668
rect -28200 -6732 -28180 -6668
rect -28284 -6748 -28180 -6732
rect -28284 -6812 -28264 -6748
rect -28200 -6812 -28180 -6748
rect -28284 -6828 -28180 -6812
rect -28284 -6892 -28264 -6828
rect -28200 -6892 -28180 -6828
rect -28284 -6908 -28180 -6892
rect -28284 -6972 -28264 -6908
rect -28200 -6972 -28180 -6908
rect -28284 -6988 -28180 -6972
rect -28284 -7052 -28264 -6988
rect -28200 -7052 -28180 -6988
rect -28284 -7068 -28180 -7052
rect -28284 -7132 -28264 -7068
rect -28200 -7132 -28180 -7068
rect -28284 -7148 -28180 -7132
rect -28284 -7212 -28264 -7148
rect -28200 -7212 -28180 -7148
rect -28284 -7228 -28180 -7212
rect -28284 -7292 -28264 -7228
rect -28200 -7292 -28180 -7228
rect -28284 -7308 -28180 -7292
rect -28284 -7372 -28264 -7308
rect -28200 -7372 -28180 -7308
rect -28284 -7388 -28180 -7372
rect -28284 -7452 -28264 -7388
rect -28200 -7452 -28180 -7388
rect -28284 -7468 -28180 -7452
rect -28284 -7532 -28264 -7468
rect -28200 -7532 -28180 -7468
rect -28284 -7548 -28180 -7532
rect -28284 -7612 -28264 -7548
rect -28200 -7612 -28180 -7548
rect -28284 -7628 -28180 -7612
rect -28284 -7692 -28264 -7628
rect -28200 -7692 -28180 -7628
rect -28284 -7708 -28180 -7692
rect -28284 -7772 -28264 -7708
rect -28200 -7772 -28180 -7708
rect -28284 -7788 -28180 -7772
rect -28284 -7852 -28264 -7788
rect -28200 -7852 -28180 -7788
rect -28284 -7868 -28180 -7852
rect -28284 -7932 -28264 -7868
rect -28200 -7932 -28180 -7868
rect -28284 -7948 -28180 -7932
rect -28284 -8012 -28264 -7948
rect -28200 -8012 -28180 -7948
rect -28284 -8028 -28180 -8012
rect -28284 -8092 -28264 -8028
rect -28200 -8092 -28180 -8028
rect -28284 -8108 -28180 -8092
rect -28284 -8172 -28264 -8108
rect -28200 -8172 -28180 -8108
rect -28284 -8188 -28180 -8172
rect -28284 -8252 -28264 -8188
rect -28200 -8252 -28180 -8188
rect -28284 -8268 -28180 -8252
rect -28284 -8332 -28264 -8268
rect -28200 -8332 -28180 -8268
rect -28284 -8348 -28180 -8332
rect -28284 -8412 -28264 -8348
rect -28200 -8412 -28180 -8348
rect -28284 -8428 -28180 -8412
rect -28284 -8492 -28264 -8428
rect -28200 -8492 -28180 -8428
rect -28284 -8508 -28180 -8492
rect -28284 -8572 -28264 -8508
rect -28200 -8572 -28180 -8508
rect -28284 -8588 -28180 -8572
rect -28284 -8652 -28264 -8588
rect -28200 -8652 -28180 -8588
rect -28284 -8668 -28180 -8652
rect -28284 -8732 -28264 -8668
rect -28200 -8732 -28180 -8668
rect -28284 -8748 -28180 -8732
rect -28284 -8812 -28264 -8748
rect -28200 -8812 -28180 -8748
rect -28284 -8828 -28180 -8812
rect -28284 -8892 -28264 -8828
rect -28200 -8892 -28180 -8828
rect -28284 -8908 -28180 -8892
rect -28284 -8972 -28264 -8908
rect -28200 -8972 -28180 -8908
rect -28284 -8988 -28180 -8972
rect -28284 -9052 -28264 -8988
rect -28200 -9052 -28180 -8988
rect -28284 -9068 -28180 -9052
rect -28284 -9132 -28264 -9068
rect -28200 -9132 -28180 -9068
rect -28284 -9148 -28180 -9132
rect -28284 -9212 -28264 -9148
rect -28200 -9212 -28180 -9148
rect -28284 -9228 -28180 -9212
rect -28284 -9292 -28264 -9228
rect -28200 -9292 -28180 -9228
rect -28284 -9308 -28180 -9292
rect -28284 -9372 -28264 -9308
rect -28200 -9372 -28180 -9308
rect -28284 -9388 -28180 -9372
rect -28284 -9452 -28264 -9388
rect -28200 -9452 -28180 -9388
rect -28284 -9468 -28180 -9452
rect -28284 -9532 -28264 -9468
rect -28200 -9532 -28180 -9468
rect -28284 -9548 -28180 -9532
rect -28284 -9612 -28264 -9548
rect -28200 -9612 -28180 -9548
rect -28284 -9628 -28180 -9612
rect -28284 -9692 -28264 -9628
rect -28200 -9692 -28180 -9628
rect -28284 -9708 -28180 -9692
rect -28284 -9772 -28264 -9708
rect -28200 -9772 -28180 -9708
rect -28284 -9788 -28180 -9772
rect -28284 -9852 -28264 -9788
rect -28200 -9852 -28180 -9788
rect -28284 -9868 -28180 -9852
rect -28284 -9932 -28264 -9868
rect -28200 -9932 -28180 -9868
rect -28284 -9948 -28180 -9932
rect -28284 -10012 -28264 -9948
rect -28200 -10012 -28180 -9948
rect -28284 -10028 -28180 -10012
rect -28284 -10092 -28264 -10028
rect -28200 -10092 -28180 -10028
rect -28284 -10108 -28180 -10092
rect -28284 -10172 -28264 -10108
rect -28200 -10172 -28180 -10108
rect -28284 -10188 -28180 -10172
rect -28284 -10252 -28264 -10188
rect -28200 -10252 -28180 -10188
rect -28284 -10268 -28180 -10252
rect -28284 -10332 -28264 -10268
rect -28200 -10332 -28180 -10268
rect -28284 -10348 -28180 -10332
rect -28284 -10412 -28264 -10348
rect -28200 -10412 -28180 -10348
rect -28284 -10428 -28180 -10412
rect -33896 -10788 -33792 -10492
rect -39085 -10868 -34163 -10839
rect -39085 -15732 -39056 -10868
rect -34192 -15732 -34163 -10868
rect -39085 -15761 -34163 -15732
rect -33896 -10852 -33876 -10788
rect -33812 -10852 -33792 -10788
rect -31064 -10839 -30960 -10441
rect -28284 -10492 -28264 -10428
rect -28200 -10492 -28180 -10428
rect -27861 -5548 -22939 -5519
rect -27861 -10412 -27832 -5548
rect -22968 -10412 -22939 -5548
rect -27861 -10441 -22939 -10412
rect -22672 -5532 -22652 -5468
rect -22588 -5532 -22568 -5468
rect -19840 -5519 -19736 -5121
rect -17060 -5172 -17040 -5108
rect -16976 -5172 -16956 -5108
rect -16637 -228 -11715 -199
rect -16637 -5092 -16608 -228
rect -11744 -5092 -11715 -228
rect -16637 -5121 -11715 -5092
rect -11448 -212 -11428 -148
rect -11364 -212 -11344 -148
rect -8616 -199 -8512 199
rect -5836 148 -5816 212
rect -5752 148 -5732 212
rect -5413 5092 -491 5121
rect -5413 228 -5384 5092
rect -520 228 -491 5092
rect -5413 199 -491 228
rect -224 5108 -204 5172
rect -140 5108 -120 5172
rect 2608 5121 2712 5519
rect 5388 5468 5408 5532
rect 5472 5468 5492 5532
rect 5811 10412 10733 10441
rect 5811 5548 5840 10412
rect 10704 5548 10733 10412
rect 5811 5519 10733 5548
rect 11000 10428 11020 10492
rect 11084 10428 11104 10492
rect 13832 10441 13936 10839
rect 16612 10788 16632 10852
rect 16696 10788 16716 10852
rect 17035 15732 21957 15761
rect 17035 10868 17064 15732
rect 21928 10868 21957 15732
rect 17035 10839 21957 10868
rect 22224 15748 22244 15812
rect 22308 15748 22328 15812
rect 25056 15761 25160 16159
rect 27836 16108 27856 16172
rect 27920 16108 27940 16172
rect 28259 21052 33181 21081
rect 28259 16188 28288 21052
rect 33152 16188 33181 21052
rect 28259 16159 33181 16188
rect 33448 21068 33468 21132
rect 33532 21068 33552 21132
rect 36280 21081 36384 21479
rect 39060 21428 39080 21492
rect 39144 21428 39164 21492
rect 39060 21132 39164 21428
rect 33448 21052 33552 21068
rect 33448 20988 33468 21052
rect 33532 20988 33552 21052
rect 33448 20972 33552 20988
rect 33448 20908 33468 20972
rect 33532 20908 33552 20972
rect 33448 20892 33552 20908
rect 33448 20828 33468 20892
rect 33532 20828 33552 20892
rect 33448 20812 33552 20828
rect 33448 20748 33468 20812
rect 33532 20748 33552 20812
rect 33448 20732 33552 20748
rect 33448 20668 33468 20732
rect 33532 20668 33552 20732
rect 33448 20652 33552 20668
rect 33448 20588 33468 20652
rect 33532 20588 33552 20652
rect 33448 20572 33552 20588
rect 33448 20508 33468 20572
rect 33532 20508 33552 20572
rect 33448 20492 33552 20508
rect 33448 20428 33468 20492
rect 33532 20428 33552 20492
rect 33448 20412 33552 20428
rect 33448 20348 33468 20412
rect 33532 20348 33552 20412
rect 33448 20332 33552 20348
rect 33448 20268 33468 20332
rect 33532 20268 33552 20332
rect 33448 20252 33552 20268
rect 33448 20188 33468 20252
rect 33532 20188 33552 20252
rect 33448 20172 33552 20188
rect 33448 20108 33468 20172
rect 33532 20108 33552 20172
rect 33448 20092 33552 20108
rect 33448 20028 33468 20092
rect 33532 20028 33552 20092
rect 33448 20012 33552 20028
rect 33448 19948 33468 20012
rect 33532 19948 33552 20012
rect 33448 19932 33552 19948
rect 33448 19868 33468 19932
rect 33532 19868 33552 19932
rect 33448 19852 33552 19868
rect 33448 19788 33468 19852
rect 33532 19788 33552 19852
rect 33448 19772 33552 19788
rect 33448 19708 33468 19772
rect 33532 19708 33552 19772
rect 33448 19692 33552 19708
rect 33448 19628 33468 19692
rect 33532 19628 33552 19692
rect 33448 19612 33552 19628
rect 33448 19548 33468 19612
rect 33532 19548 33552 19612
rect 33448 19532 33552 19548
rect 33448 19468 33468 19532
rect 33532 19468 33552 19532
rect 33448 19452 33552 19468
rect 33448 19388 33468 19452
rect 33532 19388 33552 19452
rect 33448 19372 33552 19388
rect 33448 19308 33468 19372
rect 33532 19308 33552 19372
rect 33448 19292 33552 19308
rect 33448 19228 33468 19292
rect 33532 19228 33552 19292
rect 33448 19212 33552 19228
rect 33448 19148 33468 19212
rect 33532 19148 33552 19212
rect 33448 19132 33552 19148
rect 33448 19068 33468 19132
rect 33532 19068 33552 19132
rect 33448 19052 33552 19068
rect 33448 18988 33468 19052
rect 33532 18988 33552 19052
rect 33448 18972 33552 18988
rect 33448 18908 33468 18972
rect 33532 18908 33552 18972
rect 33448 18892 33552 18908
rect 33448 18828 33468 18892
rect 33532 18828 33552 18892
rect 33448 18812 33552 18828
rect 33448 18748 33468 18812
rect 33532 18748 33552 18812
rect 33448 18732 33552 18748
rect 33448 18668 33468 18732
rect 33532 18668 33552 18732
rect 33448 18652 33552 18668
rect 33448 18588 33468 18652
rect 33532 18588 33552 18652
rect 33448 18572 33552 18588
rect 33448 18508 33468 18572
rect 33532 18508 33552 18572
rect 33448 18492 33552 18508
rect 33448 18428 33468 18492
rect 33532 18428 33552 18492
rect 33448 18412 33552 18428
rect 33448 18348 33468 18412
rect 33532 18348 33552 18412
rect 33448 18332 33552 18348
rect 33448 18268 33468 18332
rect 33532 18268 33552 18332
rect 33448 18252 33552 18268
rect 33448 18188 33468 18252
rect 33532 18188 33552 18252
rect 33448 18172 33552 18188
rect 33448 18108 33468 18172
rect 33532 18108 33552 18172
rect 33448 18092 33552 18108
rect 33448 18028 33468 18092
rect 33532 18028 33552 18092
rect 33448 18012 33552 18028
rect 33448 17948 33468 18012
rect 33532 17948 33552 18012
rect 33448 17932 33552 17948
rect 33448 17868 33468 17932
rect 33532 17868 33552 17932
rect 33448 17852 33552 17868
rect 33448 17788 33468 17852
rect 33532 17788 33552 17852
rect 33448 17772 33552 17788
rect 33448 17708 33468 17772
rect 33532 17708 33552 17772
rect 33448 17692 33552 17708
rect 33448 17628 33468 17692
rect 33532 17628 33552 17692
rect 33448 17612 33552 17628
rect 33448 17548 33468 17612
rect 33532 17548 33552 17612
rect 33448 17532 33552 17548
rect 33448 17468 33468 17532
rect 33532 17468 33552 17532
rect 33448 17452 33552 17468
rect 33448 17388 33468 17452
rect 33532 17388 33552 17452
rect 33448 17372 33552 17388
rect 33448 17308 33468 17372
rect 33532 17308 33552 17372
rect 33448 17292 33552 17308
rect 33448 17228 33468 17292
rect 33532 17228 33552 17292
rect 33448 17212 33552 17228
rect 33448 17148 33468 17212
rect 33532 17148 33552 17212
rect 33448 17132 33552 17148
rect 33448 17068 33468 17132
rect 33532 17068 33552 17132
rect 33448 17052 33552 17068
rect 33448 16988 33468 17052
rect 33532 16988 33552 17052
rect 33448 16972 33552 16988
rect 33448 16908 33468 16972
rect 33532 16908 33552 16972
rect 33448 16892 33552 16908
rect 33448 16828 33468 16892
rect 33532 16828 33552 16892
rect 33448 16812 33552 16828
rect 33448 16748 33468 16812
rect 33532 16748 33552 16812
rect 33448 16732 33552 16748
rect 33448 16668 33468 16732
rect 33532 16668 33552 16732
rect 33448 16652 33552 16668
rect 33448 16588 33468 16652
rect 33532 16588 33552 16652
rect 33448 16572 33552 16588
rect 33448 16508 33468 16572
rect 33532 16508 33552 16572
rect 33448 16492 33552 16508
rect 33448 16428 33468 16492
rect 33532 16428 33552 16492
rect 33448 16412 33552 16428
rect 33448 16348 33468 16412
rect 33532 16348 33552 16412
rect 33448 16332 33552 16348
rect 33448 16268 33468 16332
rect 33532 16268 33552 16332
rect 33448 16252 33552 16268
rect 33448 16188 33468 16252
rect 33532 16188 33552 16252
rect 33448 16172 33552 16188
rect 27836 15812 27940 16108
rect 22224 15732 22328 15748
rect 22224 15668 22244 15732
rect 22308 15668 22328 15732
rect 22224 15652 22328 15668
rect 22224 15588 22244 15652
rect 22308 15588 22328 15652
rect 22224 15572 22328 15588
rect 22224 15508 22244 15572
rect 22308 15508 22328 15572
rect 22224 15492 22328 15508
rect 22224 15428 22244 15492
rect 22308 15428 22328 15492
rect 22224 15412 22328 15428
rect 22224 15348 22244 15412
rect 22308 15348 22328 15412
rect 22224 15332 22328 15348
rect 22224 15268 22244 15332
rect 22308 15268 22328 15332
rect 22224 15252 22328 15268
rect 22224 15188 22244 15252
rect 22308 15188 22328 15252
rect 22224 15172 22328 15188
rect 22224 15108 22244 15172
rect 22308 15108 22328 15172
rect 22224 15092 22328 15108
rect 22224 15028 22244 15092
rect 22308 15028 22328 15092
rect 22224 15012 22328 15028
rect 22224 14948 22244 15012
rect 22308 14948 22328 15012
rect 22224 14932 22328 14948
rect 22224 14868 22244 14932
rect 22308 14868 22328 14932
rect 22224 14852 22328 14868
rect 22224 14788 22244 14852
rect 22308 14788 22328 14852
rect 22224 14772 22328 14788
rect 22224 14708 22244 14772
rect 22308 14708 22328 14772
rect 22224 14692 22328 14708
rect 22224 14628 22244 14692
rect 22308 14628 22328 14692
rect 22224 14612 22328 14628
rect 22224 14548 22244 14612
rect 22308 14548 22328 14612
rect 22224 14532 22328 14548
rect 22224 14468 22244 14532
rect 22308 14468 22328 14532
rect 22224 14452 22328 14468
rect 22224 14388 22244 14452
rect 22308 14388 22328 14452
rect 22224 14372 22328 14388
rect 22224 14308 22244 14372
rect 22308 14308 22328 14372
rect 22224 14292 22328 14308
rect 22224 14228 22244 14292
rect 22308 14228 22328 14292
rect 22224 14212 22328 14228
rect 22224 14148 22244 14212
rect 22308 14148 22328 14212
rect 22224 14132 22328 14148
rect 22224 14068 22244 14132
rect 22308 14068 22328 14132
rect 22224 14052 22328 14068
rect 22224 13988 22244 14052
rect 22308 13988 22328 14052
rect 22224 13972 22328 13988
rect 22224 13908 22244 13972
rect 22308 13908 22328 13972
rect 22224 13892 22328 13908
rect 22224 13828 22244 13892
rect 22308 13828 22328 13892
rect 22224 13812 22328 13828
rect 22224 13748 22244 13812
rect 22308 13748 22328 13812
rect 22224 13732 22328 13748
rect 22224 13668 22244 13732
rect 22308 13668 22328 13732
rect 22224 13652 22328 13668
rect 22224 13588 22244 13652
rect 22308 13588 22328 13652
rect 22224 13572 22328 13588
rect 22224 13508 22244 13572
rect 22308 13508 22328 13572
rect 22224 13492 22328 13508
rect 22224 13428 22244 13492
rect 22308 13428 22328 13492
rect 22224 13412 22328 13428
rect 22224 13348 22244 13412
rect 22308 13348 22328 13412
rect 22224 13332 22328 13348
rect 22224 13268 22244 13332
rect 22308 13268 22328 13332
rect 22224 13252 22328 13268
rect 22224 13188 22244 13252
rect 22308 13188 22328 13252
rect 22224 13172 22328 13188
rect 22224 13108 22244 13172
rect 22308 13108 22328 13172
rect 22224 13092 22328 13108
rect 22224 13028 22244 13092
rect 22308 13028 22328 13092
rect 22224 13012 22328 13028
rect 22224 12948 22244 13012
rect 22308 12948 22328 13012
rect 22224 12932 22328 12948
rect 22224 12868 22244 12932
rect 22308 12868 22328 12932
rect 22224 12852 22328 12868
rect 22224 12788 22244 12852
rect 22308 12788 22328 12852
rect 22224 12772 22328 12788
rect 22224 12708 22244 12772
rect 22308 12708 22328 12772
rect 22224 12692 22328 12708
rect 22224 12628 22244 12692
rect 22308 12628 22328 12692
rect 22224 12612 22328 12628
rect 22224 12548 22244 12612
rect 22308 12548 22328 12612
rect 22224 12532 22328 12548
rect 22224 12468 22244 12532
rect 22308 12468 22328 12532
rect 22224 12452 22328 12468
rect 22224 12388 22244 12452
rect 22308 12388 22328 12452
rect 22224 12372 22328 12388
rect 22224 12308 22244 12372
rect 22308 12308 22328 12372
rect 22224 12292 22328 12308
rect 22224 12228 22244 12292
rect 22308 12228 22328 12292
rect 22224 12212 22328 12228
rect 22224 12148 22244 12212
rect 22308 12148 22328 12212
rect 22224 12132 22328 12148
rect 22224 12068 22244 12132
rect 22308 12068 22328 12132
rect 22224 12052 22328 12068
rect 22224 11988 22244 12052
rect 22308 11988 22328 12052
rect 22224 11972 22328 11988
rect 22224 11908 22244 11972
rect 22308 11908 22328 11972
rect 22224 11892 22328 11908
rect 22224 11828 22244 11892
rect 22308 11828 22328 11892
rect 22224 11812 22328 11828
rect 22224 11748 22244 11812
rect 22308 11748 22328 11812
rect 22224 11732 22328 11748
rect 22224 11668 22244 11732
rect 22308 11668 22328 11732
rect 22224 11652 22328 11668
rect 22224 11588 22244 11652
rect 22308 11588 22328 11652
rect 22224 11572 22328 11588
rect 22224 11508 22244 11572
rect 22308 11508 22328 11572
rect 22224 11492 22328 11508
rect 22224 11428 22244 11492
rect 22308 11428 22328 11492
rect 22224 11412 22328 11428
rect 22224 11348 22244 11412
rect 22308 11348 22328 11412
rect 22224 11332 22328 11348
rect 22224 11268 22244 11332
rect 22308 11268 22328 11332
rect 22224 11252 22328 11268
rect 22224 11188 22244 11252
rect 22308 11188 22328 11252
rect 22224 11172 22328 11188
rect 22224 11108 22244 11172
rect 22308 11108 22328 11172
rect 22224 11092 22328 11108
rect 22224 11028 22244 11092
rect 22308 11028 22328 11092
rect 22224 11012 22328 11028
rect 22224 10948 22244 11012
rect 22308 10948 22328 11012
rect 22224 10932 22328 10948
rect 22224 10868 22244 10932
rect 22308 10868 22328 10932
rect 22224 10852 22328 10868
rect 16612 10492 16716 10788
rect 11000 10412 11104 10428
rect 11000 10348 11020 10412
rect 11084 10348 11104 10412
rect 11000 10332 11104 10348
rect 11000 10268 11020 10332
rect 11084 10268 11104 10332
rect 11000 10252 11104 10268
rect 11000 10188 11020 10252
rect 11084 10188 11104 10252
rect 11000 10172 11104 10188
rect 11000 10108 11020 10172
rect 11084 10108 11104 10172
rect 11000 10092 11104 10108
rect 11000 10028 11020 10092
rect 11084 10028 11104 10092
rect 11000 10012 11104 10028
rect 11000 9948 11020 10012
rect 11084 9948 11104 10012
rect 11000 9932 11104 9948
rect 11000 9868 11020 9932
rect 11084 9868 11104 9932
rect 11000 9852 11104 9868
rect 11000 9788 11020 9852
rect 11084 9788 11104 9852
rect 11000 9772 11104 9788
rect 11000 9708 11020 9772
rect 11084 9708 11104 9772
rect 11000 9692 11104 9708
rect 11000 9628 11020 9692
rect 11084 9628 11104 9692
rect 11000 9612 11104 9628
rect 11000 9548 11020 9612
rect 11084 9548 11104 9612
rect 11000 9532 11104 9548
rect 11000 9468 11020 9532
rect 11084 9468 11104 9532
rect 11000 9452 11104 9468
rect 11000 9388 11020 9452
rect 11084 9388 11104 9452
rect 11000 9372 11104 9388
rect 11000 9308 11020 9372
rect 11084 9308 11104 9372
rect 11000 9292 11104 9308
rect 11000 9228 11020 9292
rect 11084 9228 11104 9292
rect 11000 9212 11104 9228
rect 11000 9148 11020 9212
rect 11084 9148 11104 9212
rect 11000 9132 11104 9148
rect 11000 9068 11020 9132
rect 11084 9068 11104 9132
rect 11000 9052 11104 9068
rect 11000 8988 11020 9052
rect 11084 8988 11104 9052
rect 11000 8972 11104 8988
rect 11000 8908 11020 8972
rect 11084 8908 11104 8972
rect 11000 8892 11104 8908
rect 11000 8828 11020 8892
rect 11084 8828 11104 8892
rect 11000 8812 11104 8828
rect 11000 8748 11020 8812
rect 11084 8748 11104 8812
rect 11000 8732 11104 8748
rect 11000 8668 11020 8732
rect 11084 8668 11104 8732
rect 11000 8652 11104 8668
rect 11000 8588 11020 8652
rect 11084 8588 11104 8652
rect 11000 8572 11104 8588
rect 11000 8508 11020 8572
rect 11084 8508 11104 8572
rect 11000 8492 11104 8508
rect 11000 8428 11020 8492
rect 11084 8428 11104 8492
rect 11000 8412 11104 8428
rect 11000 8348 11020 8412
rect 11084 8348 11104 8412
rect 11000 8332 11104 8348
rect 11000 8268 11020 8332
rect 11084 8268 11104 8332
rect 11000 8252 11104 8268
rect 11000 8188 11020 8252
rect 11084 8188 11104 8252
rect 11000 8172 11104 8188
rect 11000 8108 11020 8172
rect 11084 8108 11104 8172
rect 11000 8092 11104 8108
rect 11000 8028 11020 8092
rect 11084 8028 11104 8092
rect 11000 8012 11104 8028
rect 11000 7948 11020 8012
rect 11084 7948 11104 8012
rect 11000 7932 11104 7948
rect 11000 7868 11020 7932
rect 11084 7868 11104 7932
rect 11000 7852 11104 7868
rect 11000 7788 11020 7852
rect 11084 7788 11104 7852
rect 11000 7772 11104 7788
rect 11000 7708 11020 7772
rect 11084 7708 11104 7772
rect 11000 7692 11104 7708
rect 11000 7628 11020 7692
rect 11084 7628 11104 7692
rect 11000 7612 11104 7628
rect 11000 7548 11020 7612
rect 11084 7548 11104 7612
rect 11000 7532 11104 7548
rect 11000 7468 11020 7532
rect 11084 7468 11104 7532
rect 11000 7452 11104 7468
rect 11000 7388 11020 7452
rect 11084 7388 11104 7452
rect 11000 7372 11104 7388
rect 11000 7308 11020 7372
rect 11084 7308 11104 7372
rect 11000 7292 11104 7308
rect 11000 7228 11020 7292
rect 11084 7228 11104 7292
rect 11000 7212 11104 7228
rect 11000 7148 11020 7212
rect 11084 7148 11104 7212
rect 11000 7132 11104 7148
rect 11000 7068 11020 7132
rect 11084 7068 11104 7132
rect 11000 7052 11104 7068
rect 11000 6988 11020 7052
rect 11084 6988 11104 7052
rect 11000 6972 11104 6988
rect 11000 6908 11020 6972
rect 11084 6908 11104 6972
rect 11000 6892 11104 6908
rect 11000 6828 11020 6892
rect 11084 6828 11104 6892
rect 11000 6812 11104 6828
rect 11000 6748 11020 6812
rect 11084 6748 11104 6812
rect 11000 6732 11104 6748
rect 11000 6668 11020 6732
rect 11084 6668 11104 6732
rect 11000 6652 11104 6668
rect 11000 6588 11020 6652
rect 11084 6588 11104 6652
rect 11000 6572 11104 6588
rect 11000 6508 11020 6572
rect 11084 6508 11104 6572
rect 11000 6492 11104 6508
rect 11000 6428 11020 6492
rect 11084 6428 11104 6492
rect 11000 6412 11104 6428
rect 11000 6348 11020 6412
rect 11084 6348 11104 6412
rect 11000 6332 11104 6348
rect 11000 6268 11020 6332
rect 11084 6268 11104 6332
rect 11000 6252 11104 6268
rect 11000 6188 11020 6252
rect 11084 6188 11104 6252
rect 11000 6172 11104 6188
rect 11000 6108 11020 6172
rect 11084 6108 11104 6172
rect 11000 6092 11104 6108
rect 11000 6028 11020 6092
rect 11084 6028 11104 6092
rect 11000 6012 11104 6028
rect 11000 5948 11020 6012
rect 11084 5948 11104 6012
rect 11000 5932 11104 5948
rect 11000 5868 11020 5932
rect 11084 5868 11104 5932
rect 11000 5852 11104 5868
rect 11000 5788 11020 5852
rect 11084 5788 11104 5852
rect 11000 5772 11104 5788
rect 11000 5708 11020 5772
rect 11084 5708 11104 5772
rect 11000 5692 11104 5708
rect 11000 5628 11020 5692
rect 11084 5628 11104 5692
rect 11000 5612 11104 5628
rect 11000 5548 11020 5612
rect 11084 5548 11104 5612
rect 11000 5532 11104 5548
rect 5388 5172 5492 5468
rect -224 5092 -120 5108
rect -224 5028 -204 5092
rect -140 5028 -120 5092
rect -224 5012 -120 5028
rect -224 4948 -204 5012
rect -140 4948 -120 5012
rect -224 4932 -120 4948
rect -224 4868 -204 4932
rect -140 4868 -120 4932
rect -224 4852 -120 4868
rect -224 4788 -204 4852
rect -140 4788 -120 4852
rect -224 4772 -120 4788
rect -224 4708 -204 4772
rect -140 4708 -120 4772
rect -224 4692 -120 4708
rect -224 4628 -204 4692
rect -140 4628 -120 4692
rect -224 4612 -120 4628
rect -224 4548 -204 4612
rect -140 4548 -120 4612
rect -224 4532 -120 4548
rect -224 4468 -204 4532
rect -140 4468 -120 4532
rect -224 4452 -120 4468
rect -224 4388 -204 4452
rect -140 4388 -120 4452
rect -224 4372 -120 4388
rect -224 4308 -204 4372
rect -140 4308 -120 4372
rect -224 4292 -120 4308
rect -224 4228 -204 4292
rect -140 4228 -120 4292
rect -224 4212 -120 4228
rect -224 4148 -204 4212
rect -140 4148 -120 4212
rect -224 4132 -120 4148
rect -224 4068 -204 4132
rect -140 4068 -120 4132
rect -224 4052 -120 4068
rect -224 3988 -204 4052
rect -140 3988 -120 4052
rect -224 3972 -120 3988
rect -224 3908 -204 3972
rect -140 3908 -120 3972
rect -224 3892 -120 3908
rect -224 3828 -204 3892
rect -140 3828 -120 3892
rect -224 3812 -120 3828
rect -224 3748 -204 3812
rect -140 3748 -120 3812
rect -224 3732 -120 3748
rect -224 3668 -204 3732
rect -140 3668 -120 3732
rect -224 3652 -120 3668
rect -224 3588 -204 3652
rect -140 3588 -120 3652
rect -224 3572 -120 3588
rect -224 3508 -204 3572
rect -140 3508 -120 3572
rect -224 3492 -120 3508
rect -224 3428 -204 3492
rect -140 3428 -120 3492
rect -224 3412 -120 3428
rect -224 3348 -204 3412
rect -140 3348 -120 3412
rect -224 3332 -120 3348
rect -224 3268 -204 3332
rect -140 3268 -120 3332
rect -224 3252 -120 3268
rect -224 3188 -204 3252
rect -140 3188 -120 3252
rect -224 3172 -120 3188
rect -224 3108 -204 3172
rect -140 3108 -120 3172
rect -224 3092 -120 3108
rect -224 3028 -204 3092
rect -140 3028 -120 3092
rect -224 3012 -120 3028
rect -224 2948 -204 3012
rect -140 2948 -120 3012
rect -224 2932 -120 2948
rect -224 2868 -204 2932
rect -140 2868 -120 2932
rect -224 2852 -120 2868
rect -224 2788 -204 2852
rect -140 2788 -120 2852
rect -224 2772 -120 2788
rect -224 2708 -204 2772
rect -140 2708 -120 2772
rect -224 2692 -120 2708
rect -224 2628 -204 2692
rect -140 2628 -120 2692
rect -224 2612 -120 2628
rect -224 2548 -204 2612
rect -140 2548 -120 2612
rect -224 2532 -120 2548
rect -224 2468 -204 2532
rect -140 2468 -120 2532
rect -224 2452 -120 2468
rect -224 2388 -204 2452
rect -140 2388 -120 2452
rect -224 2372 -120 2388
rect -224 2308 -204 2372
rect -140 2308 -120 2372
rect -224 2292 -120 2308
rect -224 2228 -204 2292
rect -140 2228 -120 2292
rect -224 2212 -120 2228
rect -224 2148 -204 2212
rect -140 2148 -120 2212
rect -224 2132 -120 2148
rect -224 2068 -204 2132
rect -140 2068 -120 2132
rect -224 2052 -120 2068
rect -224 1988 -204 2052
rect -140 1988 -120 2052
rect -224 1972 -120 1988
rect -224 1908 -204 1972
rect -140 1908 -120 1972
rect -224 1892 -120 1908
rect -224 1828 -204 1892
rect -140 1828 -120 1892
rect -224 1812 -120 1828
rect -224 1748 -204 1812
rect -140 1748 -120 1812
rect -224 1732 -120 1748
rect -224 1668 -204 1732
rect -140 1668 -120 1732
rect -224 1652 -120 1668
rect -224 1588 -204 1652
rect -140 1588 -120 1652
rect -224 1572 -120 1588
rect -224 1508 -204 1572
rect -140 1508 -120 1572
rect -224 1492 -120 1508
rect -224 1428 -204 1492
rect -140 1428 -120 1492
rect -224 1412 -120 1428
rect -224 1348 -204 1412
rect -140 1348 -120 1412
rect -224 1332 -120 1348
rect -224 1268 -204 1332
rect -140 1268 -120 1332
rect -224 1252 -120 1268
rect -224 1188 -204 1252
rect -140 1188 -120 1252
rect -224 1172 -120 1188
rect -224 1108 -204 1172
rect -140 1108 -120 1172
rect -224 1092 -120 1108
rect -224 1028 -204 1092
rect -140 1028 -120 1092
rect -224 1012 -120 1028
rect -224 948 -204 1012
rect -140 948 -120 1012
rect -224 932 -120 948
rect -224 868 -204 932
rect -140 868 -120 932
rect -224 852 -120 868
rect -224 788 -204 852
rect -140 788 -120 852
rect -224 772 -120 788
rect -224 708 -204 772
rect -140 708 -120 772
rect -224 692 -120 708
rect -224 628 -204 692
rect -140 628 -120 692
rect -224 612 -120 628
rect -224 548 -204 612
rect -140 548 -120 612
rect -224 532 -120 548
rect -224 468 -204 532
rect -140 468 -120 532
rect -224 452 -120 468
rect -224 388 -204 452
rect -140 388 -120 452
rect -224 372 -120 388
rect -224 308 -204 372
rect -140 308 -120 372
rect -224 292 -120 308
rect -224 228 -204 292
rect -140 228 -120 292
rect -224 212 -120 228
rect -5836 -148 -5732 148
rect -11448 -228 -11344 -212
rect -11448 -292 -11428 -228
rect -11364 -292 -11344 -228
rect -11448 -308 -11344 -292
rect -11448 -372 -11428 -308
rect -11364 -372 -11344 -308
rect -11448 -388 -11344 -372
rect -11448 -452 -11428 -388
rect -11364 -452 -11344 -388
rect -11448 -468 -11344 -452
rect -11448 -532 -11428 -468
rect -11364 -532 -11344 -468
rect -11448 -548 -11344 -532
rect -11448 -612 -11428 -548
rect -11364 -612 -11344 -548
rect -11448 -628 -11344 -612
rect -11448 -692 -11428 -628
rect -11364 -692 -11344 -628
rect -11448 -708 -11344 -692
rect -11448 -772 -11428 -708
rect -11364 -772 -11344 -708
rect -11448 -788 -11344 -772
rect -11448 -852 -11428 -788
rect -11364 -852 -11344 -788
rect -11448 -868 -11344 -852
rect -11448 -932 -11428 -868
rect -11364 -932 -11344 -868
rect -11448 -948 -11344 -932
rect -11448 -1012 -11428 -948
rect -11364 -1012 -11344 -948
rect -11448 -1028 -11344 -1012
rect -11448 -1092 -11428 -1028
rect -11364 -1092 -11344 -1028
rect -11448 -1108 -11344 -1092
rect -11448 -1172 -11428 -1108
rect -11364 -1172 -11344 -1108
rect -11448 -1188 -11344 -1172
rect -11448 -1252 -11428 -1188
rect -11364 -1252 -11344 -1188
rect -11448 -1268 -11344 -1252
rect -11448 -1332 -11428 -1268
rect -11364 -1332 -11344 -1268
rect -11448 -1348 -11344 -1332
rect -11448 -1412 -11428 -1348
rect -11364 -1412 -11344 -1348
rect -11448 -1428 -11344 -1412
rect -11448 -1492 -11428 -1428
rect -11364 -1492 -11344 -1428
rect -11448 -1508 -11344 -1492
rect -11448 -1572 -11428 -1508
rect -11364 -1572 -11344 -1508
rect -11448 -1588 -11344 -1572
rect -11448 -1652 -11428 -1588
rect -11364 -1652 -11344 -1588
rect -11448 -1668 -11344 -1652
rect -11448 -1732 -11428 -1668
rect -11364 -1732 -11344 -1668
rect -11448 -1748 -11344 -1732
rect -11448 -1812 -11428 -1748
rect -11364 -1812 -11344 -1748
rect -11448 -1828 -11344 -1812
rect -11448 -1892 -11428 -1828
rect -11364 -1892 -11344 -1828
rect -11448 -1908 -11344 -1892
rect -11448 -1972 -11428 -1908
rect -11364 -1972 -11344 -1908
rect -11448 -1988 -11344 -1972
rect -11448 -2052 -11428 -1988
rect -11364 -2052 -11344 -1988
rect -11448 -2068 -11344 -2052
rect -11448 -2132 -11428 -2068
rect -11364 -2132 -11344 -2068
rect -11448 -2148 -11344 -2132
rect -11448 -2212 -11428 -2148
rect -11364 -2212 -11344 -2148
rect -11448 -2228 -11344 -2212
rect -11448 -2292 -11428 -2228
rect -11364 -2292 -11344 -2228
rect -11448 -2308 -11344 -2292
rect -11448 -2372 -11428 -2308
rect -11364 -2372 -11344 -2308
rect -11448 -2388 -11344 -2372
rect -11448 -2452 -11428 -2388
rect -11364 -2452 -11344 -2388
rect -11448 -2468 -11344 -2452
rect -11448 -2532 -11428 -2468
rect -11364 -2532 -11344 -2468
rect -11448 -2548 -11344 -2532
rect -11448 -2612 -11428 -2548
rect -11364 -2612 -11344 -2548
rect -11448 -2628 -11344 -2612
rect -11448 -2692 -11428 -2628
rect -11364 -2692 -11344 -2628
rect -11448 -2708 -11344 -2692
rect -11448 -2772 -11428 -2708
rect -11364 -2772 -11344 -2708
rect -11448 -2788 -11344 -2772
rect -11448 -2852 -11428 -2788
rect -11364 -2852 -11344 -2788
rect -11448 -2868 -11344 -2852
rect -11448 -2932 -11428 -2868
rect -11364 -2932 -11344 -2868
rect -11448 -2948 -11344 -2932
rect -11448 -3012 -11428 -2948
rect -11364 -3012 -11344 -2948
rect -11448 -3028 -11344 -3012
rect -11448 -3092 -11428 -3028
rect -11364 -3092 -11344 -3028
rect -11448 -3108 -11344 -3092
rect -11448 -3172 -11428 -3108
rect -11364 -3172 -11344 -3108
rect -11448 -3188 -11344 -3172
rect -11448 -3252 -11428 -3188
rect -11364 -3252 -11344 -3188
rect -11448 -3268 -11344 -3252
rect -11448 -3332 -11428 -3268
rect -11364 -3332 -11344 -3268
rect -11448 -3348 -11344 -3332
rect -11448 -3412 -11428 -3348
rect -11364 -3412 -11344 -3348
rect -11448 -3428 -11344 -3412
rect -11448 -3492 -11428 -3428
rect -11364 -3492 -11344 -3428
rect -11448 -3508 -11344 -3492
rect -11448 -3572 -11428 -3508
rect -11364 -3572 -11344 -3508
rect -11448 -3588 -11344 -3572
rect -11448 -3652 -11428 -3588
rect -11364 -3652 -11344 -3588
rect -11448 -3668 -11344 -3652
rect -11448 -3732 -11428 -3668
rect -11364 -3732 -11344 -3668
rect -11448 -3748 -11344 -3732
rect -11448 -3812 -11428 -3748
rect -11364 -3812 -11344 -3748
rect -11448 -3828 -11344 -3812
rect -11448 -3892 -11428 -3828
rect -11364 -3892 -11344 -3828
rect -11448 -3908 -11344 -3892
rect -11448 -3972 -11428 -3908
rect -11364 -3972 -11344 -3908
rect -11448 -3988 -11344 -3972
rect -11448 -4052 -11428 -3988
rect -11364 -4052 -11344 -3988
rect -11448 -4068 -11344 -4052
rect -11448 -4132 -11428 -4068
rect -11364 -4132 -11344 -4068
rect -11448 -4148 -11344 -4132
rect -11448 -4212 -11428 -4148
rect -11364 -4212 -11344 -4148
rect -11448 -4228 -11344 -4212
rect -11448 -4292 -11428 -4228
rect -11364 -4292 -11344 -4228
rect -11448 -4308 -11344 -4292
rect -11448 -4372 -11428 -4308
rect -11364 -4372 -11344 -4308
rect -11448 -4388 -11344 -4372
rect -11448 -4452 -11428 -4388
rect -11364 -4452 -11344 -4388
rect -11448 -4468 -11344 -4452
rect -11448 -4532 -11428 -4468
rect -11364 -4532 -11344 -4468
rect -11448 -4548 -11344 -4532
rect -11448 -4612 -11428 -4548
rect -11364 -4612 -11344 -4548
rect -11448 -4628 -11344 -4612
rect -11448 -4692 -11428 -4628
rect -11364 -4692 -11344 -4628
rect -11448 -4708 -11344 -4692
rect -11448 -4772 -11428 -4708
rect -11364 -4772 -11344 -4708
rect -11448 -4788 -11344 -4772
rect -11448 -4852 -11428 -4788
rect -11364 -4852 -11344 -4788
rect -11448 -4868 -11344 -4852
rect -11448 -4932 -11428 -4868
rect -11364 -4932 -11344 -4868
rect -11448 -4948 -11344 -4932
rect -11448 -5012 -11428 -4948
rect -11364 -5012 -11344 -4948
rect -11448 -5028 -11344 -5012
rect -11448 -5092 -11428 -5028
rect -11364 -5092 -11344 -5028
rect -11448 -5108 -11344 -5092
rect -17060 -5468 -16956 -5172
rect -22672 -5548 -22568 -5532
rect -22672 -5612 -22652 -5548
rect -22588 -5612 -22568 -5548
rect -22672 -5628 -22568 -5612
rect -22672 -5692 -22652 -5628
rect -22588 -5692 -22568 -5628
rect -22672 -5708 -22568 -5692
rect -22672 -5772 -22652 -5708
rect -22588 -5772 -22568 -5708
rect -22672 -5788 -22568 -5772
rect -22672 -5852 -22652 -5788
rect -22588 -5852 -22568 -5788
rect -22672 -5868 -22568 -5852
rect -22672 -5932 -22652 -5868
rect -22588 -5932 -22568 -5868
rect -22672 -5948 -22568 -5932
rect -22672 -6012 -22652 -5948
rect -22588 -6012 -22568 -5948
rect -22672 -6028 -22568 -6012
rect -22672 -6092 -22652 -6028
rect -22588 -6092 -22568 -6028
rect -22672 -6108 -22568 -6092
rect -22672 -6172 -22652 -6108
rect -22588 -6172 -22568 -6108
rect -22672 -6188 -22568 -6172
rect -22672 -6252 -22652 -6188
rect -22588 -6252 -22568 -6188
rect -22672 -6268 -22568 -6252
rect -22672 -6332 -22652 -6268
rect -22588 -6332 -22568 -6268
rect -22672 -6348 -22568 -6332
rect -22672 -6412 -22652 -6348
rect -22588 -6412 -22568 -6348
rect -22672 -6428 -22568 -6412
rect -22672 -6492 -22652 -6428
rect -22588 -6492 -22568 -6428
rect -22672 -6508 -22568 -6492
rect -22672 -6572 -22652 -6508
rect -22588 -6572 -22568 -6508
rect -22672 -6588 -22568 -6572
rect -22672 -6652 -22652 -6588
rect -22588 -6652 -22568 -6588
rect -22672 -6668 -22568 -6652
rect -22672 -6732 -22652 -6668
rect -22588 -6732 -22568 -6668
rect -22672 -6748 -22568 -6732
rect -22672 -6812 -22652 -6748
rect -22588 -6812 -22568 -6748
rect -22672 -6828 -22568 -6812
rect -22672 -6892 -22652 -6828
rect -22588 -6892 -22568 -6828
rect -22672 -6908 -22568 -6892
rect -22672 -6972 -22652 -6908
rect -22588 -6972 -22568 -6908
rect -22672 -6988 -22568 -6972
rect -22672 -7052 -22652 -6988
rect -22588 -7052 -22568 -6988
rect -22672 -7068 -22568 -7052
rect -22672 -7132 -22652 -7068
rect -22588 -7132 -22568 -7068
rect -22672 -7148 -22568 -7132
rect -22672 -7212 -22652 -7148
rect -22588 -7212 -22568 -7148
rect -22672 -7228 -22568 -7212
rect -22672 -7292 -22652 -7228
rect -22588 -7292 -22568 -7228
rect -22672 -7308 -22568 -7292
rect -22672 -7372 -22652 -7308
rect -22588 -7372 -22568 -7308
rect -22672 -7388 -22568 -7372
rect -22672 -7452 -22652 -7388
rect -22588 -7452 -22568 -7388
rect -22672 -7468 -22568 -7452
rect -22672 -7532 -22652 -7468
rect -22588 -7532 -22568 -7468
rect -22672 -7548 -22568 -7532
rect -22672 -7612 -22652 -7548
rect -22588 -7612 -22568 -7548
rect -22672 -7628 -22568 -7612
rect -22672 -7692 -22652 -7628
rect -22588 -7692 -22568 -7628
rect -22672 -7708 -22568 -7692
rect -22672 -7772 -22652 -7708
rect -22588 -7772 -22568 -7708
rect -22672 -7788 -22568 -7772
rect -22672 -7852 -22652 -7788
rect -22588 -7852 -22568 -7788
rect -22672 -7868 -22568 -7852
rect -22672 -7932 -22652 -7868
rect -22588 -7932 -22568 -7868
rect -22672 -7948 -22568 -7932
rect -22672 -8012 -22652 -7948
rect -22588 -8012 -22568 -7948
rect -22672 -8028 -22568 -8012
rect -22672 -8092 -22652 -8028
rect -22588 -8092 -22568 -8028
rect -22672 -8108 -22568 -8092
rect -22672 -8172 -22652 -8108
rect -22588 -8172 -22568 -8108
rect -22672 -8188 -22568 -8172
rect -22672 -8252 -22652 -8188
rect -22588 -8252 -22568 -8188
rect -22672 -8268 -22568 -8252
rect -22672 -8332 -22652 -8268
rect -22588 -8332 -22568 -8268
rect -22672 -8348 -22568 -8332
rect -22672 -8412 -22652 -8348
rect -22588 -8412 -22568 -8348
rect -22672 -8428 -22568 -8412
rect -22672 -8492 -22652 -8428
rect -22588 -8492 -22568 -8428
rect -22672 -8508 -22568 -8492
rect -22672 -8572 -22652 -8508
rect -22588 -8572 -22568 -8508
rect -22672 -8588 -22568 -8572
rect -22672 -8652 -22652 -8588
rect -22588 -8652 -22568 -8588
rect -22672 -8668 -22568 -8652
rect -22672 -8732 -22652 -8668
rect -22588 -8732 -22568 -8668
rect -22672 -8748 -22568 -8732
rect -22672 -8812 -22652 -8748
rect -22588 -8812 -22568 -8748
rect -22672 -8828 -22568 -8812
rect -22672 -8892 -22652 -8828
rect -22588 -8892 -22568 -8828
rect -22672 -8908 -22568 -8892
rect -22672 -8972 -22652 -8908
rect -22588 -8972 -22568 -8908
rect -22672 -8988 -22568 -8972
rect -22672 -9052 -22652 -8988
rect -22588 -9052 -22568 -8988
rect -22672 -9068 -22568 -9052
rect -22672 -9132 -22652 -9068
rect -22588 -9132 -22568 -9068
rect -22672 -9148 -22568 -9132
rect -22672 -9212 -22652 -9148
rect -22588 -9212 -22568 -9148
rect -22672 -9228 -22568 -9212
rect -22672 -9292 -22652 -9228
rect -22588 -9292 -22568 -9228
rect -22672 -9308 -22568 -9292
rect -22672 -9372 -22652 -9308
rect -22588 -9372 -22568 -9308
rect -22672 -9388 -22568 -9372
rect -22672 -9452 -22652 -9388
rect -22588 -9452 -22568 -9388
rect -22672 -9468 -22568 -9452
rect -22672 -9532 -22652 -9468
rect -22588 -9532 -22568 -9468
rect -22672 -9548 -22568 -9532
rect -22672 -9612 -22652 -9548
rect -22588 -9612 -22568 -9548
rect -22672 -9628 -22568 -9612
rect -22672 -9692 -22652 -9628
rect -22588 -9692 -22568 -9628
rect -22672 -9708 -22568 -9692
rect -22672 -9772 -22652 -9708
rect -22588 -9772 -22568 -9708
rect -22672 -9788 -22568 -9772
rect -22672 -9852 -22652 -9788
rect -22588 -9852 -22568 -9788
rect -22672 -9868 -22568 -9852
rect -22672 -9932 -22652 -9868
rect -22588 -9932 -22568 -9868
rect -22672 -9948 -22568 -9932
rect -22672 -10012 -22652 -9948
rect -22588 -10012 -22568 -9948
rect -22672 -10028 -22568 -10012
rect -22672 -10092 -22652 -10028
rect -22588 -10092 -22568 -10028
rect -22672 -10108 -22568 -10092
rect -22672 -10172 -22652 -10108
rect -22588 -10172 -22568 -10108
rect -22672 -10188 -22568 -10172
rect -22672 -10252 -22652 -10188
rect -22588 -10252 -22568 -10188
rect -22672 -10268 -22568 -10252
rect -22672 -10332 -22652 -10268
rect -22588 -10332 -22568 -10268
rect -22672 -10348 -22568 -10332
rect -22672 -10412 -22652 -10348
rect -22588 -10412 -22568 -10348
rect -22672 -10428 -22568 -10412
rect -28284 -10788 -28180 -10492
rect -33896 -10868 -33792 -10852
rect -33896 -10932 -33876 -10868
rect -33812 -10932 -33792 -10868
rect -33896 -10948 -33792 -10932
rect -33896 -11012 -33876 -10948
rect -33812 -11012 -33792 -10948
rect -33896 -11028 -33792 -11012
rect -33896 -11092 -33876 -11028
rect -33812 -11092 -33792 -11028
rect -33896 -11108 -33792 -11092
rect -33896 -11172 -33876 -11108
rect -33812 -11172 -33792 -11108
rect -33896 -11188 -33792 -11172
rect -33896 -11252 -33876 -11188
rect -33812 -11252 -33792 -11188
rect -33896 -11268 -33792 -11252
rect -33896 -11332 -33876 -11268
rect -33812 -11332 -33792 -11268
rect -33896 -11348 -33792 -11332
rect -33896 -11412 -33876 -11348
rect -33812 -11412 -33792 -11348
rect -33896 -11428 -33792 -11412
rect -33896 -11492 -33876 -11428
rect -33812 -11492 -33792 -11428
rect -33896 -11508 -33792 -11492
rect -33896 -11572 -33876 -11508
rect -33812 -11572 -33792 -11508
rect -33896 -11588 -33792 -11572
rect -33896 -11652 -33876 -11588
rect -33812 -11652 -33792 -11588
rect -33896 -11668 -33792 -11652
rect -33896 -11732 -33876 -11668
rect -33812 -11732 -33792 -11668
rect -33896 -11748 -33792 -11732
rect -33896 -11812 -33876 -11748
rect -33812 -11812 -33792 -11748
rect -33896 -11828 -33792 -11812
rect -33896 -11892 -33876 -11828
rect -33812 -11892 -33792 -11828
rect -33896 -11908 -33792 -11892
rect -33896 -11972 -33876 -11908
rect -33812 -11972 -33792 -11908
rect -33896 -11988 -33792 -11972
rect -33896 -12052 -33876 -11988
rect -33812 -12052 -33792 -11988
rect -33896 -12068 -33792 -12052
rect -33896 -12132 -33876 -12068
rect -33812 -12132 -33792 -12068
rect -33896 -12148 -33792 -12132
rect -33896 -12212 -33876 -12148
rect -33812 -12212 -33792 -12148
rect -33896 -12228 -33792 -12212
rect -33896 -12292 -33876 -12228
rect -33812 -12292 -33792 -12228
rect -33896 -12308 -33792 -12292
rect -33896 -12372 -33876 -12308
rect -33812 -12372 -33792 -12308
rect -33896 -12388 -33792 -12372
rect -33896 -12452 -33876 -12388
rect -33812 -12452 -33792 -12388
rect -33896 -12468 -33792 -12452
rect -33896 -12532 -33876 -12468
rect -33812 -12532 -33792 -12468
rect -33896 -12548 -33792 -12532
rect -33896 -12612 -33876 -12548
rect -33812 -12612 -33792 -12548
rect -33896 -12628 -33792 -12612
rect -33896 -12692 -33876 -12628
rect -33812 -12692 -33792 -12628
rect -33896 -12708 -33792 -12692
rect -33896 -12772 -33876 -12708
rect -33812 -12772 -33792 -12708
rect -33896 -12788 -33792 -12772
rect -33896 -12852 -33876 -12788
rect -33812 -12852 -33792 -12788
rect -33896 -12868 -33792 -12852
rect -33896 -12932 -33876 -12868
rect -33812 -12932 -33792 -12868
rect -33896 -12948 -33792 -12932
rect -33896 -13012 -33876 -12948
rect -33812 -13012 -33792 -12948
rect -33896 -13028 -33792 -13012
rect -33896 -13092 -33876 -13028
rect -33812 -13092 -33792 -13028
rect -33896 -13108 -33792 -13092
rect -33896 -13172 -33876 -13108
rect -33812 -13172 -33792 -13108
rect -33896 -13188 -33792 -13172
rect -33896 -13252 -33876 -13188
rect -33812 -13252 -33792 -13188
rect -33896 -13268 -33792 -13252
rect -33896 -13332 -33876 -13268
rect -33812 -13332 -33792 -13268
rect -33896 -13348 -33792 -13332
rect -33896 -13412 -33876 -13348
rect -33812 -13412 -33792 -13348
rect -33896 -13428 -33792 -13412
rect -33896 -13492 -33876 -13428
rect -33812 -13492 -33792 -13428
rect -33896 -13508 -33792 -13492
rect -33896 -13572 -33876 -13508
rect -33812 -13572 -33792 -13508
rect -33896 -13588 -33792 -13572
rect -33896 -13652 -33876 -13588
rect -33812 -13652 -33792 -13588
rect -33896 -13668 -33792 -13652
rect -33896 -13732 -33876 -13668
rect -33812 -13732 -33792 -13668
rect -33896 -13748 -33792 -13732
rect -33896 -13812 -33876 -13748
rect -33812 -13812 -33792 -13748
rect -33896 -13828 -33792 -13812
rect -33896 -13892 -33876 -13828
rect -33812 -13892 -33792 -13828
rect -33896 -13908 -33792 -13892
rect -33896 -13972 -33876 -13908
rect -33812 -13972 -33792 -13908
rect -33896 -13988 -33792 -13972
rect -33896 -14052 -33876 -13988
rect -33812 -14052 -33792 -13988
rect -33896 -14068 -33792 -14052
rect -33896 -14132 -33876 -14068
rect -33812 -14132 -33792 -14068
rect -33896 -14148 -33792 -14132
rect -33896 -14212 -33876 -14148
rect -33812 -14212 -33792 -14148
rect -33896 -14228 -33792 -14212
rect -33896 -14292 -33876 -14228
rect -33812 -14292 -33792 -14228
rect -33896 -14308 -33792 -14292
rect -33896 -14372 -33876 -14308
rect -33812 -14372 -33792 -14308
rect -33896 -14388 -33792 -14372
rect -33896 -14452 -33876 -14388
rect -33812 -14452 -33792 -14388
rect -33896 -14468 -33792 -14452
rect -33896 -14532 -33876 -14468
rect -33812 -14532 -33792 -14468
rect -33896 -14548 -33792 -14532
rect -33896 -14612 -33876 -14548
rect -33812 -14612 -33792 -14548
rect -33896 -14628 -33792 -14612
rect -33896 -14692 -33876 -14628
rect -33812 -14692 -33792 -14628
rect -33896 -14708 -33792 -14692
rect -33896 -14772 -33876 -14708
rect -33812 -14772 -33792 -14708
rect -33896 -14788 -33792 -14772
rect -33896 -14852 -33876 -14788
rect -33812 -14852 -33792 -14788
rect -33896 -14868 -33792 -14852
rect -33896 -14932 -33876 -14868
rect -33812 -14932 -33792 -14868
rect -33896 -14948 -33792 -14932
rect -33896 -15012 -33876 -14948
rect -33812 -15012 -33792 -14948
rect -33896 -15028 -33792 -15012
rect -33896 -15092 -33876 -15028
rect -33812 -15092 -33792 -15028
rect -33896 -15108 -33792 -15092
rect -33896 -15172 -33876 -15108
rect -33812 -15172 -33792 -15108
rect -33896 -15188 -33792 -15172
rect -33896 -15252 -33876 -15188
rect -33812 -15252 -33792 -15188
rect -33896 -15268 -33792 -15252
rect -33896 -15332 -33876 -15268
rect -33812 -15332 -33792 -15268
rect -33896 -15348 -33792 -15332
rect -33896 -15412 -33876 -15348
rect -33812 -15412 -33792 -15348
rect -33896 -15428 -33792 -15412
rect -33896 -15492 -33876 -15428
rect -33812 -15492 -33792 -15428
rect -33896 -15508 -33792 -15492
rect -33896 -15572 -33876 -15508
rect -33812 -15572 -33792 -15508
rect -33896 -15588 -33792 -15572
rect -33896 -15652 -33876 -15588
rect -33812 -15652 -33792 -15588
rect -33896 -15668 -33792 -15652
rect -33896 -15732 -33876 -15668
rect -33812 -15732 -33792 -15668
rect -33896 -15748 -33792 -15732
rect -36676 -16159 -36572 -15761
rect -33896 -15812 -33876 -15748
rect -33812 -15812 -33792 -15748
rect -33473 -10868 -28551 -10839
rect -33473 -15732 -33444 -10868
rect -28580 -15732 -28551 -10868
rect -33473 -15761 -28551 -15732
rect -28284 -10852 -28264 -10788
rect -28200 -10852 -28180 -10788
rect -25452 -10839 -25348 -10441
rect -22672 -10492 -22652 -10428
rect -22588 -10492 -22568 -10428
rect -22249 -5548 -17327 -5519
rect -22249 -10412 -22220 -5548
rect -17356 -10412 -17327 -5548
rect -22249 -10441 -17327 -10412
rect -17060 -5532 -17040 -5468
rect -16976 -5532 -16956 -5468
rect -14228 -5519 -14124 -5121
rect -11448 -5172 -11428 -5108
rect -11364 -5172 -11344 -5108
rect -11025 -228 -6103 -199
rect -11025 -5092 -10996 -228
rect -6132 -5092 -6103 -228
rect -11025 -5121 -6103 -5092
rect -5836 -212 -5816 -148
rect -5752 -212 -5732 -148
rect -3004 -199 -2900 199
rect -224 148 -204 212
rect -140 148 -120 212
rect 199 5092 5121 5121
rect 199 228 228 5092
rect 5092 228 5121 5092
rect 199 199 5121 228
rect 5388 5108 5408 5172
rect 5472 5108 5492 5172
rect 8220 5121 8324 5519
rect 11000 5468 11020 5532
rect 11084 5468 11104 5532
rect 11423 10412 16345 10441
rect 11423 5548 11452 10412
rect 16316 5548 16345 10412
rect 11423 5519 16345 5548
rect 16612 10428 16632 10492
rect 16696 10428 16716 10492
rect 19444 10441 19548 10839
rect 22224 10788 22244 10852
rect 22308 10788 22328 10852
rect 22647 15732 27569 15761
rect 22647 10868 22676 15732
rect 27540 10868 27569 15732
rect 22647 10839 27569 10868
rect 27836 15748 27856 15812
rect 27920 15748 27940 15812
rect 30668 15761 30772 16159
rect 33448 16108 33468 16172
rect 33532 16108 33552 16172
rect 33871 21052 38793 21081
rect 33871 16188 33900 21052
rect 38764 16188 38793 21052
rect 33871 16159 38793 16188
rect 39060 21068 39080 21132
rect 39144 21068 39164 21132
rect 39060 21052 39164 21068
rect 39060 20988 39080 21052
rect 39144 20988 39164 21052
rect 39060 20972 39164 20988
rect 39060 20908 39080 20972
rect 39144 20908 39164 20972
rect 39060 20892 39164 20908
rect 39060 20828 39080 20892
rect 39144 20828 39164 20892
rect 39060 20812 39164 20828
rect 39060 20748 39080 20812
rect 39144 20748 39164 20812
rect 39060 20732 39164 20748
rect 39060 20668 39080 20732
rect 39144 20668 39164 20732
rect 39060 20652 39164 20668
rect 39060 20588 39080 20652
rect 39144 20588 39164 20652
rect 39060 20572 39164 20588
rect 39060 20508 39080 20572
rect 39144 20508 39164 20572
rect 39060 20492 39164 20508
rect 39060 20428 39080 20492
rect 39144 20428 39164 20492
rect 39060 20412 39164 20428
rect 39060 20348 39080 20412
rect 39144 20348 39164 20412
rect 39060 20332 39164 20348
rect 39060 20268 39080 20332
rect 39144 20268 39164 20332
rect 39060 20252 39164 20268
rect 39060 20188 39080 20252
rect 39144 20188 39164 20252
rect 39060 20172 39164 20188
rect 39060 20108 39080 20172
rect 39144 20108 39164 20172
rect 39060 20092 39164 20108
rect 39060 20028 39080 20092
rect 39144 20028 39164 20092
rect 39060 20012 39164 20028
rect 39060 19948 39080 20012
rect 39144 19948 39164 20012
rect 39060 19932 39164 19948
rect 39060 19868 39080 19932
rect 39144 19868 39164 19932
rect 39060 19852 39164 19868
rect 39060 19788 39080 19852
rect 39144 19788 39164 19852
rect 39060 19772 39164 19788
rect 39060 19708 39080 19772
rect 39144 19708 39164 19772
rect 39060 19692 39164 19708
rect 39060 19628 39080 19692
rect 39144 19628 39164 19692
rect 39060 19612 39164 19628
rect 39060 19548 39080 19612
rect 39144 19548 39164 19612
rect 39060 19532 39164 19548
rect 39060 19468 39080 19532
rect 39144 19468 39164 19532
rect 39060 19452 39164 19468
rect 39060 19388 39080 19452
rect 39144 19388 39164 19452
rect 39060 19372 39164 19388
rect 39060 19308 39080 19372
rect 39144 19308 39164 19372
rect 39060 19292 39164 19308
rect 39060 19228 39080 19292
rect 39144 19228 39164 19292
rect 39060 19212 39164 19228
rect 39060 19148 39080 19212
rect 39144 19148 39164 19212
rect 39060 19132 39164 19148
rect 39060 19068 39080 19132
rect 39144 19068 39164 19132
rect 39060 19052 39164 19068
rect 39060 18988 39080 19052
rect 39144 18988 39164 19052
rect 39060 18972 39164 18988
rect 39060 18908 39080 18972
rect 39144 18908 39164 18972
rect 39060 18892 39164 18908
rect 39060 18828 39080 18892
rect 39144 18828 39164 18892
rect 39060 18812 39164 18828
rect 39060 18748 39080 18812
rect 39144 18748 39164 18812
rect 39060 18732 39164 18748
rect 39060 18668 39080 18732
rect 39144 18668 39164 18732
rect 39060 18652 39164 18668
rect 39060 18588 39080 18652
rect 39144 18588 39164 18652
rect 39060 18572 39164 18588
rect 39060 18508 39080 18572
rect 39144 18508 39164 18572
rect 39060 18492 39164 18508
rect 39060 18428 39080 18492
rect 39144 18428 39164 18492
rect 39060 18412 39164 18428
rect 39060 18348 39080 18412
rect 39144 18348 39164 18412
rect 39060 18332 39164 18348
rect 39060 18268 39080 18332
rect 39144 18268 39164 18332
rect 39060 18252 39164 18268
rect 39060 18188 39080 18252
rect 39144 18188 39164 18252
rect 39060 18172 39164 18188
rect 39060 18108 39080 18172
rect 39144 18108 39164 18172
rect 39060 18092 39164 18108
rect 39060 18028 39080 18092
rect 39144 18028 39164 18092
rect 39060 18012 39164 18028
rect 39060 17948 39080 18012
rect 39144 17948 39164 18012
rect 39060 17932 39164 17948
rect 39060 17868 39080 17932
rect 39144 17868 39164 17932
rect 39060 17852 39164 17868
rect 39060 17788 39080 17852
rect 39144 17788 39164 17852
rect 39060 17772 39164 17788
rect 39060 17708 39080 17772
rect 39144 17708 39164 17772
rect 39060 17692 39164 17708
rect 39060 17628 39080 17692
rect 39144 17628 39164 17692
rect 39060 17612 39164 17628
rect 39060 17548 39080 17612
rect 39144 17548 39164 17612
rect 39060 17532 39164 17548
rect 39060 17468 39080 17532
rect 39144 17468 39164 17532
rect 39060 17452 39164 17468
rect 39060 17388 39080 17452
rect 39144 17388 39164 17452
rect 39060 17372 39164 17388
rect 39060 17308 39080 17372
rect 39144 17308 39164 17372
rect 39060 17292 39164 17308
rect 39060 17228 39080 17292
rect 39144 17228 39164 17292
rect 39060 17212 39164 17228
rect 39060 17148 39080 17212
rect 39144 17148 39164 17212
rect 39060 17132 39164 17148
rect 39060 17068 39080 17132
rect 39144 17068 39164 17132
rect 39060 17052 39164 17068
rect 39060 16988 39080 17052
rect 39144 16988 39164 17052
rect 39060 16972 39164 16988
rect 39060 16908 39080 16972
rect 39144 16908 39164 16972
rect 39060 16892 39164 16908
rect 39060 16828 39080 16892
rect 39144 16828 39164 16892
rect 39060 16812 39164 16828
rect 39060 16748 39080 16812
rect 39144 16748 39164 16812
rect 39060 16732 39164 16748
rect 39060 16668 39080 16732
rect 39144 16668 39164 16732
rect 39060 16652 39164 16668
rect 39060 16588 39080 16652
rect 39144 16588 39164 16652
rect 39060 16572 39164 16588
rect 39060 16508 39080 16572
rect 39144 16508 39164 16572
rect 39060 16492 39164 16508
rect 39060 16428 39080 16492
rect 39144 16428 39164 16492
rect 39060 16412 39164 16428
rect 39060 16348 39080 16412
rect 39144 16348 39164 16412
rect 39060 16332 39164 16348
rect 39060 16268 39080 16332
rect 39144 16268 39164 16332
rect 39060 16252 39164 16268
rect 39060 16188 39080 16252
rect 39144 16188 39164 16252
rect 39060 16172 39164 16188
rect 33448 15812 33552 16108
rect 27836 15732 27940 15748
rect 27836 15668 27856 15732
rect 27920 15668 27940 15732
rect 27836 15652 27940 15668
rect 27836 15588 27856 15652
rect 27920 15588 27940 15652
rect 27836 15572 27940 15588
rect 27836 15508 27856 15572
rect 27920 15508 27940 15572
rect 27836 15492 27940 15508
rect 27836 15428 27856 15492
rect 27920 15428 27940 15492
rect 27836 15412 27940 15428
rect 27836 15348 27856 15412
rect 27920 15348 27940 15412
rect 27836 15332 27940 15348
rect 27836 15268 27856 15332
rect 27920 15268 27940 15332
rect 27836 15252 27940 15268
rect 27836 15188 27856 15252
rect 27920 15188 27940 15252
rect 27836 15172 27940 15188
rect 27836 15108 27856 15172
rect 27920 15108 27940 15172
rect 27836 15092 27940 15108
rect 27836 15028 27856 15092
rect 27920 15028 27940 15092
rect 27836 15012 27940 15028
rect 27836 14948 27856 15012
rect 27920 14948 27940 15012
rect 27836 14932 27940 14948
rect 27836 14868 27856 14932
rect 27920 14868 27940 14932
rect 27836 14852 27940 14868
rect 27836 14788 27856 14852
rect 27920 14788 27940 14852
rect 27836 14772 27940 14788
rect 27836 14708 27856 14772
rect 27920 14708 27940 14772
rect 27836 14692 27940 14708
rect 27836 14628 27856 14692
rect 27920 14628 27940 14692
rect 27836 14612 27940 14628
rect 27836 14548 27856 14612
rect 27920 14548 27940 14612
rect 27836 14532 27940 14548
rect 27836 14468 27856 14532
rect 27920 14468 27940 14532
rect 27836 14452 27940 14468
rect 27836 14388 27856 14452
rect 27920 14388 27940 14452
rect 27836 14372 27940 14388
rect 27836 14308 27856 14372
rect 27920 14308 27940 14372
rect 27836 14292 27940 14308
rect 27836 14228 27856 14292
rect 27920 14228 27940 14292
rect 27836 14212 27940 14228
rect 27836 14148 27856 14212
rect 27920 14148 27940 14212
rect 27836 14132 27940 14148
rect 27836 14068 27856 14132
rect 27920 14068 27940 14132
rect 27836 14052 27940 14068
rect 27836 13988 27856 14052
rect 27920 13988 27940 14052
rect 27836 13972 27940 13988
rect 27836 13908 27856 13972
rect 27920 13908 27940 13972
rect 27836 13892 27940 13908
rect 27836 13828 27856 13892
rect 27920 13828 27940 13892
rect 27836 13812 27940 13828
rect 27836 13748 27856 13812
rect 27920 13748 27940 13812
rect 27836 13732 27940 13748
rect 27836 13668 27856 13732
rect 27920 13668 27940 13732
rect 27836 13652 27940 13668
rect 27836 13588 27856 13652
rect 27920 13588 27940 13652
rect 27836 13572 27940 13588
rect 27836 13508 27856 13572
rect 27920 13508 27940 13572
rect 27836 13492 27940 13508
rect 27836 13428 27856 13492
rect 27920 13428 27940 13492
rect 27836 13412 27940 13428
rect 27836 13348 27856 13412
rect 27920 13348 27940 13412
rect 27836 13332 27940 13348
rect 27836 13268 27856 13332
rect 27920 13268 27940 13332
rect 27836 13252 27940 13268
rect 27836 13188 27856 13252
rect 27920 13188 27940 13252
rect 27836 13172 27940 13188
rect 27836 13108 27856 13172
rect 27920 13108 27940 13172
rect 27836 13092 27940 13108
rect 27836 13028 27856 13092
rect 27920 13028 27940 13092
rect 27836 13012 27940 13028
rect 27836 12948 27856 13012
rect 27920 12948 27940 13012
rect 27836 12932 27940 12948
rect 27836 12868 27856 12932
rect 27920 12868 27940 12932
rect 27836 12852 27940 12868
rect 27836 12788 27856 12852
rect 27920 12788 27940 12852
rect 27836 12772 27940 12788
rect 27836 12708 27856 12772
rect 27920 12708 27940 12772
rect 27836 12692 27940 12708
rect 27836 12628 27856 12692
rect 27920 12628 27940 12692
rect 27836 12612 27940 12628
rect 27836 12548 27856 12612
rect 27920 12548 27940 12612
rect 27836 12532 27940 12548
rect 27836 12468 27856 12532
rect 27920 12468 27940 12532
rect 27836 12452 27940 12468
rect 27836 12388 27856 12452
rect 27920 12388 27940 12452
rect 27836 12372 27940 12388
rect 27836 12308 27856 12372
rect 27920 12308 27940 12372
rect 27836 12292 27940 12308
rect 27836 12228 27856 12292
rect 27920 12228 27940 12292
rect 27836 12212 27940 12228
rect 27836 12148 27856 12212
rect 27920 12148 27940 12212
rect 27836 12132 27940 12148
rect 27836 12068 27856 12132
rect 27920 12068 27940 12132
rect 27836 12052 27940 12068
rect 27836 11988 27856 12052
rect 27920 11988 27940 12052
rect 27836 11972 27940 11988
rect 27836 11908 27856 11972
rect 27920 11908 27940 11972
rect 27836 11892 27940 11908
rect 27836 11828 27856 11892
rect 27920 11828 27940 11892
rect 27836 11812 27940 11828
rect 27836 11748 27856 11812
rect 27920 11748 27940 11812
rect 27836 11732 27940 11748
rect 27836 11668 27856 11732
rect 27920 11668 27940 11732
rect 27836 11652 27940 11668
rect 27836 11588 27856 11652
rect 27920 11588 27940 11652
rect 27836 11572 27940 11588
rect 27836 11508 27856 11572
rect 27920 11508 27940 11572
rect 27836 11492 27940 11508
rect 27836 11428 27856 11492
rect 27920 11428 27940 11492
rect 27836 11412 27940 11428
rect 27836 11348 27856 11412
rect 27920 11348 27940 11412
rect 27836 11332 27940 11348
rect 27836 11268 27856 11332
rect 27920 11268 27940 11332
rect 27836 11252 27940 11268
rect 27836 11188 27856 11252
rect 27920 11188 27940 11252
rect 27836 11172 27940 11188
rect 27836 11108 27856 11172
rect 27920 11108 27940 11172
rect 27836 11092 27940 11108
rect 27836 11028 27856 11092
rect 27920 11028 27940 11092
rect 27836 11012 27940 11028
rect 27836 10948 27856 11012
rect 27920 10948 27940 11012
rect 27836 10932 27940 10948
rect 27836 10868 27856 10932
rect 27920 10868 27940 10932
rect 27836 10852 27940 10868
rect 22224 10492 22328 10788
rect 16612 10412 16716 10428
rect 16612 10348 16632 10412
rect 16696 10348 16716 10412
rect 16612 10332 16716 10348
rect 16612 10268 16632 10332
rect 16696 10268 16716 10332
rect 16612 10252 16716 10268
rect 16612 10188 16632 10252
rect 16696 10188 16716 10252
rect 16612 10172 16716 10188
rect 16612 10108 16632 10172
rect 16696 10108 16716 10172
rect 16612 10092 16716 10108
rect 16612 10028 16632 10092
rect 16696 10028 16716 10092
rect 16612 10012 16716 10028
rect 16612 9948 16632 10012
rect 16696 9948 16716 10012
rect 16612 9932 16716 9948
rect 16612 9868 16632 9932
rect 16696 9868 16716 9932
rect 16612 9852 16716 9868
rect 16612 9788 16632 9852
rect 16696 9788 16716 9852
rect 16612 9772 16716 9788
rect 16612 9708 16632 9772
rect 16696 9708 16716 9772
rect 16612 9692 16716 9708
rect 16612 9628 16632 9692
rect 16696 9628 16716 9692
rect 16612 9612 16716 9628
rect 16612 9548 16632 9612
rect 16696 9548 16716 9612
rect 16612 9532 16716 9548
rect 16612 9468 16632 9532
rect 16696 9468 16716 9532
rect 16612 9452 16716 9468
rect 16612 9388 16632 9452
rect 16696 9388 16716 9452
rect 16612 9372 16716 9388
rect 16612 9308 16632 9372
rect 16696 9308 16716 9372
rect 16612 9292 16716 9308
rect 16612 9228 16632 9292
rect 16696 9228 16716 9292
rect 16612 9212 16716 9228
rect 16612 9148 16632 9212
rect 16696 9148 16716 9212
rect 16612 9132 16716 9148
rect 16612 9068 16632 9132
rect 16696 9068 16716 9132
rect 16612 9052 16716 9068
rect 16612 8988 16632 9052
rect 16696 8988 16716 9052
rect 16612 8972 16716 8988
rect 16612 8908 16632 8972
rect 16696 8908 16716 8972
rect 16612 8892 16716 8908
rect 16612 8828 16632 8892
rect 16696 8828 16716 8892
rect 16612 8812 16716 8828
rect 16612 8748 16632 8812
rect 16696 8748 16716 8812
rect 16612 8732 16716 8748
rect 16612 8668 16632 8732
rect 16696 8668 16716 8732
rect 16612 8652 16716 8668
rect 16612 8588 16632 8652
rect 16696 8588 16716 8652
rect 16612 8572 16716 8588
rect 16612 8508 16632 8572
rect 16696 8508 16716 8572
rect 16612 8492 16716 8508
rect 16612 8428 16632 8492
rect 16696 8428 16716 8492
rect 16612 8412 16716 8428
rect 16612 8348 16632 8412
rect 16696 8348 16716 8412
rect 16612 8332 16716 8348
rect 16612 8268 16632 8332
rect 16696 8268 16716 8332
rect 16612 8252 16716 8268
rect 16612 8188 16632 8252
rect 16696 8188 16716 8252
rect 16612 8172 16716 8188
rect 16612 8108 16632 8172
rect 16696 8108 16716 8172
rect 16612 8092 16716 8108
rect 16612 8028 16632 8092
rect 16696 8028 16716 8092
rect 16612 8012 16716 8028
rect 16612 7948 16632 8012
rect 16696 7948 16716 8012
rect 16612 7932 16716 7948
rect 16612 7868 16632 7932
rect 16696 7868 16716 7932
rect 16612 7852 16716 7868
rect 16612 7788 16632 7852
rect 16696 7788 16716 7852
rect 16612 7772 16716 7788
rect 16612 7708 16632 7772
rect 16696 7708 16716 7772
rect 16612 7692 16716 7708
rect 16612 7628 16632 7692
rect 16696 7628 16716 7692
rect 16612 7612 16716 7628
rect 16612 7548 16632 7612
rect 16696 7548 16716 7612
rect 16612 7532 16716 7548
rect 16612 7468 16632 7532
rect 16696 7468 16716 7532
rect 16612 7452 16716 7468
rect 16612 7388 16632 7452
rect 16696 7388 16716 7452
rect 16612 7372 16716 7388
rect 16612 7308 16632 7372
rect 16696 7308 16716 7372
rect 16612 7292 16716 7308
rect 16612 7228 16632 7292
rect 16696 7228 16716 7292
rect 16612 7212 16716 7228
rect 16612 7148 16632 7212
rect 16696 7148 16716 7212
rect 16612 7132 16716 7148
rect 16612 7068 16632 7132
rect 16696 7068 16716 7132
rect 16612 7052 16716 7068
rect 16612 6988 16632 7052
rect 16696 6988 16716 7052
rect 16612 6972 16716 6988
rect 16612 6908 16632 6972
rect 16696 6908 16716 6972
rect 16612 6892 16716 6908
rect 16612 6828 16632 6892
rect 16696 6828 16716 6892
rect 16612 6812 16716 6828
rect 16612 6748 16632 6812
rect 16696 6748 16716 6812
rect 16612 6732 16716 6748
rect 16612 6668 16632 6732
rect 16696 6668 16716 6732
rect 16612 6652 16716 6668
rect 16612 6588 16632 6652
rect 16696 6588 16716 6652
rect 16612 6572 16716 6588
rect 16612 6508 16632 6572
rect 16696 6508 16716 6572
rect 16612 6492 16716 6508
rect 16612 6428 16632 6492
rect 16696 6428 16716 6492
rect 16612 6412 16716 6428
rect 16612 6348 16632 6412
rect 16696 6348 16716 6412
rect 16612 6332 16716 6348
rect 16612 6268 16632 6332
rect 16696 6268 16716 6332
rect 16612 6252 16716 6268
rect 16612 6188 16632 6252
rect 16696 6188 16716 6252
rect 16612 6172 16716 6188
rect 16612 6108 16632 6172
rect 16696 6108 16716 6172
rect 16612 6092 16716 6108
rect 16612 6028 16632 6092
rect 16696 6028 16716 6092
rect 16612 6012 16716 6028
rect 16612 5948 16632 6012
rect 16696 5948 16716 6012
rect 16612 5932 16716 5948
rect 16612 5868 16632 5932
rect 16696 5868 16716 5932
rect 16612 5852 16716 5868
rect 16612 5788 16632 5852
rect 16696 5788 16716 5852
rect 16612 5772 16716 5788
rect 16612 5708 16632 5772
rect 16696 5708 16716 5772
rect 16612 5692 16716 5708
rect 16612 5628 16632 5692
rect 16696 5628 16716 5692
rect 16612 5612 16716 5628
rect 16612 5548 16632 5612
rect 16696 5548 16716 5612
rect 16612 5532 16716 5548
rect 11000 5172 11104 5468
rect 5388 5092 5492 5108
rect 5388 5028 5408 5092
rect 5472 5028 5492 5092
rect 5388 5012 5492 5028
rect 5388 4948 5408 5012
rect 5472 4948 5492 5012
rect 5388 4932 5492 4948
rect 5388 4868 5408 4932
rect 5472 4868 5492 4932
rect 5388 4852 5492 4868
rect 5388 4788 5408 4852
rect 5472 4788 5492 4852
rect 5388 4772 5492 4788
rect 5388 4708 5408 4772
rect 5472 4708 5492 4772
rect 5388 4692 5492 4708
rect 5388 4628 5408 4692
rect 5472 4628 5492 4692
rect 5388 4612 5492 4628
rect 5388 4548 5408 4612
rect 5472 4548 5492 4612
rect 5388 4532 5492 4548
rect 5388 4468 5408 4532
rect 5472 4468 5492 4532
rect 5388 4452 5492 4468
rect 5388 4388 5408 4452
rect 5472 4388 5492 4452
rect 5388 4372 5492 4388
rect 5388 4308 5408 4372
rect 5472 4308 5492 4372
rect 5388 4292 5492 4308
rect 5388 4228 5408 4292
rect 5472 4228 5492 4292
rect 5388 4212 5492 4228
rect 5388 4148 5408 4212
rect 5472 4148 5492 4212
rect 5388 4132 5492 4148
rect 5388 4068 5408 4132
rect 5472 4068 5492 4132
rect 5388 4052 5492 4068
rect 5388 3988 5408 4052
rect 5472 3988 5492 4052
rect 5388 3972 5492 3988
rect 5388 3908 5408 3972
rect 5472 3908 5492 3972
rect 5388 3892 5492 3908
rect 5388 3828 5408 3892
rect 5472 3828 5492 3892
rect 5388 3812 5492 3828
rect 5388 3748 5408 3812
rect 5472 3748 5492 3812
rect 5388 3732 5492 3748
rect 5388 3668 5408 3732
rect 5472 3668 5492 3732
rect 5388 3652 5492 3668
rect 5388 3588 5408 3652
rect 5472 3588 5492 3652
rect 5388 3572 5492 3588
rect 5388 3508 5408 3572
rect 5472 3508 5492 3572
rect 5388 3492 5492 3508
rect 5388 3428 5408 3492
rect 5472 3428 5492 3492
rect 5388 3412 5492 3428
rect 5388 3348 5408 3412
rect 5472 3348 5492 3412
rect 5388 3332 5492 3348
rect 5388 3268 5408 3332
rect 5472 3268 5492 3332
rect 5388 3252 5492 3268
rect 5388 3188 5408 3252
rect 5472 3188 5492 3252
rect 5388 3172 5492 3188
rect 5388 3108 5408 3172
rect 5472 3108 5492 3172
rect 5388 3092 5492 3108
rect 5388 3028 5408 3092
rect 5472 3028 5492 3092
rect 5388 3012 5492 3028
rect 5388 2948 5408 3012
rect 5472 2948 5492 3012
rect 5388 2932 5492 2948
rect 5388 2868 5408 2932
rect 5472 2868 5492 2932
rect 5388 2852 5492 2868
rect 5388 2788 5408 2852
rect 5472 2788 5492 2852
rect 5388 2772 5492 2788
rect 5388 2708 5408 2772
rect 5472 2708 5492 2772
rect 5388 2692 5492 2708
rect 5388 2628 5408 2692
rect 5472 2628 5492 2692
rect 5388 2612 5492 2628
rect 5388 2548 5408 2612
rect 5472 2548 5492 2612
rect 5388 2532 5492 2548
rect 5388 2468 5408 2532
rect 5472 2468 5492 2532
rect 5388 2452 5492 2468
rect 5388 2388 5408 2452
rect 5472 2388 5492 2452
rect 5388 2372 5492 2388
rect 5388 2308 5408 2372
rect 5472 2308 5492 2372
rect 5388 2292 5492 2308
rect 5388 2228 5408 2292
rect 5472 2228 5492 2292
rect 5388 2212 5492 2228
rect 5388 2148 5408 2212
rect 5472 2148 5492 2212
rect 5388 2132 5492 2148
rect 5388 2068 5408 2132
rect 5472 2068 5492 2132
rect 5388 2052 5492 2068
rect 5388 1988 5408 2052
rect 5472 1988 5492 2052
rect 5388 1972 5492 1988
rect 5388 1908 5408 1972
rect 5472 1908 5492 1972
rect 5388 1892 5492 1908
rect 5388 1828 5408 1892
rect 5472 1828 5492 1892
rect 5388 1812 5492 1828
rect 5388 1748 5408 1812
rect 5472 1748 5492 1812
rect 5388 1732 5492 1748
rect 5388 1668 5408 1732
rect 5472 1668 5492 1732
rect 5388 1652 5492 1668
rect 5388 1588 5408 1652
rect 5472 1588 5492 1652
rect 5388 1572 5492 1588
rect 5388 1508 5408 1572
rect 5472 1508 5492 1572
rect 5388 1492 5492 1508
rect 5388 1428 5408 1492
rect 5472 1428 5492 1492
rect 5388 1412 5492 1428
rect 5388 1348 5408 1412
rect 5472 1348 5492 1412
rect 5388 1332 5492 1348
rect 5388 1268 5408 1332
rect 5472 1268 5492 1332
rect 5388 1252 5492 1268
rect 5388 1188 5408 1252
rect 5472 1188 5492 1252
rect 5388 1172 5492 1188
rect 5388 1108 5408 1172
rect 5472 1108 5492 1172
rect 5388 1092 5492 1108
rect 5388 1028 5408 1092
rect 5472 1028 5492 1092
rect 5388 1012 5492 1028
rect 5388 948 5408 1012
rect 5472 948 5492 1012
rect 5388 932 5492 948
rect 5388 868 5408 932
rect 5472 868 5492 932
rect 5388 852 5492 868
rect 5388 788 5408 852
rect 5472 788 5492 852
rect 5388 772 5492 788
rect 5388 708 5408 772
rect 5472 708 5492 772
rect 5388 692 5492 708
rect 5388 628 5408 692
rect 5472 628 5492 692
rect 5388 612 5492 628
rect 5388 548 5408 612
rect 5472 548 5492 612
rect 5388 532 5492 548
rect 5388 468 5408 532
rect 5472 468 5492 532
rect 5388 452 5492 468
rect 5388 388 5408 452
rect 5472 388 5492 452
rect 5388 372 5492 388
rect 5388 308 5408 372
rect 5472 308 5492 372
rect 5388 292 5492 308
rect 5388 228 5408 292
rect 5472 228 5492 292
rect 5388 212 5492 228
rect -224 -148 -120 148
rect -5836 -228 -5732 -212
rect -5836 -292 -5816 -228
rect -5752 -292 -5732 -228
rect -5836 -308 -5732 -292
rect -5836 -372 -5816 -308
rect -5752 -372 -5732 -308
rect -5836 -388 -5732 -372
rect -5836 -452 -5816 -388
rect -5752 -452 -5732 -388
rect -5836 -468 -5732 -452
rect -5836 -532 -5816 -468
rect -5752 -532 -5732 -468
rect -5836 -548 -5732 -532
rect -5836 -612 -5816 -548
rect -5752 -612 -5732 -548
rect -5836 -628 -5732 -612
rect -5836 -692 -5816 -628
rect -5752 -692 -5732 -628
rect -5836 -708 -5732 -692
rect -5836 -772 -5816 -708
rect -5752 -772 -5732 -708
rect -5836 -788 -5732 -772
rect -5836 -852 -5816 -788
rect -5752 -852 -5732 -788
rect -5836 -868 -5732 -852
rect -5836 -932 -5816 -868
rect -5752 -932 -5732 -868
rect -5836 -948 -5732 -932
rect -5836 -1012 -5816 -948
rect -5752 -1012 -5732 -948
rect -5836 -1028 -5732 -1012
rect -5836 -1092 -5816 -1028
rect -5752 -1092 -5732 -1028
rect -5836 -1108 -5732 -1092
rect -5836 -1172 -5816 -1108
rect -5752 -1172 -5732 -1108
rect -5836 -1188 -5732 -1172
rect -5836 -1252 -5816 -1188
rect -5752 -1252 -5732 -1188
rect -5836 -1268 -5732 -1252
rect -5836 -1332 -5816 -1268
rect -5752 -1332 -5732 -1268
rect -5836 -1348 -5732 -1332
rect -5836 -1412 -5816 -1348
rect -5752 -1412 -5732 -1348
rect -5836 -1428 -5732 -1412
rect -5836 -1492 -5816 -1428
rect -5752 -1492 -5732 -1428
rect -5836 -1508 -5732 -1492
rect -5836 -1572 -5816 -1508
rect -5752 -1572 -5732 -1508
rect -5836 -1588 -5732 -1572
rect -5836 -1652 -5816 -1588
rect -5752 -1652 -5732 -1588
rect -5836 -1668 -5732 -1652
rect -5836 -1732 -5816 -1668
rect -5752 -1732 -5732 -1668
rect -5836 -1748 -5732 -1732
rect -5836 -1812 -5816 -1748
rect -5752 -1812 -5732 -1748
rect -5836 -1828 -5732 -1812
rect -5836 -1892 -5816 -1828
rect -5752 -1892 -5732 -1828
rect -5836 -1908 -5732 -1892
rect -5836 -1972 -5816 -1908
rect -5752 -1972 -5732 -1908
rect -5836 -1988 -5732 -1972
rect -5836 -2052 -5816 -1988
rect -5752 -2052 -5732 -1988
rect -5836 -2068 -5732 -2052
rect -5836 -2132 -5816 -2068
rect -5752 -2132 -5732 -2068
rect -5836 -2148 -5732 -2132
rect -5836 -2212 -5816 -2148
rect -5752 -2212 -5732 -2148
rect -5836 -2228 -5732 -2212
rect -5836 -2292 -5816 -2228
rect -5752 -2292 -5732 -2228
rect -5836 -2308 -5732 -2292
rect -5836 -2372 -5816 -2308
rect -5752 -2372 -5732 -2308
rect -5836 -2388 -5732 -2372
rect -5836 -2452 -5816 -2388
rect -5752 -2452 -5732 -2388
rect -5836 -2468 -5732 -2452
rect -5836 -2532 -5816 -2468
rect -5752 -2532 -5732 -2468
rect -5836 -2548 -5732 -2532
rect -5836 -2612 -5816 -2548
rect -5752 -2612 -5732 -2548
rect -5836 -2628 -5732 -2612
rect -5836 -2692 -5816 -2628
rect -5752 -2692 -5732 -2628
rect -5836 -2708 -5732 -2692
rect -5836 -2772 -5816 -2708
rect -5752 -2772 -5732 -2708
rect -5836 -2788 -5732 -2772
rect -5836 -2852 -5816 -2788
rect -5752 -2852 -5732 -2788
rect -5836 -2868 -5732 -2852
rect -5836 -2932 -5816 -2868
rect -5752 -2932 -5732 -2868
rect -5836 -2948 -5732 -2932
rect -5836 -3012 -5816 -2948
rect -5752 -3012 -5732 -2948
rect -5836 -3028 -5732 -3012
rect -5836 -3092 -5816 -3028
rect -5752 -3092 -5732 -3028
rect -5836 -3108 -5732 -3092
rect -5836 -3172 -5816 -3108
rect -5752 -3172 -5732 -3108
rect -5836 -3188 -5732 -3172
rect -5836 -3252 -5816 -3188
rect -5752 -3252 -5732 -3188
rect -5836 -3268 -5732 -3252
rect -5836 -3332 -5816 -3268
rect -5752 -3332 -5732 -3268
rect -5836 -3348 -5732 -3332
rect -5836 -3412 -5816 -3348
rect -5752 -3412 -5732 -3348
rect -5836 -3428 -5732 -3412
rect -5836 -3492 -5816 -3428
rect -5752 -3492 -5732 -3428
rect -5836 -3508 -5732 -3492
rect -5836 -3572 -5816 -3508
rect -5752 -3572 -5732 -3508
rect -5836 -3588 -5732 -3572
rect -5836 -3652 -5816 -3588
rect -5752 -3652 -5732 -3588
rect -5836 -3668 -5732 -3652
rect -5836 -3732 -5816 -3668
rect -5752 -3732 -5732 -3668
rect -5836 -3748 -5732 -3732
rect -5836 -3812 -5816 -3748
rect -5752 -3812 -5732 -3748
rect -5836 -3828 -5732 -3812
rect -5836 -3892 -5816 -3828
rect -5752 -3892 -5732 -3828
rect -5836 -3908 -5732 -3892
rect -5836 -3972 -5816 -3908
rect -5752 -3972 -5732 -3908
rect -5836 -3988 -5732 -3972
rect -5836 -4052 -5816 -3988
rect -5752 -4052 -5732 -3988
rect -5836 -4068 -5732 -4052
rect -5836 -4132 -5816 -4068
rect -5752 -4132 -5732 -4068
rect -5836 -4148 -5732 -4132
rect -5836 -4212 -5816 -4148
rect -5752 -4212 -5732 -4148
rect -5836 -4228 -5732 -4212
rect -5836 -4292 -5816 -4228
rect -5752 -4292 -5732 -4228
rect -5836 -4308 -5732 -4292
rect -5836 -4372 -5816 -4308
rect -5752 -4372 -5732 -4308
rect -5836 -4388 -5732 -4372
rect -5836 -4452 -5816 -4388
rect -5752 -4452 -5732 -4388
rect -5836 -4468 -5732 -4452
rect -5836 -4532 -5816 -4468
rect -5752 -4532 -5732 -4468
rect -5836 -4548 -5732 -4532
rect -5836 -4612 -5816 -4548
rect -5752 -4612 -5732 -4548
rect -5836 -4628 -5732 -4612
rect -5836 -4692 -5816 -4628
rect -5752 -4692 -5732 -4628
rect -5836 -4708 -5732 -4692
rect -5836 -4772 -5816 -4708
rect -5752 -4772 -5732 -4708
rect -5836 -4788 -5732 -4772
rect -5836 -4852 -5816 -4788
rect -5752 -4852 -5732 -4788
rect -5836 -4868 -5732 -4852
rect -5836 -4932 -5816 -4868
rect -5752 -4932 -5732 -4868
rect -5836 -4948 -5732 -4932
rect -5836 -5012 -5816 -4948
rect -5752 -5012 -5732 -4948
rect -5836 -5028 -5732 -5012
rect -5836 -5092 -5816 -5028
rect -5752 -5092 -5732 -5028
rect -5836 -5108 -5732 -5092
rect -11448 -5468 -11344 -5172
rect -17060 -5548 -16956 -5532
rect -17060 -5612 -17040 -5548
rect -16976 -5612 -16956 -5548
rect -17060 -5628 -16956 -5612
rect -17060 -5692 -17040 -5628
rect -16976 -5692 -16956 -5628
rect -17060 -5708 -16956 -5692
rect -17060 -5772 -17040 -5708
rect -16976 -5772 -16956 -5708
rect -17060 -5788 -16956 -5772
rect -17060 -5852 -17040 -5788
rect -16976 -5852 -16956 -5788
rect -17060 -5868 -16956 -5852
rect -17060 -5932 -17040 -5868
rect -16976 -5932 -16956 -5868
rect -17060 -5948 -16956 -5932
rect -17060 -6012 -17040 -5948
rect -16976 -6012 -16956 -5948
rect -17060 -6028 -16956 -6012
rect -17060 -6092 -17040 -6028
rect -16976 -6092 -16956 -6028
rect -17060 -6108 -16956 -6092
rect -17060 -6172 -17040 -6108
rect -16976 -6172 -16956 -6108
rect -17060 -6188 -16956 -6172
rect -17060 -6252 -17040 -6188
rect -16976 -6252 -16956 -6188
rect -17060 -6268 -16956 -6252
rect -17060 -6332 -17040 -6268
rect -16976 -6332 -16956 -6268
rect -17060 -6348 -16956 -6332
rect -17060 -6412 -17040 -6348
rect -16976 -6412 -16956 -6348
rect -17060 -6428 -16956 -6412
rect -17060 -6492 -17040 -6428
rect -16976 -6492 -16956 -6428
rect -17060 -6508 -16956 -6492
rect -17060 -6572 -17040 -6508
rect -16976 -6572 -16956 -6508
rect -17060 -6588 -16956 -6572
rect -17060 -6652 -17040 -6588
rect -16976 -6652 -16956 -6588
rect -17060 -6668 -16956 -6652
rect -17060 -6732 -17040 -6668
rect -16976 -6732 -16956 -6668
rect -17060 -6748 -16956 -6732
rect -17060 -6812 -17040 -6748
rect -16976 -6812 -16956 -6748
rect -17060 -6828 -16956 -6812
rect -17060 -6892 -17040 -6828
rect -16976 -6892 -16956 -6828
rect -17060 -6908 -16956 -6892
rect -17060 -6972 -17040 -6908
rect -16976 -6972 -16956 -6908
rect -17060 -6988 -16956 -6972
rect -17060 -7052 -17040 -6988
rect -16976 -7052 -16956 -6988
rect -17060 -7068 -16956 -7052
rect -17060 -7132 -17040 -7068
rect -16976 -7132 -16956 -7068
rect -17060 -7148 -16956 -7132
rect -17060 -7212 -17040 -7148
rect -16976 -7212 -16956 -7148
rect -17060 -7228 -16956 -7212
rect -17060 -7292 -17040 -7228
rect -16976 -7292 -16956 -7228
rect -17060 -7308 -16956 -7292
rect -17060 -7372 -17040 -7308
rect -16976 -7372 -16956 -7308
rect -17060 -7388 -16956 -7372
rect -17060 -7452 -17040 -7388
rect -16976 -7452 -16956 -7388
rect -17060 -7468 -16956 -7452
rect -17060 -7532 -17040 -7468
rect -16976 -7532 -16956 -7468
rect -17060 -7548 -16956 -7532
rect -17060 -7612 -17040 -7548
rect -16976 -7612 -16956 -7548
rect -17060 -7628 -16956 -7612
rect -17060 -7692 -17040 -7628
rect -16976 -7692 -16956 -7628
rect -17060 -7708 -16956 -7692
rect -17060 -7772 -17040 -7708
rect -16976 -7772 -16956 -7708
rect -17060 -7788 -16956 -7772
rect -17060 -7852 -17040 -7788
rect -16976 -7852 -16956 -7788
rect -17060 -7868 -16956 -7852
rect -17060 -7932 -17040 -7868
rect -16976 -7932 -16956 -7868
rect -17060 -7948 -16956 -7932
rect -17060 -8012 -17040 -7948
rect -16976 -8012 -16956 -7948
rect -17060 -8028 -16956 -8012
rect -17060 -8092 -17040 -8028
rect -16976 -8092 -16956 -8028
rect -17060 -8108 -16956 -8092
rect -17060 -8172 -17040 -8108
rect -16976 -8172 -16956 -8108
rect -17060 -8188 -16956 -8172
rect -17060 -8252 -17040 -8188
rect -16976 -8252 -16956 -8188
rect -17060 -8268 -16956 -8252
rect -17060 -8332 -17040 -8268
rect -16976 -8332 -16956 -8268
rect -17060 -8348 -16956 -8332
rect -17060 -8412 -17040 -8348
rect -16976 -8412 -16956 -8348
rect -17060 -8428 -16956 -8412
rect -17060 -8492 -17040 -8428
rect -16976 -8492 -16956 -8428
rect -17060 -8508 -16956 -8492
rect -17060 -8572 -17040 -8508
rect -16976 -8572 -16956 -8508
rect -17060 -8588 -16956 -8572
rect -17060 -8652 -17040 -8588
rect -16976 -8652 -16956 -8588
rect -17060 -8668 -16956 -8652
rect -17060 -8732 -17040 -8668
rect -16976 -8732 -16956 -8668
rect -17060 -8748 -16956 -8732
rect -17060 -8812 -17040 -8748
rect -16976 -8812 -16956 -8748
rect -17060 -8828 -16956 -8812
rect -17060 -8892 -17040 -8828
rect -16976 -8892 -16956 -8828
rect -17060 -8908 -16956 -8892
rect -17060 -8972 -17040 -8908
rect -16976 -8972 -16956 -8908
rect -17060 -8988 -16956 -8972
rect -17060 -9052 -17040 -8988
rect -16976 -9052 -16956 -8988
rect -17060 -9068 -16956 -9052
rect -17060 -9132 -17040 -9068
rect -16976 -9132 -16956 -9068
rect -17060 -9148 -16956 -9132
rect -17060 -9212 -17040 -9148
rect -16976 -9212 -16956 -9148
rect -17060 -9228 -16956 -9212
rect -17060 -9292 -17040 -9228
rect -16976 -9292 -16956 -9228
rect -17060 -9308 -16956 -9292
rect -17060 -9372 -17040 -9308
rect -16976 -9372 -16956 -9308
rect -17060 -9388 -16956 -9372
rect -17060 -9452 -17040 -9388
rect -16976 -9452 -16956 -9388
rect -17060 -9468 -16956 -9452
rect -17060 -9532 -17040 -9468
rect -16976 -9532 -16956 -9468
rect -17060 -9548 -16956 -9532
rect -17060 -9612 -17040 -9548
rect -16976 -9612 -16956 -9548
rect -17060 -9628 -16956 -9612
rect -17060 -9692 -17040 -9628
rect -16976 -9692 -16956 -9628
rect -17060 -9708 -16956 -9692
rect -17060 -9772 -17040 -9708
rect -16976 -9772 -16956 -9708
rect -17060 -9788 -16956 -9772
rect -17060 -9852 -17040 -9788
rect -16976 -9852 -16956 -9788
rect -17060 -9868 -16956 -9852
rect -17060 -9932 -17040 -9868
rect -16976 -9932 -16956 -9868
rect -17060 -9948 -16956 -9932
rect -17060 -10012 -17040 -9948
rect -16976 -10012 -16956 -9948
rect -17060 -10028 -16956 -10012
rect -17060 -10092 -17040 -10028
rect -16976 -10092 -16956 -10028
rect -17060 -10108 -16956 -10092
rect -17060 -10172 -17040 -10108
rect -16976 -10172 -16956 -10108
rect -17060 -10188 -16956 -10172
rect -17060 -10252 -17040 -10188
rect -16976 -10252 -16956 -10188
rect -17060 -10268 -16956 -10252
rect -17060 -10332 -17040 -10268
rect -16976 -10332 -16956 -10268
rect -17060 -10348 -16956 -10332
rect -17060 -10412 -17040 -10348
rect -16976 -10412 -16956 -10348
rect -17060 -10428 -16956 -10412
rect -22672 -10788 -22568 -10492
rect -28284 -10868 -28180 -10852
rect -28284 -10932 -28264 -10868
rect -28200 -10932 -28180 -10868
rect -28284 -10948 -28180 -10932
rect -28284 -11012 -28264 -10948
rect -28200 -11012 -28180 -10948
rect -28284 -11028 -28180 -11012
rect -28284 -11092 -28264 -11028
rect -28200 -11092 -28180 -11028
rect -28284 -11108 -28180 -11092
rect -28284 -11172 -28264 -11108
rect -28200 -11172 -28180 -11108
rect -28284 -11188 -28180 -11172
rect -28284 -11252 -28264 -11188
rect -28200 -11252 -28180 -11188
rect -28284 -11268 -28180 -11252
rect -28284 -11332 -28264 -11268
rect -28200 -11332 -28180 -11268
rect -28284 -11348 -28180 -11332
rect -28284 -11412 -28264 -11348
rect -28200 -11412 -28180 -11348
rect -28284 -11428 -28180 -11412
rect -28284 -11492 -28264 -11428
rect -28200 -11492 -28180 -11428
rect -28284 -11508 -28180 -11492
rect -28284 -11572 -28264 -11508
rect -28200 -11572 -28180 -11508
rect -28284 -11588 -28180 -11572
rect -28284 -11652 -28264 -11588
rect -28200 -11652 -28180 -11588
rect -28284 -11668 -28180 -11652
rect -28284 -11732 -28264 -11668
rect -28200 -11732 -28180 -11668
rect -28284 -11748 -28180 -11732
rect -28284 -11812 -28264 -11748
rect -28200 -11812 -28180 -11748
rect -28284 -11828 -28180 -11812
rect -28284 -11892 -28264 -11828
rect -28200 -11892 -28180 -11828
rect -28284 -11908 -28180 -11892
rect -28284 -11972 -28264 -11908
rect -28200 -11972 -28180 -11908
rect -28284 -11988 -28180 -11972
rect -28284 -12052 -28264 -11988
rect -28200 -12052 -28180 -11988
rect -28284 -12068 -28180 -12052
rect -28284 -12132 -28264 -12068
rect -28200 -12132 -28180 -12068
rect -28284 -12148 -28180 -12132
rect -28284 -12212 -28264 -12148
rect -28200 -12212 -28180 -12148
rect -28284 -12228 -28180 -12212
rect -28284 -12292 -28264 -12228
rect -28200 -12292 -28180 -12228
rect -28284 -12308 -28180 -12292
rect -28284 -12372 -28264 -12308
rect -28200 -12372 -28180 -12308
rect -28284 -12388 -28180 -12372
rect -28284 -12452 -28264 -12388
rect -28200 -12452 -28180 -12388
rect -28284 -12468 -28180 -12452
rect -28284 -12532 -28264 -12468
rect -28200 -12532 -28180 -12468
rect -28284 -12548 -28180 -12532
rect -28284 -12612 -28264 -12548
rect -28200 -12612 -28180 -12548
rect -28284 -12628 -28180 -12612
rect -28284 -12692 -28264 -12628
rect -28200 -12692 -28180 -12628
rect -28284 -12708 -28180 -12692
rect -28284 -12772 -28264 -12708
rect -28200 -12772 -28180 -12708
rect -28284 -12788 -28180 -12772
rect -28284 -12852 -28264 -12788
rect -28200 -12852 -28180 -12788
rect -28284 -12868 -28180 -12852
rect -28284 -12932 -28264 -12868
rect -28200 -12932 -28180 -12868
rect -28284 -12948 -28180 -12932
rect -28284 -13012 -28264 -12948
rect -28200 -13012 -28180 -12948
rect -28284 -13028 -28180 -13012
rect -28284 -13092 -28264 -13028
rect -28200 -13092 -28180 -13028
rect -28284 -13108 -28180 -13092
rect -28284 -13172 -28264 -13108
rect -28200 -13172 -28180 -13108
rect -28284 -13188 -28180 -13172
rect -28284 -13252 -28264 -13188
rect -28200 -13252 -28180 -13188
rect -28284 -13268 -28180 -13252
rect -28284 -13332 -28264 -13268
rect -28200 -13332 -28180 -13268
rect -28284 -13348 -28180 -13332
rect -28284 -13412 -28264 -13348
rect -28200 -13412 -28180 -13348
rect -28284 -13428 -28180 -13412
rect -28284 -13492 -28264 -13428
rect -28200 -13492 -28180 -13428
rect -28284 -13508 -28180 -13492
rect -28284 -13572 -28264 -13508
rect -28200 -13572 -28180 -13508
rect -28284 -13588 -28180 -13572
rect -28284 -13652 -28264 -13588
rect -28200 -13652 -28180 -13588
rect -28284 -13668 -28180 -13652
rect -28284 -13732 -28264 -13668
rect -28200 -13732 -28180 -13668
rect -28284 -13748 -28180 -13732
rect -28284 -13812 -28264 -13748
rect -28200 -13812 -28180 -13748
rect -28284 -13828 -28180 -13812
rect -28284 -13892 -28264 -13828
rect -28200 -13892 -28180 -13828
rect -28284 -13908 -28180 -13892
rect -28284 -13972 -28264 -13908
rect -28200 -13972 -28180 -13908
rect -28284 -13988 -28180 -13972
rect -28284 -14052 -28264 -13988
rect -28200 -14052 -28180 -13988
rect -28284 -14068 -28180 -14052
rect -28284 -14132 -28264 -14068
rect -28200 -14132 -28180 -14068
rect -28284 -14148 -28180 -14132
rect -28284 -14212 -28264 -14148
rect -28200 -14212 -28180 -14148
rect -28284 -14228 -28180 -14212
rect -28284 -14292 -28264 -14228
rect -28200 -14292 -28180 -14228
rect -28284 -14308 -28180 -14292
rect -28284 -14372 -28264 -14308
rect -28200 -14372 -28180 -14308
rect -28284 -14388 -28180 -14372
rect -28284 -14452 -28264 -14388
rect -28200 -14452 -28180 -14388
rect -28284 -14468 -28180 -14452
rect -28284 -14532 -28264 -14468
rect -28200 -14532 -28180 -14468
rect -28284 -14548 -28180 -14532
rect -28284 -14612 -28264 -14548
rect -28200 -14612 -28180 -14548
rect -28284 -14628 -28180 -14612
rect -28284 -14692 -28264 -14628
rect -28200 -14692 -28180 -14628
rect -28284 -14708 -28180 -14692
rect -28284 -14772 -28264 -14708
rect -28200 -14772 -28180 -14708
rect -28284 -14788 -28180 -14772
rect -28284 -14852 -28264 -14788
rect -28200 -14852 -28180 -14788
rect -28284 -14868 -28180 -14852
rect -28284 -14932 -28264 -14868
rect -28200 -14932 -28180 -14868
rect -28284 -14948 -28180 -14932
rect -28284 -15012 -28264 -14948
rect -28200 -15012 -28180 -14948
rect -28284 -15028 -28180 -15012
rect -28284 -15092 -28264 -15028
rect -28200 -15092 -28180 -15028
rect -28284 -15108 -28180 -15092
rect -28284 -15172 -28264 -15108
rect -28200 -15172 -28180 -15108
rect -28284 -15188 -28180 -15172
rect -28284 -15252 -28264 -15188
rect -28200 -15252 -28180 -15188
rect -28284 -15268 -28180 -15252
rect -28284 -15332 -28264 -15268
rect -28200 -15332 -28180 -15268
rect -28284 -15348 -28180 -15332
rect -28284 -15412 -28264 -15348
rect -28200 -15412 -28180 -15348
rect -28284 -15428 -28180 -15412
rect -28284 -15492 -28264 -15428
rect -28200 -15492 -28180 -15428
rect -28284 -15508 -28180 -15492
rect -28284 -15572 -28264 -15508
rect -28200 -15572 -28180 -15508
rect -28284 -15588 -28180 -15572
rect -28284 -15652 -28264 -15588
rect -28200 -15652 -28180 -15588
rect -28284 -15668 -28180 -15652
rect -28284 -15732 -28264 -15668
rect -28200 -15732 -28180 -15668
rect -28284 -15748 -28180 -15732
rect -33896 -16108 -33792 -15812
rect -39085 -16188 -34163 -16159
rect -39085 -21052 -39056 -16188
rect -34192 -21052 -34163 -16188
rect -39085 -21081 -34163 -21052
rect -33896 -16172 -33876 -16108
rect -33812 -16172 -33792 -16108
rect -31064 -16159 -30960 -15761
rect -28284 -15812 -28264 -15748
rect -28200 -15812 -28180 -15748
rect -27861 -10868 -22939 -10839
rect -27861 -15732 -27832 -10868
rect -22968 -15732 -22939 -10868
rect -27861 -15761 -22939 -15732
rect -22672 -10852 -22652 -10788
rect -22588 -10852 -22568 -10788
rect -19840 -10839 -19736 -10441
rect -17060 -10492 -17040 -10428
rect -16976 -10492 -16956 -10428
rect -16637 -5548 -11715 -5519
rect -16637 -10412 -16608 -5548
rect -11744 -10412 -11715 -5548
rect -16637 -10441 -11715 -10412
rect -11448 -5532 -11428 -5468
rect -11364 -5532 -11344 -5468
rect -8616 -5519 -8512 -5121
rect -5836 -5172 -5816 -5108
rect -5752 -5172 -5732 -5108
rect -5413 -228 -491 -199
rect -5413 -5092 -5384 -228
rect -520 -5092 -491 -228
rect -5413 -5121 -491 -5092
rect -224 -212 -204 -148
rect -140 -212 -120 -148
rect 2608 -199 2712 199
rect 5388 148 5408 212
rect 5472 148 5492 212
rect 5811 5092 10733 5121
rect 5811 228 5840 5092
rect 10704 228 10733 5092
rect 5811 199 10733 228
rect 11000 5108 11020 5172
rect 11084 5108 11104 5172
rect 13832 5121 13936 5519
rect 16612 5468 16632 5532
rect 16696 5468 16716 5532
rect 17035 10412 21957 10441
rect 17035 5548 17064 10412
rect 21928 5548 21957 10412
rect 17035 5519 21957 5548
rect 22224 10428 22244 10492
rect 22308 10428 22328 10492
rect 25056 10441 25160 10839
rect 27836 10788 27856 10852
rect 27920 10788 27940 10852
rect 28259 15732 33181 15761
rect 28259 10868 28288 15732
rect 33152 10868 33181 15732
rect 28259 10839 33181 10868
rect 33448 15748 33468 15812
rect 33532 15748 33552 15812
rect 36280 15761 36384 16159
rect 39060 16108 39080 16172
rect 39144 16108 39164 16172
rect 39060 15812 39164 16108
rect 33448 15732 33552 15748
rect 33448 15668 33468 15732
rect 33532 15668 33552 15732
rect 33448 15652 33552 15668
rect 33448 15588 33468 15652
rect 33532 15588 33552 15652
rect 33448 15572 33552 15588
rect 33448 15508 33468 15572
rect 33532 15508 33552 15572
rect 33448 15492 33552 15508
rect 33448 15428 33468 15492
rect 33532 15428 33552 15492
rect 33448 15412 33552 15428
rect 33448 15348 33468 15412
rect 33532 15348 33552 15412
rect 33448 15332 33552 15348
rect 33448 15268 33468 15332
rect 33532 15268 33552 15332
rect 33448 15252 33552 15268
rect 33448 15188 33468 15252
rect 33532 15188 33552 15252
rect 33448 15172 33552 15188
rect 33448 15108 33468 15172
rect 33532 15108 33552 15172
rect 33448 15092 33552 15108
rect 33448 15028 33468 15092
rect 33532 15028 33552 15092
rect 33448 15012 33552 15028
rect 33448 14948 33468 15012
rect 33532 14948 33552 15012
rect 33448 14932 33552 14948
rect 33448 14868 33468 14932
rect 33532 14868 33552 14932
rect 33448 14852 33552 14868
rect 33448 14788 33468 14852
rect 33532 14788 33552 14852
rect 33448 14772 33552 14788
rect 33448 14708 33468 14772
rect 33532 14708 33552 14772
rect 33448 14692 33552 14708
rect 33448 14628 33468 14692
rect 33532 14628 33552 14692
rect 33448 14612 33552 14628
rect 33448 14548 33468 14612
rect 33532 14548 33552 14612
rect 33448 14532 33552 14548
rect 33448 14468 33468 14532
rect 33532 14468 33552 14532
rect 33448 14452 33552 14468
rect 33448 14388 33468 14452
rect 33532 14388 33552 14452
rect 33448 14372 33552 14388
rect 33448 14308 33468 14372
rect 33532 14308 33552 14372
rect 33448 14292 33552 14308
rect 33448 14228 33468 14292
rect 33532 14228 33552 14292
rect 33448 14212 33552 14228
rect 33448 14148 33468 14212
rect 33532 14148 33552 14212
rect 33448 14132 33552 14148
rect 33448 14068 33468 14132
rect 33532 14068 33552 14132
rect 33448 14052 33552 14068
rect 33448 13988 33468 14052
rect 33532 13988 33552 14052
rect 33448 13972 33552 13988
rect 33448 13908 33468 13972
rect 33532 13908 33552 13972
rect 33448 13892 33552 13908
rect 33448 13828 33468 13892
rect 33532 13828 33552 13892
rect 33448 13812 33552 13828
rect 33448 13748 33468 13812
rect 33532 13748 33552 13812
rect 33448 13732 33552 13748
rect 33448 13668 33468 13732
rect 33532 13668 33552 13732
rect 33448 13652 33552 13668
rect 33448 13588 33468 13652
rect 33532 13588 33552 13652
rect 33448 13572 33552 13588
rect 33448 13508 33468 13572
rect 33532 13508 33552 13572
rect 33448 13492 33552 13508
rect 33448 13428 33468 13492
rect 33532 13428 33552 13492
rect 33448 13412 33552 13428
rect 33448 13348 33468 13412
rect 33532 13348 33552 13412
rect 33448 13332 33552 13348
rect 33448 13268 33468 13332
rect 33532 13268 33552 13332
rect 33448 13252 33552 13268
rect 33448 13188 33468 13252
rect 33532 13188 33552 13252
rect 33448 13172 33552 13188
rect 33448 13108 33468 13172
rect 33532 13108 33552 13172
rect 33448 13092 33552 13108
rect 33448 13028 33468 13092
rect 33532 13028 33552 13092
rect 33448 13012 33552 13028
rect 33448 12948 33468 13012
rect 33532 12948 33552 13012
rect 33448 12932 33552 12948
rect 33448 12868 33468 12932
rect 33532 12868 33552 12932
rect 33448 12852 33552 12868
rect 33448 12788 33468 12852
rect 33532 12788 33552 12852
rect 33448 12772 33552 12788
rect 33448 12708 33468 12772
rect 33532 12708 33552 12772
rect 33448 12692 33552 12708
rect 33448 12628 33468 12692
rect 33532 12628 33552 12692
rect 33448 12612 33552 12628
rect 33448 12548 33468 12612
rect 33532 12548 33552 12612
rect 33448 12532 33552 12548
rect 33448 12468 33468 12532
rect 33532 12468 33552 12532
rect 33448 12452 33552 12468
rect 33448 12388 33468 12452
rect 33532 12388 33552 12452
rect 33448 12372 33552 12388
rect 33448 12308 33468 12372
rect 33532 12308 33552 12372
rect 33448 12292 33552 12308
rect 33448 12228 33468 12292
rect 33532 12228 33552 12292
rect 33448 12212 33552 12228
rect 33448 12148 33468 12212
rect 33532 12148 33552 12212
rect 33448 12132 33552 12148
rect 33448 12068 33468 12132
rect 33532 12068 33552 12132
rect 33448 12052 33552 12068
rect 33448 11988 33468 12052
rect 33532 11988 33552 12052
rect 33448 11972 33552 11988
rect 33448 11908 33468 11972
rect 33532 11908 33552 11972
rect 33448 11892 33552 11908
rect 33448 11828 33468 11892
rect 33532 11828 33552 11892
rect 33448 11812 33552 11828
rect 33448 11748 33468 11812
rect 33532 11748 33552 11812
rect 33448 11732 33552 11748
rect 33448 11668 33468 11732
rect 33532 11668 33552 11732
rect 33448 11652 33552 11668
rect 33448 11588 33468 11652
rect 33532 11588 33552 11652
rect 33448 11572 33552 11588
rect 33448 11508 33468 11572
rect 33532 11508 33552 11572
rect 33448 11492 33552 11508
rect 33448 11428 33468 11492
rect 33532 11428 33552 11492
rect 33448 11412 33552 11428
rect 33448 11348 33468 11412
rect 33532 11348 33552 11412
rect 33448 11332 33552 11348
rect 33448 11268 33468 11332
rect 33532 11268 33552 11332
rect 33448 11252 33552 11268
rect 33448 11188 33468 11252
rect 33532 11188 33552 11252
rect 33448 11172 33552 11188
rect 33448 11108 33468 11172
rect 33532 11108 33552 11172
rect 33448 11092 33552 11108
rect 33448 11028 33468 11092
rect 33532 11028 33552 11092
rect 33448 11012 33552 11028
rect 33448 10948 33468 11012
rect 33532 10948 33552 11012
rect 33448 10932 33552 10948
rect 33448 10868 33468 10932
rect 33532 10868 33552 10932
rect 33448 10852 33552 10868
rect 27836 10492 27940 10788
rect 22224 10412 22328 10428
rect 22224 10348 22244 10412
rect 22308 10348 22328 10412
rect 22224 10332 22328 10348
rect 22224 10268 22244 10332
rect 22308 10268 22328 10332
rect 22224 10252 22328 10268
rect 22224 10188 22244 10252
rect 22308 10188 22328 10252
rect 22224 10172 22328 10188
rect 22224 10108 22244 10172
rect 22308 10108 22328 10172
rect 22224 10092 22328 10108
rect 22224 10028 22244 10092
rect 22308 10028 22328 10092
rect 22224 10012 22328 10028
rect 22224 9948 22244 10012
rect 22308 9948 22328 10012
rect 22224 9932 22328 9948
rect 22224 9868 22244 9932
rect 22308 9868 22328 9932
rect 22224 9852 22328 9868
rect 22224 9788 22244 9852
rect 22308 9788 22328 9852
rect 22224 9772 22328 9788
rect 22224 9708 22244 9772
rect 22308 9708 22328 9772
rect 22224 9692 22328 9708
rect 22224 9628 22244 9692
rect 22308 9628 22328 9692
rect 22224 9612 22328 9628
rect 22224 9548 22244 9612
rect 22308 9548 22328 9612
rect 22224 9532 22328 9548
rect 22224 9468 22244 9532
rect 22308 9468 22328 9532
rect 22224 9452 22328 9468
rect 22224 9388 22244 9452
rect 22308 9388 22328 9452
rect 22224 9372 22328 9388
rect 22224 9308 22244 9372
rect 22308 9308 22328 9372
rect 22224 9292 22328 9308
rect 22224 9228 22244 9292
rect 22308 9228 22328 9292
rect 22224 9212 22328 9228
rect 22224 9148 22244 9212
rect 22308 9148 22328 9212
rect 22224 9132 22328 9148
rect 22224 9068 22244 9132
rect 22308 9068 22328 9132
rect 22224 9052 22328 9068
rect 22224 8988 22244 9052
rect 22308 8988 22328 9052
rect 22224 8972 22328 8988
rect 22224 8908 22244 8972
rect 22308 8908 22328 8972
rect 22224 8892 22328 8908
rect 22224 8828 22244 8892
rect 22308 8828 22328 8892
rect 22224 8812 22328 8828
rect 22224 8748 22244 8812
rect 22308 8748 22328 8812
rect 22224 8732 22328 8748
rect 22224 8668 22244 8732
rect 22308 8668 22328 8732
rect 22224 8652 22328 8668
rect 22224 8588 22244 8652
rect 22308 8588 22328 8652
rect 22224 8572 22328 8588
rect 22224 8508 22244 8572
rect 22308 8508 22328 8572
rect 22224 8492 22328 8508
rect 22224 8428 22244 8492
rect 22308 8428 22328 8492
rect 22224 8412 22328 8428
rect 22224 8348 22244 8412
rect 22308 8348 22328 8412
rect 22224 8332 22328 8348
rect 22224 8268 22244 8332
rect 22308 8268 22328 8332
rect 22224 8252 22328 8268
rect 22224 8188 22244 8252
rect 22308 8188 22328 8252
rect 22224 8172 22328 8188
rect 22224 8108 22244 8172
rect 22308 8108 22328 8172
rect 22224 8092 22328 8108
rect 22224 8028 22244 8092
rect 22308 8028 22328 8092
rect 22224 8012 22328 8028
rect 22224 7948 22244 8012
rect 22308 7948 22328 8012
rect 22224 7932 22328 7948
rect 22224 7868 22244 7932
rect 22308 7868 22328 7932
rect 22224 7852 22328 7868
rect 22224 7788 22244 7852
rect 22308 7788 22328 7852
rect 22224 7772 22328 7788
rect 22224 7708 22244 7772
rect 22308 7708 22328 7772
rect 22224 7692 22328 7708
rect 22224 7628 22244 7692
rect 22308 7628 22328 7692
rect 22224 7612 22328 7628
rect 22224 7548 22244 7612
rect 22308 7548 22328 7612
rect 22224 7532 22328 7548
rect 22224 7468 22244 7532
rect 22308 7468 22328 7532
rect 22224 7452 22328 7468
rect 22224 7388 22244 7452
rect 22308 7388 22328 7452
rect 22224 7372 22328 7388
rect 22224 7308 22244 7372
rect 22308 7308 22328 7372
rect 22224 7292 22328 7308
rect 22224 7228 22244 7292
rect 22308 7228 22328 7292
rect 22224 7212 22328 7228
rect 22224 7148 22244 7212
rect 22308 7148 22328 7212
rect 22224 7132 22328 7148
rect 22224 7068 22244 7132
rect 22308 7068 22328 7132
rect 22224 7052 22328 7068
rect 22224 6988 22244 7052
rect 22308 6988 22328 7052
rect 22224 6972 22328 6988
rect 22224 6908 22244 6972
rect 22308 6908 22328 6972
rect 22224 6892 22328 6908
rect 22224 6828 22244 6892
rect 22308 6828 22328 6892
rect 22224 6812 22328 6828
rect 22224 6748 22244 6812
rect 22308 6748 22328 6812
rect 22224 6732 22328 6748
rect 22224 6668 22244 6732
rect 22308 6668 22328 6732
rect 22224 6652 22328 6668
rect 22224 6588 22244 6652
rect 22308 6588 22328 6652
rect 22224 6572 22328 6588
rect 22224 6508 22244 6572
rect 22308 6508 22328 6572
rect 22224 6492 22328 6508
rect 22224 6428 22244 6492
rect 22308 6428 22328 6492
rect 22224 6412 22328 6428
rect 22224 6348 22244 6412
rect 22308 6348 22328 6412
rect 22224 6332 22328 6348
rect 22224 6268 22244 6332
rect 22308 6268 22328 6332
rect 22224 6252 22328 6268
rect 22224 6188 22244 6252
rect 22308 6188 22328 6252
rect 22224 6172 22328 6188
rect 22224 6108 22244 6172
rect 22308 6108 22328 6172
rect 22224 6092 22328 6108
rect 22224 6028 22244 6092
rect 22308 6028 22328 6092
rect 22224 6012 22328 6028
rect 22224 5948 22244 6012
rect 22308 5948 22328 6012
rect 22224 5932 22328 5948
rect 22224 5868 22244 5932
rect 22308 5868 22328 5932
rect 22224 5852 22328 5868
rect 22224 5788 22244 5852
rect 22308 5788 22328 5852
rect 22224 5772 22328 5788
rect 22224 5708 22244 5772
rect 22308 5708 22328 5772
rect 22224 5692 22328 5708
rect 22224 5628 22244 5692
rect 22308 5628 22328 5692
rect 22224 5612 22328 5628
rect 22224 5548 22244 5612
rect 22308 5548 22328 5612
rect 22224 5532 22328 5548
rect 16612 5172 16716 5468
rect 11000 5092 11104 5108
rect 11000 5028 11020 5092
rect 11084 5028 11104 5092
rect 11000 5012 11104 5028
rect 11000 4948 11020 5012
rect 11084 4948 11104 5012
rect 11000 4932 11104 4948
rect 11000 4868 11020 4932
rect 11084 4868 11104 4932
rect 11000 4852 11104 4868
rect 11000 4788 11020 4852
rect 11084 4788 11104 4852
rect 11000 4772 11104 4788
rect 11000 4708 11020 4772
rect 11084 4708 11104 4772
rect 11000 4692 11104 4708
rect 11000 4628 11020 4692
rect 11084 4628 11104 4692
rect 11000 4612 11104 4628
rect 11000 4548 11020 4612
rect 11084 4548 11104 4612
rect 11000 4532 11104 4548
rect 11000 4468 11020 4532
rect 11084 4468 11104 4532
rect 11000 4452 11104 4468
rect 11000 4388 11020 4452
rect 11084 4388 11104 4452
rect 11000 4372 11104 4388
rect 11000 4308 11020 4372
rect 11084 4308 11104 4372
rect 11000 4292 11104 4308
rect 11000 4228 11020 4292
rect 11084 4228 11104 4292
rect 11000 4212 11104 4228
rect 11000 4148 11020 4212
rect 11084 4148 11104 4212
rect 11000 4132 11104 4148
rect 11000 4068 11020 4132
rect 11084 4068 11104 4132
rect 11000 4052 11104 4068
rect 11000 3988 11020 4052
rect 11084 3988 11104 4052
rect 11000 3972 11104 3988
rect 11000 3908 11020 3972
rect 11084 3908 11104 3972
rect 11000 3892 11104 3908
rect 11000 3828 11020 3892
rect 11084 3828 11104 3892
rect 11000 3812 11104 3828
rect 11000 3748 11020 3812
rect 11084 3748 11104 3812
rect 11000 3732 11104 3748
rect 11000 3668 11020 3732
rect 11084 3668 11104 3732
rect 11000 3652 11104 3668
rect 11000 3588 11020 3652
rect 11084 3588 11104 3652
rect 11000 3572 11104 3588
rect 11000 3508 11020 3572
rect 11084 3508 11104 3572
rect 11000 3492 11104 3508
rect 11000 3428 11020 3492
rect 11084 3428 11104 3492
rect 11000 3412 11104 3428
rect 11000 3348 11020 3412
rect 11084 3348 11104 3412
rect 11000 3332 11104 3348
rect 11000 3268 11020 3332
rect 11084 3268 11104 3332
rect 11000 3252 11104 3268
rect 11000 3188 11020 3252
rect 11084 3188 11104 3252
rect 11000 3172 11104 3188
rect 11000 3108 11020 3172
rect 11084 3108 11104 3172
rect 11000 3092 11104 3108
rect 11000 3028 11020 3092
rect 11084 3028 11104 3092
rect 11000 3012 11104 3028
rect 11000 2948 11020 3012
rect 11084 2948 11104 3012
rect 11000 2932 11104 2948
rect 11000 2868 11020 2932
rect 11084 2868 11104 2932
rect 11000 2852 11104 2868
rect 11000 2788 11020 2852
rect 11084 2788 11104 2852
rect 11000 2772 11104 2788
rect 11000 2708 11020 2772
rect 11084 2708 11104 2772
rect 11000 2692 11104 2708
rect 11000 2628 11020 2692
rect 11084 2628 11104 2692
rect 11000 2612 11104 2628
rect 11000 2548 11020 2612
rect 11084 2548 11104 2612
rect 11000 2532 11104 2548
rect 11000 2468 11020 2532
rect 11084 2468 11104 2532
rect 11000 2452 11104 2468
rect 11000 2388 11020 2452
rect 11084 2388 11104 2452
rect 11000 2372 11104 2388
rect 11000 2308 11020 2372
rect 11084 2308 11104 2372
rect 11000 2292 11104 2308
rect 11000 2228 11020 2292
rect 11084 2228 11104 2292
rect 11000 2212 11104 2228
rect 11000 2148 11020 2212
rect 11084 2148 11104 2212
rect 11000 2132 11104 2148
rect 11000 2068 11020 2132
rect 11084 2068 11104 2132
rect 11000 2052 11104 2068
rect 11000 1988 11020 2052
rect 11084 1988 11104 2052
rect 11000 1972 11104 1988
rect 11000 1908 11020 1972
rect 11084 1908 11104 1972
rect 11000 1892 11104 1908
rect 11000 1828 11020 1892
rect 11084 1828 11104 1892
rect 11000 1812 11104 1828
rect 11000 1748 11020 1812
rect 11084 1748 11104 1812
rect 11000 1732 11104 1748
rect 11000 1668 11020 1732
rect 11084 1668 11104 1732
rect 11000 1652 11104 1668
rect 11000 1588 11020 1652
rect 11084 1588 11104 1652
rect 11000 1572 11104 1588
rect 11000 1508 11020 1572
rect 11084 1508 11104 1572
rect 11000 1492 11104 1508
rect 11000 1428 11020 1492
rect 11084 1428 11104 1492
rect 11000 1412 11104 1428
rect 11000 1348 11020 1412
rect 11084 1348 11104 1412
rect 11000 1332 11104 1348
rect 11000 1268 11020 1332
rect 11084 1268 11104 1332
rect 11000 1252 11104 1268
rect 11000 1188 11020 1252
rect 11084 1188 11104 1252
rect 11000 1172 11104 1188
rect 11000 1108 11020 1172
rect 11084 1108 11104 1172
rect 11000 1092 11104 1108
rect 11000 1028 11020 1092
rect 11084 1028 11104 1092
rect 11000 1012 11104 1028
rect 11000 948 11020 1012
rect 11084 948 11104 1012
rect 11000 932 11104 948
rect 11000 868 11020 932
rect 11084 868 11104 932
rect 11000 852 11104 868
rect 11000 788 11020 852
rect 11084 788 11104 852
rect 11000 772 11104 788
rect 11000 708 11020 772
rect 11084 708 11104 772
rect 11000 692 11104 708
rect 11000 628 11020 692
rect 11084 628 11104 692
rect 11000 612 11104 628
rect 11000 548 11020 612
rect 11084 548 11104 612
rect 11000 532 11104 548
rect 11000 468 11020 532
rect 11084 468 11104 532
rect 11000 452 11104 468
rect 11000 388 11020 452
rect 11084 388 11104 452
rect 11000 372 11104 388
rect 11000 308 11020 372
rect 11084 308 11104 372
rect 11000 292 11104 308
rect 11000 228 11020 292
rect 11084 228 11104 292
rect 11000 212 11104 228
rect 5388 -148 5492 148
rect -224 -228 -120 -212
rect -224 -292 -204 -228
rect -140 -292 -120 -228
rect -224 -308 -120 -292
rect -224 -372 -204 -308
rect -140 -372 -120 -308
rect -224 -388 -120 -372
rect -224 -452 -204 -388
rect -140 -452 -120 -388
rect -224 -468 -120 -452
rect -224 -532 -204 -468
rect -140 -532 -120 -468
rect -224 -548 -120 -532
rect -224 -612 -204 -548
rect -140 -612 -120 -548
rect -224 -628 -120 -612
rect -224 -692 -204 -628
rect -140 -692 -120 -628
rect -224 -708 -120 -692
rect -224 -772 -204 -708
rect -140 -772 -120 -708
rect -224 -788 -120 -772
rect -224 -852 -204 -788
rect -140 -852 -120 -788
rect -224 -868 -120 -852
rect -224 -932 -204 -868
rect -140 -932 -120 -868
rect -224 -948 -120 -932
rect -224 -1012 -204 -948
rect -140 -1012 -120 -948
rect -224 -1028 -120 -1012
rect -224 -1092 -204 -1028
rect -140 -1092 -120 -1028
rect -224 -1108 -120 -1092
rect -224 -1172 -204 -1108
rect -140 -1172 -120 -1108
rect -224 -1188 -120 -1172
rect -224 -1252 -204 -1188
rect -140 -1252 -120 -1188
rect -224 -1268 -120 -1252
rect -224 -1332 -204 -1268
rect -140 -1332 -120 -1268
rect -224 -1348 -120 -1332
rect -224 -1412 -204 -1348
rect -140 -1412 -120 -1348
rect -224 -1428 -120 -1412
rect -224 -1492 -204 -1428
rect -140 -1492 -120 -1428
rect -224 -1508 -120 -1492
rect -224 -1572 -204 -1508
rect -140 -1572 -120 -1508
rect -224 -1588 -120 -1572
rect -224 -1652 -204 -1588
rect -140 -1652 -120 -1588
rect -224 -1668 -120 -1652
rect -224 -1732 -204 -1668
rect -140 -1732 -120 -1668
rect -224 -1748 -120 -1732
rect -224 -1812 -204 -1748
rect -140 -1812 -120 -1748
rect -224 -1828 -120 -1812
rect -224 -1892 -204 -1828
rect -140 -1892 -120 -1828
rect -224 -1908 -120 -1892
rect -224 -1972 -204 -1908
rect -140 -1972 -120 -1908
rect -224 -1988 -120 -1972
rect -224 -2052 -204 -1988
rect -140 -2052 -120 -1988
rect -224 -2068 -120 -2052
rect -224 -2132 -204 -2068
rect -140 -2132 -120 -2068
rect -224 -2148 -120 -2132
rect -224 -2212 -204 -2148
rect -140 -2212 -120 -2148
rect -224 -2228 -120 -2212
rect -224 -2292 -204 -2228
rect -140 -2292 -120 -2228
rect -224 -2308 -120 -2292
rect -224 -2372 -204 -2308
rect -140 -2372 -120 -2308
rect -224 -2388 -120 -2372
rect -224 -2452 -204 -2388
rect -140 -2452 -120 -2388
rect -224 -2468 -120 -2452
rect -224 -2532 -204 -2468
rect -140 -2532 -120 -2468
rect -224 -2548 -120 -2532
rect -224 -2612 -204 -2548
rect -140 -2612 -120 -2548
rect -224 -2628 -120 -2612
rect -224 -2692 -204 -2628
rect -140 -2692 -120 -2628
rect -224 -2708 -120 -2692
rect -224 -2772 -204 -2708
rect -140 -2772 -120 -2708
rect -224 -2788 -120 -2772
rect -224 -2852 -204 -2788
rect -140 -2852 -120 -2788
rect -224 -2868 -120 -2852
rect -224 -2932 -204 -2868
rect -140 -2932 -120 -2868
rect -224 -2948 -120 -2932
rect -224 -3012 -204 -2948
rect -140 -3012 -120 -2948
rect -224 -3028 -120 -3012
rect -224 -3092 -204 -3028
rect -140 -3092 -120 -3028
rect -224 -3108 -120 -3092
rect -224 -3172 -204 -3108
rect -140 -3172 -120 -3108
rect -224 -3188 -120 -3172
rect -224 -3252 -204 -3188
rect -140 -3252 -120 -3188
rect -224 -3268 -120 -3252
rect -224 -3332 -204 -3268
rect -140 -3332 -120 -3268
rect -224 -3348 -120 -3332
rect -224 -3412 -204 -3348
rect -140 -3412 -120 -3348
rect -224 -3428 -120 -3412
rect -224 -3492 -204 -3428
rect -140 -3492 -120 -3428
rect -224 -3508 -120 -3492
rect -224 -3572 -204 -3508
rect -140 -3572 -120 -3508
rect -224 -3588 -120 -3572
rect -224 -3652 -204 -3588
rect -140 -3652 -120 -3588
rect -224 -3668 -120 -3652
rect -224 -3732 -204 -3668
rect -140 -3732 -120 -3668
rect -224 -3748 -120 -3732
rect -224 -3812 -204 -3748
rect -140 -3812 -120 -3748
rect -224 -3828 -120 -3812
rect -224 -3892 -204 -3828
rect -140 -3892 -120 -3828
rect -224 -3908 -120 -3892
rect -224 -3972 -204 -3908
rect -140 -3972 -120 -3908
rect -224 -3988 -120 -3972
rect -224 -4052 -204 -3988
rect -140 -4052 -120 -3988
rect -224 -4068 -120 -4052
rect -224 -4132 -204 -4068
rect -140 -4132 -120 -4068
rect -224 -4148 -120 -4132
rect -224 -4212 -204 -4148
rect -140 -4212 -120 -4148
rect -224 -4228 -120 -4212
rect -224 -4292 -204 -4228
rect -140 -4292 -120 -4228
rect -224 -4308 -120 -4292
rect -224 -4372 -204 -4308
rect -140 -4372 -120 -4308
rect -224 -4388 -120 -4372
rect -224 -4452 -204 -4388
rect -140 -4452 -120 -4388
rect -224 -4468 -120 -4452
rect -224 -4532 -204 -4468
rect -140 -4532 -120 -4468
rect -224 -4548 -120 -4532
rect -224 -4612 -204 -4548
rect -140 -4612 -120 -4548
rect -224 -4628 -120 -4612
rect -224 -4692 -204 -4628
rect -140 -4692 -120 -4628
rect -224 -4708 -120 -4692
rect -224 -4772 -204 -4708
rect -140 -4772 -120 -4708
rect -224 -4788 -120 -4772
rect -224 -4852 -204 -4788
rect -140 -4852 -120 -4788
rect -224 -4868 -120 -4852
rect -224 -4932 -204 -4868
rect -140 -4932 -120 -4868
rect -224 -4948 -120 -4932
rect -224 -5012 -204 -4948
rect -140 -5012 -120 -4948
rect -224 -5028 -120 -5012
rect -224 -5092 -204 -5028
rect -140 -5092 -120 -5028
rect -224 -5108 -120 -5092
rect -5836 -5468 -5732 -5172
rect -11448 -5548 -11344 -5532
rect -11448 -5612 -11428 -5548
rect -11364 -5612 -11344 -5548
rect -11448 -5628 -11344 -5612
rect -11448 -5692 -11428 -5628
rect -11364 -5692 -11344 -5628
rect -11448 -5708 -11344 -5692
rect -11448 -5772 -11428 -5708
rect -11364 -5772 -11344 -5708
rect -11448 -5788 -11344 -5772
rect -11448 -5852 -11428 -5788
rect -11364 -5852 -11344 -5788
rect -11448 -5868 -11344 -5852
rect -11448 -5932 -11428 -5868
rect -11364 -5932 -11344 -5868
rect -11448 -5948 -11344 -5932
rect -11448 -6012 -11428 -5948
rect -11364 -6012 -11344 -5948
rect -11448 -6028 -11344 -6012
rect -11448 -6092 -11428 -6028
rect -11364 -6092 -11344 -6028
rect -11448 -6108 -11344 -6092
rect -11448 -6172 -11428 -6108
rect -11364 -6172 -11344 -6108
rect -11448 -6188 -11344 -6172
rect -11448 -6252 -11428 -6188
rect -11364 -6252 -11344 -6188
rect -11448 -6268 -11344 -6252
rect -11448 -6332 -11428 -6268
rect -11364 -6332 -11344 -6268
rect -11448 -6348 -11344 -6332
rect -11448 -6412 -11428 -6348
rect -11364 -6412 -11344 -6348
rect -11448 -6428 -11344 -6412
rect -11448 -6492 -11428 -6428
rect -11364 -6492 -11344 -6428
rect -11448 -6508 -11344 -6492
rect -11448 -6572 -11428 -6508
rect -11364 -6572 -11344 -6508
rect -11448 -6588 -11344 -6572
rect -11448 -6652 -11428 -6588
rect -11364 -6652 -11344 -6588
rect -11448 -6668 -11344 -6652
rect -11448 -6732 -11428 -6668
rect -11364 -6732 -11344 -6668
rect -11448 -6748 -11344 -6732
rect -11448 -6812 -11428 -6748
rect -11364 -6812 -11344 -6748
rect -11448 -6828 -11344 -6812
rect -11448 -6892 -11428 -6828
rect -11364 -6892 -11344 -6828
rect -11448 -6908 -11344 -6892
rect -11448 -6972 -11428 -6908
rect -11364 -6972 -11344 -6908
rect -11448 -6988 -11344 -6972
rect -11448 -7052 -11428 -6988
rect -11364 -7052 -11344 -6988
rect -11448 -7068 -11344 -7052
rect -11448 -7132 -11428 -7068
rect -11364 -7132 -11344 -7068
rect -11448 -7148 -11344 -7132
rect -11448 -7212 -11428 -7148
rect -11364 -7212 -11344 -7148
rect -11448 -7228 -11344 -7212
rect -11448 -7292 -11428 -7228
rect -11364 -7292 -11344 -7228
rect -11448 -7308 -11344 -7292
rect -11448 -7372 -11428 -7308
rect -11364 -7372 -11344 -7308
rect -11448 -7388 -11344 -7372
rect -11448 -7452 -11428 -7388
rect -11364 -7452 -11344 -7388
rect -11448 -7468 -11344 -7452
rect -11448 -7532 -11428 -7468
rect -11364 -7532 -11344 -7468
rect -11448 -7548 -11344 -7532
rect -11448 -7612 -11428 -7548
rect -11364 -7612 -11344 -7548
rect -11448 -7628 -11344 -7612
rect -11448 -7692 -11428 -7628
rect -11364 -7692 -11344 -7628
rect -11448 -7708 -11344 -7692
rect -11448 -7772 -11428 -7708
rect -11364 -7772 -11344 -7708
rect -11448 -7788 -11344 -7772
rect -11448 -7852 -11428 -7788
rect -11364 -7852 -11344 -7788
rect -11448 -7868 -11344 -7852
rect -11448 -7932 -11428 -7868
rect -11364 -7932 -11344 -7868
rect -11448 -7948 -11344 -7932
rect -11448 -8012 -11428 -7948
rect -11364 -8012 -11344 -7948
rect -11448 -8028 -11344 -8012
rect -11448 -8092 -11428 -8028
rect -11364 -8092 -11344 -8028
rect -11448 -8108 -11344 -8092
rect -11448 -8172 -11428 -8108
rect -11364 -8172 -11344 -8108
rect -11448 -8188 -11344 -8172
rect -11448 -8252 -11428 -8188
rect -11364 -8252 -11344 -8188
rect -11448 -8268 -11344 -8252
rect -11448 -8332 -11428 -8268
rect -11364 -8332 -11344 -8268
rect -11448 -8348 -11344 -8332
rect -11448 -8412 -11428 -8348
rect -11364 -8412 -11344 -8348
rect -11448 -8428 -11344 -8412
rect -11448 -8492 -11428 -8428
rect -11364 -8492 -11344 -8428
rect -11448 -8508 -11344 -8492
rect -11448 -8572 -11428 -8508
rect -11364 -8572 -11344 -8508
rect -11448 -8588 -11344 -8572
rect -11448 -8652 -11428 -8588
rect -11364 -8652 -11344 -8588
rect -11448 -8668 -11344 -8652
rect -11448 -8732 -11428 -8668
rect -11364 -8732 -11344 -8668
rect -11448 -8748 -11344 -8732
rect -11448 -8812 -11428 -8748
rect -11364 -8812 -11344 -8748
rect -11448 -8828 -11344 -8812
rect -11448 -8892 -11428 -8828
rect -11364 -8892 -11344 -8828
rect -11448 -8908 -11344 -8892
rect -11448 -8972 -11428 -8908
rect -11364 -8972 -11344 -8908
rect -11448 -8988 -11344 -8972
rect -11448 -9052 -11428 -8988
rect -11364 -9052 -11344 -8988
rect -11448 -9068 -11344 -9052
rect -11448 -9132 -11428 -9068
rect -11364 -9132 -11344 -9068
rect -11448 -9148 -11344 -9132
rect -11448 -9212 -11428 -9148
rect -11364 -9212 -11344 -9148
rect -11448 -9228 -11344 -9212
rect -11448 -9292 -11428 -9228
rect -11364 -9292 -11344 -9228
rect -11448 -9308 -11344 -9292
rect -11448 -9372 -11428 -9308
rect -11364 -9372 -11344 -9308
rect -11448 -9388 -11344 -9372
rect -11448 -9452 -11428 -9388
rect -11364 -9452 -11344 -9388
rect -11448 -9468 -11344 -9452
rect -11448 -9532 -11428 -9468
rect -11364 -9532 -11344 -9468
rect -11448 -9548 -11344 -9532
rect -11448 -9612 -11428 -9548
rect -11364 -9612 -11344 -9548
rect -11448 -9628 -11344 -9612
rect -11448 -9692 -11428 -9628
rect -11364 -9692 -11344 -9628
rect -11448 -9708 -11344 -9692
rect -11448 -9772 -11428 -9708
rect -11364 -9772 -11344 -9708
rect -11448 -9788 -11344 -9772
rect -11448 -9852 -11428 -9788
rect -11364 -9852 -11344 -9788
rect -11448 -9868 -11344 -9852
rect -11448 -9932 -11428 -9868
rect -11364 -9932 -11344 -9868
rect -11448 -9948 -11344 -9932
rect -11448 -10012 -11428 -9948
rect -11364 -10012 -11344 -9948
rect -11448 -10028 -11344 -10012
rect -11448 -10092 -11428 -10028
rect -11364 -10092 -11344 -10028
rect -11448 -10108 -11344 -10092
rect -11448 -10172 -11428 -10108
rect -11364 -10172 -11344 -10108
rect -11448 -10188 -11344 -10172
rect -11448 -10252 -11428 -10188
rect -11364 -10252 -11344 -10188
rect -11448 -10268 -11344 -10252
rect -11448 -10332 -11428 -10268
rect -11364 -10332 -11344 -10268
rect -11448 -10348 -11344 -10332
rect -11448 -10412 -11428 -10348
rect -11364 -10412 -11344 -10348
rect -11448 -10428 -11344 -10412
rect -17060 -10788 -16956 -10492
rect -22672 -10868 -22568 -10852
rect -22672 -10932 -22652 -10868
rect -22588 -10932 -22568 -10868
rect -22672 -10948 -22568 -10932
rect -22672 -11012 -22652 -10948
rect -22588 -11012 -22568 -10948
rect -22672 -11028 -22568 -11012
rect -22672 -11092 -22652 -11028
rect -22588 -11092 -22568 -11028
rect -22672 -11108 -22568 -11092
rect -22672 -11172 -22652 -11108
rect -22588 -11172 -22568 -11108
rect -22672 -11188 -22568 -11172
rect -22672 -11252 -22652 -11188
rect -22588 -11252 -22568 -11188
rect -22672 -11268 -22568 -11252
rect -22672 -11332 -22652 -11268
rect -22588 -11332 -22568 -11268
rect -22672 -11348 -22568 -11332
rect -22672 -11412 -22652 -11348
rect -22588 -11412 -22568 -11348
rect -22672 -11428 -22568 -11412
rect -22672 -11492 -22652 -11428
rect -22588 -11492 -22568 -11428
rect -22672 -11508 -22568 -11492
rect -22672 -11572 -22652 -11508
rect -22588 -11572 -22568 -11508
rect -22672 -11588 -22568 -11572
rect -22672 -11652 -22652 -11588
rect -22588 -11652 -22568 -11588
rect -22672 -11668 -22568 -11652
rect -22672 -11732 -22652 -11668
rect -22588 -11732 -22568 -11668
rect -22672 -11748 -22568 -11732
rect -22672 -11812 -22652 -11748
rect -22588 -11812 -22568 -11748
rect -22672 -11828 -22568 -11812
rect -22672 -11892 -22652 -11828
rect -22588 -11892 -22568 -11828
rect -22672 -11908 -22568 -11892
rect -22672 -11972 -22652 -11908
rect -22588 -11972 -22568 -11908
rect -22672 -11988 -22568 -11972
rect -22672 -12052 -22652 -11988
rect -22588 -12052 -22568 -11988
rect -22672 -12068 -22568 -12052
rect -22672 -12132 -22652 -12068
rect -22588 -12132 -22568 -12068
rect -22672 -12148 -22568 -12132
rect -22672 -12212 -22652 -12148
rect -22588 -12212 -22568 -12148
rect -22672 -12228 -22568 -12212
rect -22672 -12292 -22652 -12228
rect -22588 -12292 -22568 -12228
rect -22672 -12308 -22568 -12292
rect -22672 -12372 -22652 -12308
rect -22588 -12372 -22568 -12308
rect -22672 -12388 -22568 -12372
rect -22672 -12452 -22652 -12388
rect -22588 -12452 -22568 -12388
rect -22672 -12468 -22568 -12452
rect -22672 -12532 -22652 -12468
rect -22588 -12532 -22568 -12468
rect -22672 -12548 -22568 -12532
rect -22672 -12612 -22652 -12548
rect -22588 -12612 -22568 -12548
rect -22672 -12628 -22568 -12612
rect -22672 -12692 -22652 -12628
rect -22588 -12692 -22568 -12628
rect -22672 -12708 -22568 -12692
rect -22672 -12772 -22652 -12708
rect -22588 -12772 -22568 -12708
rect -22672 -12788 -22568 -12772
rect -22672 -12852 -22652 -12788
rect -22588 -12852 -22568 -12788
rect -22672 -12868 -22568 -12852
rect -22672 -12932 -22652 -12868
rect -22588 -12932 -22568 -12868
rect -22672 -12948 -22568 -12932
rect -22672 -13012 -22652 -12948
rect -22588 -13012 -22568 -12948
rect -22672 -13028 -22568 -13012
rect -22672 -13092 -22652 -13028
rect -22588 -13092 -22568 -13028
rect -22672 -13108 -22568 -13092
rect -22672 -13172 -22652 -13108
rect -22588 -13172 -22568 -13108
rect -22672 -13188 -22568 -13172
rect -22672 -13252 -22652 -13188
rect -22588 -13252 -22568 -13188
rect -22672 -13268 -22568 -13252
rect -22672 -13332 -22652 -13268
rect -22588 -13332 -22568 -13268
rect -22672 -13348 -22568 -13332
rect -22672 -13412 -22652 -13348
rect -22588 -13412 -22568 -13348
rect -22672 -13428 -22568 -13412
rect -22672 -13492 -22652 -13428
rect -22588 -13492 -22568 -13428
rect -22672 -13508 -22568 -13492
rect -22672 -13572 -22652 -13508
rect -22588 -13572 -22568 -13508
rect -22672 -13588 -22568 -13572
rect -22672 -13652 -22652 -13588
rect -22588 -13652 -22568 -13588
rect -22672 -13668 -22568 -13652
rect -22672 -13732 -22652 -13668
rect -22588 -13732 -22568 -13668
rect -22672 -13748 -22568 -13732
rect -22672 -13812 -22652 -13748
rect -22588 -13812 -22568 -13748
rect -22672 -13828 -22568 -13812
rect -22672 -13892 -22652 -13828
rect -22588 -13892 -22568 -13828
rect -22672 -13908 -22568 -13892
rect -22672 -13972 -22652 -13908
rect -22588 -13972 -22568 -13908
rect -22672 -13988 -22568 -13972
rect -22672 -14052 -22652 -13988
rect -22588 -14052 -22568 -13988
rect -22672 -14068 -22568 -14052
rect -22672 -14132 -22652 -14068
rect -22588 -14132 -22568 -14068
rect -22672 -14148 -22568 -14132
rect -22672 -14212 -22652 -14148
rect -22588 -14212 -22568 -14148
rect -22672 -14228 -22568 -14212
rect -22672 -14292 -22652 -14228
rect -22588 -14292 -22568 -14228
rect -22672 -14308 -22568 -14292
rect -22672 -14372 -22652 -14308
rect -22588 -14372 -22568 -14308
rect -22672 -14388 -22568 -14372
rect -22672 -14452 -22652 -14388
rect -22588 -14452 -22568 -14388
rect -22672 -14468 -22568 -14452
rect -22672 -14532 -22652 -14468
rect -22588 -14532 -22568 -14468
rect -22672 -14548 -22568 -14532
rect -22672 -14612 -22652 -14548
rect -22588 -14612 -22568 -14548
rect -22672 -14628 -22568 -14612
rect -22672 -14692 -22652 -14628
rect -22588 -14692 -22568 -14628
rect -22672 -14708 -22568 -14692
rect -22672 -14772 -22652 -14708
rect -22588 -14772 -22568 -14708
rect -22672 -14788 -22568 -14772
rect -22672 -14852 -22652 -14788
rect -22588 -14852 -22568 -14788
rect -22672 -14868 -22568 -14852
rect -22672 -14932 -22652 -14868
rect -22588 -14932 -22568 -14868
rect -22672 -14948 -22568 -14932
rect -22672 -15012 -22652 -14948
rect -22588 -15012 -22568 -14948
rect -22672 -15028 -22568 -15012
rect -22672 -15092 -22652 -15028
rect -22588 -15092 -22568 -15028
rect -22672 -15108 -22568 -15092
rect -22672 -15172 -22652 -15108
rect -22588 -15172 -22568 -15108
rect -22672 -15188 -22568 -15172
rect -22672 -15252 -22652 -15188
rect -22588 -15252 -22568 -15188
rect -22672 -15268 -22568 -15252
rect -22672 -15332 -22652 -15268
rect -22588 -15332 -22568 -15268
rect -22672 -15348 -22568 -15332
rect -22672 -15412 -22652 -15348
rect -22588 -15412 -22568 -15348
rect -22672 -15428 -22568 -15412
rect -22672 -15492 -22652 -15428
rect -22588 -15492 -22568 -15428
rect -22672 -15508 -22568 -15492
rect -22672 -15572 -22652 -15508
rect -22588 -15572 -22568 -15508
rect -22672 -15588 -22568 -15572
rect -22672 -15652 -22652 -15588
rect -22588 -15652 -22568 -15588
rect -22672 -15668 -22568 -15652
rect -22672 -15732 -22652 -15668
rect -22588 -15732 -22568 -15668
rect -22672 -15748 -22568 -15732
rect -28284 -16108 -28180 -15812
rect -33896 -16188 -33792 -16172
rect -33896 -16252 -33876 -16188
rect -33812 -16252 -33792 -16188
rect -33896 -16268 -33792 -16252
rect -33896 -16332 -33876 -16268
rect -33812 -16332 -33792 -16268
rect -33896 -16348 -33792 -16332
rect -33896 -16412 -33876 -16348
rect -33812 -16412 -33792 -16348
rect -33896 -16428 -33792 -16412
rect -33896 -16492 -33876 -16428
rect -33812 -16492 -33792 -16428
rect -33896 -16508 -33792 -16492
rect -33896 -16572 -33876 -16508
rect -33812 -16572 -33792 -16508
rect -33896 -16588 -33792 -16572
rect -33896 -16652 -33876 -16588
rect -33812 -16652 -33792 -16588
rect -33896 -16668 -33792 -16652
rect -33896 -16732 -33876 -16668
rect -33812 -16732 -33792 -16668
rect -33896 -16748 -33792 -16732
rect -33896 -16812 -33876 -16748
rect -33812 -16812 -33792 -16748
rect -33896 -16828 -33792 -16812
rect -33896 -16892 -33876 -16828
rect -33812 -16892 -33792 -16828
rect -33896 -16908 -33792 -16892
rect -33896 -16972 -33876 -16908
rect -33812 -16972 -33792 -16908
rect -33896 -16988 -33792 -16972
rect -33896 -17052 -33876 -16988
rect -33812 -17052 -33792 -16988
rect -33896 -17068 -33792 -17052
rect -33896 -17132 -33876 -17068
rect -33812 -17132 -33792 -17068
rect -33896 -17148 -33792 -17132
rect -33896 -17212 -33876 -17148
rect -33812 -17212 -33792 -17148
rect -33896 -17228 -33792 -17212
rect -33896 -17292 -33876 -17228
rect -33812 -17292 -33792 -17228
rect -33896 -17308 -33792 -17292
rect -33896 -17372 -33876 -17308
rect -33812 -17372 -33792 -17308
rect -33896 -17388 -33792 -17372
rect -33896 -17452 -33876 -17388
rect -33812 -17452 -33792 -17388
rect -33896 -17468 -33792 -17452
rect -33896 -17532 -33876 -17468
rect -33812 -17532 -33792 -17468
rect -33896 -17548 -33792 -17532
rect -33896 -17612 -33876 -17548
rect -33812 -17612 -33792 -17548
rect -33896 -17628 -33792 -17612
rect -33896 -17692 -33876 -17628
rect -33812 -17692 -33792 -17628
rect -33896 -17708 -33792 -17692
rect -33896 -17772 -33876 -17708
rect -33812 -17772 -33792 -17708
rect -33896 -17788 -33792 -17772
rect -33896 -17852 -33876 -17788
rect -33812 -17852 -33792 -17788
rect -33896 -17868 -33792 -17852
rect -33896 -17932 -33876 -17868
rect -33812 -17932 -33792 -17868
rect -33896 -17948 -33792 -17932
rect -33896 -18012 -33876 -17948
rect -33812 -18012 -33792 -17948
rect -33896 -18028 -33792 -18012
rect -33896 -18092 -33876 -18028
rect -33812 -18092 -33792 -18028
rect -33896 -18108 -33792 -18092
rect -33896 -18172 -33876 -18108
rect -33812 -18172 -33792 -18108
rect -33896 -18188 -33792 -18172
rect -33896 -18252 -33876 -18188
rect -33812 -18252 -33792 -18188
rect -33896 -18268 -33792 -18252
rect -33896 -18332 -33876 -18268
rect -33812 -18332 -33792 -18268
rect -33896 -18348 -33792 -18332
rect -33896 -18412 -33876 -18348
rect -33812 -18412 -33792 -18348
rect -33896 -18428 -33792 -18412
rect -33896 -18492 -33876 -18428
rect -33812 -18492 -33792 -18428
rect -33896 -18508 -33792 -18492
rect -33896 -18572 -33876 -18508
rect -33812 -18572 -33792 -18508
rect -33896 -18588 -33792 -18572
rect -33896 -18652 -33876 -18588
rect -33812 -18652 -33792 -18588
rect -33896 -18668 -33792 -18652
rect -33896 -18732 -33876 -18668
rect -33812 -18732 -33792 -18668
rect -33896 -18748 -33792 -18732
rect -33896 -18812 -33876 -18748
rect -33812 -18812 -33792 -18748
rect -33896 -18828 -33792 -18812
rect -33896 -18892 -33876 -18828
rect -33812 -18892 -33792 -18828
rect -33896 -18908 -33792 -18892
rect -33896 -18972 -33876 -18908
rect -33812 -18972 -33792 -18908
rect -33896 -18988 -33792 -18972
rect -33896 -19052 -33876 -18988
rect -33812 -19052 -33792 -18988
rect -33896 -19068 -33792 -19052
rect -33896 -19132 -33876 -19068
rect -33812 -19132 -33792 -19068
rect -33896 -19148 -33792 -19132
rect -33896 -19212 -33876 -19148
rect -33812 -19212 -33792 -19148
rect -33896 -19228 -33792 -19212
rect -33896 -19292 -33876 -19228
rect -33812 -19292 -33792 -19228
rect -33896 -19308 -33792 -19292
rect -33896 -19372 -33876 -19308
rect -33812 -19372 -33792 -19308
rect -33896 -19388 -33792 -19372
rect -33896 -19452 -33876 -19388
rect -33812 -19452 -33792 -19388
rect -33896 -19468 -33792 -19452
rect -33896 -19532 -33876 -19468
rect -33812 -19532 -33792 -19468
rect -33896 -19548 -33792 -19532
rect -33896 -19612 -33876 -19548
rect -33812 -19612 -33792 -19548
rect -33896 -19628 -33792 -19612
rect -33896 -19692 -33876 -19628
rect -33812 -19692 -33792 -19628
rect -33896 -19708 -33792 -19692
rect -33896 -19772 -33876 -19708
rect -33812 -19772 -33792 -19708
rect -33896 -19788 -33792 -19772
rect -33896 -19852 -33876 -19788
rect -33812 -19852 -33792 -19788
rect -33896 -19868 -33792 -19852
rect -33896 -19932 -33876 -19868
rect -33812 -19932 -33792 -19868
rect -33896 -19948 -33792 -19932
rect -33896 -20012 -33876 -19948
rect -33812 -20012 -33792 -19948
rect -33896 -20028 -33792 -20012
rect -33896 -20092 -33876 -20028
rect -33812 -20092 -33792 -20028
rect -33896 -20108 -33792 -20092
rect -33896 -20172 -33876 -20108
rect -33812 -20172 -33792 -20108
rect -33896 -20188 -33792 -20172
rect -33896 -20252 -33876 -20188
rect -33812 -20252 -33792 -20188
rect -33896 -20268 -33792 -20252
rect -33896 -20332 -33876 -20268
rect -33812 -20332 -33792 -20268
rect -33896 -20348 -33792 -20332
rect -33896 -20412 -33876 -20348
rect -33812 -20412 -33792 -20348
rect -33896 -20428 -33792 -20412
rect -33896 -20492 -33876 -20428
rect -33812 -20492 -33792 -20428
rect -33896 -20508 -33792 -20492
rect -33896 -20572 -33876 -20508
rect -33812 -20572 -33792 -20508
rect -33896 -20588 -33792 -20572
rect -33896 -20652 -33876 -20588
rect -33812 -20652 -33792 -20588
rect -33896 -20668 -33792 -20652
rect -33896 -20732 -33876 -20668
rect -33812 -20732 -33792 -20668
rect -33896 -20748 -33792 -20732
rect -33896 -20812 -33876 -20748
rect -33812 -20812 -33792 -20748
rect -33896 -20828 -33792 -20812
rect -33896 -20892 -33876 -20828
rect -33812 -20892 -33792 -20828
rect -33896 -20908 -33792 -20892
rect -33896 -20972 -33876 -20908
rect -33812 -20972 -33792 -20908
rect -33896 -20988 -33792 -20972
rect -33896 -21052 -33876 -20988
rect -33812 -21052 -33792 -20988
rect -33896 -21068 -33792 -21052
rect -36676 -21479 -36572 -21081
rect -33896 -21132 -33876 -21068
rect -33812 -21132 -33792 -21068
rect -33473 -16188 -28551 -16159
rect -33473 -21052 -33444 -16188
rect -28580 -21052 -28551 -16188
rect -33473 -21081 -28551 -21052
rect -28284 -16172 -28264 -16108
rect -28200 -16172 -28180 -16108
rect -25452 -16159 -25348 -15761
rect -22672 -15812 -22652 -15748
rect -22588 -15812 -22568 -15748
rect -22249 -10868 -17327 -10839
rect -22249 -15732 -22220 -10868
rect -17356 -15732 -17327 -10868
rect -22249 -15761 -17327 -15732
rect -17060 -10852 -17040 -10788
rect -16976 -10852 -16956 -10788
rect -14228 -10839 -14124 -10441
rect -11448 -10492 -11428 -10428
rect -11364 -10492 -11344 -10428
rect -11025 -5548 -6103 -5519
rect -11025 -10412 -10996 -5548
rect -6132 -10412 -6103 -5548
rect -11025 -10441 -6103 -10412
rect -5836 -5532 -5816 -5468
rect -5752 -5532 -5732 -5468
rect -3004 -5519 -2900 -5121
rect -224 -5172 -204 -5108
rect -140 -5172 -120 -5108
rect 199 -228 5121 -199
rect 199 -5092 228 -228
rect 5092 -5092 5121 -228
rect 199 -5121 5121 -5092
rect 5388 -212 5408 -148
rect 5472 -212 5492 -148
rect 8220 -199 8324 199
rect 11000 148 11020 212
rect 11084 148 11104 212
rect 11423 5092 16345 5121
rect 11423 228 11452 5092
rect 16316 228 16345 5092
rect 11423 199 16345 228
rect 16612 5108 16632 5172
rect 16696 5108 16716 5172
rect 19444 5121 19548 5519
rect 22224 5468 22244 5532
rect 22308 5468 22328 5532
rect 22647 10412 27569 10441
rect 22647 5548 22676 10412
rect 27540 5548 27569 10412
rect 22647 5519 27569 5548
rect 27836 10428 27856 10492
rect 27920 10428 27940 10492
rect 30668 10441 30772 10839
rect 33448 10788 33468 10852
rect 33532 10788 33552 10852
rect 33871 15732 38793 15761
rect 33871 10868 33900 15732
rect 38764 10868 38793 15732
rect 33871 10839 38793 10868
rect 39060 15748 39080 15812
rect 39144 15748 39164 15812
rect 39060 15732 39164 15748
rect 39060 15668 39080 15732
rect 39144 15668 39164 15732
rect 39060 15652 39164 15668
rect 39060 15588 39080 15652
rect 39144 15588 39164 15652
rect 39060 15572 39164 15588
rect 39060 15508 39080 15572
rect 39144 15508 39164 15572
rect 39060 15492 39164 15508
rect 39060 15428 39080 15492
rect 39144 15428 39164 15492
rect 39060 15412 39164 15428
rect 39060 15348 39080 15412
rect 39144 15348 39164 15412
rect 39060 15332 39164 15348
rect 39060 15268 39080 15332
rect 39144 15268 39164 15332
rect 39060 15252 39164 15268
rect 39060 15188 39080 15252
rect 39144 15188 39164 15252
rect 39060 15172 39164 15188
rect 39060 15108 39080 15172
rect 39144 15108 39164 15172
rect 39060 15092 39164 15108
rect 39060 15028 39080 15092
rect 39144 15028 39164 15092
rect 39060 15012 39164 15028
rect 39060 14948 39080 15012
rect 39144 14948 39164 15012
rect 39060 14932 39164 14948
rect 39060 14868 39080 14932
rect 39144 14868 39164 14932
rect 39060 14852 39164 14868
rect 39060 14788 39080 14852
rect 39144 14788 39164 14852
rect 39060 14772 39164 14788
rect 39060 14708 39080 14772
rect 39144 14708 39164 14772
rect 39060 14692 39164 14708
rect 39060 14628 39080 14692
rect 39144 14628 39164 14692
rect 39060 14612 39164 14628
rect 39060 14548 39080 14612
rect 39144 14548 39164 14612
rect 39060 14532 39164 14548
rect 39060 14468 39080 14532
rect 39144 14468 39164 14532
rect 39060 14452 39164 14468
rect 39060 14388 39080 14452
rect 39144 14388 39164 14452
rect 39060 14372 39164 14388
rect 39060 14308 39080 14372
rect 39144 14308 39164 14372
rect 39060 14292 39164 14308
rect 39060 14228 39080 14292
rect 39144 14228 39164 14292
rect 39060 14212 39164 14228
rect 39060 14148 39080 14212
rect 39144 14148 39164 14212
rect 39060 14132 39164 14148
rect 39060 14068 39080 14132
rect 39144 14068 39164 14132
rect 39060 14052 39164 14068
rect 39060 13988 39080 14052
rect 39144 13988 39164 14052
rect 39060 13972 39164 13988
rect 39060 13908 39080 13972
rect 39144 13908 39164 13972
rect 39060 13892 39164 13908
rect 39060 13828 39080 13892
rect 39144 13828 39164 13892
rect 39060 13812 39164 13828
rect 39060 13748 39080 13812
rect 39144 13748 39164 13812
rect 39060 13732 39164 13748
rect 39060 13668 39080 13732
rect 39144 13668 39164 13732
rect 39060 13652 39164 13668
rect 39060 13588 39080 13652
rect 39144 13588 39164 13652
rect 39060 13572 39164 13588
rect 39060 13508 39080 13572
rect 39144 13508 39164 13572
rect 39060 13492 39164 13508
rect 39060 13428 39080 13492
rect 39144 13428 39164 13492
rect 39060 13412 39164 13428
rect 39060 13348 39080 13412
rect 39144 13348 39164 13412
rect 39060 13332 39164 13348
rect 39060 13268 39080 13332
rect 39144 13268 39164 13332
rect 39060 13252 39164 13268
rect 39060 13188 39080 13252
rect 39144 13188 39164 13252
rect 39060 13172 39164 13188
rect 39060 13108 39080 13172
rect 39144 13108 39164 13172
rect 39060 13092 39164 13108
rect 39060 13028 39080 13092
rect 39144 13028 39164 13092
rect 39060 13012 39164 13028
rect 39060 12948 39080 13012
rect 39144 12948 39164 13012
rect 39060 12932 39164 12948
rect 39060 12868 39080 12932
rect 39144 12868 39164 12932
rect 39060 12852 39164 12868
rect 39060 12788 39080 12852
rect 39144 12788 39164 12852
rect 39060 12772 39164 12788
rect 39060 12708 39080 12772
rect 39144 12708 39164 12772
rect 39060 12692 39164 12708
rect 39060 12628 39080 12692
rect 39144 12628 39164 12692
rect 39060 12612 39164 12628
rect 39060 12548 39080 12612
rect 39144 12548 39164 12612
rect 39060 12532 39164 12548
rect 39060 12468 39080 12532
rect 39144 12468 39164 12532
rect 39060 12452 39164 12468
rect 39060 12388 39080 12452
rect 39144 12388 39164 12452
rect 39060 12372 39164 12388
rect 39060 12308 39080 12372
rect 39144 12308 39164 12372
rect 39060 12292 39164 12308
rect 39060 12228 39080 12292
rect 39144 12228 39164 12292
rect 39060 12212 39164 12228
rect 39060 12148 39080 12212
rect 39144 12148 39164 12212
rect 39060 12132 39164 12148
rect 39060 12068 39080 12132
rect 39144 12068 39164 12132
rect 39060 12052 39164 12068
rect 39060 11988 39080 12052
rect 39144 11988 39164 12052
rect 39060 11972 39164 11988
rect 39060 11908 39080 11972
rect 39144 11908 39164 11972
rect 39060 11892 39164 11908
rect 39060 11828 39080 11892
rect 39144 11828 39164 11892
rect 39060 11812 39164 11828
rect 39060 11748 39080 11812
rect 39144 11748 39164 11812
rect 39060 11732 39164 11748
rect 39060 11668 39080 11732
rect 39144 11668 39164 11732
rect 39060 11652 39164 11668
rect 39060 11588 39080 11652
rect 39144 11588 39164 11652
rect 39060 11572 39164 11588
rect 39060 11508 39080 11572
rect 39144 11508 39164 11572
rect 39060 11492 39164 11508
rect 39060 11428 39080 11492
rect 39144 11428 39164 11492
rect 39060 11412 39164 11428
rect 39060 11348 39080 11412
rect 39144 11348 39164 11412
rect 39060 11332 39164 11348
rect 39060 11268 39080 11332
rect 39144 11268 39164 11332
rect 39060 11252 39164 11268
rect 39060 11188 39080 11252
rect 39144 11188 39164 11252
rect 39060 11172 39164 11188
rect 39060 11108 39080 11172
rect 39144 11108 39164 11172
rect 39060 11092 39164 11108
rect 39060 11028 39080 11092
rect 39144 11028 39164 11092
rect 39060 11012 39164 11028
rect 39060 10948 39080 11012
rect 39144 10948 39164 11012
rect 39060 10932 39164 10948
rect 39060 10868 39080 10932
rect 39144 10868 39164 10932
rect 39060 10852 39164 10868
rect 33448 10492 33552 10788
rect 27836 10412 27940 10428
rect 27836 10348 27856 10412
rect 27920 10348 27940 10412
rect 27836 10332 27940 10348
rect 27836 10268 27856 10332
rect 27920 10268 27940 10332
rect 27836 10252 27940 10268
rect 27836 10188 27856 10252
rect 27920 10188 27940 10252
rect 27836 10172 27940 10188
rect 27836 10108 27856 10172
rect 27920 10108 27940 10172
rect 27836 10092 27940 10108
rect 27836 10028 27856 10092
rect 27920 10028 27940 10092
rect 27836 10012 27940 10028
rect 27836 9948 27856 10012
rect 27920 9948 27940 10012
rect 27836 9932 27940 9948
rect 27836 9868 27856 9932
rect 27920 9868 27940 9932
rect 27836 9852 27940 9868
rect 27836 9788 27856 9852
rect 27920 9788 27940 9852
rect 27836 9772 27940 9788
rect 27836 9708 27856 9772
rect 27920 9708 27940 9772
rect 27836 9692 27940 9708
rect 27836 9628 27856 9692
rect 27920 9628 27940 9692
rect 27836 9612 27940 9628
rect 27836 9548 27856 9612
rect 27920 9548 27940 9612
rect 27836 9532 27940 9548
rect 27836 9468 27856 9532
rect 27920 9468 27940 9532
rect 27836 9452 27940 9468
rect 27836 9388 27856 9452
rect 27920 9388 27940 9452
rect 27836 9372 27940 9388
rect 27836 9308 27856 9372
rect 27920 9308 27940 9372
rect 27836 9292 27940 9308
rect 27836 9228 27856 9292
rect 27920 9228 27940 9292
rect 27836 9212 27940 9228
rect 27836 9148 27856 9212
rect 27920 9148 27940 9212
rect 27836 9132 27940 9148
rect 27836 9068 27856 9132
rect 27920 9068 27940 9132
rect 27836 9052 27940 9068
rect 27836 8988 27856 9052
rect 27920 8988 27940 9052
rect 27836 8972 27940 8988
rect 27836 8908 27856 8972
rect 27920 8908 27940 8972
rect 27836 8892 27940 8908
rect 27836 8828 27856 8892
rect 27920 8828 27940 8892
rect 27836 8812 27940 8828
rect 27836 8748 27856 8812
rect 27920 8748 27940 8812
rect 27836 8732 27940 8748
rect 27836 8668 27856 8732
rect 27920 8668 27940 8732
rect 27836 8652 27940 8668
rect 27836 8588 27856 8652
rect 27920 8588 27940 8652
rect 27836 8572 27940 8588
rect 27836 8508 27856 8572
rect 27920 8508 27940 8572
rect 27836 8492 27940 8508
rect 27836 8428 27856 8492
rect 27920 8428 27940 8492
rect 27836 8412 27940 8428
rect 27836 8348 27856 8412
rect 27920 8348 27940 8412
rect 27836 8332 27940 8348
rect 27836 8268 27856 8332
rect 27920 8268 27940 8332
rect 27836 8252 27940 8268
rect 27836 8188 27856 8252
rect 27920 8188 27940 8252
rect 27836 8172 27940 8188
rect 27836 8108 27856 8172
rect 27920 8108 27940 8172
rect 27836 8092 27940 8108
rect 27836 8028 27856 8092
rect 27920 8028 27940 8092
rect 27836 8012 27940 8028
rect 27836 7948 27856 8012
rect 27920 7948 27940 8012
rect 27836 7932 27940 7948
rect 27836 7868 27856 7932
rect 27920 7868 27940 7932
rect 27836 7852 27940 7868
rect 27836 7788 27856 7852
rect 27920 7788 27940 7852
rect 27836 7772 27940 7788
rect 27836 7708 27856 7772
rect 27920 7708 27940 7772
rect 27836 7692 27940 7708
rect 27836 7628 27856 7692
rect 27920 7628 27940 7692
rect 27836 7612 27940 7628
rect 27836 7548 27856 7612
rect 27920 7548 27940 7612
rect 27836 7532 27940 7548
rect 27836 7468 27856 7532
rect 27920 7468 27940 7532
rect 27836 7452 27940 7468
rect 27836 7388 27856 7452
rect 27920 7388 27940 7452
rect 27836 7372 27940 7388
rect 27836 7308 27856 7372
rect 27920 7308 27940 7372
rect 27836 7292 27940 7308
rect 27836 7228 27856 7292
rect 27920 7228 27940 7292
rect 27836 7212 27940 7228
rect 27836 7148 27856 7212
rect 27920 7148 27940 7212
rect 27836 7132 27940 7148
rect 27836 7068 27856 7132
rect 27920 7068 27940 7132
rect 27836 7052 27940 7068
rect 27836 6988 27856 7052
rect 27920 6988 27940 7052
rect 27836 6972 27940 6988
rect 27836 6908 27856 6972
rect 27920 6908 27940 6972
rect 27836 6892 27940 6908
rect 27836 6828 27856 6892
rect 27920 6828 27940 6892
rect 27836 6812 27940 6828
rect 27836 6748 27856 6812
rect 27920 6748 27940 6812
rect 27836 6732 27940 6748
rect 27836 6668 27856 6732
rect 27920 6668 27940 6732
rect 27836 6652 27940 6668
rect 27836 6588 27856 6652
rect 27920 6588 27940 6652
rect 27836 6572 27940 6588
rect 27836 6508 27856 6572
rect 27920 6508 27940 6572
rect 27836 6492 27940 6508
rect 27836 6428 27856 6492
rect 27920 6428 27940 6492
rect 27836 6412 27940 6428
rect 27836 6348 27856 6412
rect 27920 6348 27940 6412
rect 27836 6332 27940 6348
rect 27836 6268 27856 6332
rect 27920 6268 27940 6332
rect 27836 6252 27940 6268
rect 27836 6188 27856 6252
rect 27920 6188 27940 6252
rect 27836 6172 27940 6188
rect 27836 6108 27856 6172
rect 27920 6108 27940 6172
rect 27836 6092 27940 6108
rect 27836 6028 27856 6092
rect 27920 6028 27940 6092
rect 27836 6012 27940 6028
rect 27836 5948 27856 6012
rect 27920 5948 27940 6012
rect 27836 5932 27940 5948
rect 27836 5868 27856 5932
rect 27920 5868 27940 5932
rect 27836 5852 27940 5868
rect 27836 5788 27856 5852
rect 27920 5788 27940 5852
rect 27836 5772 27940 5788
rect 27836 5708 27856 5772
rect 27920 5708 27940 5772
rect 27836 5692 27940 5708
rect 27836 5628 27856 5692
rect 27920 5628 27940 5692
rect 27836 5612 27940 5628
rect 27836 5548 27856 5612
rect 27920 5548 27940 5612
rect 27836 5532 27940 5548
rect 22224 5172 22328 5468
rect 16612 5092 16716 5108
rect 16612 5028 16632 5092
rect 16696 5028 16716 5092
rect 16612 5012 16716 5028
rect 16612 4948 16632 5012
rect 16696 4948 16716 5012
rect 16612 4932 16716 4948
rect 16612 4868 16632 4932
rect 16696 4868 16716 4932
rect 16612 4852 16716 4868
rect 16612 4788 16632 4852
rect 16696 4788 16716 4852
rect 16612 4772 16716 4788
rect 16612 4708 16632 4772
rect 16696 4708 16716 4772
rect 16612 4692 16716 4708
rect 16612 4628 16632 4692
rect 16696 4628 16716 4692
rect 16612 4612 16716 4628
rect 16612 4548 16632 4612
rect 16696 4548 16716 4612
rect 16612 4532 16716 4548
rect 16612 4468 16632 4532
rect 16696 4468 16716 4532
rect 16612 4452 16716 4468
rect 16612 4388 16632 4452
rect 16696 4388 16716 4452
rect 16612 4372 16716 4388
rect 16612 4308 16632 4372
rect 16696 4308 16716 4372
rect 16612 4292 16716 4308
rect 16612 4228 16632 4292
rect 16696 4228 16716 4292
rect 16612 4212 16716 4228
rect 16612 4148 16632 4212
rect 16696 4148 16716 4212
rect 16612 4132 16716 4148
rect 16612 4068 16632 4132
rect 16696 4068 16716 4132
rect 16612 4052 16716 4068
rect 16612 3988 16632 4052
rect 16696 3988 16716 4052
rect 16612 3972 16716 3988
rect 16612 3908 16632 3972
rect 16696 3908 16716 3972
rect 16612 3892 16716 3908
rect 16612 3828 16632 3892
rect 16696 3828 16716 3892
rect 16612 3812 16716 3828
rect 16612 3748 16632 3812
rect 16696 3748 16716 3812
rect 16612 3732 16716 3748
rect 16612 3668 16632 3732
rect 16696 3668 16716 3732
rect 16612 3652 16716 3668
rect 16612 3588 16632 3652
rect 16696 3588 16716 3652
rect 16612 3572 16716 3588
rect 16612 3508 16632 3572
rect 16696 3508 16716 3572
rect 16612 3492 16716 3508
rect 16612 3428 16632 3492
rect 16696 3428 16716 3492
rect 16612 3412 16716 3428
rect 16612 3348 16632 3412
rect 16696 3348 16716 3412
rect 16612 3332 16716 3348
rect 16612 3268 16632 3332
rect 16696 3268 16716 3332
rect 16612 3252 16716 3268
rect 16612 3188 16632 3252
rect 16696 3188 16716 3252
rect 16612 3172 16716 3188
rect 16612 3108 16632 3172
rect 16696 3108 16716 3172
rect 16612 3092 16716 3108
rect 16612 3028 16632 3092
rect 16696 3028 16716 3092
rect 16612 3012 16716 3028
rect 16612 2948 16632 3012
rect 16696 2948 16716 3012
rect 16612 2932 16716 2948
rect 16612 2868 16632 2932
rect 16696 2868 16716 2932
rect 16612 2852 16716 2868
rect 16612 2788 16632 2852
rect 16696 2788 16716 2852
rect 16612 2772 16716 2788
rect 16612 2708 16632 2772
rect 16696 2708 16716 2772
rect 16612 2692 16716 2708
rect 16612 2628 16632 2692
rect 16696 2628 16716 2692
rect 16612 2612 16716 2628
rect 16612 2548 16632 2612
rect 16696 2548 16716 2612
rect 16612 2532 16716 2548
rect 16612 2468 16632 2532
rect 16696 2468 16716 2532
rect 16612 2452 16716 2468
rect 16612 2388 16632 2452
rect 16696 2388 16716 2452
rect 16612 2372 16716 2388
rect 16612 2308 16632 2372
rect 16696 2308 16716 2372
rect 16612 2292 16716 2308
rect 16612 2228 16632 2292
rect 16696 2228 16716 2292
rect 16612 2212 16716 2228
rect 16612 2148 16632 2212
rect 16696 2148 16716 2212
rect 16612 2132 16716 2148
rect 16612 2068 16632 2132
rect 16696 2068 16716 2132
rect 16612 2052 16716 2068
rect 16612 1988 16632 2052
rect 16696 1988 16716 2052
rect 16612 1972 16716 1988
rect 16612 1908 16632 1972
rect 16696 1908 16716 1972
rect 16612 1892 16716 1908
rect 16612 1828 16632 1892
rect 16696 1828 16716 1892
rect 16612 1812 16716 1828
rect 16612 1748 16632 1812
rect 16696 1748 16716 1812
rect 16612 1732 16716 1748
rect 16612 1668 16632 1732
rect 16696 1668 16716 1732
rect 16612 1652 16716 1668
rect 16612 1588 16632 1652
rect 16696 1588 16716 1652
rect 16612 1572 16716 1588
rect 16612 1508 16632 1572
rect 16696 1508 16716 1572
rect 16612 1492 16716 1508
rect 16612 1428 16632 1492
rect 16696 1428 16716 1492
rect 16612 1412 16716 1428
rect 16612 1348 16632 1412
rect 16696 1348 16716 1412
rect 16612 1332 16716 1348
rect 16612 1268 16632 1332
rect 16696 1268 16716 1332
rect 16612 1252 16716 1268
rect 16612 1188 16632 1252
rect 16696 1188 16716 1252
rect 16612 1172 16716 1188
rect 16612 1108 16632 1172
rect 16696 1108 16716 1172
rect 16612 1092 16716 1108
rect 16612 1028 16632 1092
rect 16696 1028 16716 1092
rect 16612 1012 16716 1028
rect 16612 948 16632 1012
rect 16696 948 16716 1012
rect 16612 932 16716 948
rect 16612 868 16632 932
rect 16696 868 16716 932
rect 16612 852 16716 868
rect 16612 788 16632 852
rect 16696 788 16716 852
rect 16612 772 16716 788
rect 16612 708 16632 772
rect 16696 708 16716 772
rect 16612 692 16716 708
rect 16612 628 16632 692
rect 16696 628 16716 692
rect 16612 612 16716 628
rect 16612 548 16632 612
rect 16696 548 16716 612
rect 16612 532 16716 548
rect 16612 468 16632 532
rect 16696 468 16716 532
rect 16612 452 16716 468
rect 16612 388 16632 452
rect 16696 388 16716 452
rect 16612 372 16716 388
rect 16612 308 16632 372
rect 16696 308 16716 372
rect 16612 292 16716 308
rect 16612 228 16632 292
rect 16696 228 16716 292
rect 16612 212 16716 228
rect 11000 -148 11104 148
rect 5388 -228 5492 -212
rect 5388 -292 5408 -228
rect 5472 -292 5492 -228
rect 5388 -308 5492 -292
rect 5388 -372 5408 -308
rect 5472 -372 5492 -308
rect 5388 -388 5492 -372
rect 5388 -452 5408 -388
rect 5472 -452 5492 -388
rect 5388 -468 5492 -452
rect 5388 -532 5408 -468
rect 5472 -532 5492 -468
rect 5388 -548 5492 -532
rect 5388 -612 5408 -548
rect 5472 -612 5492 -548
rect 5388 -628 5492 -612
rect 5388 -692 5408 -628
rect 5472 -692 5492 -628
rect 5388 -708 5492 -692
rect 5388 -772 5408 -708
rect 5472 -772 5492 -708
rect 5388 -788 5492 -772
rect 5388 -852 5408 -788
rect 5472 -852 5492 -788
rect 5388 -868 5492 -852
rect 5388 -932 5408 -868
rect 5472 -932 5492 -868
rect 5388 -948 5492 -932
rect 5388 -1012 5408 -948
rect 5472 -1012 5492 -948
rect 5388 -1028 5492 -1012
rect 5388 -1092 5408 -1028
rect 5472 -1092 5492 -1028
rect 5388 -1108 5492 -1092
rect 5388 -1172 5408 -1108
rect 5472 -1172 5492 -1108
rect 5388 -1188 5492 -1172
rect 5388 -1252 5408 -1188
rect 5472 -1252 5492 -1188
rect 5388 -1268 5492 -1252
rect 5388 -1332 5408 -1268
rect 5472 -1332 5492 -1268
rect 5388 -1348 5492 -1332
rect 5388 -1412 5408 -1348
rect 5472 -1412 5492 -1348
rect 5388 -1428 5492 -1412
rect 5388 -1492 5408 -1428
rect 5472 -1492 5492 -1428
rect 5388 -1508 5492 -1492
rect 5388 -1572 5408 -1508
rect 5472 -1572 5492 -1508
rect 5388 -1588 5492 -1572
rect 5388 -1652 5408 -1588
rect 5472 -1652 5492 -1588
rect 5388 -1668 5492 -1652
rect 5388 -1732 5408 -1668
rect 5472 -1732 5492 -1668
rect 5388 -1748 5492 -1732
rect 5388 -1812 5408 -1748
rect 5472 -1812 5492 -1748
rect 5388 -1828 5492 -1812
rect 5388 -1892 5408 -1828
rect 5472 -1892 5492 -1828
rect 5388 -1908 5492 -1892
rect 5388 -1972 5408 -1908
rect 5472 -1972 5492 -1908
rect 5388 -1988 5492 -1972
rect 5388 -2052 5408 -1988
rect 5472 -2052 5492 -1988
rect 5388 -2068 5492 -2052
rect 5388 -2132 5408 -2068
rect 5472 -2132 5492 -2068
rect 5388 -2148 5492 -2132
rect 5388 -2212 5408 -2148
rect 5472 -2212 5492 -2148
rect 5388 -2228 5492 -2212
rect 5388 -2292 5408 -2228
rect 5472 -2292 5492 -2228
rect 5388 -2308 5492 -2292
rect 5388 -2372 5408 -2308
rect 5472 -2372 5492 -2308
rect 5388 -2388 5492 -2372
rect 5388 -2452 5408 -2388
rect 5472 -2452 5492 -2388
rect 5388 -2468 5492 -2452
rect 5388 -2532 5408 -2468
rect 5472 -2532 5492 -2468
rect 5388 -2548 5492 -2532
rect 5388 -2612 5408 -2548
rect 5472 -2612 5492 -2548
rect 5388 -2628 5492 -2612
rect 5388 -2692 5408 -2628
rect 5472 -2692 5492 -2628
rect 5388 -2708 5492 -2692
rect 5388 -2772 5408 -2708
rect 5472 -2772 5492 -2708
rect 5388 -2788 5492 -2772
rect 5388 -2852 5408 -2788
rect 5472 -2852 5492 -2788
rect 5388 -2868 5492 -2852
rect 5388 -2932 5408 -2868
rect 5472 -2932 5492 -2868
rect 5388 -2948 5492 -2932
rect 5388 -3012 5408 -2948
rect 5472 -3012 5492 -2948
rect 5388 -3028 5492 -3012
rect 5388 -3092 5408 -3028
rect 5472 -3092 5492 -3028
rect 5388 -3108 5492 -3092
rect 5388 -3172 5408 -3108
rect 5472 -3172 5492 -3108
rect 5388 -3188 5492 -3172
rect 5388 -3252 5408 -3188
rect 5472 -3252 5492 -3188
rect 5388 -3268 5492 -3252
rect 5388 -3332 5408 -3268
rect 5472 -3332 5492 -3268
rect 5388 -3348 5492 -3332
rect 5388 -3412 5408 -3348
rect 5472 -3412 5492 -3348
rect 5388 -3428 5492 -3412
rect 5388 -3492 5408 -3428
rect 5472 -3492 5492 -3428
rect 5388 -3508 5492 -3492
rect 5388 -3572 5408 -3508
rect 5472 -3572 5492 -3508
rect 5388 -3588 5492 -3572
rect 5388 -3652 5408 -3588
rect 5472 -3652 5492 -3588
rect 5388 -3668 5492 -3652
rect 5388 -3732 5408 -3668
rect 5472 -3732 5492 -3668
rect 5388 -3748 5492 -3732
rect 5388 -3812 5408 -3748
rect 5472 -3812 5492 -3748
rect 5388 -3828 5492 -3812
rect 5388 -3892 5408 -3828
rect 5472 -3892 5492 -3828
rect 5388 -3908 5492 -3892
rect 5388 -3972 5408 -3908
rect 5472 -3972 5492 -3908
rect 5388 -3988 5492 -3972
rect 5388 -4052 5408 -3988
rect 5472 -4052 5492 -3988
rect 5388 -4068 5492 -4052
rect 5388 -4132 5408 -4068
rect 5472 -4132 5492 -4068
rect 5388 -4148 5492 -4132
rect 5388 -4212 5408 -4148
rect 5472 -4212 5492 -4148
rect 5388 -4228 5492 -4212
rect 5388 -4292 5408 -4228
rect 5472 -4292 5492 -4228
rect 5388 -4308 5492 -4292
rect 5388 -4372 5408 -4308
rect 5472 -4372 5492 -4308
rect 5388 -4388 5492 -4372
rect 5388 -4452 5408 -4388
rect 5472 -4452 5492 -4388
rect 5388 -4468 5492 -4452
rect 5388 -4532 5408 -4468
rect 5472 -4532 5492 -4468
rect 5388 -4548 5492 -4532
rect 5388 -4612 5408 -4548
rect 5472 -4612 5492 -4548
rect 5388 -4628 5492 -4612
rect 5388 -4692 5408 -4628
rect 5472 -4692 5492 -4628
rect 5388 -4708 5492 -4692
rect 5388 -4772 5408 -4708
rect 5472 -4772 5492 -4708
rect 5388 -4788 5492 -4772
rect 5388 -4852 5408 -4788
rect 5472 -4852 5492 -4788
rect 5388 -4868 5492 -4852
rect 5388 -4932 5408 -4868
rect 5472 -4932 5492 -4868
rect 5388 -4948 5492 -4932
rect 5388 -5012 5408 -4948
rect 5472 -5012 5492 -4948
rect 5388 -5028 5492 -5012
rect 5388 -5092 5408 -5028
rect 5472 -5092 5492 -5028
rect 5388 -5108 5492 -5092
rect -224 -5468 -120 -5172
rect -5836 -5548 -5732 -5532
rect -5836 -5612 -5816 -5548
rect -5752 -5612 -5732 -5548
rect -5836 -5628 -5732 -5612
rect -5836 -5692 -5816 -5628
rect -5752 -5692 -5732 -5628
rect -5836 -5708 -5732 -5692
rect -5836 -5772 -5816 -5708
rect -5752 -5772 -5732 -5708
rect -5836 -5788 -5732 -5772
rect -5836 -5852 -5816 -5788
rect -5752 -5852 -5732 -5788
rect -5836 -5868 -5732 -5852
rect -5836 -5932 -5816 -5868
rect -5752 -5932 -5732 -5868
rect -5836 -5948 -5732 -5932
rect -5836 -6012 -5816 -5948
rect -5752 -6012 -5732 -5948
rect -5836 -6028 -5732 -6012
rect -5836 -6092 -5816 -6028
rect -5752 -6092 -5732 -6028
rect -5836 -6108 -5732 -6092
rect -5836 -6172 -5816 -6108
rect -5752 -6172 -5732 -6108
rect -5836 -6188 -5732 -6172
rect -5836 -6252 -5816 -6188
rect -5752 -6252 -5732 -6188
rect -5836 -6268 -5732 -6252
rect -5836 -6332 -5816 -6268
rect -5752 -6332 -5732 -6268
rect -5836 -6348 -5732 -6332
rect -5836 -6412 -5816 -6348
rect -5752 -6412 -5732 -6348
rect -5836 -6428 -5732 -6412
rect -5836 -6492 -5816 -6428
rect -5752 -6492 -5732 -6428
rect -5836 -6508 -5732 -6492
rect -5836 -6572 -5816 -6508
rect -5752 -6572 -5732 -6508
rect -5836 -6588 -5732 -6572
rect -5836 -6652 -5816 -6588
rect -5752 -6652 -5732 -6588
rect -5836 -6668 -5732 -6652
rect -5836 -6732 -5816 -6668
rect -5752 -6732 -5732 -6668
rect -5836 -6748 -5732 -6732
rect -5836 -6812 -5816 -6748
rect -5752 -6812 -5732 -6748
rect -5836 -6828 -5732 -6812
rect -5836 -6892 -5816 -6828
rect -5752 -6892 -5732 -6828
rect -5836 -6908 -5732 -6892
rect -5836 -6972 -5816 -6908
rect -5752 -6972 -5732 -6908
rect -5836 -6988 -5732 -6972
rect -5836 -7052 -5816 -6988
rect -5752 -7052 -5732 -6988
rect -5836 -7068 -5732 -7052
rect -5836 -7132 -5816 -7068
rect -5752 -7132 -5732 -7068
rect -5836 -7148 -5732 -7132
rect -5836 -7212 -5816 -7148
rect -5752 -7212 -5732 -7148
rect -5836 -7228 -5732 -7212
rect -5836 -7292 -5816 -7228
rect -5752 -7292 -5732 -7228
rect -5836 -7308 -5732 -7292
rect -5836 -7372 -5816 -7308
rect -5752 -7372 -5732 -7308
rect -5836 -7388 -5732 -7372
rect -5836 -7452 -5816 -7388
rect -5752 -7452 -5732 -7388
rect -5836 -7468 -5732 -7452
rect -5836 -7532 -5816 -7468
rect -5752 -7532 -5732 -7468
rect -5836 -7548 -5732 -7532
rect -5836 -7612 -5816 -7548
rect -5752 -7612 -5732 -7548
rect -5836 -7628 -5732 -7612
rect -5836 -7692 -5816 -7628
rect -5752 -7692 -5732 -7628
rect -5836 -7708 -5732 -7692
rect -5836 -7772 -5816 -7708
rect -5752 -7772 -5732 -7708
rect -5836 -7788 -5732 -7772
rect -5836 -7852 -5816 -7788
rect -5752 -7852 -5732 -7788
rect -5836 -7868 -5732 -7852
rect -5836 -7932 -5816 -7868
rect -5752 -7932 -5732 -7868
rect -5836 -7948 -5732 -7932
rect -5836 -8012 -5816 -7948
rect -5752 -8012 -5732 -7948
rect -5836 -8028 -5732 -8012
rect -5836 -8092 -5816 -8028
rect -5752 -8092 -5732 -8028
rect -5836 -8108 -5732 -8092
rect -5836 -8172 -5816 -8108
rect -5752 -8172 -5732 -8108
rect -5836 -8188 -5732 -8172
rect -5836 -8252 -5816 -8188
rect -5752 -8252 -5732 -8188
rect -5836 -8268 -5732 -8252
rect -5836 -8332 -5816 -8268
rect -5752 -8332 -5732 -8268
rect -5836 -8348 -5732 -8332
rect -5836 -8412 -5816 -8348
rect -5752 -8412 -5732 -8348
rect -5836 -8428 -5732 -8412
rect -5836 -8492 -5816 -8428
rect -5752 -8492 -5732 -8428
rect -5836 -8508 -5732 -8492
rect -5836 -8572 -5816 -8508
rect -5752 -8572 -5732 -8508
rect -5836 -8588 -5732 -8572
rect -5836 -8652 -5816 -8588
rect -5752 -8652 -5732 -8588
rect -5836 -8668 -5732 -8652
rect -5836 -8732 -5816 -8668
rect -5752 -8732 -5732 -8668
rect -5836 -8748 -5732 -8732
rect -5836 -8812 -5816 -8748
rect -5752 -8812 -5732 -8748
rect -5836 -8828 -5732 -8812
rect -5836 -8892 -5816 -8828
rect -5752 -8892 -5732 -8828
rect -5836 -8908 -5732 -8892
rect -5836 -8972 -5816 -8908
rect -5752 -8972 -5732 -8908
rect -5836 -8988 -5732 -8972
rect -5836 -9052 -5816 -8988
rect -5752 -9052 -5732 -8988
rect -5836 -9068 -5732 -9052
rect -5836 -9132 -5816 -9068
rect -5752 -9132 -5732 -9068
rect -5836 -9148 -5732 -9132
rect -5836 -9212 -5816 -9148
rect -5752 -9212 -5732 -9148
rect -5836 -9228 -5732 -9212
rect -5836 -9292 -5816 -9228
rect -5752 -9292 -5732 -9228
rect -5836 -9308 -5732 -9292
rect -5836 -9372 -5816 -9308
rect -5752 -9372 -5732 -9308
rect -5836 -9388 -5732 -9372
rect -5836 -9452 -5816 -9388
rect -5752 -9452 -5732 -9388
rect -5836 -9468 -5732 -9452
rect -5836 -9532 -5816 -9468
rect -5752 -9532 -5732 -9468
rect -5836 -9548 -5732 -9532
rect -5836 -9612 -5816 -9548
rect -5752 -9612 -5732 -9548
rect -5836 -9628 -5732 -9612
rect -5836 -9692 -5816 -9628
rect -5752 -9692 -5732 -9628
rect -5836 -9708 -5732 -9692
rect -5836 -9772 -5816 -9708
rect -5752 -9772 -5732 -9708
rect -5836 -9788 -5732 -9772
rect -5836 -9852 -5816 -9788
rect -5752 -9852 -5732 -9788
rect -5836 -9868 -5732 -9852
rect -5836 -9932 -5816 -9868
rect -5752 -9932 -5732 -9868
rect -5836 -9948 -5732 -9932
rect -5836 -10012 -5816 -9948
rect -5752 -10012 -5732 -9948
rect -5836 -10028 -5732 -10012
rect -5836 -10092 -5816 -10028
rect -5752 -10092 -5732 -10028
rect -5836 -10108 -5732 -10092
rect -5836 -10172 -5816 -10108
rect -5752 -10172 -5732 -10108
rect -5836 -10188 -5732 -10172
rect -5836 -10252 -5816 -10188
rect -5752 -10252 -5732 -10188
rect -5836 -10268 -5732 -10252
rect -5836 -10332 -5816 -10268
rect -5752 -10332 -5732 -10268
rect -5836 -10348 -5732 -10332
rect -5836 -10412 -5816 -10348
rect -5752 -10412 -5732 -10348
rect -5836 -10428 -5732 -10412
rect -11448 -10788 -11344 -10492
rect -17060 -10868 -16956 -10852
rect -17060 -10932 -17040 -10868
rect -16976 -10932 -16956 -10868
rect -17060 -10948 -16956 -10932
rect -17060 -11012 -17040 -10948
rect -16976 -11012 -16956 -10948
rect -17060 -11028 -16956 -11012
rect -17060 -11092 -17040 -11028
rect -16976 -11092 -16956 -11028
rect -17060 -11108 -16956 -11092
rect -17060 -11172 -17040 -11108
rect -16976 -11172 -16956 -11108
rect -17060 -11188 -16956 -11172
rect -17060 -11252 -17040 -11188
rect -16976 -11252 -16956 -11188
rect -17060 -11268 -16956 -11252
rect -17060 -11332 -17040 -11268
rect -16976 -11332 -16956 -11268
rect -17060 -11348 -16956 -11332
rect -17060 -11412 -17040 -11348
rect -16976 -11412 -16956 -11348
rect -17060 -11428 -16956 -11412
rect -17060 -11492 -17040 -11428
rect -16976 -11492 -16956 -11428
rect -17060 -11508 -16956 -11492
rect -17060 -11572 -17040 -11508
rect -16976 -11572 -16956 -11508
rect -17060 -11588 -16956 -11572
rect -17060 -11652 -17040 -11588
rect -16976 -11652 -16956 -11588
rect -17060 -11668 -16956 -11652
rect -17060 -11732 -17040 -11668
rect -16976 -11732 -16956 -11668
rect -17060 -11748 -16956 -11732
rect -17060 -11812 -17040 -11748
rect -16976 -11812 -16956 -11748
rect -17060 -11828 -16956 -11812
rect -17060 -11892 -17040 -11828
rect -16976 -11892 -16956 -11828
rect -17060 -11908 -16956 -11892
rect -17060 -11972 -17040 -11908
rect -16976 -11972 -16956 -11908
rect -17060 -11988 -16956 -11972
rect -17060 -12052 -17040 -11988
rect -16976 -12052 -16956 -11988
rect -17060 -12068 -16956 -12052
rect -17060 -12132 -17040 -12068
rect -16976 -12132 -16956 -12068
rect -17060 -12148 -16956 -12132
rect -17060 -12212 -17040 -12148
rect -16976 -12212 -16956 -12148
rect -17060 -12228 -16956 -12212
rect -17060 -12292 -17040 -12228
rect -16976 -12292 -16956 -12228
rect -17060 -12308 -16956 -12292
rect -17060 -12372 -17040 -12308
rect -16976 -12372 -16956 -12308
rect -17060 -12388 -16956 -12372
rect -17060 -12452 -17040 -12388
rect -16976 -12452 -16956 -12388
rect -17060 -12468 -16956 -12452
rect -17060 -12532 -17040 -12468
rect -16976 -12532 -16956 -12468
rect -17060 -12548 -16956 -12532
rect -17060 -12612 -17040 -12548
rect -16976 -12612 -16956 -12548
rect -17060 -12628 -16956 -12612
rect -17060 -12692 -17040 -12628
rect -16976 -12692 -16956 -12628
rect -17060 -12708 -16956 -12692
rect -17060 -12772 -17040 -12708
rect -16976 -12772 -16956 -12708
rect -17060 -12788 -16956 -12772
rect -17060 -12852 -17040 -12788
rect -16976 -12852 -16956 -12788
rect -17060 -12868 -16956 -12852
rect -17060 -12932 -17040 -12868
rect -16976 -12932 -16956 -12868
rect -17060 -12948 -16956 -12932
rect -17060 -13012 -17040 -12948
rect -16976 -13012 -16956 -12948
rect -17060 -13028 -16956 -13012
rect -17060 -13092 -17040 -13028
rect -16976 -13092 -16956 -13028
rect -17060 -13108 -16956 -13092
rect -17060 -13172 -17040 -13108
rect -16976 -13172 -16956 -13108
rect -17060 -13188 -16956 -13172
rect -17060 -13252 -17040 -13188
rect -16976 -13252 -16956 -13188
rect -17060 -13268 -16956 -13252
rect -17060 -13332 -17040 -13268
rect -16976 -13332 -16956 -13268
rect -17060 -13348 -16956 -13332
rect -17060 -13412 -17040 -13348
rect -16976 -13412 -16956 -13348
rect -17060 -13428 -16956 -13412
rect -17060 -13492 -17040 -13428
rect -16976 -13492 -16956 -13428
rect -17060 -13508 -16956 -13492
rect -17060 -13572 -17040 -13508
rect -16976 -13572 -16956 -13508
rect -17060 -13588 -16956 -13572
rect -17060 -13652 -17040 -13588
rect -16976 -13652 -16956 -13588
rect -17060 -13668 -16956 -13652
rect -17060 -13732 -17040 -13668
rect -16976 -13732 -16956 -13668
rect -17060 -13748 -16956 -13732
rect -17060 -13812 -17040 -13748
rect -16976 -13812 -16956 -13748
rect -17060 -13828 -16956 -13812
rect -17060 -13892 -17040 -13828
rect -16976 -13892 -16956 -13828
rect -17060 -13908 -16956 -13892
rect -17060 -13972 -17040 -13908
rect -16976 -13972 -16956 -13908
rect -17060 -13988 -16956 -13972
rect -17060 -14052 -17040 -13988
rect -16976 -14052 -16956 -13988
rect -17060 -14068 -16956 -14052
rect -17060 -14132 -17040 -14068
rect -16976 -14132 -16956 -14068
rect -17060 -14148 -16956 -14132
rect -17060 -14212 -17040 -14148
rect -16976 -14212 -16956 -14148
rect -17060 -14228 -16956 -14212
rect -17060 -14292 -17040 -14228
rect -16976 -14292 -16956 -14228
rect -17060 -14308 -16956 -14292
rect -17060 -14372 -17040 -14308
rect -16976 -14372 -16956 -14308
rect -17060 -14388 -16956 -14372
rect -17060 -14452 -17040 -14388
rect -16976 -14452 -16956 -14388
rect -17060 -14468 -16956 -14452
rect -17060 -14532 -17040 -14468
rect -16976 -14532 -16956 -14468
rect -17060 -14548 -16956 -14532
rect -17060 -14612 -17040 -14548
rect -16976 -14612 -16956 -14548
rect -17060 -14628 -16956 -14612
rect -17060 -14692 -17040 -14628
rect -16976 -14692 -16956 -14628
rect -17060 -14708 -16956 -14692
rect -17060 -14772 -17040 -14708
rect -16976 -14772 -16956 -14708
rect -17060 -14788 -16956 -14772
rect -17060 -14852 -17040 -14788
rect -16976 -14852 -16956 -14788
rect -17060 -14868 -16956 -14852
rect -17060 -14932 -17040 -14868
rect -16976 -14932 -16956 -14868
rect -17060 -14948 -16956 -14932
rect -17060 -15012 -17040 -14948
rect -16976 -15012 -16956 -14948
rect -17060 -15028 -16956 -15012
rect -17060 -15092 -17040 -15028
rect -16976 -15092 -16956 -15028
rect -17060 -15108 -16956 -15092
rect -17060 -15172 -17040 -15108
rect -16976 -15172 -16956 -15108
rect -17060 -15188 -16956 -15172
rect -17060 -15252 -17040 -15188
rect -16976 -15252 -16956 -15188
rect -17060 -15268 -16956 -15252
rect -17060 -15332 -17040 -15268
rect -16976 -15332 -16956 -15268
rect -17060 -15348 -16956 -15332
rect -17060 -15412 -17040 -15348
rect -16976 -15412 -16956 -15348
rect -17060 -15428 -16956 -15412
rect -17060 -15492 -17040 -15428
rect -16976 -15492 -16956 -15428
rect -17060 -15508 -16956 -15492
rect -17060 -15572 -17040 -15508
rect -16976 -15572 -16956 -15508
rect -17060 -15588 -16956 -15572
rect -17060 -15652 -17040 -15588
rect -16976 -15652 -16956 -15588
rect -17060 -15668 -16956 -15652
rect -17060 -15732 -17040 -15668
rect -16976 -15732 -16956 -15668
rect -17060 -15748 -16956 -15732
rect -22672 -16108 -22568 -15812
rect -28284 -16188 -28180 -16172
rect -28284 -16252 -28264 -16188
rect -28200 -16252 -28180 -16188
rect -28284 -16268 -28180 -16252
rect -28284 -16332 -28264 -16268
rect -28200 -16332 -28180 -16268
rect -28284 -16348 -28180 -16332
rect -28284 -16412 -28264 -16348
rect -28200 -16412 -28180 -16348
rect -28284 -16428 -28180 -16412
rect -28284 -16492 -28264 -16428
rect -28200 -16492 -28180 -16428
rect -28284 -16508 -28180 -16492
rect -28284 -16572 -28264 -16508
rect -28200 -16572 -28180 -16508
rect -28284 -16588 -28180 -16572
rect -28284 -16652 -28264 -16588
rect -28200 -16652 -28180 -16588
rect -28284 -16668 -28180 -16652
rect -28284 -16732 -28264 -16668
rect -28200 -16732 -28180 -16668
rect -28284 -16748 -28180 -16732
rect -28284 -16812 -28264 -16748
rect -28200 -16812 -28180 -16748
rect -28284 -16828 -28180 -16812
rect -28284 -16892 -28264 -16828
rect -28200 -16892 -28180 -16828
rect -28284 -16908 -28180 -16892
rect -28284 -16972 -28264 -16908
rect -28200 -16972 -28180 -16908
rect -28284 -16988 -28180 -16972
rect -28284 -17052 -28264 -16988
rect -28200 -17052 -28180 -16988
rect -28284 -17068 -28180 -17052
rect -28284 -17132 -28264 -17068
rect -28200 -17132 -28180 -17068
rect -28284 -17148 -28180 -17132
rect -28284 -17212 -28264 -17148
rect -28200 -17212 -28180 -17148
rect -28284 -17228 -28180 -17212
rect -28284 -17292 -28264 -17228
rect -28200 -17292 -28180 -17228
rect -28284 -17308 -28180 -17292
rect -28284 -17372 -28264 -17308
rect -28200 -17372 -28180 -17308
rect -28284 -17388 -28180 -17372
rect -28284 -17452 -28264 -17388
rect -28200 -17452 -28180 -17388
rect -28284 -17468 -28180 -17452
rect -28284 -17532 -28264 -17468
rect -28200 -17532 -28180 -17468
rect -28284 -17548 -28180 -17532
rect -28284 -17612 -28264 -17548
rect -28200 -17612 -28180 -17548
rect -28284 -17628 -28180 -17612
rect -28284 -17692 -28264 -17628
rect -28200 -17692 -28180 -17628
rect -28284 -17708 -28180 -17692
rect -28284 -17772 -28264 -17708
rect -28200 -17772 -28180 -17708
rect -28284 -17788 -28180 -17772
rect -28284 -17852 -28264 -17788
rect -28200 -17852 -28180 -17788
rect -28284 -17868 -28180 -17852
rect -28284 -17932 -28264 -17868
rect -28200 -17932 -28180 -17868
rect -28284 -17948 -28180 -17932
rect -28284 -18012 -28264 -17948
rect -28200 -18012 -28180 -17948
rect -28284 -18028 -28180 -18012
rect -28284 -18092 -28264 -18028
rect -28200 -18092 -28180 -18028
rect -28284 -18108 -28180 -18092
rect -28284 -18172 -28264 -18108
rect -28200 -18172 -28180 -18108
rect -28284 -18188 -28180 -18172
rect -28284 -18252 -28264 -18188
rect -28200 -18252 -28180 -18188
rect -28284 -18268 -28180 -18252
rect -28284 -18332 -28264 -18268
rect -28200 -18332 -28180 -18268
rect -28284 -18348 -28180 -18332
rect -28284 -18412 -28264 -18348
rect -28200 -18412 -28180 -18348
rect -28284 -18428 -28180 -18412
rect -28284 -18492 -28264 -18428
rect -28200 -18492 -28180 -18428
rect -28284 -18508 -28180 -18492
rect -28284 -18572 -28264 -18508
rect -28200 -18572 -28180 -18508
rect -28284 -18588 -28180 -18572
rect -28284 -18652 -28264 -18588
rect -28200 -18652 -28180 -18588
rect -28284 -18668 -28180 -18652
rect -28284 -18732 -28264 -18668
rect -28200 -18732 -28180 -18668
rect -28284 -18748 -28180 -18732
rect -28284 -18812 -28264 -18748
rect -28200 -18812 -28180 -18748
rect -28284 -18828 -28180 -18812
rect -28284 -18892 -28264 -18828
rect -28200 -18892 -28180 -18828
rect -28284 -18908 -28180 -18892
rect -28284 -18972 -28264 -18908
rect -28200 -18972 -28180 -18908
rect -28284 -18988 -28180 -18972
rect -28284 -19052 -28264 -18988
rect -28200 -19052 -28180 -18988
rect -28284 -19068 -28180 -19052
rect -28284 -19132 -28264 -19068
rect -28200 -19132 -28180 -19068
rect -28284 -19148 -28180 -19132
rect -28284 -19212 -28264 -19148
rect -28200 -19212 -28180 -19148
rect -28284 -19228 -28180 -19212
rect -28284 -19292 -28264 -19228
rect -28200 -19292 -28180 -19228
rect -28284 -19308 -28180 -19292
rect -28284 -19372 -28264 -19308
rect -28200 -19372 -28180 -19308
rect -28284 -19388 -28180 -19372
rect -28284 -19452 -28264 -19388
rect -28200 -19452 -28180 -19388
rect -28284 -19468 -28180 -19452
rect -28284 -19532 -28264 -19468
rect -28200 -19532 -28180 -19468
rect -28284 -19548 -28180 -19532
rect -28284 -19612 -28264 -19548
rect -28200 -19612 -28180 -19548
rect -28284 -19628 -28180 -19612
rect -28284 -19692 -28264 -19628
rect -28200 -19692 -28180 -19628
rect -28284 -19708 -28180 -19692
rect -28284 -19772 -28264 -19708
rect -28200 -19772 -28180 -19708
rect -28284 -19788 -28180 -19772
rect -28284 -19852 -28264 -19788
rect -28200 -19852 -28180 -19788
rect -28284 -19868 -28180 -19852
rect -28284 -19932 -28264 -19868
rect -28200 -19932 -28180 -19868
rect -28284 -19948 -28180 -19932
rect -28284 -20012 -28264 -19948
rect -28200 -20012 -28180 -19948
rect -28284 -20028 -28180 -20012
rect -28284 -20092 -28264 -20028
rect -28200 -20092 -28180 -20028
rect -28284 -20108 -28180 -20092
rect -28284 -20172 -28264 -20108
rect -28200 -20172 -28180 -20108
rect -28284 -20188 -28180 -20172
rect -28284 -20252 -28264 -20188
rect -28200 -20252 -28180 -20188
rect -28284 -20268 -28180 -20252
rect -28284 -20332 -28264 -20268
rect -28200 -20332 -28180 -20268
rect -28284 -20348 -28180 -20332
rect -28284 -20412 -28264 -20348
rect -28200 -20412 -28180 -20348
rect -28284 -20428 -28180 -20412
rect -28284 -20492 -28264 -20428
rect -28200 -20492 -28180 -20428
rect -28284 -20508 -28180 -20492
rect -28284 -20572 -28264 -20508
rect -28200 -20572 -28180 -20508
rect -28284 -20588 -28180 -20572
rect -28284 -20652 -28264 -20588
rect -28200 -20652 -28180 -20588
rect -28284 -20668 -28180 -20652
rect -28284 -20732 -28264 -20668
rect -28200 -20732 -28180 -20668
rect -28284 -20748 -28180 -20732
rect -28284 -20812 -28264 -20748
rect -28200 -20812 -28180 -20748
rect -28284 -20828 -28180 -20812
rect -28284 -20892 -28264 -20828
rect -28200 -20892 -28180 -20828
rect -28284 -20908 -28180 -20892
rect -28284 -20972 -28264 -20908
rect -28200 -20972 -28180 -20908
rect -28284 -20988 -28180 -20972
rect -28284 -21052 -28264 -20988
rect -28200 -21052 -28180 -20988
rect -28284 -21068 -28180 -21052
rect -33896 -21428 -33792 -21132
rect -39085 -21508 -34163 -21479
rect -39085 -26372 -39056 -21508
rect -34192 -26372 -34163 -21508
rect -39085 -26401 -34163 -26372
rect -33896 -21492 -33876 -21428
rect -33812 -21492 -33792 -21428
rect -31064 -21479 -30960 -21081
rect -28284 -21132 -28264 -21068
rect -28200 -21132 -28180 -21068
rect -27861 -16188 -22939 -16159
rect -27861 -21052 -27832 -16188
rect -22968 -21052 -22939 -16188
rect -27861 -21081 -22939 -21052
rect -22672 -16172 -22652 -16108
rect -22588 -16172 -22568 -16108
rect -19840 -16159 -19736 -15761
rect -17060 -15812 -17040 -15748
rect -16976 -15812 -16956 -15748
rect -16637 -10868 -11715 -10839
rect -16637 -15732 -16608 -10868
rect -11744 -15732 -11715 -10868
rect -16637 -15761 -11715 -15732
rect -11448 -10852 -11428 -10788
rect -11364 -10852 -11344 -10788
rect -8616 -10839 -8512 -10441
rect -5836 -10492 -5816 -10428
rect -5752 -10492 -5732 -10428
rect -5413 -5548 -491 -5519
rect -5413 -10412 -5384 -5548
rect -520 -10412 -491 -5548
rect -5413 -10441 -491 -10412
rect -224 -5532 -204 -5468
rect -140 -5532 -120 -5468
rect 2608 -5519 2712 -5121
rect 5388 -5172 5408 -5108
rect 5472 -5172 5492 -5108
rect 5811 -228 10733 -199
rect 5811 -5092 5840 -228
rect 10704 -5092 10733 -228
rect 5811 -5121 10733 -5092
rect 11000 -212 11020 -148
rect 11084 -212 11104 -148
rect 13832 -199 13936 199
rect 16612 148 16632 212
rect 16696 148 16716 212
rect 17035 5092 21957 5121
rect 17035 228 17064 5092
rect 21928 228 21957 5092
rect 17035 199 21957 228
rect 22224 5108 22244 5172
rect 22308 5108 22328 5172
rect 25056 5121 25160 5519
rect 27836 5468 27856 5532
rect 27920 5468 27940 5532
rect 28259 10412 33181 10441
rect 28259 5548 28288 10412
rect 33152 5548 33181 10412
rect 28259 5519 33181 5548
rect 33448 10428 33468 10492
rect 33532 10428 33552 10492
rect 36280 10441 36384 10839
rect 39060 10788 39080 10852
rect 39144 10788 39164 10852
rect 39060 10492 39164 10788
rect 33448 10412 33552 10428
rect 33448 10348 33468 10412
rect 33532 10348 33552 10412
rect 33448 10332 33552 10348
rect 33448 10268 33468 10332
rect 33532 10268 33552 10332
rect 33448 10252 33552 10268
rect 33448 10188 33468 10252
rect 33532 10188 33552 10252
rect 33448 10172 33552 10188
rect 33448 10108 33468 10172
rect 33532 10108 33552 10172
rect 33448 10092 33552 10108
rect 33448 10028 33468 10092
rect 33532 10028 33552 10092
rect 33448 10012 33552 10028
rect 33448 9948 33468 10012
rect 33532 9948 33552 10012
rect 33448 9932 33552 9948
rect 33448 9868 33468 9932
rect 33532 9868 33552 9932
rect 33448 9852 33552 9868
rect 33448 9788 33468 9852
rect 33532 9788 33552 9852
rect 33448 9772 33552 9788
rect 33448 9708 33468 9772
rect 33532 9708 33552 9772
rect 33448 9692 33552 9708
rect 33448 9628 33468 9692
rect 33532 9628 33552 9692
rect 33448 9612 33552 9628
rect 33448 9548 33468 9612
rect 33532 9548 33552 9612
rect 33448 9532 33552 9548
rect 33448 9468 33468 9532
rect 33532 9468 33552 9532
rect 33448 9452 33552 9468
rect 33448 9388 33468 9452
rect 33532 9388 33552 9452
rect 33448 9372 33552 9388
rect 33448 9308 33468 9372
rect 33532 9308 33552 9372
rect 33448 9292 33552 9308
rect 33448 9228 33468 9292
rect 33532 9228 33552 9292
rect 33448 9212 33552 9228
rect 33448 9148 33468 9212
rect 33532 9148 33552 9212
rect 33448 9132 33552 9148
rect 33448 9068 33468 9132
rect 33532 9068 33552 9132
rect 33448 9052 33552 9068
rect 33448 8988 33468 9052
rect 33532 8988 33552 9052
rect 33448 8972 33552 8988
rect 33448 8908 33468 8972
rect 33532 8908 33552 8972
rect 33448 8892 33552 8908
rect 33448 8828 33468 8892
rect 33532 8828 33552 8892
rect 33448 8812 33552 8828
rect 33448 8748 33468 8812
rect 33532 8748 33552 8812
rect 33448 8732 33552 8748
rect 33448 8668 33468 8732
rect 33532 8668 33552 8732
rect 33448 8652 33552 8668
rect 33448 8588 33468 8652
rect 33532 8588 33552 8652
rect 33448 8572 33552 8588
rect 33448 8508 33468 8572
rect 33532 8508 33552 8572
rect 33448 8492 33552 8508
rect 33448 8428 33468 8492
rect 33532 8428 33552 8492
rect 33448 8412 33552 8428
rect 33448 8348 33468 8412
rect 33532 8348 33552 8412
rect 33448 8332 33552 8348
rect 33448 8268 33468 8332
rect 33532 8268 33552 8332
rect 33448 8252 33552 8268
rect 33448 8188 33468 8252
rect 33532 8188 33552 8252
rect 33448 8172 33552 8188
rect 33448 8108 33468 8172
rect 33532 8108 33552 8172
rect 33448 8092 33552 8108
rect 33448 8028 33468 8092
rect 33532 8028 33552 8092
rect 33448 8012 33552 8028
rect 33448 7948 33468 8012
rect 33532 7948 33552 8012
rect 33448 7932 33552 7948
rect 33448 7868 33468 7932
rect 33532 7868 33552 7932
rect 33448 7852 33552 7868
rect 33448 7788 33468 7852
rect 33532 7788 33552 7852
rect 33448 7772 33552 7788
rect 33448 7708 33468 7772
rect 33532 7708 33552 7772
rect 33448 7692 33552 7708
rect 33448 7628 33468 7692
rect 33532 7628 33552 7692
rect 33448 7612 33552 7628
rect 33448 7548 33468 7612
rect 33532 7548 33552 7612
rect 33448 7532 33552 7548
rect 33448 7468 33468 7532
rect 33532 7468 33552 7532
rect 33448 7452 33552 7468
rect 33448 7388 33468 7452
rect 33532 7388 33552 7452
rect 33448 7372 33552 7388
rect 33448 7308 33468 7372
rect 33532 7308 33552 7372
rect 33448 7292 33552 7308
rect 33448 7228 33468 7292
rect 33532 7228 33552 7292
rect 33448 7212 33552 7228
rect 33448 7148 33468 7212
rect 33532 7148 33552 7212
rect 33448 7132 33552 7148
rect 33448 7068 33468 7132
rect 33532 7068 33552 7132
rect 33448 7052 33552 7068
rect 33448 6988 33468 7052
rect 33532 6988 33552 7052
rect 33448 6972 33552 6988
rect 33448 6908 33468 6972
rect 33532 6908 33552 6972
rect 33448 6892 33552 6908
rect 33448 6828 33468 6892
rect 33532 6828 33552 6892
rect 33448 6812 33552 6828
rect 33448 6748 33468 6812
rect 33532 6748 33552 6812
rect 33448 6732 33552 6748
rect 33448 6668 33468 6732
rect 33532 6668 33552 6732
rect 33448 6652 33552 6668
rect 33448 6588 33468 6652
rect 33532 6588 33552 6652
rect 33448 6572 33552 6588
rect 33448 6508 33468 6572
rect 33532 6508 33552 6572
rect 33448 6492 33552 6508
rect 33448 6428 33468 6492
rect 33532 6428 33552 6492
rect 33448 6412 33552 6428
rect 33448 6348 33468 6412
rect 33532 6348 33552 6412
rect 33448 6332 33552 6348
rect 33448 6268 33468 6332
rect 33532 6268 33552 6332
rect 33448 6252 33552 6268
rect 33448 6188 33468 6252
rect 33532 6188 33552 6252
rect 33448 6172 33552 6188
rect 33448 6108 33468 6172
rect 33532 6108 33552 6172
rect 33448 6092 33552 6108
rect 33448 6028 33468 6092
rect 33532 6028 33552 6092
rect 33448 6012 33552 6028
rect 33448 5948 33468 6012
rect 33532 5948 33552 6012
rect 33448 5932 33552 5948
rect 33448 5868 33468 5932
rect 33532 5868 33552 5932
rect 33448 5852 33552 5868
rect 33448 5788 33468 5852
rect 33532 5788 33552 5852
rect 33448 5772 33552 5788
rect 33448 5708 33468 5772
rect 33532 5708 33552 5772
rect 33448 5692 33552 5708
rect 33448 5628 33468 5692
rect 33532 5628 33552 5692
rect 33448 5612 33552 5628
rect 33448 5548 33468 5612
rect 33532 5548 33552 5612
rect 33448 5532 33552 5548
rect 27836 5172 27940 5468
rect 22224 5092 22328 5108
rect 22224 5028 22244 5092
rect 22308 5028 22328 5092
rect 22224 5012 22328 5028
rect 22224 4948 22244 5012
rect 22308 4948 22328 5012
rect 22224 4932 22328 4948
rect 22224 4868 22244 4932
rect 22308 4868 22328 4932
rect 22224 4852 22328 4868
rect 22224 4788 22244 4852
rect 22308 4788 22328 4852
rect 22224 4772 22328 4788
rect 22224 4708 22244 4772
rect 22308 4708 22328 4772
rect 22224 4692 22328 4708
rect 22224 4628 22244 4692
rect 22308 4628 22328 4692
rect 22224 4612 22328 4628
rect 22224 4548 22244 4612
rect 22308 4548 22328 4612
rect 22224 4532 22328 4548
rect 22224 4468 22244 4532
rect 22308 4468 22328 4532
rect 22224 4452 22328 4468
rect 22224 4388 22244 4452
rect 22308 4388 22328 4452
rect 22224 4372 22328 4388
rect 22224 4308 22244 4372
rect 22308 4308 22328 4372
rect 22224 4292 22328 4308
rect 22224 4228 22244 4292
rect 22308 4228 22328 4292
rect 22224 4212 22328 4228
rect 22224 4148 22244 4212
rect 22308 4148 22328 4212
rect 22224 4132 22328 4148
rect 22224 4068 22244 4132
rect 22308 4068 22328 4132
rect 22224 4052 22328 4068
rect 22224 3988 22244 4052
rect 22308 3988 22328 4052
rect 22224 3972 22328 3988
rect 22224 3908 22244 3972
rect 22308 3908 22328 3972
rect 22224 3892 22328 3908
rect 22224 3828 22244 3892
rect 22308 3828 22328 3892
rect 22224 3812 22328 3828
rect 22224 3748 22244 3812
rect 22308 3748 22328 3812
rect 22224 3732 22328 3748
rect 22224 3668 22244 3732
rect 22308 3668 22328 3732
rect 22224 3652 22328 3668
rect 22224 3588 22244 3652
rect 22308 3588 22328 3652
rect 22224 3572 22328 3588
rect 22224 3508 22244 3572
rect 22308 3508 22328 3572
rect 22224 3492 22328 3508
rect 22224 3428 22244 3492
rect 22308 3428 22328 3492
rect 22224 3412 22328 3428
rect 22224 3348 22244 3412
rect 22308 3348 22328 3412
rect 22224 3332 22328 3348
rect 22224 3268 22244 3332
rect 22308 3268 22328 3332
rect 22224 3252 22328 3268
rect 22224 3188 22244 3252
rect 22308 3188 22328 3252
rect 22224 3172 22328 3188
rect 22224 3108 22244 3172
rect 22308 3108 22328 3172
rect 22224 3092 22328 3108
rect 22224 3028 22244 3092
rect 22308 3028 22328 3092
rect 22224 3012 22328 3028
rect 22224 2948 22244 3012
rect 22308 2948 22328 3012
rect 22224 2932 22328 2948
rect 22224 2868 22244 2932
rect 22308 2868 22328 2932
rect 22224 2852 22328 2868
rect 22224 2788 22244 2852
rect 22308 2788 22328 2852
rect 22224 2772 22328 2788
rect 22224 2708 22244 2772
rect 22308 2708 22328 2772
rect 22224 2692 22328 2708
rect 22224 2628 22244 2692
rect 22308 2628 22328 2692
rect 22224 2612 22328 2628
rect 22224 2548 22244 2612
rect 22308 2548 22328 2612
rect 22224 2532 22328 2548
rect 22224 2468 22244 2532
rect 22308 2468 22328 2532
rect 22224 2452 22328 2468
rect 22224 2388 22244 2452
rect 22308 2388 22328 2452
rect 22224 2372 22328 2388
rect 22224 2308 22244 2372
rect 22308 2308 22328 2372
rect 22224 2292 22328 2308
rect 22224 2228 22244 2292
rect 22308 2228 22328 2292
rect 22224 2212 22328 2228
rect 22224 2148 22244 2212
rect 22308 2148 22328 2212
rect 22224 2132 22328 2148
rect 22224 2068 22244 2132
rect 22308 2068 22328 2132
rect 22224 2052 22328 2068
rect 22224 1988 22244 2052
rect 22308 1988 22328 2052
rect 22224 1972 22328 1988
rect 22224 1908 22244 1972
rect 22308 1908 22328 1972
rect 22224 1892 22328 1908
rect 22224 1828 22244 1892
rect 22308 1828 22328 1892
rect 22224 1812 22328 1828
rect 22224 1748 22244 1812
rect 22308 1748 22328 1812
rect 22224 1732 22328 1748
rect 22224 1668 22244 1732
rect 22308 1668 22328 1732
rect 22224 1652 22328 1668
rect 22224 1588 22244 1652
rect 22308 1588 22328 1652
rect 22224 1572 22328 1588
rect 22224 1508 22244 1572
rect 22308 1508 22328 1572
rect 22224 1492 22328 1508
rect 22224 1428 22244 1492
rect 22308 1428 22328 1492
rect 22224 1412 22328 1428
rect 22224 1348 22244 1412
rect 22308 1348 22328 1412
rect 22224 1332 22328 1348
rect 22224 1268 22244 1332
rect 22308 1268 22328 1332
rect 22224 1252 22328 1268
rect 22224 1188 22244 1252
rect 22308 1188 22328 1252
rect 22224 1172 22328 1188
rect 22224 1108 22244 1172
rect 22308 1108 22328 1172
rect 22224 1092 22328 1108
rect 22224 1028 22244 1092
rect 22308 1028 22328 1092
rect 22224 1012 22328 1028
rect 22224 948 22244 1012
rect 22308 948 22328 1012
rect 22224 932 22328 948
rect 22224 868 22244 932
rect 22308 868 22328 932
rect 22224 852 22328 868
rect 22224 788 22244 852
rect 22308 788 22328 852
rect 22224 772 22328 788
rect 22224 708 22244 772
rect 22308 708 22328 772
rect 22224 692 22328 708
rect 22224 628 22244 692
rect 22308 628 22328 692
rect 22224 612 22328 628
rect 22224 548 22244 612
rect 22308 548 22328 612
rect 22224 532 22328 548
rect 22224 468 22244 532
rect 22308 468 22328 532
rect 22224 452 22328 468
rect 22224 388 22244 452
rect 22308 388 22328 452
rect 22224 372 22328 388
rect 22224 308 22244 372
rect 22308 308 22328 372
rect 22224 292 22328 308
rect 22224 228 22244 292
rect 22308 228 22328 292
rect 22224 212 22328 228
rect 16612 -148 16716 148
rect 11000 -228 11104 -212
rect 11000 -292 11020 -228
rect 11084 -292 11104 -228
rect 11000 -308 11104 -292
rect 11000 -372 11020 -308
rect 11084 -372 11104 -308
rect 11000 -388 11104 -372
rect 11000 -452 11020 -388
rect 11084 -452 11104 -388
rect 11000 -468 11104 -452
rect 11000 -532 11020 -468
rect 11084 -532 11104 -468
rect 11000 -548 11104 -532
rect 11000 -612 11020 -548
rect 11084 -612 11104 -548
rect 11000 -628 11104 -612
rect 11000 -692 11020 -628
rect 11084 -692 11104 -628
rect 11000 -708 11104 -692
rect 11000 -772 11020 -708
rect 11084 -772 11104 -708
rect 11000 -788 11104 -772
rect 11000 -852 11020 -788
rect 11084 -852 11104 -788
rect 11000 -868 11104 -852
rect 11000 -932 11020 -868
rect 11084 -932 11104 -868
rect 11000 -948 11104 -932
rect 11000 -1012 11020 -948
rect 11084 -1012 11104 -948
rect 11000 -1028 11104 -1012
rect 11000 -1092 11020 -1028
rect 11084 -1092 11104 -1028
rect 11000 -1108 11104 -1092
rect 11000 -1172 11020 -1108
rect 11084 -1172 11104 -1108
rect 11000 -1188 11104 -1172
rect 11000 -1252 11020 -1188
rect 11084 -1252 11104 -1188
rect 11000 -1268 11104 -1252
rect 11000 -1332 11020 -1268
rect 11084 -1332 11104 -1268
rect 11000 -1348 11104 -1332
rect 11000 -1412 11020 -1348
rect 11084 -1412 11104 -1348
rect 11000 -1428 11104 -1412
rect 11000 -1492 11020 -1428
rect 11084 -1492 11104 -1428
rect 11000 -1508 11104 -1492
rect 11000 -1572 11020 -1508
rect 11084 -1572 11104 -1508
rect 11000 -1588 11104 -1572
rect 11000 -1652 11020 -1588
rect 11084 -1652 11104 -1588
rect 11000 -1668 11104 -1652
rect 11000 -1732 11020 -1668
rect 11084 -1732 11104 -1668
rect 11000 -1748 11104 -1732
rect 11000 -1812 11020 -1748
rect 11084 -1812 11104 -1748
rect 11000 -1828 11104 -1812
rect 11000 -1892 11020 -1828
rect 11084 -1892 11104 -1828
rect 11000 -1908 11104 -1892
rect 11000 -1972 11020 -1908
rect 11084 -1972 11104 -1908
rect 11000 -1988 11104 -1972
rect 11000 -2052 11020 -1988
rect 11084 -2052 11104 -1988
rect 11000 -2068 11104 -2052
rect 11000 -2132 11020 -2068
rect 11084 -2132 11104 -2068
rect 11000 -2148 11104 -2132
rect 11000 -2212 11020 -2148
rect 11084 -2212 11104 -2148
rect 11000 -2228 11104 -2212
rect 11000 -2292 11020 -2228
rect 11084 -2292 11104 -2228
rect 11000 -2308 11104 -2292
rect 11000 -2372 11020 -2308
rect 11084 -2372 11104 -2308
rect 11000 -2388 11104 -2372
rect 11000 -2452 11020 -2388
rect 11084 -2452 11104 -2388
rect 11000 -2468 11104 -2452
rect 11000 -2532 11020 -2468
rect 11084 -2532 11104 -2468
rect 11000 -2548 11104 -2532
rect 11000 -2612 11020 -2548
rect 11084 -2612 11104 -2548
rect 11000 -2628 11104 -2612
rect 11000 -2692 11020 -2628
rect 11084 -2692 11104 -2628
rect 11000 -2708 11104 -2692
rect 11000 -2772 11020 -2708
rect 11084 -2772 11104 -2708
rect 11000 -2788 11104 -2772
rect 11000 -2852 11020 -2788
rect 11084 -2852 11104 -2788
rect 11000 -2868 11104 -2852
rect 11000 -2932 11020 -2868
rect 11084 -2932 11104 -2868
rect 11000 -2948 11104 -2932
rect 11000 -3012 11020 -2948
rect 11084 -3012 11104 -2948
rect 11000 -3028 11104 -3012
rect 11000 -3092 11020 -3028
rect 11084 -3092 11104 -3028
rect 11000 -3108 11104 -3092
rect 11000 -3172 11020 -3108
rect 11084 -3172 11104 -3108
rect 11000 -3188 11104 -3172
rect 11000 -3252 11020 -3188
rect 11084 -3252 11104 -3188
rect 11000 -3268 11104 -3252
rect 11000 -3332 11020 -3268
rect 11084 -3332 11104 -3268
rect 11000 -3348 11104 -3332
rect 11000 -3412 11020 -3348
rect 11084 -3412 11104 -3348
rect 11000 -3428 11104 -3412
rect 11000 -3492 11020 -3428
rect 11084 -3492 11104 -3428
rect 11000 -3508 11104 -3492
rect 11000 -3572 11020 -3508
rect 11084 -3572 11104 -3508
rect 11000 -3588 11104 -3572
rect 11000 -3652 11020 -3588
rect 11084 -3652 11104 -3588
rect 11000 -3668 11104 -3652
rect 11000 -3732 11020 -3668
rect 11084 -3732 11104 -3668
rect 11000 -3748 11104 -3732
rect 11000 -3812 11020 -3748
rect 11084 -3812 11104 -3748
rect 11000 -3828 11104 -3812
rect 11000 -3892 11020 -3828
rect 11084 -3892 11104 -3828
rect 11000 -3908 11104 -3892
rect 11000 -3972 11020 -3908
rect 11084 -3972 11104 -3908
rect 11000 -3988 11104 -3972
rect 11000 -4052 11020 -3988
rect 11084 -4052 11104 -3988
rect 11000 -4068 11104 -4052
rect 11000 -4132 11020 -4068
rect 11084 -4132 11104 -4068
rect 11000 -4148 11104 -4132
rect 11000 -4212 11020 -4148
rect 11084 -4212 11104 -4148
rect 11000 -4228 11104 -4212
rect 11000 -4292 11020 -4228
rect 11084 -4292 11104 -4228
rect 11000 -4308 11104 -4292
rect 11000 -4372 11020 -4308
rect 11084 -4372 11104 -4308
rect 11000 -4388 11104 -4372
rect 11000 -4452 11020 -4388
rect 11084 -4452 11104 -4388
rect 11000 -4468 11104 -4452
rect 11000 -4532 11020 -4468
rect 11084 -4532 11104 -4468
rect 11000 -4548 11104 -4532
rect 11000 -4612 11020 -4548
rect 11084 -4612 11104 -4548
rect 11000 -4628 11104 -4612
rect 11000 -4692 11020 -4628
rect 11084 -4692 11104 -4628
rect 11000 -4708 11104 -4692
rect 11000 -4772 11020 -4708
rect 11084 -4772 11104 -4708
rect 11000 -4788 11104 -4772
rect 11000 -4852 11020 -4788
rect 11084 -4852 11104 -4788
rect 11000 -4868 11104 -4852
rect 11000 -4932 11020 -4868
rect 11084 -4932 11104 -4868
rect 11000 -4948 11104 -4932
rect 11000 -5012 11020 -4948
rect 11084 -5012 11104 -4948
rect 11000 -5028 11104 -5012
rect 11000 -5092 11020 -5028
rect 11084 -5092 11104 -5028
rect 11000 -5108 11104 -5092
rect 5388 -5468 5492 -5172
rect -224 -5548 -120 -5532
rect -224 -5612 -204 -5548
rect -140 -5612 -120 -5548
rect -224 -5628 -120 -5612
rect -224 -5692 -204 -5628
rect -140 -5692 -120 -5628
rect -224 -5708 -120 -5692
rect -224 -5772 -204 -5708
rect -140 -5772 -120 -5708
rect -224 -5788 -120 -5772
rect -224 -5852 -204 -5788
rect -140 -5852 -120 -5788
rect -224 -5868 -120 -5852
rect -224 -5932 -204 -5868
rect -140 -5932 -120 -5868
rect -224 -5948 -120 -5932
rect -224 -6012 -204 -5948
rect -140 -6012 -120 -5948
rect -224 -6028 -120 -6012
rect -224 -6092 -204 -6028
rect -140 -6092 -120 -6028
rect -224 -6108 -120 -6092
rect -224 -6172 -204 -6108
rect -140 -6172 -120 -6108
rect -224 -6188 -120 -6172
rect -224 -6252 -204 -6188
rect -140 -6252 -120 -6188
rect -224 -6268 -120 -6252
rect -224 -6332 -204 -6268
rect -140 -6332 -120 -6268
rect -224 -6348 -120 -6332
rect -224 -6412 -204 -6348
rect -140 -6412 -120 -6348
rect -224 -6428 -120 -6412
rect -224 -6492 -204 -6428
rect -140 -6492 -120 -6428
rect -224 -6508 -120 -6492
rect -224 -6572 -204 -6508
rect -140 -6572 -120 -6508
rect -224 -6588 -120 -6572
rect -224 -6652 -204 -6588
rect -140 -6652 -120 -6588
rect -224 -6668 -120 -6652
rect -224 -6732 -204 -6668
rect -140 -6732 -120 -6668
rect -224 -6748 -120 -6732
rect -224 -6812 -204 -6748
rect -140 -6812 -120 -6748
rect -224 -6828 -120 -6812
rect -224 -6892 -204 -6828
rect -140 -6892 -120 -6828
rect -224 -6908 -120 -6892
rect -224 -6972 -204 -6908
rect -140 -6972 -120 -6908
rect -224 -6988 -120 -6972
rect -224 -7052 -204 -6988
rect -140 -7052 -120 -6988
rect -224 -7068 -120 -7052
rect -224 -7132 -204 -7068
rect -140 -7132 -120 -7068
rect -224 -7148 -120 -7132
rect -224 -7212 -204 -7148
rect -140 -7212 -120 -7148
rect -224 -7228 -120 -7212
rect -224 -7292 -204 -7228
rect -140 -7292 -120 -7228
rect -224 -7308 -120 -7292
rect -224 -7372 -204 -7308
rect -140 -7372 -120 -7308
rect -224 -7388 -120 -7372
rect -224 -7452 -204 -7388
rect -140 -7452 -120 -7388
rect -224 -7468 -120 -7452
rect -224 -7532 -204 -7468
rect -140 -7532 -120 -7468
rect -224 -7548 -120 -7532
rect -224 -7612 -204 -7548
rect -140 -7612 -120 -7548
rect -224 -7628 -120 -7612
rect -224 -7692 -204 -7628
rect -140 -7692 -120 -7628
rect -224 -7708 -120 -7692
rect -224 -7772 -204 -7708
rect -140 -7772 -120 -7708
rect -224 -7788 -120 -7772
rect -224 -7852 -204 -7788
rect -140 -7852 -120 -7788
rect -224 -7868 -120 -7852
rect -224 -7932 -204 -7868
rect -140 -7932 -120 -7868
rect -224 -7948 -120 -7932
rect -224 -8012 -204 -7948
rect -140 -8012 -120 -7948
rect -224 -8028 -120 -8012
rect -224 -8092 -204 -8028
rect -140 -8092 -120 -8028
rect -224 -8108 -120 -8092
rect -224 -8172 -204 -8108
rect -140 -8172 -120 -8108
rect -224 -8188 -120 -8172
rect -224 -8252 -204 -8188
rect -140 -8252 -120 -8188
rect -224 -8268 -120 -8252
rect -224 -8332 -204 -8268
rect -140 -8332 -120 -8268
rect -224 -8348 -120 -8332
rect -224 -8412 -204 -8348
rect -140 -8412 -120 -8348
rect -224 -8428 -120 -8412
rect -224 -8492 -204 -8428
rect -140 -8492 -120 -8428
rect -224 -8508 -120 -8492
rect -224 -8572 -204 -8508
rect -140 -8572 -120 -8508
rect -224 -8588 -120 -8572
rect -224 -8652 -204 -8588
rect -140 -8652 -120 -8588
rect -224 -8668 -120 -8652
rect -224 -8732 -204 -8668
rect -140 -8732 -120 -8668
rect -224 -8748 -120 -8732
rect -224 -8812 -204 -8748
rect -140 -8812 -120 -8748
rect -224 -8828 -120 -8812
rect -224 -8892 -204 -8828
rect -140 -8892 -120 -8828
rect -224 -8908 -120 -8892
rect -224 -8972 -204 -8908
rect -140 -8972 -120 -8908
rect -224 -8988 -120 -8972
rect -224 -9052 -204 -8988
rect -140 -9052 -120 -8988
rect -224 -9068 -120 -9052
rect -224 -9132 -204 -9068
rect -140 -9132 -120 -9068
rect -224 -9148 -120 -9132
rect -224 -9212 -204 -9148
rect -140 -9212 -120 -9148
rect -224 -9228 -120 -9212
rect -224 -9292 -204 -9228
rect -140 -9292 -120 -9228
rect -224 -9308 -120 -9292
rect -224 -9372 -204 -9308
rect -140 -9372 -120 -9308
rect -224 -9388 -120 -9372
rect -224 -9452 -204 -9388
rect -140 -9452 -120 -9388
rect -224 -9468 -120 -9452
rect -224 -9532 -204 -9468
rect -140 -9532 -120 -9468
rect -224 -9548 -120 -9532
rect -224 -9612 -204 -9548
rect -140 -9612 -120 -9548
rect -224 -9628 -120 -9612
rect -224 -9692 -204 -9628
rect -140 -9692 -120 -9628
rect -224 -9708 -120 -9692
rect -224 -9772 -204 -9708
rect -140 -9772 -120 -9708
rect -224 -9788 -120 -9772
rect -224 -9852 -204 -9788
rect -140 -9852 -120 -9788
rect -224 -9868 -120 -9852
rect -224 -9932 -204 -9868
rect -140 -9932 -120 -9868
rect -224 -9948 -120 -9932
rect -224 -10012 -204 -9948
rect -140 -10012 -120 -9948
rect -224 -10028 -120 -10012
rect -224 -10092 -204 -10028
rect -140 -10092 -120 -10028
rect -224 -10108 -120 -10092
rect -224 -10172 -204 -10108
rect -140 -10172 -120 -10108
rect -224 -10188 -120 -10172
rect -224 -10252 -204 -10188
rect -140 -10252 -120 -10188
rect -224 -10268 -120 -10252
rect -224 -10332 -204 -10268
rect -140 -10332 -120 -10268
rect -224 -10348 -120 -10332
rect -224 -10412 -204 -10348
rect -140 -10412 -120 -10348
rect -224 -10428 -120 -10412
rect -5836 -10788 -5732 -10492
rect -11448 -10868 -11344 -10852
rect -11448 -10932 -11428 -10868
rect -11364 -10932 -11344 -10868
rect -11448 -10948 -11344 -10932
rect -11448 -11012 -11428 -10948
rect -11364 -11012 -11344 -10948
rect -11448 -11028 -11344 -11012
rect -11448 -11092 -11428 -11028
rect -11364 -11092 -11344 -11028
rect -11448 -11108 -11344 -11092
rect -11448 -11172 -11428 -11108
rect -11364 -11172 -11344 -11108
rect -11448 -11188 -11344 -11172
rect -11448 -11252 -11428 -11188
rect -11364 -11252 -11344 -11188
rect -11448 -11268 -11344 -11252
rect -11448 -11332 -11428 -11268
rect -11364 -11332 -11344 -11268
rect -11448 -11348 -11344 -11332
rect -11448 -11412 -11428 -11348
rect -11364 -11412 -11344 -11348
rect -11448 -11428 -11344 -11412
rect -11448 -11492 -11428 -11428
rect -11364 -11492 -11344 -11428
rect -11448 -11508 -11344 -11492
rect -11448 -11572 -11428 -11508
rect -11364 -11572 -11344 -11508
rect -11448 -11588 -11344 -11572
rect -11448 -11652 -11428 -11588
rect -11364 -11652 -11344 -11588
rect -11448 -11668 -11344 -11652
rect -11448 -11732 -11428 -11668
rect -11364 -11732 -11344 -11668
rect -11448 -11748 -11344 -11732
rect -11448 -11812 -11428 -11748
rect -11364 -11812 -11344 -11748
rect -11448 -11828 -11344 -11812
rect -11448 -11892 -11428 -11828
rect -11364 -11892 -11344 -11828
rect -11448 -11908 -11344 -11892
rect -11448 -11972 -11428 -11908
rect -11364 -11972 -11344 -11908
rect -11448 -11988 -11344 -11972
rect -11448 -12052 -11428 -11988
rect -11364 -12052 -11344 -11988
rect -11448 -12068 -11344 -12052
rect -11448 -12132 -11428 -12068
rect -11364 -12132 -11344 -12068
rect -11448 -12148 -11344 -12132
rect -11448 -12212 -11428 -12148
rect -11364 -12212 -11344 -12148
rect -11448 -12228 -11344 -12212
rect -11448 -12292 -11428 -12228
rect -11364 -12292 -11344 -12228
rect -11448 -12308 -11344 -12292
rect -11448 -12372 -11428 -12308
rect -11364 -12372 -11344 -12308
rect -11448 -12388 -11344 -12372
rect -11448 -12452 -11428 -12388
rect -11364 -12452 -11344 -12388
rect -11448 -12468 -11344 -12452
rect -11448 -12532 -11428 -12468
rect -11364 -12532 -11344 -12468
rect -11448 -12548 -11344 -12532
rect -11448 -12612 -11428 -12548
rect -11364 -12612 -11344 -12548
rect -11448 -12628 -11344 -12612
rect -11448 -12692 -11428 -12628
rect -11364 -12692 -11344 -12628
rect -11448 -12708 -11344 -12692
rect -11448 -12772 -11428 -12708
rect -11364 -12772 -11344 -12708
rect -11448 -12788 -11344 -12772
rect -11448 -12852 -11428 -12788
rect -11364 -12852 -11344 -12788
rect -11448 -12868 -11344 -12852
rect -11448 -12932 -11428 -12868
rect -11364 -12932 -11344 -12868
rect -11448 -12948 -11344 -12932
rect -11448 -13012 -11428 -12948
rect -11364 -13012 -11344 -12948
rect -11448 -13028 -11344 -13012
rect -11448 -13092 -11428 -13028
rect -11364 -13092 -11344 -13028
rect -11448 -13108 -11344 -13092
rect -11448 -13172 -11428 -13108
rect -11364 -13172 -11344 -13108
rect -11448 -13188 -11344 -13172
rect -11448 -13252 -11428 -13188
rect -11364 -13252 -11344 -13188
rect -11448 -13268 -11344 -13252
rect -11448 -13332 -11428 -13268
rect -11364 -13332 -11344 -13268
rect -11448 -13348 -11344 -13332
rect -11448 -13412 -11428 -13348
rect -11364 -13412 -11344 -13348
rect -11448 -13428 -11344 -13412
rect -11448 -13492 -11428 -13428
rect -11364 -13492 -11344 -13428
rect -11448 -13508 -11344 -13492
rect -11448 -13572 -11428 -13508
rect -11364 -13572 -11344 -13508
rect -11448 -13588 -11344 -13572
rect -11448 -13652 -11428 -13588
rect -11364 -13652 -11344 -13588
rect -11448 -13668 -11344 -13652
rect -11448 -13732 -11428 -13668
rect -11364 -13732 -11344 -13668
rect -11448 -13748 -11344 -13732
rect -11448 -13812 -11428 -13748
rect -11364 -13812 -11344 -13748
rect -11448 -13828 -11344 -13812
rect -11448 -13892 -11428 -13828
rect -11364 -13892 -11344 -13828
rect -11448 -13908 -11344 -13892
rect -11448 -13972 -11428 -13908
rect -11364 -13972 -11344 -13908
rect -11448 -13988 -11344 -13972
rect -11448 -14052 -11428 -13988
rect -11364 -14052 -11344 -13988
rect -11448 -14068 -11344 -14052
rect -11448 -14132 -11428 -14068
rect -11364 -14132 -11344 -14068
rect -11448 -14148 -11344 -14132
rect -11448 -14212 -11428 -14148
rect -11364 -14212 -11344 -14148
rect -11448 -14228 -11344 -14212
rect -11448 -14292 -11428 -14228
rect -11364 -14292 -11344 -14228
rect -11448 -14308 -11344 -14292
rect -11448 -14372 -11428 -14308
rect -11364 -14372 -11344 -14308
rect -11448 -14388 -11344 -14372
rect -11448 -14452 -11428 -14388
rect -11364 -14452 -11344 -14388
rect -11448 -14468 -11344 -14452
rect -11448 -14532 -11428 -14468
rect -11364 -14532 -11344 -14468
rect -11448 -14548 -11344 -14532
rect -11448 -14612 -11428 -14548
rect -11364 -14612 -11344 -14548
rect -11448 -14628 -11344 -14612
rect -11448 -14692 -11428 -14628
rect -11364 -14692 -11344 -14628
rect -11448 -14708 -11344 -14692
rect -11448 -14772 -11428 -14708
rect -11364 -14772 -11344 -14708
rect -11448 -14788 -11344 -14772
rect -11448 -14852 -11428 -14788
rect -11364 -14852 -11344 -14788
rect -11448 -14868 -11344 -14852
rect -11448 -14932 -11428 -14868
rect -11364 -14932 -11344 -14868
rect -11448 -14948 -11344 -14932
rect -11448 -15012 -11428 -14948
rect -11364 -15012 -11344 -14948
rect -11448 -15028 -11344 -15012
rect -11448 -15092 -11428 -15028
rect -11364 -15092 -11344 -15028
rect -11448 -15108 -11344 -15092
rect -11448 -15172 -11428 -15108
rect -11364 -15172 -11344 -15108
rect -11448 -15188 -11344 -15172
rect -11448 -15252 -11428 -15188
rect -11364 -15252 -11344 -15188
rect -11448 -15268 -11344 -15252
rect -11448 -15332 -11428 -15268
rect -11364 -15332 -11344 -15268
rect -11448 -15348 -11344 -15332
rect -11448 -15412 -11428 -15348
rect -11364 -15412 -11344 -15348
rect -11448 -15428 -11344 -15412
rect -11448 -15492 -11428 -15428
rect -11364 -15492 -11344 -15428
rect -11448 -15508 -11344 -15492
rect -11448 -15572 -11428 -15508
rect -11364 -15572 -11344 -15508
rect -11448 -15588 -11344 -15572
rect -11448 -15652 -11428 -15588
rect -11364 -15652 -11344 -15588
rect -11448 -15668 -11344 -15652
rect -11448 -15732 -11428 -15668
rect -11364 -15732 -11344 -15668
rect -11448 -15748 -11344 -15732
rect -17060 -16108 -16956 -15812
rect -22672 -16188 -22568 -16172
rect -22672 -16252 -22652 -16188
rect -22588 -16252 -22568 -16188
rect -22672 -16268 -22568 -16252
rect -22672 -16332 -22652 -16268
rect -22588 -16332 -22568 -16268
rect -22672 -16348 -22568 -16332
rect -22672 -16412 -22652 -16348
rect -22588 -16412 -22568 -16348
rect -22672 -16428 -22568 -16412
rect -22672 -16492 -22652 -16428
rect -22588 -16492 -22568 -16428
rect -22672 -16508 -22568 -16492
rect -22672 -16572 -22652 -16508
rect -22588 -16572 -22568 -16508
rect -22672 -16588 -22568 -16572
rect -22672 -16652 -22652 -16588
rect -22588 -16652 -22568 -16588
rect -22672 -16668 -22568 -16652
rect -22672 -16732 -22652 -16668
rect -22588 -16732 -22568 -16668
rect -22672 -16748 -22568 -16732
rect -22672 -16812 -22652 -16748
rect -22588 -16812 -22568 -16748
rect -22672 -16828 -22568 -16812
rect -22672 -16892 -22652 -16828
rect -22588 -16892 -22568 -16828
rect -22672 -16908 -22568 -16892
rect -22672 -16972 -22652 -16908
rect -22588 -16972 -22568 -16908
rect -22672 -16988 -22568 -16972
rect -22672 -17052 -22652 -16988
rect -22588 -17052 -22568 -16988
rect -22672 -17068 -22568 -17052
rect -22672 -17132 -22652 -17068
rect -22588 -17132 -22568 -17068
rect -22672 -17148 -22568 -17132
rect -22672 -17212 -22652 -17148
rect -22588 -17212 -22568 -17148
rect -22672 -17228 -22568 -17212
rect -22672 -17292 -22652 -17228
rect -22588 -17292 -22568 -17228
rect -22672 -17308 -22568 -17292
rect -22672 -17372 -22652 -17308
rect -22588 -17372 -22568 -17308
rect -22672 -17388 -22568 -17372
rect -22672 -17452 -22652 -17388
rect -22588 -17452 -22568 -17388
rect -22672 -17468 -22568 -17452
rect -22672 -17532 -22652 -17468
rect -22588 -17532 -22568 -17468
rect -22672 -17548 -22568 -17532
rect -22672 -17612 -22652 -17548
rect -22588 -17612 -22568 -17548
rect -22672 -17628 -22568 -17612
rect -22672 -17692 -22652 -17628
rect -22588 -17692 -22568 -17628
rect -22672 -17708 -22568 -17692
rect -22672 -17772 -22652 -17708
rect -22588 -17772 -22568 -17708
rect -22672 -17788 -22568 -17772
rect -22672 -17852 -22652 -17788
rect -22588 -17852 -22568 -17788
rect -22672 -17868 -22568 -17852
rect -22672 -17932 -22652 -17868
rect -22588 -17932 -22568 -17868
rect -22672 -17948 -22568 -17932
rect -22672 -18012 -22652 -17948
rect -22588 -18012 -22568 -17948
rect -22672 -18028 -22568 -18012
rect -22672 -18092 -22652 -18028
rect -22588 -18092 -22568 -18028
rect -22672 -18108 -22568 -18092
rect -22672 -18172 -22652 -18108
rect -22588 -18172 -22568 -18108
rect -22672 -18188 -22568 -18172
rect -22672 -18252 -22652 -18188
rect -22588 -18252 -22568 -18188
rect -22672 -18268 -22568 -18252
rect -22672 -18332 -22652 -18268
rect -22588 -18332 -22568 -18268
rect -22672 -18348 -22568 -18332
rect -22672 -18412 -22652 -18348
rect -22588 -18412 -22568 -18348
rect -22672 -18428 -22568 -18412
rect -22672 -18492 -22652 -18428
rect -22588 -18492 -22568 -18428
rect -22672 -18508 -22568 -18492
rect -22672 -18572 -22652 -18508
rect -22588 -18572 -22568 -18508
rect -22672 -18588 -22568 -18572
rect -22672 -18652 -22652 -18588
rect -22588 -18652 -22568 -18588
rect -22672 -18668 -22568 -18652
rect -22672 -18732 -22652 -18668
rect -22588 -18732 -22568 -18668
rect -22672 -18748 -22568 -18732
rect -22672 -18812 -22652 -18748
rect -22588 -18812 -22568 -18748
rect -22672 -18828 -22568 -18812
rect -22672 -18892 -22652 -18828
rect -22588 -18892 -22568 -18828
rect -22672 -18908 -22568 -18892
rect -22672 -18972 -22652 -18908
rect -22588 -18972 -22568 -18908
rect -22672 -18988 -22568 -18972
rect -22672 -19052 -22652 -18988
rect -22588 -19052 -22568 -18988
rect -22672 -19068 -22568 -19052
rect -22672 -19132 -22652 -19068
rect -22588 -19132 -22568 -19068
rect -22672 -19148 -22568 -19132
rect -22672 -19212 -22652 -19148
rect -22588 -19212 -22568 -19148
rect -22672 -19228 -22568 -19212
rect -22672 -19292 -22652 -19228
rect -22588 -19292 -22568 -19228
rect -22672 -19308 -22568 -19292
rect -22672 -19372 -22652 -19308
rect -22588 -19372 -22568 -19308
rect -22672 -19388 -22568 -19372
rect -22672 -19452 -22652 -19388
rect -22588 -19452 -22568 -19388
rect -22672 -19468 -22568 -19452
rect -22672 -19532 -22652 -19468
rect -22588 -19532 -22568 -19468
rect -22672 -19548 -22568 -19532
rect -22672 -19612 -22652 -19548
rect -22588 -19612 -22568 -19548
rect -22672 -19628 -22568 -19612
rect -22672 -19692 -22652 -19628
rect -22588 -19692 -22568 -19628
rect -22672 -19708 -22568 -19692
rect -22672 -19772 -22652 -19708
rect -22588 -19772 -22568 -19708
rect -22672 -19788 -22568 -19772
rect -22672 -19852 -22652 -19788
rect -22588 -19852 -22568 -19788
rect -22672 -19868 -22568 -19852
rect -22672 -19932 -22652 -19868
rect -22588 -19932 -22568 -19868
rect -22672 -19948 -22568 -19932
rect -22672 -20012 -22652 -19948
rect -22588 -20012 -22568 -19948
rect -22672 -20028 -22568 -20012
rect -22672 -20092 -22652 -20028
rect -22588 -20092 -22568 -20028
rect -22672 -20108 -22568 -20092
rect -22672 -20172 -22652 -20108
rect -22588 -20172 -22568 -20108
rect -22672 -20188 -22568 -20172
rect -22672 -20252 -22652 -20188
rect -22588 -20252 -22568 -20188
rect -22672 -20268 -22568 -20252
rect -22672 -20332 -22652 -20268
rect -22588 -20332 -22568 -20268
rect -22672 -20348 -22568 -20332
rect -22672 -20412 -22652 -20348
rect -22588 -20412 -22568 -20348
rect -22672 -20428 -22568 -20412
rect -22672 -20492 -22652 -20428
rect -22588 -20492 -22568 -20428
rect -22672 -20508 -22568 -20492
rect -22672 -20572 -22652 -20508
rect -22588 -20572 -22568 -20508
rect -22672 -20588 -22568 -20572
rect -22672 -20652 -22652 -20588
rect -22588 -20652 -22568 -20588
rect -22672 -20668 -22568 -20652
rect -22672 -20732 -22652 -20668
rect -22588 -20732 -22568 -20668
rect -22672 -20748 -22568 -20732
rect -22672 -20812 -22652 -20748
rect -22588 -20812 -22568 -20748
rect -22672 -20828 -22568 -20812
rect -22672 -20892 -22652 -20828
rect -22588 -20892 -22568 -20828
rect -22672 -20908 -22568 -20892
rect -22672 -20972 -22652 -20908
rect -22588 -20972 -22568 -20908
rect -22672 -20988 -22568 -20972
rect -22672 -21052 -22652 -20988
rect -22588 -21052 -22568 -20988
rect -22672 -21068 -22568 -21052
rect -28284 -21428 -28180 -21132
rect -33896 -21508 -33792 -21492
rect -33896 -21572 -33876 -21508
rect -33812 -21572 -33792 -21508
rect -33896 -21588 -33792 -21572
rect -33896 -21652 -33876 -21588
rect -33812 -21652 -33792 -21588
rect -33896 -21668 -33792 -21652
rect -33896 -21732 -33876 -21668
rect -33812 -21732 -33792 -21668
rect -33896 -21748 -33792 -21732
rect -33896 -21812 -33876 -21748
rect -33812 -21812 -33792 -21748
rect -33896 -21828 -33792 -21812
rect -33896 -21892 -33876 -21828
rect -33812 -21892 -33792 -21828
rect -33896 -21908 -33792 -21892
rect -33896 -21972 -33876 -21908
rect -33812 -21972 -33792 -21908
rect -33896 -21988 -33792 -21972
rect -33896 -22052 -33876 -21988
rect -33812 -22052 -33792 -21988
rect -33896 -22068 -33792 -22052
rect -33896 -22132 -33876 -22068
rect -33812 -22132 -33792 -22068
rect -33896 -22148 -33792 -22132
rect -33896 -22212 -33876 -22148
rect -33812 -22212 -33792 -22148
rect -33896 -22228 -33792 -22212
rect -33896 -22292 -33876 -22228
rect -33812 -22292 -33792 -22228
rect -33896 -22308 -33792 -22292
rect -33896 -22372 -33876 -22308
rect -33812 -22372 -33792 -22308
rect -33896 -22388 -33792 -22372
rect -33896 -22452 -33876 -22388
rect -33812 -22452 -33792 -22388
rect -33896 -22468 -33792 -22452
rect -33896 -22532 -33876 -22468
rect -33812 -22532 -33792 -22468
rect -33896 -22548 -33792 -22532
rect -33896 -22612 -33876 -22548
rect -33812 -22612 -33792 -22548
rect -33896 -22628 -33792 -22612
rect -33896 -22692 -33876 -22628
rect -33812 -22692 -33792 -22628
rect -33896 -22708 -33792 -22692
rect -33896 -22772 -33876 -22708
rect -33812 -22772 -33792 -22708
rect -33896 -22788 -33792 -22772
rect -33896 -22852 -33876 -22788
rect -33812 -22852 -33792 -22788
rect -33896 -22868 -33792 -22852
rect -33896 -22932 -33876 -22868
rect -33812 -22932 -33792 -22868
rect -33896 -22948 -33792 -22932
rect -33896 -23012 -33876 -22948
rect -33812 -23012 -33792 -22948
rect -33896 -23028 -33792 -23012
rect -33896 -23092 -33876 -23028
rect -33812 -23092 -33792 -23028
rect -33896 -23108 -33792 -23092
rect -33896 -23172 -33876 -23108
rect -33812 -23172 -33792 -23108
rect -33896 -23188 -33792 -23172
rect -33896 -23252 -33876 -23188
rect -33812 -23252 -33792 -23188
rect -33896 -23268 -33792 -23252
rect -33896 -23332 -33876 -23268
rect -33812 -23332 -33792 -23268
rect -33896 -23348 -33792 -23332
rect -33896 -23412 -33876 -23348
rect -33812 -23412 -33792 -23348
rect -33896 -23428 -33792 -23412
rect -33896 -23492 -33876 -23428
rect -33812 -23492 -33792 -23428
rect -33896 -23508 -33792 -23492
rect -33896 -23572 -33876 -23508
rect -33812 -23572 -33792 -23508
rect -33896 -23588 -33792 -23572
rect -33896 -23652 -33876 -23588
rect -33812 -23652 -33792 -23588
rect -33896 -23668 -33792 -23652
rect -33896 -23732 -33876 -23668
rect -33812 -23732 -33792 -23668
rect -33896 -23748 -33792 -23732
rect -33896 -23812 -33876 -23748
rect -33812 -23812 -33792 -23748
rect -33896 -23828 -33792 -23812
rect -33896 -23892 -33876 -23828
rect -33812 -23892 -33792 -23828
rect -33896 -23908 -33792 -23892
rect -33896 -23972 -33876 -23908
rect -33812 -23972 -33792 -23908
rect -33896 -23988 -33792 -23972
rect -33896 -24052 -33876 -23988
rect -33812 -24052 -33792 -23988
rect -33896 -24068 -33792 -24052
rect -33896 -24132 -33876 -24068
rect -33812 -24132 -33792 -24068
rect -33896 -24148 -33792 -24132
rect -33896 -24212 -33876 -24148
rect -33812 -24212 -33792 -24148
rect -33896 -24228 -33792 -24212
rect -33896 -24292 -33876 -24228
rect -33812 -24292 -33792 -24228
rect -33896 -24308 -33792 -24292
rect -33896 -24372 -33876 -24308
rect -33812 -24372 -33792 -24308
rect -33896 -24388 -33792 -24372
rect -33896 -24452 -33876 -24388
rect -33812 -24452 -33792 -24388
rect -33896 -24468 -33792 -24452
rect -33896 -24532 -33876 -24468
rect -33812 -24532 -33792 -24468
rect -33896 -24548 -33792 -24532
rect -33896 -24612 -33876 -24548
rect -33812 -24612 -33792 -24548
rect -33896 -24628 -33792 -24612
rect -33896 -24692 -33876 -24628
rect -33812 -24692 -33792 -24628
rect -33896 -24708 -33792 -24692
rect -33896 -24772 -33876 -24708
rect -33812 -24772 -33792 -24708
rect -33896 -24788 -33792 -24772
rect -33896 -24852 -33876 -24788
rect -33812 -24852 -33792 -24788
rect -33896 -24868 -33792 -24852
rect -33896 -24932 -33876 -24868
rect -33812 -24932 -33792 -24868
rect -33896 -24948 -33792 -24932
rect -33896 -25012 -33876 -24948
rect -33812 -25012 -33792 -24948
rect -33896 -25028 -33792 -25012
rect -33896 -25092 -33876 -25028
rect -33812 -25092 -33792 -25028
rect -33896 -25108 -33792 -25092
rect -33896 -25172 -33876 -25108
rect -33812 -25172 -33792 -25108
rect -33896 -25188 -33792 -25172
rect -33896 -25252 -33876 -25188
rect -33812 -25252 -33792 -25188
rect -33896 -25268 -33792 -25252
rect -33896 -25332 -33876 -25268
rect -33812 -25332 -33792 -25268
rect -33896 -25348 -33792 -25332
rect -33896 -25412 -33876 -25348
rect -33812 -25412 -33792 -25348
rect -33896 -25428 -33792 -25412
rect -33896 -25492 -33876 -25428
rect -33812 -25492 -33792 -25428
rect -33896 -25508 -33792 -25492
rect -33896 -25572 -33876 -25508
rect -33812 -25572 -33792 -25508
rect -33896 -25588 -33792 -25572
rect -33896 -25652 -33876 -25588
rect -33812 -25652 -33792 -25588
rect -33896 -25668 -33792 -25652
rect -33896 -25732 -33876 -25668
rect -33812 -25732 -33792 -25668
rect -33896 -25748 -33792 -25732
rect -33896 -25812 -33876 -25748
rect -33812 -25812 -33792 -25748
rect -33896 -25828 -33792 -25812
rect -33896 -25892 -33876 -25828
rect -33812 -25892 -33792 -25828
rect -33896 -25908 -33792 -25892
rect -33896 -25972 -33876 -25908
rect -33812 -25972 -33792 -25908
rect -33896 -25988 -33792 -25972
rect -33896 -26052 -33876 -25988
rect -33812 -26052 -33792 -25988
rect -33896 -26068 -33792 -26052
rect -33896 -26132 -33876 -26068
rect -33812 -26132 -33792 -26068
rect -33896 -26148 -33792 -26132
rect -33896 -26212 -33876 -26148
rect -33812 -26212 -33792 -26148
rect -33896 -26228 -33792 -26212
rect -33896 -26292 -33876 -26228
rect -33812 -26292 -33792 -26228
rect -33896 -26308 -33792 -26292
rect -33896 -26372 -33876 -26308
rect -33812 -26372 -33792 -26308
rect -33896 -26388 -33792 -26372
rect -36676 -26799 -36572 -26401
rect -33896 -26452 -33876 -26388
rect -33812 -26452 -33792 -26388
rect -33473 -21508 -28551 -21479
rect -33473 -26372 -33444 -21508
rect -28580 -26372 -28551 -21508
rect -33473 -26401 -28551 -26372
rect -28284 -21492 -28264 -21428
rect -28200 -21492 -28180 -21428
rect -25452 -21479 -25348 -21081
rect -22672 -21132 -22652 -21068
rect -22588 -21132 -22568 -21068
rect -22249 -16188 -17327 -16159
rect -22249 -21052 -22220 -16188
rect -17356 -21052 -17327 -16188
rect -22249 -21081 -17327 -21052
rect -17060 -16172 -17040 -16108
rect -16976 -16172 -16956 -16108
rect -14228 -16159 -14124 -15761
rect -11448 -15812 -11428 -15748
rect -11364 -15812 -11344 -15748
rect -11025 -10868 -6103 -10839
rect -11025 -15732 -10996 -10868
rect -6132 -15732 -6103 -10868
rect -11025 -15761 -6103 -15732
rect -5836 -10852 -5816 -10788
rect -5752 -10852 -5732 -10788
rect -3004 -10839 -2900 -10441
rect -224 -10492 -204 -10428
rect -140 -10492 -120 -10428
rect 199 -5548 5121 -5519
rect 199 -10412 228 -5548
rect 5092 -10412 5121 -5548
rect 199 -10441 5121 -10412
rect 5388 -5532 5408 -5468
rect 5472 -5532 5492 -5468
rect 8220 -5519 8324 -5121
rect 11000 -5172 11020 -5108
rect 11084 -5172 11104 -5108
rect 11423 -228 16345 -199
rect 11423 -5092 11452 -228
rect 16316 -5092 16345 -228
rect 11423 -5121 16345 -5092
rect 16612 -212 16632 -148
rect 16696 -212 16716 -148
rect 19444 -199 19548 199
rect 22224 148 22244 212
rect 22308 148 22328 212
rect 22647 5092 27569 5121
rect 22647 228 22676 5092
rect 27540 228 27569 5092
rect 22647 199 27569 228
rect 27836 5108 27856 5172
rect 27920 5108 27940 5172
rect 30668 5121 30772 5519
rect 33448 5468 33468 5532
rect 33532 5468 33552 5532
rect 33871 10412 38793 10441
rect 33871 5548 33900 10412
rect 38764 5548 38793 10412
rect 33871 5519 38793 5548
rect 39060 10428 39080 10492
rect 39144 10428 39164 10492
rect 39060 10412 39164 10428
rect 39060 10348 39080 10412
rect 39144 10348 39164 10412
rect 39060 10332 39164 10348
rect 39060 10268 39080 10332
rect 39144 10268 39164 10332
rect 39060 10252 39164 10268
rect 39060 10188 39080 10252
rect 39144 10188 39164 10252
rect 39060 10172 39164 10188
rect 39060 10108 39080 10172
rect 39144 10108 39164 10172
rect 39060 10092 39164 10108
rect 39060 10028 39080 10092
rect 39144 10028 39164 10092
rect 39060 10012 39164 10028
rect 39060 9948 39080 10012
rect 39144 9948 39164 10012
rect 39060 9932 39164 9948
rect 39060 9868 39080 9932
rect 39144 9868 39164 9932
rect 39060 9852 39164 9868
rect 39060 9788 39080 9852
rect 39144 9788 39164 9852
rect 39060 9772 39164 9788
rect 39060 9708 39080 9772
rect 39144 9708 39164 9772
rect 39060 9692 39164 9708
rect 39060 9628 39080 9692
rect 39144 9628 39164 9692
rect 39060 9612 39164 9628
rect 39060 9548 39080 9612
rect 39144 9548 39164 9612
rect 39060 9532 39164 9548
rect 39060 9468 39080 9532
rect 39144 9468 39164 9532
rect 39060 9452 39164 9468
rect 39060 9388 39080 9452
rect 39144 9388 39164 9452
rect 39060 9372 39164 9388
rect 39060 9308 39080 9372
rect 39144 9308 39164 9372
rect 39060 9292 39164 9308
rect 39060 9228 39080 9292
rect 39144 9228 39164 9292
rect 39060 9212 39164 9228
rect 39060 9148 39080 9212
rect 39144 9148 39164 9212
rect 39060 9132 39164 9148
rect 39060 9068 39080 9132
rect 39144 9068 39164 9132
rect 39060 9052 39164 9068
rect 39060 8988 39080 9052
rect 39144 8988 39164 9052
rect 39060 8972 39164 8988
rect 39060 8908 39080 8972
rect 39144 8908 39164 8972
rect 39060 8892 39164 8908
rect 39060 8828 39080 8892
rect 39144 8828 39164 8892
rect 39060 8812 39164 8828
rect 39060 8748 39080 8812
rect 39144 8748 39164 8812
rect 39060 8732 39164 8748
rect 39060 8668 39080 8732
rect 39144 8668 39164 8732
rect 39060 8652 39164 8668
rect 39060 8588 39080 8652
rect 39144 8588 39164 8652
rect 39060 8572 39164 8588
rect 39060 8508 39080 8572
rect 39144 8508 39164 8572
rect 39060 8492 39164 8508
rect 39060 8428 39080 8492
rect 39144 8428 39164 8492
rect 39060 8412 39164 8428
rect 39060 8348 39080 8412
rect 39144 8348 39164 8412
rect 39060 8332 39164 8348
rect 39060 8268 39080 8332
rect 39144 8268 39164 8332
rect 39060 8252 39164 8268
rect 39060 8188 39080 8252
rect 39144 8188 39164 8252
rect 39060 8172 39164 8188
rect 39060 8108 39080 8172
rect 39144 8108 39164 8172
rect 39060 8092 39164 8108
rect 39060 8028 39080 8092
rect 39144 8028 39164 8092
rect 39060 8012 39164 8028
rect 39060 7948 39080 8012
rect 39144 7948 39164 8012
rect 39060 7932 39164 7948
rect 39060 7868 39080 7932
rect 39144 7868 39164 7932
rect 39060 7852 39164 7868
rect 39060 7788 39080 7852
rect 39144 7788 39164 7852
rect 39060 7772 39164 7788
rect 39060 7708 39080 7772
rect 39144 7708 39164 7772
rect 39060 7692 39164 7708
rect 39060 7628 39080 7692
rect 39144 7628 39164 7692
rect 39060 7612 39164 7628
rect 39060 7548 39080 7612
rect 39144 7548 39164 7612
rect 39060 7532 39164 7548
rect 39060 7468 39080 7532
rect 39144 7468 39164 7532
rect 39060 7452 39164 7468
rect 39060 7388 39080 7452
rect 39144 7388 39164 7452
rect 39060 7372 39164 7388
rect 39060 7308 39080 7372
rect 39144 7308 39164 7372
rect 39060 7292 39164 7308
rect 39060 7228 39080 7292
rect 39144 7228 39164 7292
rect 39060 7212 39164 7228
rect 39060 7148 39080 7212
rect 39144 7148 39164 7212
rect 39060 7132 39164 7148
rect 39060 7068 39080 7132
rect 39144 7068 39164 7132
rect 39060 7052 39164 7068
rect 39060 6988 39080 7052
rect 39144 6988 39164 7052
rect 39060 6972 39164 6988
rect 39060 6908 39080 6972
rect 39144 6908 39164 6972
rect 39060 6892 39164 6908
rect 39060 6828 39080 6892
rect 39144 6828 39164 6892
rect 39060 6812 39164 6828
rect 39060 6748 39080 6812
rect 39144 6748 39164 6812
rect 39060 6732 39164 6748
rect 39060 6668 39080 6732
rect 39144 6668 39164 6732
rect 39060 6652 39164 6668
rect 39060 6588 39080 6652
rect 39144 6588 39164 6652
rect 39060 6572 39164 6588
rect 39060 6508 39080 6572
rect 39144 6508 39164 6572
rect 39060 6492 39164 6508
rect 39060 6428 39080 6492
rect 39144 6428 39164 6492
rect 39060 6412 39164 6428
rect 39060 6348 39080 6412
rect 39144 6348 39164 6412
rect 39060 6332 39164 6348
rect 39060 6268 39080 6332
rect 39144 6268 39164 6332
rect 39060 6252 39164 6268
rect 39060 6188 39080 6252
rect 39144 6188 39164 6252
rect 39060 6172 39164 6188
rect 39060 6108 39080 6172
rect 39144 6108 39164 6172
rect 39060 6092 39164 6108
rect 39060 6028 39080 6092
rect 39144 6028 39164 6092
rect 39060 6012 39164 6028
rect 39060 5948 39080 6012
rect 39144 5948 39164 6012
rect 39060 5932 39164 5948
rect 39060 5868 39080 5932
rect 39144 5868 39164 5932
rect 39060 5852 39164 5868
rect 39060 5788 39080 5852
rect 39144 5788 39164 5852
rect 39060 5772 39164 5788
rect 39060 5708 39080 5772
rect 39144 5708 39164 5772
rect 39060 5692 39164 5708
rect 39060 5628 39080 5692
rect 39144 5628 39164 5692
rect 39060 5612 39164 5628
rect 39060 5548 39080 5612
rect 39144 5548 39164 5612
rect 39060 5532 39164 5548
rect 33448 5172 33552 5468
rect 27836 5092 27940 5108
rect 27836 5028 27856 5092
rect 27920 5028 27940 5092
rect 27836 5012 27940 5028
rect 27836 4948 27856 5012
rect 27920 4948 27940 5012
rect 27836 4932 27940 4948
rect 27836 4868 27856 4932
rect 27920 4868 27940 4932
rect 27836 4852 27940 4868
rect 27836 4788 27856 4852
rect 27920 4788 27940 4852
rect 27836 4772 27940 4788
rect 27836 4708 27856 4772
rect 27920 4708 27940 4772
rect 27836 4692 27940 4708
rect 27836 4628 27856 4692
rect 27920 4628 27940 4692
rect 27836 4612 27940 4628
rect 27836 4548 27856 4612
rect 27920 4548 27940 4612
rect 27836 4532 27940 4548
rect 27836 4468 27856 4532
rect 27920 4468 27940 4532
rect 27836 4452 27940 4468
rect 27836 4388 27856 4452
rect 27920 4388 27940 4452
rect 27836 4372 27940 4388
rect 27836 4308 27856 4372
rect 27920 4308 27940 4372
rect 27836 4292 27940 4308
rect 27836 4228 27856 4292
rect 27920 4228 27940 4292
rect 27836 4212 27940 4228
rect 27836 4148 27856 4212
rect 27920 4148 27940 4212
rect 27836 4132 27940 4148
rect 27836 4068 27856 4132
rect 27920 4068 27940 4132
rect 27836 4052 27940 4068
rect 27836 3988 27856 4052
rect 27920 3988 27940 4052
rect 27836 3972 27940 3988
rect 27836 3908 27856 3972
rect 27920 3908 27940 3972
rect 27836 3892 27940 3908
rect 27836 3828 27856 3892
rect 27920 3828 27940 3892
rect 27836 3812 27940 3828
rect 27836 3748 27856 3812
rect 27920 3748 27940 3812
rect 27836 3732 27940 3748
rect 27836 3668 27856 3732
rect 27920 3668 27940 3732
rect 27836 3652 27940 3668
rect 27836 3588 27856 3652
rect 27920 3588 27940 3652
rect 27836 3572 27940 3588
rect 27836 3508 27856 3572
rect 27920 3508 27940 3572
rect 27836 3492 27940 3508
rect 27836 3428 27856 3492
rect 27920 3428 27940 3492
rect 27836 3412 27940 3428
rect 27836 3348 27856 3412
rect 27920 3348 27940 3412
rect 27836 3332 27940 3348
rect 27836 3268 27856 3332
rect 27920 3268 27940 3332
rect 27836 3252 27940 3268
rect 27836 3188 27856 3252
rect 27920 3188 27940 3252
rect 27836 3172 27940 3188
rect 27836 3108 27856 3172
rect 27920 3108 27940 3172
rect 27836 3092 27940 3108
rect 27836 3028 27856 3092
rect 27920 3028 27940 3092
rect 27836 3012 27940 3028
rect 27836 2948 27856 3012
rect 27920 2948 27940 3012
rect 27836 2932 27940 2948
rect 27836 2868 27856 2932
rect 27920 2868 27940 2932
rect 27836 2852 27940 2868
rect 27836 2788 27856 2852
rect 27920 2788 27940 2852
rect 27836 2772 27940 2788
rect 27836 2708 27856 2772
rect 27920 2708 27940 2772
rect 27836 2692 27940 2708
rect 27836 2628 27856 2692
rect 27920 2628 27940 2692
rect 27836 2612 27940 2628
rect 27836 2548 27856 2612
rect 27920 2548 27940 2612
rect 27836 2532 27940 2548
rect 27836 2468 27856 2532
rect 27920 2468 27940 2532
rect 27836 2452 27940 2468
rect 27836 2388 27856 2452
rect 27920 2388 27940 2452
rect 27836 2372 27940 2388
rect 27836 2308 27856 2372
rect 27920 2308 27940 2372
rect 27836 2292 27940 2308
rect 27836 2228 27856 2292
rect 27920 2228 27940 2292
rect 27836 2212 27940 2228
rect 27836 2148 27856 2212
rect 27920 2148 27940 2212
rect 27836 2132 27940 2148
rect 27836 2068 27856 2132
rect 27920 2068 27940 2132
rect 27836 2052 27940 2068
rect 27836 1988 27856 2052
rect 27920 1988 27940 2052
rect 27836 1972 27940 1988
rect 27836 1908 27856 1972
rect 27920 1908 27940 1972
rect 27836 1892 27940 1908
rect 27836 1828 27856 1892
rect 27920 1828 27940 1892
rect 27836 1812 27940 1828
rect 27836 1748 27856 1812
rect 27920 1748 27940 1812
rect 27836 1732 27940 1748
rect 27836 1668 27856 1732
rect 27920 1668 27940 1732
rect 27836 1652 27940 1668
rect 27836 1588 27856 1652
rect 27920 1588 27940 1652
rect 27836 1572 27940 1588
rect 27836 1508 27856 1572
rect 27920 1508 27940 1572
rect 27836 1492 27940 1508
rect 27836 1428 27856 1492
rect 27920 1428 27940 1492
rect 27836 1412 27940 1428
rect 27836 1348 27856 1412
rect 27920 1348 27940 1412
rect 27836 1332 27940 1348
rect 27836 1268 27856 1332
rect 27920 1268 27940 1332
rect 27836 1252 27940 1268
rect 27836 1188 27856 1252
rect 27920 1188 27940 1252
rect 27836 1172 27940 1188
rect 27836 1108 27856 1172
rect 27920 1108 27940 1172
rect 27836 1092 27940 1108
rect 27836 1028 27856 1092
rect 27920 1028 27940 1092
rect 27836 1012 27940 1028
rect 27836 948 27856 1012
rect 27920 948 27940 1012
rect 27836 932 27940 948
rect 27836 868 27856 932
rect 27920 868 27940 932
rect 27836 852 27940 868
rect 27836 788 27856 852
rect 27920 788 27940 852
rect 27836 772 27940 788
rect 27836 708 27856 772
rect 27920 708 27940 772
rect 27836 692 27940 708
rect 27836 628 27856 692
rect 27920 628 27940 692
rect 27836 612 27940 628
rect 27836 548 27856 612
rect 27920 548 27940 612
rect 27836 532 27940 548
rect 27836 468 27856 532
rect 27920 468 27940 532
rect 27836 452 27940 468
rect 27836 388 27856 452
rect 27920 388 27940 452
rect 27836 372 27940 388
rect 27836 308 27856 372
rect 27920 308 27940 372
rect 27836 292 27940 308
rect 27836 228 27856 292
rect 27920 228 27940 292
rect 27836 212 27940 228
rect 22224 -148 22328 148
rect 16612 -228 16716 -212
rect 16612 -292 16632 -228
rect 16696 -292 16716 -228
rect 16612 -308 16716 -292
rect 16612 -372 16632 -308
rect 16696 -372 16716 -308
rect 16612 -388 16716 -372
rect 16612 -452 16632 -388
rect 16696 -452 16716 -388
rect 16612 -468 16716 -452
rect 16612 -532 16632 -468
rect 16696 -532 16716 -468
rect 16612 -548 16716 -532
rect 16612 -612 16632 -548
rect 16696 -612 16716 -548
rect 16612 -628 16716 -612
rect 16612 -692 16632 -628
rect 16696 -692 16716 -628
rect 16612 -708 16716 -692
rect 16612 -772 16632 -708
rect 16696 -772 16716 -708
rect 16612 -788 16716 -772
rect 16612 -852 16632 -788
rect 16696 -852 16716 -788
rect 16612 -868 16716 -852
rect 16612 -932 16632 -868
rect 16696 -932 16716 -868
rect 16612 -948 16716 -932
rect 16612 -1012 16632 -948
rect 16696 -1012 16716 -948
rect 16612 -1028 16716 -1012
rect 16612 -1092 16632 -1028
rect 16696 -1092 16716 -1028
rect 16612 -1108 16716 -1092
rect 16612 -1172 16632 -1108
rect 16696 -1172 16716 -1108
rect 16612 -1188 16716 -1172
rect 16612 -1252 16632 -1188
rect 16696 -1252 16716 -1188
rect 16612 -1268 16716 -1252
rect 16612 -1332 16632 -1268
rect 16696 -1332 16716 -1268
rect 16612 -1348 16716 -1332
rect 16612 -1412 16632 -1348
rect 16696 -1412 16716 -1348
rect 16612 -1428 16716 -1412
rect 16612 -1492 16632 -1428
rect 16696 -1492 16716 -1428
rect 16612 -1508 16716 -1492
rect 16612 -1572 16632 -1508
rect 16696 -1572 16716 -1508
rect 16612 -1588 16716 -1572
rect 16612 -1652 16632 -1588
rect 16696 -1652 16716 -1588
rect 16612 -1668 16716 -1652
rect 16612 -1732 16632 -1668
rect 16696 -1732 16716 -1668
rect 16612 -1748 16716 -1732
rect 16612 -1812 16632 -1748
rect 16696 -1812 16716 -1748
rect 16612 -1828 16716 -1812
rect 16612 -1892 16632 -1828
rect 16696 -1892 16716 -1828
rect 16612 -1908 16716 -1892
rect 16612 -1972 16632 -1908
rect 16696 -1972 16716 -1908
rect 16612 -1988 16716 -1972
rect 16612 -2052 16632 -1988
rect 16696 -2052 16716 -1988
rect 16612 -2068 16716 -2052
rect 16612 -2132 16632 -2068
rect 16696 -2132 16716 -2068
rect 16612 -2148 16716 -2132
rect 16612 -2212 16632 -2148
rect 16696 -2212 16716 -2148
rect 16612 -2228 16716 -2212
rect 16612 -2292 16632 -2228
rect 16696 -2292 16716 -2228
rect 16612 -2308 16716 -2292
rect 16612 -2372 16632 -2308
rect 16696 -2372 16716 -2308
rect 16612 -2388 16716 -2372
rect 16612 -2452 16632 -2388
rect 16696 -2452 16716 -2388
rect 16612 -2468 16716 -2452
rect 16612 -2532 16632 -2468
rect 16696 -2532 16716 -2468
rect 16612 -2548 16716 -2532
rect 16612 -2612 16632 -2548
rect 16696 -2612 16716 -2548
rect 16612 -2628 16716 -2612
rect 16612 -2692 16632 -2628
rect 16696 -2692 16716 -2628
rect 16612 -2708 16716 -2692
rect 16612 -2772 16632 -2708
rect 16696 -2772 16716 -2708
rect 16612 -2788 16716 -2772
rect 16612 -2852 16632 -2788
rect 16696 -2852 16716 -2788
rect 16612 -2868 16716 -2852
rect 16612 -2932 16632 -2868
rect 16696 -2932 16716 -2868
rect 16612 -2948 16716 -2932
rect 16612 -3012 16632 -2948
rect 16696 -3012 16716 -2948
rect 16612 -3028 16716 -3012
rect 16612 -3092 16632 -3028
rect 16696 -3092 16716 -3028
rect 16612 -3108 16716 -3092
rect 16612 -3172 16632 -3108
rect 16696 -3172 16716 -3108
rect 16612 -3188 16716 -3172
rect 16612 -3252 16632 -3188
rect 16696 -3252 16716 -3188
rect 16612 -3268 16716 -3252
rect 16612 -3332 16632 -3268
rect 16696 -3332 16716 -3268
rect 16612 -3348 16716 -3332
rect 16612 -3412 16632 -3348
rect 16696 -3412 16716 -3348
rect 16612 -3428 16716 -3412
rect 16612 -3492 16632 -3428
rect 16696 -3492 16716 -3428
rect 16612 -3508 16716 -3492
rect 16612 -3572 16632 -3508
rect 16696 -3572 16716 -3508
rect 16612 -3588 16716 -3572
rect 16612 -3652 16632 -3588
rect 16696 -3652 16716 -3588
rect 16612 -3668 16716 -3652
rect 16612 -3732 16632 -3668
rect 16696 -3732 16716 -3668
rect 16612 -3748 16716 -3732
rect 16612 -3812 16632 -3748
rect 16696 -3812 16716 -3748
rect 16612 -3828 16716 -3812
rect 16612 -3892 16632 -3828
rect 16696 -3892 16716 -3828
rect 16612 -3908 16716 -3892
rect 16612 -3972 16632 -3908
rect 16696 -3972 16716 -3908
rect 16612 -3988 16716 -3972
rect 16612 -4052 16632 -3988
rect 16696 -4052 16716 -3988
rect 16612 -4068 16716 -4052
rect 16612 -4132 16632 -4068
rect 16696 -4132 16716 -4068
rect 16612 -4148 16716 -4132
rect 16612 -4212 16632 -4148
rect 16696 -4212 16716 -4148
rect 16612 -4228 16716 -4212
rect 16612 -4292 16632 -4228
rect 16696 -4292 16716 -4228
rect 16612 -4308 16716 -4292
rect 16612 -4372 16632 -4308
rect 16696 -4372 16716 -4308
rect 16612 -4388 16716 -4372
rect 16612 -4452 16632 -4388
rect 16696 -4452 16716 -4388
rect 16612 -4468 16716 -4452
rect 16612 -4532 16632 -4468
rect 16696 -4532 16716 -4468
rect 16612 -4548 16716 -4532
rect 16612 -4612 16632 -4548
rect 16696 -4612 16716 -4548
rect 16612 -4628 16716 -4612
rect 16612 -4692 16632 -4628
rect 16696 -4692 16716 -4628
rect 16612 -4708 16716 -4692
rect 16612 -4772 16632 -4708
rect 16696 -4772 16716 -4708
rect 16612 -4788 16716 -4772
rect 16612 -4852 16632 -4788
rect 16696 -4852 16716 -4788
rect 16612 -4868 16716 -4852
rect 16612 -4932 16632 -4868
rect 16696 -4932 16716 -4868
rect 16612 -4948 16716 -4932
rect 16612 -5012 16632 -4948
rect 16696 -5012 16716 -4948
rect 16612 -5028 16716 -5012
rect 16612 -5092 16632 -5028
rect 16696 -5092 16716 -5028
rect 16612 -5108 16716 -5092
rect 11000 -5468 11104 -5172
rect 5388 -5548 5492 -5532
rect 5388 -5612 5408 -5548
rect 5472 -5612 5492 -5548
rect 5388 -5628 5492 -5612
rect 5388 -5692 5408 -5628
rect 5472 -5692 5492 -5628
rect 5388 -5708 5492 -5692
rect 5388 -5772 5408 -5708
rect 5472 -5772 5492 -5708
rect 5388 -5788 5492 -5772
rect 5388 -5852 5408 -5788
rect 5472 -5852 5492 -5788
rect 5388 -5868 5492 -5852
rect 5388 -5932 5408 -5868
rect 5472 -5932 5492 -5868
rect 5388 -5948 5492 -5932
rect 5388 -6012 5408 -5948
rect 5472 -6012 5492 -5948
rect 5388 -6028 5492 -6012
rect 5388 -6092 5408 -6028
rect 5472 -6092 5492 -6028
rect 5388 -6108 5492 -6092
rect 5388 -6172 5408 -6108
rect 5472 -6172 5492 -6108
rect 5388 -6188 5492 -6172
rect 5388 -6252 5408 -6188
rect 5472 -6252 5492 -6188
rect 5388 -6268 5492 -6252
rect 5388 -6332 5408 -6268
rect 5472 -6332 5492 -6268
rect 5388 -6348 5492 -6332
rect 5388 -6412 5408 -6348
rect 5472 -6412 5492 -6348
rect 5388 -6428 5492 -6412
rect 5388 -6492 5408 -6428
rect 5472 -6492 5492 -6428
rect 5388 -6508 5492 -6492
rect 5388 -6572 5408 -6508
rect 5472 -6572 5492 -6508
rect 5388 -6588 5492 -6572
rect 5388 -6652 5408 -6588
rect 5472 -6652 5492 -6588
rect 5388 -6668 5492 -6652
rect 5388 -6732 5408 -6668
rect 5472 -6732 5492 -6668
rect 5388 -6748 5492 -6732
rect 5388 -6812 5408 -6748
rect 5472 -6812 5492 -6748
rect 5388 -6828 5492 -6812
rect 5388 -6892 5408 -6828
rect 5472 -6892 5492 -6828
rect 5388 -6908 5492 -6892
rect 5388 -6972 5408 -6908
rect 5472 -6972 5492 -6908
rect 5388 -6988 5492 -6972
rect 5388 -7052 5408 -6988
rect 5472 -7052 5492 -6988
rect 5388 -7068 5492 -7052
rect 5388 -7132 5408 -7068
rect 5472 -7132 5492 -7068
rect 5388 -7148 5492 -7132
rect 5388 -7212 5408 -7148
rect 5472 -7212 5492 -7148
rect 5388 -7228 5492 -7212
rect 5388 -7292 5408 -7228
rect 5472 -7292 5492 -7228
rect 5388 -7308 5492 -7292
rect 5388 -7372 5408 -7308
rect 5472 -7372 5492 -7308
rect 5388 -7388 5492 -7372
rect 5388 -7452 5408 -7388
rect 5472 -7452 5492 -7388
rect 5388 -7468 5492 -7452
rect 5388 -7532 5408 -7468
rect 5472 -7532 5492 -7468
rect 5388 -7548 5492 -7532
rect 5388 -7612 5408 -7548
rect 5472 -7612 5492 -7548
rect 5388 -7628 5492 -7612
rect 5388 -7692 5408 -7628
rect 5472 -7692 5492 -7628
rect 5388 -7708 5492 -7692
rect 5388 -7772 5408 -7708
rect 5472 -7772 5492 -7708
rect 5388 -7788 5492 -7772
rect 5388 -7852 5408 -7788
rect 5472 -7852 5492 -7788
rect 5388 -7868 5492 -7852
rect 5388 -7932 5408 -7868
rect 5472 -7932 5492 -7868
rect 5388 -7948 5492 -7932
rect 5388 -8012 5408 -7948
rect 5472 -8012 5492 -7948
rect 5388 -8028 5492 -8012
rect 5388 -8092 5408 -8028
rect 5472 -8092 5492 -8028
rect 5388 -8108 5492 -8092
rect 5388 -8172 5408 -8108
rect 5472 -8172 5492 -8108
rect 5388 -8188 5492 -8172
rect 5388 -8252 5408 -8188
rect 5472 -8252 5492 -8188
rect 5388 -8268 5492 -8252
rect 5388 -8332 5408 -8268
rect 5472 -8332 5492 -8268
rect 5388 -8348 5492 -8332
rect 5388 -8412 5408 -8348
rect 5472 -8412 5492 -8348
rect 5388 -8428 5492 -8412
rect 5388 -8492 5408 -8428
rect 5472 -8492 5492 -8428
rect 5388 -8508 5492 -8492
rect 5388 -8572 5408 -8508
rect 5472 -8572 5492 -8508
rect 5388 -8588 5492 -8572
rect 5388 -8652 5408 -8588
rect 5472 -8652 5492 -8588
rect 5388 -8668 5492 -8652
rect 5388 -8732 5408 -8668
rect 5472 -8732 5492 -8668
rect 5388 -8748 5492 -8732
rect 5388 -8812 5408 -8748
rect 5472 -8812 5492 -8748
rect 5388 -8828 5492 -8812
rect 5388 -8892 5408 -8828
rect 5472 -8892 5492 -8828
rect 5388 -8908 5492 -8892
rect 5388 -8972 5408 -8908
rect 5472 -8972 5492 -8908
rect 5388 -8988 5492 -8972
rect 5388 -9052 5408 -8988
rect 5472 -9052 5492 -8988
rect 5388 -9068 5492 -9052
rect 5388 -9132 5408 -9068
rect 5472 -9132 5492 -9068
rect 5388 -9148 5492 -9132
rect 5388 -9212 5408 -9148
rect 5472 -9212 5492 -9148
rect 5388 -9228 5492 -9212
rect 5388 -9292 5408 -9228
rect 5472 -9292 5492 -9228
rect 5388 -9308 5492 -9292
rect 5388 -9372 5408 -9308
rect 5472 -9372 5492 -9308
rect 5388 -9388 5492 -9372
rect 5388 -9452 5408 -9388
rect 5472 -9452 5492 -9388
rect 5388 -9468 5492 -9452
rect 5388 -9532 5408 -9468
rect 5472 -9532 5492 -9468
rect 5388 -9548 5492 -9532
rect 5388 -9612 5408 -9548
rect 5472 -9612 5492 -9548
rect 5388 -9628 5492 -9612
rect 5388 -9692 5408 -9628
rect 5472 -9692 5492 -9628
rect 5388 -9708 5492 -9692
rect 5388 -9772 5408 -9708
rect 5472 -9772 5492 -9708
rect 5388 -9788 5492 -9772
rect 5388 -9852 5408 -9788
rect 5472 -9852 5492 -9788
rect 5388 -9868 5492 -9852
rect 5388 -9932 5408 -9868
rect 5472 -9932 5492 -9868
rect 5388 -9948 5492 -9932
rect 5388 -10012 5408 -9948
rect 5472 -10012 5492 -9948
rect 5388 -10028 5492 -10012
rect 5388 -10092 5408 -10028
rect 5472 -10092 5492 -10028
rect 5388 -10108 5492 -10092
rect 5388 -10172 5408 -10108
rect 5472 -10172 5492 -10108
rect 5388 -10188 5492 -10172
rect 5388 -10252 5408 -10188
rect 5472 -10252 5492 -10188
rect 5388 -10268 5492 -10252
rect 5388 -10332 5408 -10268
rect 5472 -10332 5492 -10268
rect 5388 -10348 5492 -10332
rect 5388 -10412 5408 -10348
rect 5472 -10412 5492 -10348
rect 5388 -10428 5492 -10412
rect -224 -10788 -120 -10492
rect -5836 -10868 -5732 -10852
rect -5836 -10932 -5816 -10868
rect -5752 -10932 -5732 -10868
rect -5836 -10948 -5732 -10932
rect -5836 -11012 -5816 -10948
rect -5752 -11012 -5732 -10948
rect -5836 -11028 -5732 -11012
rect -5836 -11092 -5816 -11028
rect -5752 -11092 -5732 -11028
rect -5836 -11108 -5732 -11092
rect -5836 -11172 -5816 -11108
rect -5752 -11172 -5732 -11108
rect -5836 -11188 -5732 -11172
rect -5836 -11252 -5816 -11188
rect -5752 -11252 -5732 -11188
rect -5836 -11268 -5732 -11252
rect -5836 -11332 -5816 -11268
rect -5752 -11332 -5732 -11268
rect -5836 -11348 -5732 -11332
rect -5836 -11412 -5816 -11348
rect -5752 -11412 -5732 -11348
rect -5836 -11428 -5732 -11412
rect -5836 -11492 -5816 -11428
rect -5752 -11492 -5732 -11428
rect -5836 -11508 -5732 -11492
rect -5836 -11572 -5816 -11508
rect -5752 -11572 -5732 -11508
rect -5836 -11588 -5732 -11572
rect -5836 -11652 -5816 -11588
rect -5752 -11652 -5732 -11588
rect -5836 -11668 -5732 -11652
rect -5836 -11732 -5816 -11668
rect -5752 -11732 -5732 -11668
rect -5836 -11748 -5732 -11732
rect -5836 -11812 -5816 -11748
rect -5752 -11812 -5732 -11748
rect -5836 -11828 -5732 -11812
rect -5836 -11892 -5816 -11828
rect -5752 -11892 -5732 -11828
rect -5836 -11908 -5732 -11892
rect -5836 -11972 -5816 -11908
rect -5752 -11972 -5732 -11908
rect -5836 -11988 -5732 -11972
rect -5836 -12052 -5816 -11988
rect -5752 -12052 -5732 -11988
rect -5836 -12068 -5732 -12052
rect -5836 -12132 -5816 -12068
rect -5752 -12132 -5732 -12068
rect -5836 -12148 -5732 -12132
rect -5836 -12212 -5816 -12148
rect -5752 -12212 -5732 -12148
rect -5836 -12228 -5732 -12212
rect -5836 -12292 -5816 -12228
rect -5752 -12292 -5732 -12228
rect -5836 -12308 -5732 -12292
rect -5836 -12372 -5816 -12308
rect -5752 -12372 -5732 -12308
rect -5836 -12388 -5732 -12372
rect -5836 -12452 -5816 -12388
rect -5752 -12452 -5732 -12388
rect -5836 -12468 -5732 -12452
rect -5836 -12532 -5816 -12468
rect -5752 -12532 -5732 -12468
rect -5836 -12548 -5732 -12532
rect -5836 -12612 -5816 -12548
rect -5752 -12612 -5732 -12548
rect -5836 -12628 -5732 -12612
rect -5836 -12692 -5816 -12628
rect -5752 -12692 -5732 -12628
rect -5836 -12708 -5732 -12692
rect -5836 -12772 -5816 -12708
rect -5752 -12772 -5732 -12708
rect -5836 -12788 -5732 -12772
rect -5836 -12852 -5816 -12788
rect -5752 -12852 -5732 -12788
rect -5836 -12868 -5732 -12852
rect -5836 -12932 -5816 -12868
rect -5752 -12932 -5732 -12868
rect -5836 -12948 -5732 -12932
rect -5836 -13012 -5816 -12948
rect -5752 -13012 -5732 -12948
rect -5836 -13028 -5732 -13012
rect -5836 -13092 -5816 -13028
rect -5752 -13092 -5732 -13028
rect -5836 -13108 -5732 -13092
rect -5836 -13172 -5816 -13108
rect -5752 -13172 -5732 -13108
rect -5836 -13188 -5732 -13172
rect -5836 -13252 -5816 -13188
rect -5752 -13252 -5732 -13188
rect -5836 -13268 -5732 -13252
rect -5836 -13332 -5816 -13268
rect -5752 -13332 -5732 -13268
rect -5836 -13348 -5732 -13332
rect -5836 -13412 -5816 -13348
rect -5752 -13412 -5732 -13348
rect -5836 -13428 -5732 -13412
rect -5836 -13492 -5816 -13428
rect -5752 -13492 -5732 -13428
rect -5836 -13508 -5732 -13492
rect -5836 -13572 -5816 -13508
rect -5752 -13572 -5732 -13508
rect -5836 -13588 -5732 -13572
rect -5836 -13652 -5816 -13588
rect -5752 -13652 -5732 -13588
rect -5836 -13668 -5732 -13652
rect -5836 -13732 -5816 -13668
rect -5752 -13732 -5732 -13668
rect -5836 -13748 -5732 -13732
rect -5836 -13812 -5816 -13748
rect -5752 -13812 -5732 -13748
rect -5836 -13828 -5732 -13812
rect -5836 -13892 -5816 -13828
rect -5752 -13892 -5732 -13828
rect -5836 -13908 -5732 -13892
rect -5836 -13972 -5816 -13908
rect -5752 -13972 -5732 -13908
rect -5836 -13988 -5732 -13972
rect -5836 -14052 -5816 -13988
rect -5752 -14052 -5732 -13988
rect -5836 -14068 -5732 -14052
rect -5836 -14132 -5816 -14068
rect -5752 -14132 -5732 -14068
rect -5836 -14148 -5732 -14132
rect -5836 -14212 -5816 -14148
rect -5752 -14212 -5732 -14148
rect -5836 -14228 -5732 -14212
rect -5836 -14292 -5816 -14228
rect -5752 -14292 -5732 -14228
rect -5836 -14308 -5732 -14292
rect -5836 -14372 -5816 -14308
rect -5752 -14372 -5732 -14308
rect -5836 -14388 -5732 -14372
rect -5836 -14452 -5816 -14388
rect -5752 -14452 -5732 -14388
rect -5836 -14468 -5732 -14452
rect -5836 -14532 -5816 -14468
rect -5752 -14532 -5732 -14468
rect -5836 -14548 -5732 -14532
rect -5836 -14612 -5816 -14548
rect -5752 -14612 -5732 -14548
rect -5836 -14628 -5732 -14612
rect -5836 -14692 -5816 -14628
rect -5752 -14692 -5732 -14628
rect -5836 -14708 -5732 -14692
rect -5836 -14772 -5816 -14708
rect -5752 -14772 -5732 -14708
rect -5836 -14788 -5732 -14772
rect -5836 -14852 -5816 -14788
rect -5752 -14852 -5732 -14788
rect -5836 -14868 -5732 -14852
rect -5836 -14932 -5816 -14868
rect -5752 -14932 -5732 -14868
rect -5836 -14948 -5732 -14932
rect -5836 -15012 -5816 -14948
rect -5752 -15012 -5732 -14948
rect -5836 -15028 -5732 -15012
rect -5836 -15092 -5816 -15028
rect -5752 -15092 -5732 -15028
rect -5836 -15108 -5732 -15092
rect -5836 -15172 -5816 -15108
rect -5752 -15172 -5732 -15108
rect -5836 -15188 -5732 -15172
rect -5836 -15252 -5816 -15188
rect -5752 -15252 -5732 -15188
rect -5836 -15268 -5732 -15252
rect -5836 -15332 -5816 -15268
rect -5752 -15332 -5732 -15268
rect -5836 -15348 -5732 -15332
rect -5836 -15412 -5816 -15348
rect -5752 -15412 -5732 -15348
rect -5836 -15428 -5732 -15412
rect -5836 -15492 -5816 -15428
rect -5752 -15492 -5732 -15428
rect -5836 -15508 -5732 -15492
rect -5836 -15572 -5816 -15508
rect -5752 -15572 -5732 -15508
rect -5836 -15588 -5732 -15572
rect -5836 -15652 -5816 -15588
rect -5752 -15652 -5732 -15588
rect -5836 -15668 -5732 -15652
rect -5836 -15732 -5816 -15668
rect -5752 -15732 -5732 -15668
rect -5836 -15748 -5732 -15732
rect -11448 -16108 -11344 -15812
rect -17060 -16188 -16956 -16172
rect -17060 -16252 -17040 -16188
rect -16976 -16252 -16956 -16188
rect -17060 -16268 -16956 -16252
rect -17060 -16332 -17040 -16268
rect -16976 -16332 -16956 -16268
rect -17060 -16348 -16956 -16332
rect -17060 -16412 -17040 -16348
rect -16976 -16412 -16956 -16348
rect -17060 -16428 -16956 -16412
rect -17060 -16492 -17040 -16428
rect -16976 -16492 -16956 -16428
rect -17060 -16508 -16956 -16492
rect -17060 -16572 -17040 -16508
rect -16976 -16572 -16956 -16508
rect -17060 -16588 -16956 -16572
rect -17060 -16652 -17040 -16588
rect -16976 -16652 -16956 -16588
rect -17060 -16668 -16956 -16652
rect -17060 -16732 -17040 -16668
rect -16976 -16732 -16956 -16668
rect -17060 -16748 -16956 -16732
rect -17060 -16812 -17040 -16748
rect -16976 -16812 -16956 -16748
rect -17060 -16828 -16956 -16812
rect -17060 -16892 -17040 -16828
rect -16976 -16892 -16956 -16828
rect -17060 -16908 -16956 -16892
rect -17060 -16972 -17040 -16908
rect -16976 -16972 -16956 -16908
rect -17060 -16988 -16956 -16972
rect -17060 -17052 -17040 -16988
rect -16976 -17052 -16956 -16988
rect -17060 -17068 -16956 -17052
rect -17060 -17132 -17040 -17068
rect -16976 -17132 -16956 -17068
rect -17060 -17148 -16956 -17132
rect -17060 -17212 -17040 -17148
rect -16976 -17212 -16956 -17148
rect -17060 -17228 -16956 -17212
rect -17060 -17292 -17040 -17228
rect -16976 -17292 -16956 -17228
rect -17060 -17308 -16956 -17292
rect -17060 -17372 -17040 -17308
rect -16976 -17372 -16956 -17308
rect -17060 -17388 -16956 -17372
rect -17060 -17452 -17040 -17388
rect -16976 -17452 -16956 -17388
rect -17060 -17468 -16956 -17452
rect -17060 -17532 -17040 -17468
rect -16976 -17532 -16956 -17468
rect -17060 -17548 -16956 -17532
rect -17060 -17612 -17040 -17548
rect -16976 -17612 -16956 -17548
rect -17060 -17628 -16956 -17612
rect -17060 -17692 -17040 -17628
rect -16976 -17692 -16956 -17628
rect -17060 -17708 -16956 -17692
rect -17060 -17772 -17040 -17708
rect -16976 -17772 -16956 -17708
rect -17060 -17788 -16956 -17772
rect -17060 -17852 -17040 -17788
rect -16976 -17852 -16956 -17788
rect -17060 -17868 -16956 -17852
rect -17060 -17932 -17040 -17868
rect -16976 -17932 -16956 -17868
rect -17060 -17948 -16956 -17932
rect -17060 -18012 -17040 -17948
rect -16976 -18012 -16956 -17948
rect -17060 -18028 -16956 -18012
rect -17060 -18092 -17040 -18028
rect -16976 -18092 -16956 -18028
rect -17060 -18108 -16956 -18092
rect -17060 -18172 -17040 -18108
rect -16976 -18172 -16956 -18108
rect -17060 -18188 -16956 -18172
rect -17060 -18252 -17040 -18188
rect -16976 -18252 -16956 -18188
rect -17060 -18268 -16956 -18252
rect -17060 -18332 -17040 -18268
rect -16976 -18332 -16956 -18268
rect -17060 -18348 -16956 -18332
rect -17060 -18412 -17040 -18348
rect -16976 -18412 -16956 -18348
rect -17060 -18428 -16956 -18412
rect -17060 -18492 -17040 -18428
rect -16976 -18492 -16956 -18428
rect -17060 -18508 -16956 -18492
rect -17060 -18572 -17040 -18508
rect -16976 -18572 -16956 -18508
rect -17060 -18588 -16956 -18572
rect -17060 -18652 -17040 -18588
rect -16976 -18652 -16956 -18588
rect -17060 -18668 -16956 -18652
rect -17060 -18732 -17040 -18668
rect -16976 -18732 -16956 -18668
rect -17060 -18748 -16956 -18732
rect -17060 -18812 -17040 -18748
rect -16976 -18812 -16956 -18748
rect -17060 -18828 -16956 -18812
rect -17060 -18892 -17040 -18828
rect -16976 -18892 -16956 -18828
rect -17060 -18908 -16956 -18892
rect -17060 -18972 -17040 -18908
rect -16976 -18972 -16956 -18908
rect -17060 -18988 -16956 -18972
rect -17060 -19052 -17040 -18988
rect -16976 -19052 -16956 -18988
rect -17060 -19068 -16956 -19052
rect -17060 -19132 -17040 -19068
rect -16976 -19132 -16956 -19068
rect -17060 -19148 -16956 -19132
rect -17060 -19212 -17040 -19148
rect -16976 -19212 -16956 -19148
rect -17060 -19228 -16956 -19212
rect -17060 -19292 -17040 -19228
rect -16976 -19292 -16956 -19228
rect -17060 -19308 -16956 -19292
rect -17060 -19372 -17040 -19308
rect -16976 -19372 -16956 -19308
rect -17060 -19388 -16956 -19372
rect -17060 -19452 -17040 -19388
rect -16976 -19452 -16956 -19388
rect -17060 -19468 -16956 -19452
rect -17060 -19532 -17040 -19468
rect -16976 -19532 -16956 -19468
rect -17060 -19548 -16956 -19532
rect -17060 -19612 -17040 -19548
rect -16976 -19612 -16956 -19548
rect -17060 -19628 -16956 -19612
rect -17060 -19692 -17040 -19628
rect -16976 -19692 -16956 -19628
rect -17060 -19708 -16956 -19692
rect -17060 -19772 -17040 -19708
rect -16976 -19772 -16956 -19708
rect -17060 -19788 -16956 -19772
rect -17060 -19852 -17040 -19788
rect -16976 -19852 -16956 -19788
rect -17060 -19868 -16956 -19852
rect -17060 -19932 -17040 -19868
rect -16976 -19932 -16956 -19868
rect -17060 -19948 -16956 -19932
rect -17060 -20012 -17040 -19948
rect -16976 -20012 -16956 -19948
rect -17060 -20028 -16956 -20012
rect -17060 -20092 -17040 -20028
rect -16976 -20092 -16956 -20028
rect -17060 -20108 -16956 -20092
rect -17060 -20172 -17040 -20108
rect -16976 -20172 -16956 -20108
rect -17060 -20188 -16956 -20172
rect -17060 -20252 -17040 -20188
rect -16976 -20252 -16956 -20188
rect -17060 -20268 -16956 -20252
rect -17060 -20332 -17040 -20268
rect -16976 -20332 -16956 -20268
rect -17060 -20348 -16956 -20332
rect -17060 -20412 -17040 -20348
rect -16976 -20412 -16956 -20348
rect -17060 -20428 -16956 -20412
rect -17060 -20492 -17040 -20428
rect -16976 -20492 -16956 -20428
rect -17060 -20508 -16956 -20492
rect -17060 -20572 -17040 -20508
rect -16976 -20572 -16956 -20508
rect -17060 -20588 -16956 -20572
rect -17060 -20652 -17040 -20588
rect -16976 -20652 -16956 -20588
rect -17060 -20668 -16956 -20652
rect -17060 -20732 -17040 -20668
rect -16976 -20732 -16956 -20668
rect -17060 -20748 -16956 -20732
rect -17060 -20812 -17040 -20748
rect -16976 -20812 -16956 -20748
rect -17060 -20828 -16956 -20812
rect -17060 -20892 -17040 -20828
rect -16976 -20892 -16956 -20828
rect -17060 -20908 -16956 -20892
rect -17060 -20972 -17040 -20908
rect -16976 -20972 -16956 -20908
rect -17060 -20988 -16956 -20972
rect -17060 -21052 -17040 -20988
rect -16976 -21052 -16956 -20988
rect -17060 -21068 -16956 -21052
rect -22672 -21428 -22568 -21132
rect -28284 -21508 -28180 -21492
rect -28284 -21572 -28264 -21508
rect -28200 -21572 -28180 -21508
rect -28284 -21588 -28180 -21572
rect -28284 -21652 -28264 -21588
rect -28200 -21652 -28180 -21588
rect -28284 -21668 -28180 -21652
rect -28284 -21732 -28264 -21668
rect -28200 -21732 -28180 -21668
rect -28284 -21748 -28180 -21732
rect -28284 -21812 -28264 -21748
rect -28200 -21812 -28180 -21748
rect -28284 -21828 -28180 -21812
rect -28284 -21892 -28264 -21828
rect -28200 -21892 -28180 -21828
rect -28284 -21908 -28180 -21892
rect -28284 -21972 -28264 -21908
rect -28200 -21972 -28180 -21908
rect -28284 -21988 -28180 -21972
rect -28284 -22052 -28264 -21988
rect -28200 -22052 -28180 -21988
rect -28284 -22068 -28180 -22052
rect -28284 -22132 -28264 -22068
rect -28200 -22132 -28180 -22068
rect -28284 -22148 -28180 -22132
rect -28284 -22212 -28264 -22148
rect -28200 -22212 -28180 -22148
rect -28284 -22228 -28180 -22212
rect -28284 -22292 -28264 -22228
rect -28200 -22292 -28180 -22228
rect -28284 -22308 -28180 -22292
rect -28284 -22372 -28264 -22308
rect -28200 -22372 -28180 -22308
rect -28284 -22388 -28180 -22372
rect -28284 -22452 -28264 -22388
rect -28200 -22452 -28180 -22388
rect -28284 -22468 -28180 -22452
rect -28284 -22532 -28264 -22468
rect -28200 -22532 -28180 -22468
rect -28284 -22548 -28180 -22532
rect -28284 -22612 -28264 -22548
rect -28200 -22612 -28180 -22548
rect -28284 -22628 -28180 -22612
rect -28284 -22692 -28264 -22628
rect -28200 -22692 -28180 -22628
rect -28284 -22708 -28180 -22692
rect -28284 -22772 -28264 -22708
rect -28200 -22772 -28180 -22708
rect -28284 -22788 -28180 -22772
rect -28284 -22852 -28264 -22788
rect -28200 -22852 -28180 -22788
rect -28284 -22868 -28180 -22852
rect -28284 -22932 -28264 -22868
rect -28200 -22932 -28180 -22868
rect -28284 -22948 -28180 -22932
rect -28284 -23012 -28264 -22948
rect -28200 -23012 -28180 -22948
rect -28284 -23028 -28180 -23012
rect -28284 -23092 -28264 -23028
rect -28200 -23092 -28180 -23028
rect -28284 -23108 -28180 -23092
rect -28284 -23172 -28264 -23108
rect -28200 -23172 -28180 -23108
rect -28284 -23188 -28180 -23172
rect -28284 -23252 -28264 -23188
rect -28200 -23252 -28180 -23188
rect -28284 -23268 -28180 -23252
rect -28284 -23332 -28264 -23268
rect -28200 -23332 -28180 -23268
rect -28284 -23348 -28180 -23332
rect -28284 -23412 -28264 -23348
rect -28200 -23412 -28180 -23348
rect -28284 -23428 -28180 -23412
rect -28284 -23492 -28264 -23428
rect -28200 -23492 -28180 -23428
rect -28284 -23508 -28180 -23492
rect -28284 -23572 -28264 -23508
rect -28200 -23572 -28180 -23508
rect -28284 -23588 -28180 -23572
rect -28284 -23652 -28264 -23588
rect -28200 -23652 -28180 -23588
rect -28284 -23668 -28180 -23652
rect -28284 -23732 -28264 -23668
rect -28200 -23732 -28180 -23668
rect -28284 -23748 -28180 -23732
rect -28284 -23812 -28264 -23748
rect -28200 -23812 -28180 -23748
rect -28284 -23828 -28180 -23812
rect -28284 -23892 -28264 -23828
rect -28200 -23892 -28180 -23828
rect -28284 -23908 -28180 -23892
rect -28284 -23972 -28264 -23908
rect -28200 -23972 -28180 -23908
rect -28284 -23988 -28180 -23972
rect -28284 -24052 -28264 -23988
rect -28200 -24052 -28180 -23988
rect -28284 -24068 -28180 -24052
rect -28284 -24132 -28264 -24068
rect -28200 -24132 -28180 -24068
rect -28284 -24148 -28180 -24132
rect -28284 -24212 -28264 -24148
rect -28200 -24212 -28180 -24148
rect -28284 -24228 -28180 -24212
rect -28284 -24292 -28264 -24228
rect -28200 -24292 -28180 -24228
rect -28284 -24308 -28180 -24292
rect -28284 -24372 -28264 -24308
rect -28200 -24372 -28180 -24308
rect -28284 -24388 -28180 -24372
rect -28284 -24452 -28264 -24388
rect -28200 -24452 -28180 -24388
rect -28284 -24468 -28180 -24452
rect -28284 -24532 -28264 -24468
rect -28200 -24532 -28180 -24468
rect -28284 -24548 -28180 -24532
rect -28284 -24612 -28264 -24548
rect -28200 -24612 -28180 -24548
rect -28284 -24628 -28180 -24612
rect -28284 -24692 -28264 -24628
rect -28200 -24692 -28180 -24628
rect -28284 -24708 -28180 -24692
rect -28284 -24772 -28264 -24708
rect -28200 -24772 -28180 -24708
rect -28284 -24788 -28180 -24772
rect -28284 -24852 -28264 -24788
rect -28200 -24852 -28180 -24788
rect -28284 -24868 -28180 -24852
rect -28284 -24932 -28264 -24868
rect -28200 -24932 -28180 -24868
rect -28284 -24948 -28180 -24932
rect -28284 -25012 -28264 -24948
rect -28200 -25012 -28180 -24948
rect -28284 -25028 -28180 -25012
rect -28284 -25092 -28264 -25028
rect -28200 -25092 -28180 -25028
rect -28284 -25108 -28180 -25092
rect -28284 -25172 -28264 -25108
rect -28200 -25172 -28180 -25108
rect -28284 -25188 -28180 -25172
rect -28284 -25252 -28264 -25188
rect -28200 -25252 -28180 -25188
rect -28284 -25268 -28180 -25252
rect -28284 -25332 -28264 -25268
rect -28200 -25332 -28180 -25268
rect -28284 -25348 -28180 -25332
rect -28284 -25412 -28264 -25348
rect -28200 -25412 -28180 -25348
rect -28284 -25428 -28180 -25412
rect -28284 -25492 -28264 -25428
rect -28200 -25492 -28180 -25428
rect -28284 -25508 -28180 -25492
rect -28284 -25572 -28264 -25508
rect -28200 -25572 -28180 -25508
rect -28284 -25588 -28180 -25572
rect -28284 -25652 -28264 -25588
rect -28200 -25652 -28180 -25588
rect -28284 -25668 -28180 -25652
rect -28284 -25732 -28264 -25668
rect -28200 -25732 -28180 -25668
rect -28284 -25748 -28180 -25732
rect -28284 -25812 -28264 -25748
rect -28200 -25812 -28180 -25748
rect -28284 -25828 -28180 -25812
rect -28284 -25892 -28264 -25828
rect -28200 -25892 -28180 -25828
rect -28284 -25908 -28180 -25892
rect -28284 -25972 -28264 -25908
rect -28200 -25972 -28180 -25908
rect -28284 -25988 -28180 -25972
rect -28284 -26052 -28264 -25988
rect -28200 -26052 -28180 -25988
rect -28284 -26068 -28180 -26052
rect -28284 -26132 -28264 -26068
rect -28200 -26132 -28180 -26068
rect -28284 -26148 -28180 -26132
rect -28284 -26212 -28264 -26148
rect -28200 -26212 -28180 -26148
rect -28284 -26228 -28180 -26212
rect -28284 -26292 -28264 -26228
rect -28200 -26292 -28180 -26228
rect -28284 -26308 -28180 -26292
rect -28284 -26372 -28264 -26308
rect -28200 -26372 -28180 -26308
rect -28284 -26388 -28180 -26372
rect -33896 -26748 -33792 -26452
rect -39085 -26828 -34163 -26799
rect -39085 -31692 -39056 -26828
rect -34192 -31692 -34163 -26828
rect -39085 -31721 -34163 -31692
rect -33896 -26812 -33876 -26748
rect -33812 -26812 -33792 -26748
rect -31064 -26799 -30960 -26401
rect -28284 -26452 -28264 -26388
rect -28200 -26452 -28180 -26388
rect -27861 -21508 -22939 -21479
rect -27861 -26372 -27832 -21508
rect -22968 -26372 -22939 -21508
rect -27861 -26401 -22939 -26372
rect -22672 -21492 -22652 -21428
rect -22588 -21492 -22568 -21428
rect -19840 -21479 -19736 -21081
rect -17060 -21132 -17040 -21068
rect -16976 -21132 -16956 -21068
rect -16637 -16188 -11715 -16159
rect -16637 -21052 -16608 -16188
rect -11744 -21052 -11715 -16188
rect -16637 -21081 -11715 -21052
rect -11448 -16172 -11428 -16108
rect -11364 -16172 -11344 -16108
rect -8616 -16159 -8512 -15761
rect -5836 -15812 -5816 -15748
rect -5752 -15812 -5732 -15748
rect -5413 -10868 -491 -10839
rect -5413 -15732 -5384 -10868
rect -520 -15732 -491 -10868
rect -5413 -15761 -491 -15732
rect -224 -10852 -204 -10788
rect -140 -10852 -120 -10788
rect 2608 -10839 2712 -10441
rect 5388 -10492 5408 -10428
rect 5472 -10492 5492 -10428
rect 5811 -5548 10733 -5519
rect 5811 -10412 5840 -5548
rect 10704 -10412 10733 -5548
rect 5811 -10441 10733 -10412
rect 11000 -5532 11020 -5468
rect 11084 -5532 11104 -5468
rect 13832 -5519 13936 -5121
rect 16612 -5172 16632 -5108
rect 16696 -5172 16716 -5108
rect 17035 -228 21957 -199
rect 17035 -5092 17064 -228
rect 21928 -5092 21957 -228
rect 17035 -5121 21957 -5092
rect 22224 -212 22244 -148
rect 22308 -212 22328 -148
rect 25056 -199 25160 199
rect 27836 148 27856 212
rect 27920 148 27940 212
rect 28259 5092 33181 5121
rect 28259 228 28288 5092
rect 33152 228 33181 5092
rect 28259 199 33181 228
rect 33448 5108 33468 5172
rect 33532 5108 33552 5172
rect 36280 5121 36384 5519
rect 39060 5468 39080 5532
rect 39144 5468 39164 5532
rect 39060 5172 39164 5468
rect 33448 5092 33552 5108
rect 33448 5028 33468 5092
rect 33532 5028 33552 5092
rect 33448 5012 33552 5028
rect 33448 4948 33468 5012
rect 33532 4948 33552 5012
rect 33448 4932 33552 4948
rect 33448 4868 33468 4932
rect 33532 4868 33552 4932
rect 33448 4852 33552 4868
rect 33448 4788 33468 4852
rect 33532 4788 33552 4852
rect 33448 4772 33552 4788
rect 33448 4708 33468 4772
rect 33532 4708 33552 4772
rect 33448 4692 33552 4708
rect 33448 4628 33468 4692
rect 33532 4628 33552 4692
rect 33448 4612 33552 4628
rect 33448 4548 33468 4612
rect 33532 4548 33552 4612
rect 33448 4532 33552 4548
rect 33448 4468 33468 4532
rect 33532 4468 33552 4532
rect 33448 4452 33552 4468
rect 33448 4388 33468 4452
rect 33532 4388 33552 4452
rect 33448 4372 33552 4388
rect 33448 4308 33468 4372
rect 33532 4308 33552 4372
rect 33448 4292 33552 4308
rect 33448 4228 33468 4292
rect 33532 4228 33552 4292
rect 33448 4212 33552 4228
rect 33448 4148 33468 4212
rect 33532 4148 33552 4212
rect 33448 4132 33552 4148
rect 33448 4068 33468 4132
rect 33532 4068 33552 4132
rect 33448 4052 33552 4068
rect 33448 3988 33468 4052
rect 33532 3988 33552 4052
rect 33448 3972 33552 3988
rect 33448 3908 33468 3972
rect 33532 3908 33552 3972
rect 33448 3892 33552 3908
rect 33448 3828 33468 3892
rect 33532 3828 33552 3892
rect 33448 3812 33552 3828
rect 33448 3748 33468 3812
rect 33532 3748 33552 3812
rect 33448 3732 33552 3748
rect 33448 3668 33468 3732
rect 33532 3668 33552 3732
rect 33448 3652 33552 3668
rect 33448 3588 33468 3652
rect 33532 3588 33552 3652
rect 33448 3572 33552 3588
rect 33448 3508 33468 3572
rect 33532 3508 33552 3572
rect 33448 3492 33552 3508
rect 33448 3428 33468 3492
rect 33532 3428 33552 3492
rect 33448 3412 33552 3428
rect 33448 3348 33468 3412
rect 33532 3348 33552 3412
rect 33448 3332 33552 3348
rect 33448 3268 33468 3332
rect 33532 3268 33552 3332
rect 33448 3252 33552 3268
rect 33448 3188 33468 3252
rect 33532 3188 33552 3252
rect 33448 3172 33552 3188
rect 33448 3108 33468 3172
rect 33532 3108 33552 3172
rect 33448 3092 33552 3108
rect 33448 3028 33468 3092
rect 33532 3028 33552 3092
rect 33448 3012 33552 3028
rect 33448 2948 33468 3012
rect 33532 2948 33552 3012
rect 33448 2932 33552 2948
rect 33448 2868 33468 2932
rect 33532 2868 33552 2932
rect 33448 2852 33552 2868
rect 33448 2788 33468 2852
rect 33532 2788 33552 2852
rect 33448 2772 33552 2788
rect 33448 2708 33468 2772
rect 33532 2708 33552 2772
rect 33448 2692 33552 2708
rect 33448 2628 33468 2692
rect 33532 2628 33552 2692
rect 33448 2612 33552 2628
rect 33448 2548 33468 2612
rect 33532 2548 33552 2612
rect 33448 2532 33552 2548
rect 33448 2468 33468 2532
rect 33532 2468 33552 2532
rect 33448 2452 33552 2468
rect 33448 2388 33468 2452
rect 33532 2388 33552 2452
rect 33448 2372 33552 2388
rect 33448 2308 33468 2372
rect 33532 2308 33552 2372
rect 33448 2292 33552 2308
rect 33448 2228 33468 2292
rect 33532 2228 33552 2292
rect 33448 2212 33552 2228
rect 33448 2148 33468 2212
rect 33532 2148 33552 2212
rect 33448 2132 33552 2148
rect 33448 2068 33468 2132
rect 33532 2068 33552 2132
rect 33448 2052 33552 2068
rect 33448 1988 33468 2052
rect 33532 1988 33552 2052
rect 33448 1972 33552 1988
rect 33448 1908 33468 1972
rect 33532 1908 33552 1972
rect 33448 1892 33552 1908
rect 33448 1828 33468 1892
rect 33532 1828 33552 1892
rect 33448 1812 33552 1828
rect 33448 1748 33468 1812
rect 33532 1748 33552 1812
rect 33448 1732 33552 1748
rect 33448 1668 33468 1732
rect 33532 1668 33552 1732
rect 33448 1652 33552 1668
rect 33448 1588 33468 1652
rect 33532 1588 33552 1652
rect 33448 1572 33552 1588
rect 33448 1508 33468 1572
rect 33532 1508 33552 1572
rect 33448 1492 33552 1508
rect 33448 1428 33468 1492
rect 33532 1428 33552 1492
rect 33448 1412 33552 1428
rect 33448 1348 33468 1412
rect 33532 1348 33552 1412
rect 33448 1332 33552 1348
rect 33448 1268 33468 1332
rect 33532 1268 33552 1332
rect 33448 1252 33552 1268
rect 33448 1188 33468 1252
rect 33532 1188 33552 1252
rect 33448 1172 33552 1188
rect 33448 1108 33468 1172
rect 33532 1108 33552 1172
rect 33448 1092 33552 1108
rect 33448 1028 33468 1092
rect 33532 1028 33552 1092
rect 33448 1012 33552 1028
rect 33448 948 33468 1012
rect 33532 948 33552 1012
rect 33448 932 33552 948
rect 33448 868 33468 932
rect 33532 868 33552 932
rect 33448 852 33552 868
rect 33448 788 33468 852
rect 33532 788 33552 852
rect 33448 772 33552 788
rect 33448 708 33468 772
rect 33532 708 33552 772
rect 33448 692 33552 708
rect 33448 628 33468 692
rect 33532 628 33552 692
rect 33448 612 33552 628
rect 33448 548 33468 612
rect 33532 548 33552 612
rect 33448 532 33552 548
rect 33448 468 33468 532
rect 33532 468 33552 532
rect 33448 452 33552 468
rect 33448 388 33468 452
rect 33532 388 33552 452
rect 33448 372 33552 388
rect 33448 308 33468 372
rect 33532 308 33552 372
rect 33448 292 33552 308
rect 33448 228 33468 292
rect 33532 228 33552 292
rect 33448 212 33552 228
rect 27836 -148 27940 148
rect 22224 -228 22328 -212
rect 22224 -292 22244 -228
rect 22308 -292 22328 -228
rect 22224 -308 22328 -292
rect 22224 -372 22244 -308
rect 22308 -372 22328 -308
rect 22224 -388 22328 -372
rect 22224 -452 22244 -388
rect 22308 -452 22328 -388
rect 22224 -468 22328 -452
rect 22224 -532 22244 -468
rect 22308 -532 22328 -468
rect 22224 -548 22328 -532
rect 22224 -612 22244 -548
rect 22308 -612 22328 -548
rect 22224 -628 22328 -612
rect 22224 -692 22244 -628
rect 22308 -692 22328 -628
rect 22224 -708 22328 -692
rect 22224 -772 22244 -708
rect 22308 -772 22328 -708
rect 22224 -788 22328 -772
rect 22224 -852 22244 -788
rect 22308 -852 22328 -788
rect 22224 -868 22328 -852
rect 22224 -932 22244 -868
rect 22308 -932 22328 -868
rect 22224 -948 22328 -932
rect 22224 -1012 22244 -948
rect 22308 -1012 22328 -948
rect 22224 -1028 22328 -1012
rect 22224 -1092 22244 -1028
rect 22308 -1092 22328 -1028
rect 22224 -1108 22328 -1092
rect 22224 -1172 22244 -1108
rect 22308 -1172 22328 -1108
rect 22224 -1188 22328 -1172
rect 22224 -1252 22244 -1188
rect 22308 -1252 22328 -1188
rect 22224 -1268 22328 -1252
rect 22224 -1332 22244 -1268
rect 22308 -1332 22328 -1268
rect 22224 -1348 22328 -1332
rect 22224 -1412 22244 -1348
rect 22308 -1412 22328 -1348
rect 22224 -1428 22328 -1412
rect 22224 -1492 22244 -1428
rect 22308 -1492 22328 -1428
rect 22224 -1508 22328 -1492
rect 22224 -1572 22244 -1508
rect 22308 -1572 22328 -1508
rect 22224 -1588 22328 -1572
rect 22224 -1652 22244 -1588
rect 22308 -1652 22328 -1588
rect 22224 -1668 22328 -1652
rect 22224 -1732 22244 -1668
rect 22308 -1732 22328 -1668
rect 22224 -1748 22328 -1732
rect 22224 -1812 22244 -1748
rect 22308 -1812 22328 -1748
rect 22224 -1828 22328 -1812
rect 22224 -1892 22244 -1828
rect 22308 -1892 22328 -1828
rect 22224 -1908 22328 -1892
rect 22224 -1972 22244 -1908
rect 22308 -1972 22328 -1908
rect 22224 -1988 22328 -1972
rect 22224 -2052 22244 -1988
rect 22308 -2052 22328 -1988
rect 22224 -2068 22328 -2052
rect 22224 -2132 22244 -2068
rect 22308 -2132 22328 -2068
rect 22224 -2148 22328 -2132
rect 22224 -2212 22244 -2148
rect 22308 -2212 22328 -2148
rect 22224 -2228 22328 -2212
rect 22224 -2292 22244 -2228
rect 22308 -2292 22328 -2228
rect 22224 -2308 22328 -2292
rect 22224 -2372 22244 -2308
rect 22308 -2372 22328 -2308
rect 22224 -2388 22328 -2372
rect 22224 -2452 22244 -2388
rect 22308 -2452 22328 -2388
rect 22224 -2468 22328 -2452
rect 22224 -2532 22244 -2468
rect 22308 -2532 22328 -2468
rect 22224 -2548 22328 -2532
rect 22224 -2612 22244 -2548
rect 22308 -2612 22328 -2548
rect 22224 -2628 22328 -2612
rect 22224 -2692 22244 -2628
rect 22308 -2692 22328 -2628
rect 22224 -2708 22328 -2692
rect 22224 -2772 22244 -2708
rect 22308 -2772 22328 -2708
rect 22224 -2788 22328 -2772
rect 22224 -2852 22244 -2788
rect 22308 -2852 22328 -2788
rect 22224 -2868 22328 -2852
rect 22224 -2932 22244 -2868
rect 22308 -2932 22328 -2868
rect 22224 -2948 22328 -2932
rect 22224 -3012 22244 -2948
rect 22308 -3012 22328 -2948
rect 22224 -3028 22328 -3012
rect 22224 -3092 22244 -3028
rect 22308 -3092 22328 -3028
rect 22224 -3108 22328 -3092
rect 22224 -3172 22244 -3108
rect 22308 -3172 22328 -3108
rect 22224 -3188 22328 -3172
rect 22224 -3252 22244 -3188
rect 22308 -3252 22328 -3188
rect 22224 -3268 22328 -3252
rect 22224 -3332 22244 -3268
rect 22308 -3332 22328 -3268
rect 22224 -3348 22328 -3332
rect 22224 -3412 22244 -3348
rect 22308 -3412 22328 -3348
rect 22224 -3428 22328 -3412
rect 22224 -3492 22244 -3428
rect 22308 -3492 22328 -3428
rect 22224 -3508 22328 -3492
rect 22224 -3572 22244 -3508
rect 22308 -3572 22328 -3508
rect 22224 -3588 22328 -3572
rect 22224 -3652 22244 -3588
rect 22308 -3652 22328 -3588
rect 22224 -3668 22328 -3652
rect 22224 -3732 22244 -3668
rect 22308 -3732 22328 -3668
rect 22224 -3748 22328 -3732
rect 22224 -3812 22244 -3748
rect 22308 -3812 22328 -3748
rect 22224 -3828 22328 -3812
rect 22224 -3892 22244 -3828
rect 22308 -3892 22328 -3828
rect 22224 -3908 22328 -3892
rect 22224 -3972 22244 -3908
rect 22308 -3972 22328 -3908
rect 22224 -3988 22328 -3972
rect 22224 -4052 22244 -3988
rect 22308 -4052 22328 -3988
rect 22224 -4068 22328 -4052
rect 22224 -4132 22244 -4068
rect 22308 -4132 22328 -4068
rect 22224 -4148 22328 -4132
rect 22224 -4212 22244 -4148
rect 22308 -4212 22328 -4148
rect 22224 -4228 22328 -4212
rect 22224 -4292 22244 -4228
rect 22308 -4292 22328 -4228
rect 22224 -4308 22328 -4292
rect 22224 -4372 22244 -4308
rect 22308 -4372 22328 -4308
rect 22224 -4388 22328 -4372
rect 22224 -4452 22244 -4388
rect 22308 -4452 22328 -4388
rect 22224 -4468 22328 -4452
rect 22224 -4532 22244 -4468
rect 22308 -4532 22328 -4468
rect 22224 -4548 22328 -4532
rect 22224 -4612 22244 -4548
rect 22308 -4612 22328 -4548
rect 22224 -4628 22328 -4612
rect 22224 -4692 22244 -4628
rect 22308 -4692 22328 -4628
rect 22224 -4708 22328 -4692
rect 22224 -4772 22244 -4708
rect 22308 -4772 22328 -4708
rect 22224 -4788 22328 -4772
rect 22224 -4852 22244 -4788
rect 22308 -4852 22328 -4788
rect 22224 -4868 22328 -4852
rect 22224 -4932 22244 -4868
rect 22308 -4932 22328 -4868
rect 22224 -4948 22328 -4932
rect 22224 -5012 22244 -4948
rect 22308 -5012 22328 -4948
rect 22224 -5028 22328 -5012
rect 22224 -5092 22244 -5028
rect 22308 -5092 22328 -5028
rect 22224 -5108 22328 -5092
rect 16612 -5468 16716 -5172
rect 11000 -5548 11104 -5532
rect 11000 -5612 11020 -5548
rect 11084 -5612 11104 -5548
rect 11000 -5628 11104 -5612
rect 11000 -5692 11020 -5628
rect 11084 -5692 11104 -5628
rect 11000 -5708 11104 -5692
rect 11000 -5772 11020 -5708
rect 11084 -5772 11104 -5708
rect 11000 -5788 11104 -5772
rect 11000 -5852 11020 -5788
rect 11084 -5852 11104 -5788
rect 11000 -5868 11104 -5852
rect 11000 -5932 11020 -5868
rect 11084 -5932 11104 -5868
rect 11000 -5948 11104 -5932
rect 11000 -6012 11020 -5948
rect 11084 -6012 11104 -5948
rect 11000 -6028 11104 -6012
rect 11000 -6092 11020 -6028
rect 11084 -6092 11104 -6028
rect 11000 -6108 11104 -6092
rect 11000 -6172 11020 -6108
rect 11084 -6172 11104 -6108
rect 11000 -6188 11104 -6172
rect 11000 -6252 11020 -6188
rect 11084 -6252 11104 -6188
rect 11000 -6268 11104 -6252
rect 11000 -6332 11020 -6268
rect 11084 -6332 11104 -6268
rect 11000 -6348 11104 -6332
rect 11000 -6412 11020 -6348
rect 11084 -6412 11104 -6348
rect 11000 -6428 11104 -6412
rect 11000 -6492 11020 -6428
rect 11084 -6492 11104 -6428
rect 11000 -6508 11104 -6492
rect 11000 -6572 11020 -6508
rect 11084 -6572 11104 -6508
rect 11000 -6588 11104 -6572
rect 11000 -6652 11020 -6588
rect 11084 -6652 11104 -6588
rect 11000 -6668 11104 -6652
rect 11000 -6732 11020 -6668
rect 11084 -6732 11104 -6668
rect 11000 -6748 11104 -6732
rect 11000 -6812 11020 -6748
rect 11084 -6812 11104 -6748
rect 11000 -6828 11104 -6812
rect 11000 -6892 11020 -6828
rect 11084 -6892 11104 -6828
rect 11000 -6908 11104 -6892
rect 11000 -6972 11020 -6908
rect 11084 -6972 11104 -6908
rect 11000 -6988 11104 -6972
rect 11000 -7052 11020 -6988
rect 11084 -7052 11104 -6988
rect 11000 -7068 11104 -7052
rect 11000 -7132 11020 -7068
rect 11084 -7132 11104 -7068
rect 11000 -7148 11104 -7132
rect 11000 -7212 11020 -7148
rect 11084 -7212 11104 -7148
rect 11000 -7228 11104 -7212
rect 11000 -7292 11020 -7228
rect 11084 -7292 11104 -7228
rect 11000 -7308 11104 -7292
rect 11000 -7372 11020 -7308
rect 11084 -7372 11104 -7308
rect 11000 -7388 11104 -7372
rect 11000 -7452 11020 -7388
rect 11084 -7452 11104 -7388
rect 11000 -7468 11104 -7452
rect 11000 -7532 11020 -7468
rect 11084 -7532 11104 -7468
rect 11000 -7548 11104 -7532
rect 11000 -7612 11020 -7548
rect 11084 -7612 11104 -7548
rect 11000 -7628 11104 -7612
rect 11000 -7692 11020 -7628
rect 11084 -7692 11104 -7628
rect 11000 -7708 11104 -7692
rect 11000 -7772 11020 -7708
rect 11084 -7772 11104 -7708
rect 11000 -7788 11104 -7772
rect 11000 -7852 11020 -7788
rect 11084 -7852 11104 -7788
rect 11000 -7868 11104 -7852
rect 11000 -7932 11020 -7868
rect 11084 -7932 11104 -7868
rect 11000 -7948 11104 -7932
rect 11000 -8012 11020 -7948
rect 11084 -8012 11104 -7948
rect 11000 -8028 11104 -8012
rect 11000 -8092 11020 -8028
rect 11084 -8092 11104 -8028
rect 11000 -8108 11104 -8092
rect 11000 -8172 11020 -8108
rect 11084 -8172 11104 -8108
rect 11000 -8188 11104 -8172
rect 11000 -8252 11020 -8188
rect 11084 -8252 11104 -8188
rect 11000 -8268 11104 -8252
rect 11000 -8332 11020 -8268
rect 11084 -8332 11104 -8268
rect 11000 -8348 11104 -8332
rect 11000 -8412 11020 -8348
rect 11084 -8412 11104 -8348
rect 11000 -8428 11104 -8412
rect 11000 -8492 11020 -8428
rect 11084 -8492 11104 -8428
rect 11000 -8508 11104 -8492
rect 11000 -8572 11020 -8508
rect 11084 -8572 11104 -8508
rect 11000 -8588 11104 -8572
rect 11000 -8652 11020 -8588
rect 11084 -8652 11104 -8588
rect 11000 -8668 11104 -8652
rect 11000 -8732 11020 -8668
rect 11084 -8732 11104 -8668
rect 11000 -8748 11104 -8732
rect 11000 -8812 11020 -8748
rect 11084 -8812 11104 -8748
rect 11000 -8828 11104 -8812
rect 11000 -8892 11020 -8828
rect 11084 -8892 11104 -8828
rect 11000 -8908 11104 -8892
rect 11000 -8972 11020 -8908
rect 11084 -8972 11104 -8908
rect 11000 -8988 11104 -8972
rect 11000 -9052 11020 -8988
rect 11084 -9052 11104 -8988
rect 11000 -9068 11104 -9052
rect 11000 -9132 11020 -9068
rect 11084 -9132 11104 -9068
rect 11000 -9148 11104 -9132
rect 11000 -9212 11020 -9148
rect 11084 -9212 11104 -9148
rect 11000 -9228 11104 -9212
rect 11000 -9292 11020 -9228
rect 11084 -9292 11104 -9228
rect 11000 -9308 11104 -9292
rect 11000 -9372 11020 -9308
rect 11084 -9372 11104 -9308
rect 11000 -9388 11104 -9372
rect 11000 -9452 11020 -9388
rect 11084 -9452 11104 -9388
rect 11000 -9468 11104 -9452
rect 11000 -9532 11020 -9468
rect 11084 -9532 11104 -9468
rect 11000 -9548 11104 -9532
rect 11000 -9612 11020 -9548
rect 11084 -9612 11104 -9548
rect 11000 -9628 11104 -9612
rect 11000 -9692 11020 -9628
rect 11084 -9692 11104 -9628
rect 11000 -9708 11104 -9692
rect 11000 -9772 11020 -9708
rect 11084 -9772 11104 -9708
rect 11000 -9788 11104 -9772
rect 11000 -9852 11020 -9788
rect 11084 -9852 11104 -9788
rect 11000 -9868 11104 -9852
rect 11000 -9932 11020 -9868
rect 11084 -9932 11104 -9868
rect 11000 -9948 11104 -9932
rect 11000 -10012 11020 -9948
rect 11084 -10012 11104 -9948
rect 11000 -10028 11104 -10012
rect 11000 -10092 11020 -10028
rect 11084 -10092 11104 -10028
rect 11000 -10108 11104 -10092
rect 11000 -10172 11020 -10108
rect 11084 -10172 11104 -10108
rect 11000 -10188 11104 -10172
rect 11000 -10252 11020 -10188
rect 11084 -10252 11104 -10188
rect 11000 -10268 11104 -10252
rect 11000 -10332 11020 -10268
rect 11084 -10332 11104 -10268
rect 11000 -10348 11104 -10332
rect 11000 -10412 11020 -10348
rect 11084 -10412 11104 -10348
rect 11000 -10428 11104 -10412
rect 5388 -10788 5492 -10492
rect -224 -10868 -120 -10852
rect -224 -10932 -204 -10868
rect -140 -10932 -120 -10868
rect -224 -10948 -120 -10932
rect -224 -11012 -204 -10948
rect -140 -11012 -120 -10948
rect -224 -11028 -120 -11012
rect -224 -11092 -204 -11028
rect -140 -11092 -120 -11028
rect -224 -11108 -120 -11092
rect -224 -11172 -204 -11108
rect -140 -11172 -120 -11108
rect -224 -11188 -120 -11172
rect -224 -11252 -204 -11188
rect -140 -11252 -120 -11188
rect -224 -11268 -120 -11252
rect -224 -11332 -204 -11268
rect -140 -11332 -120 -11268
rect -224 -11348 -120 -11332
rect -224 -11412 -204 -11348
rect -140 -11412 -120 -11348
rect -224 -11428 -120 -11412
rect -224 -11492 -204 -11428
rect -140 -11492 -120 -11428
rect -224 -11508 -120 -11492
rect -224 -11572 -204 -11508
rect -140 -11572 -120 -11508
rect -224 -11588 -120 -11572
rect -224 -11652 -204 -11588
rect -140 -11652 -120 -11588
rect -224 -11668 -120 -11652
rect -224 -11732 -204 -11668
rect -140 -11732 -120 -11668
rect -224 -11748 -120 -11732
rect -224 -11812 -204 -11748
rect -140 -11812 -120 -11748
rect -224 -11828 -120 -11812
rect -224 -11892 -204 -11828
rect -140 -11892 -120 -11828
rect -224 -11908 -120 -11892
rect -224 -11972 -204 -11908
rect -140 -11972 -120 -11908
rect -224 -11988 -120 -11972
rect -224 -12052 -204 -11988
rect -140 -12052 -120 -11988
rect -224 -12068 -120 -12052
rect -224 -12132 -204 -12068
rect -140 -12132 -120 -12068
rect -224 -12148 -120 -12132
rect -224 -12212 -204 -12148
rect -140 -12212 -120 -12148
rect -224 -12228 -120 -12212
rect -224 -12292 -204 -12228
rect -140 -12292 -120 -12228
rect -224 -12308 -120 -12292
rect -224 -12372 -204 -12308
rect -140 -12372 -120 -12308
rect -224 -12388 -120 -12372
rect -224 -12452 -204 -12388
rect -140 -12452 -120 -12388
rect -224 -12468 -120 -12452
rect -224 -12532 -204 -12468
rect -140 -12532 -120 -12468
rect -224 -12548 -120 -12532
rect -224 -12612 -204 -12548
rect -140 -12612 -120 -12548
rect -224 -12628 -120 -12612
rect -224 -12692 -204 -12628
rect -140 -12692 -120 -12628
rect -224 -12708 -120 -12692
rect -224 -12772 -204 -12708
rect -140 -12772 -120 -12708
rect -224 -12788 -120 -12772
rect -224 -12852 -204 -12788
rect -140 -12852 -120 -12788
rect -224 -12868 -120 -12852
rect -224 -12932 -204 -12868
rect -140 -12932 -120 -12868
rect -224 -12948 -120 -12932
rect -224 -13012 -204 -12948
rect -140 -13012 -120 -12948
rect -224 -13028 -120 -13012
rect -224 -13092 -204 -13028
rect -140 -13092 -120 -13028
rect -224 -13108 -120 -13092
rect -224 -13172 -204 -13108
rect -140 -13172 -120 -13108
rect -224 -13188 -120 -13172
rect -224 -13252 -204 -13188
rect -140 -13252 -120 -13188
rect -224 -13268 -120 -13252
rect -224 -13332 -204 -13268
rect -140 -13332 -120 -13268
rect -224 -13348 -120 -13332
rect -224 -13412 -204 -13348
rect -140 -13412 -120 -13348
rect -224 -13428 -120 -13412
rect -224 -13492 -204 -13428
rect -140 -13492 -120 -13428
rect -224 -13508 -120 -13492
rect -224 -13572 -204 -13508
rect -140 -13572 -120 -13508
rect -224 -13588 -120 -13572
rect -224 -13652 -204 -13588
rect -140 -13652 -120 -13588
rect -224 -13668 -120 -13652
rect -224 -13732 -204 -13668
rect -140 -13732 -120 -13668
rect -224 -13748 -120 -13732
rect -224 -13812 -204 -13748
rect -140 -13812 -120 -13748
rect -224 -13828 -120 -13812
rect -224 -13892 -204 -13828
rect -140 -13892 -120 -13828
rect -224 -13908 -120 -13892
rect -224 -13972 -204 -13908
rect -140 -13972 -120 -13908
rect -224 -13988 -120 -13972
rect -224 -14052 -204 -13988
rect -140 -14052 -120 -13988
rect -224 -14068 -120 -14052
rect -224 -14132 -204 -14068
rect -140 -14132 -120 -14068
rect -224 -14148 -120 -14132
rect -224 -14212 -204 -14148
rect -140 -14212 -120 -14148
rect -224 -14228 -120 -14212
rect -224 -14292 -204 -14228
rect -140 -14292 -120 -14228
rect -224 -14308 -120 -14292
rect -224 -14372 -204 -14308
rect -140 -14372 -120 -14308
rect -224 -14388 -120 -14372
rect -224 -14452 -204 -14388
rect -140 -14452 -120 -14388
rect -224 -14468 -120 -14452
rect -224 -14532 -204 -14468
rect -140 -14532 -120 -14468
rect -224 -14548 -120 -14532
rect -224 -14612 -204 -14548
rect -140 -14612 -120 -14548
rect -224 -14628 -120 -14612
rect -224 -14692 -204 -14628
rect -140 -14692 -120 -14628
rect -224 -14708 -120 -14692
rect -224 -14772 -204 -14708
rect -140 -14772 -120 -14708
rect -224 -14788 -120 -14772
rect -224 -14852 -204 -14788
rect -140 -14852 -120 -14788
rect -224 -14868 -120 -14852
rect -224 -14932 -204 -14868
rect -140 -14932 -120 -14868
rect -224 -14948 -120 -14932
rect -224 -15012 -204 -14948
rect -140 -15012 -120 -14948
rect -224 -15028 -120 -15012
rect -224 -15092 -204 -15028
rect -140 -15092 -120 -15028
rect -224 -15108 -120 -15092
rect -224 -15172 -204 -15108
rect -140 -15172 -120 -15108
rect -224 -15188 -120 -15172
rect -224 -15252 -204 -15188
rect -140 -15252 -120 -15188
rect -224 -15268 -120 -15252
rect -224 -15332 -204 -15268
rect -140 -15332 -120 -15268
rect -224 -15348 -120 -15332
rect -224 -15412 -204 -15348
rect -140 -15412 -120 -15348
rect -224 -15428 -120 -15412
rect -224 -15492 -204 -15428
rect -140 -15492 -120 -15428
rect -224 -15508 -120 -15492
rect -224 -15572 -204 -15508
rect -140 -15572 -120 -15508
rect -224 -15588 -120 -15572
rect -224 -15652 -204 -15588
rect -140 -15652 -120 -15588
rect -224 -15668 -120 -15652
rect -224 -15732 -204 -15668
rect -140 -15732 -120 -15668
rect -224 -15748 -120 -15732
rect -5836 -16108 -5732 -15812
rect -11448 -16188 -11344 -16172
rect -11448 -16252 -11428 -16188
rect -11364 -16252 -11344 -16188
rect -11448 -16268 -11344 -16252
rect -11448 -16332 -11428 -16268
rect -11364 -16332 -11344 -16268
rect -11448 -16348 -11344 -16332
rect -11448 -16412 -11428 -16348
rect -11364 -16412 -11344 -16348
rect -11448 -16428 -11344 -16412
rect -11448 -16492 -11428 -16428
rect -11364 -16492 -11344 -16428
rect -11448 -16508 -11344 -16492
rect -11448 -16572 -11428 -16508
rect -11364 -16572 -11344 -16508
rect -11448 -16588 -11344 -16572
rect -11448 -16652 -11428 -16588
rect -11364 -16652 -11344 -16588
rect -11448 -16668 -11344 -16652
rect -11448 -16732 -11428 -16668
rect -11364 -16732 -11344 -16668
rect -11448 -16748 -11344 -16732
rect -11448 -16812 -11428 -16748
rect -11364 -16812 -11344 -16748
rect -11448 -16828 -11344 -16812
rect -11448 -16892 -11428 -16828
rect -11364 -16892 -11344 -16828
rect -11448 -16908 -11344 -16892
rect -11448 -16972 -11428 -16908
rect -11364 -16972 -11344 -16908
rect -11448 -16988 -11344 -16972
rect -11448 -17052 -11428 -16988
rect -11364 -17052 -11344 -16988
rect -11448 -17068 -11344 -17052
rect -11448 -17132 -11428 -17068
rect -11364 -17132 -11344 -17068
rect -11448 -17148 -11344 -17132
rect -11448 -17212 -11428 -17148
rect -11364 -17212 -11344 -17148
rect -11448 -17228 -11344 -17212
rect -11448 -17292 -11428 -17228
rect -11364 -17292 -11344 -17228
rect -11448 -17308 -11344 -17292
rect -11448 -17372 -11428 -17308
rect -11364 -17372 -11344 -17308
rect -11448 -17388 -11344 -17372
rect -11448 -17452 -11428 -17388
rect -11364 -17452 -11344 -17388
rect -11448 -17468 -11344 -17452
rect -11448 -17532 -11428 -17468
rect -11364 -17532 -11344 -17468
rect -11448 -17548 -11344 -17532
rect -11448 -17612 -11428 -17548
rect -11364 -17612 -11344 -17548
rect -11448 -17628 -11344 -17612
rect -11448 -17692 -11428 -17628
rect -11364 -17692 -11344 -17628
rect -11448 -17708 -11344 -17692
rect -11448 -17772 -11428 -17708
rect -11364 -17772 -11344 -17708
rect -11448 -17788 -11344 -17772
rect -11448 -17852 -11428 -17788
rect -11364 -17852 -11344 -17788
rect -11448 -17868 -11344 -17852
rect -11448 -17932 -11428 -17868
rect -11364 -17932 -11344 -17868
rect -11448 -17948 -11344 -17932
rect -11448 -18012 -11428 -17948
rect -11364 -18012 -11344 -17948
rect -11448 -18028 -11344 -18012
rect -11448 -18092 -11428 -18028
rect -11364 -18092 -11344 -18028
rect -11448 -18108 -11344 -18092
rect -11448 -18172 -11428 -18108
rect -11364 -18172 -11344 -18108
rect -11448 -18188 -11344 -18172
rect -11448 -18252 -11428 -18188
rect -11364 -18252 -11344 -18188
rect -11448 -18268 -11344 -18252
rect -11448 -18332 -11428 -18268
rect -11364 -18332 -11344 -18268
rect -11448 -18348 -11344 -18332
rect -11448 -18412 -11428 -18348
rect -11364 -18412 -11344 -18348
rect -11448 -18428 -11344 -18412
rect -11448 -18492 -11428 -18428
rect -11364 -18492 -11344 -18428
rect -11448 -18508 -11344 -18492
rect -11448 -18572 -11428 -18508
rect -11364 -18572 -11344 -18508
rect -11448 -18588 -11344 -18572
rect -11448 -18652 -11428 -18588
rect -11364 -18652 -11344 -18588
rect -11448 -18668 -11344 -18652
rect -11448 -18732 -11428 -18668
rect -11364 -18732 -11344 -18668
rect -11448 -18748 -11344 -18732
rect -11448 -18812 -11428 -18748
rect -11364 -18812 -11344 -18748
rect -11448 -18828 -11344 -18812
rect -11448 -18892 -11428 -18828
rect -11364 -18892 -11344 -18828
rect -11448 -18908 -11344 -18892
rect -11448 -18972 -11428 -18908
rect -11364 -18972 -11344 -18908
rect -11448 -18988 -11344 -18972
rect -11448 -19052 -11428 -18988
rect -11364 -19052 -11344 -18988
rect -11448 -19068 -11344 -19052
rect -11448 -19132 -11428 -19068
rect -11364 -19132 -11344 -19068
rect -11448 -19148 -11344 -19132
rect -11448 -19212 -11428 -19148
rect -11364 -19212 -11344 -19148
rect -11448 -19228 -11344 -19212
rect -11448 -19292 -11428 -19228
rect -11364 -19292 -11344 -19228
rect -11448 -19308 -11344 -19292
rect -11448 -19372 -11428 -19308
rect -11364 -19372 -11344 -19308
rect -11448 -19388 -11344 -19372
rect -11448 -19452 -11428 -19388
rect -11364 -19452 -11344 -19388
rect -11448 -19468 -11344 -19452
rect -11448 -19532 -11428 -19468
rect -11364 -19532 -11344 -19468
rect -11448 -19548 -11344 -19532
rect -11448 -19612 -11428 -19548
rect -11364 -19612 -11344 -19548
rect -11448 -19628 -11344 -19612
rect -11448 -19692 -11428 -19628
rect -11364 -19692 -11344 -19628
rect -11448 -19708 -11344 -19692
rect -11448 -19772 -11428 -19708
rect -11364 -19772 -11344 -19708
rect -11448 -19788 -11344 -19772
rect -11448 -19852 -11428 -19788
rect -11364 -19852 -11344 -19788
rect -11448 -19868 -11344 -19852
rect -11448 -19932 -11428 -19868
rect -11364 -19932 -11344 -19868
rect -11448 -19948 -11344 -19932
rect -11448 -20012 -11428 -19948
rect -11364 -20012 -11344 -19948
rect -11448 -20028 -11344 -20012
rect -11448 -20092 -11428 -20028
rect -11364 -20092 -11344 -20028
rect -11448 -20108 -11344 -20092
rect -11448 -20172 -11428 -20108
rect -11364 -20172 -11344 -20108
rect -11448 -20188 -11344 -20172
rect -11448 -20252 -11428 -20188
rect -11364 -20252 -11344 -20188
rect -11448 -20268 -11344 -20252
rect -11448 -20332 -11428 -20268
rect -11364 -20332 -11344 -20268
rect -11448 -20348 -11344 -20332
rect -11448 -20412 -11428 -20348
rect -11364 -20412 -11344 -20348
rect -11448 -20428 -11344 -20412
rect -11448 -20492 -11428 -20428
rect -11364 -20492 -11344 -20428
rect -11448 -20508 -11344 -20492
rect -11448 -20572 -11428 -20508
rect -11364 -20572 -11344 -20508
rect -11448 -20588 -11344 -20572
rect -11448 -20652 -11428 -20588
rect -11364 -20652 -11344 -20588
rect -11448 -20668 -11344 -20652
rect -11448 -20732 -11428 -20668
rect -11364 -20732 -11344 -20668
rect -11448 -20748 -11344 -20732
rect -11448 -20812 -11428 -20748
rect -11364 -20812 -11344 -20748
rect -11448 -20828 -11344 -20812
rect -11448 -20892 -11428 -20828
rect -11364 -20892 -11344 -20828
rect -11448 -20908 -11344 -20892
rect -11448 -20972 -11428 -20908
rect -11364 -20972 -11344 -20908
rect -11448 -20988 -11344 -20972
rect -11448 -21052 -11428 -20988
rect -11364 -21052 -11344 -20988
rect -11448 -21068 -11344 -21052
rect -17060 -21428 -16956 -21132
rect -22672 -21508 -22568 -21492
rect -22672 -21572 -22652 -21508
rect -22588 -21572 -22568 -21508
rect -22672 -21588 -22568 -21572
rect -22672 -21652 -22652 -21588
rect -22588 -21652 -22568 -21588
rect -22672 -21668 -22568 -21652
rect -22672 -21732 -22652 -21668
rect -22588 -21732 -22568 -21668
rect -22672 -21748 -22568 -21732
rect -22672 -21812 -22652 -21748
rect -22588 -21812 -22568 -21748
rect -22672 -21828 -22568 -21812
rect -22672 -21892 -22652 -21828
rect -22588 -21892 -22568 -21828
rect -22672 -21908 -22568 -21892
rect -22672 -21972 -22652 -21908
rect -22588 -21972 -22568 -21908
rect -22672 -21988 -22568 -21972
rect -22672 -22052 -22652 -21988
rect -22588 -22052 -22568 -21988
rect -22672 -22068 -22568 -22052
rect -22672 -22132 -22652 -22068
rect -22588 -22132 -22568 -22068
rect -22672 -22148 -22568 -22132
rect -22672 -22212 -22652 -22148
rect -22588 -22212 -22568 -22148
rect -22672 -22228 -22568 -22212
rect -22672 -22292 -22652 -22228
rect -22588 -22292 -22568 -22228
rect -22672 -22308 -22568 -22292
rect -22672 -22372 -22652 -22308
rect -22588 -22372 -22568 -22308
rect -22672 -22388 -22568 -22372
rect -22672 -22452 -22652 -22388
rect -22588 -22452 -22568 -22388
rect -22672 -22468 -22568 -22452
rect -22672 -22532 -22652 -22468
rect -22588 -22532 -22568 -22468
rect -22672 -22548 -22568 -22532
rect -22672 -22612 -22652 -22548
rect -22588 -22612 -22568 -22548
rect -22672 -22628 -22568 -22612
rect -22672 -22692 -22652 -22628
rect -22588 -22692 -22568 -22628
rect -22672 -22708 -22568 -22692
rect -22672 -22772 -22652 -22708
rect -22588 -22772 -22568 -22708
rect -22672 -22788 -22568 -22772
rect -22672 -22852 -22652 -22788
rect -22588 -22852 -22568 -22788
rect -22672 -22868 -22568 -22852
rect -22672 -22932 -22652 -22868
rect -22588 -22932 -22568 -22868
rect -22672 -22948 -22568 -22932
rect -22672 -23012 -22652 -22948
rect -22588 -23012 -22568 -22948
rect -22672 -23028 -22568 -23012
rect -22672 -23092 -22652 -23028
rect -22588 -23092 -22568 -23028
rect -22672 -23108 -22568 -23092
rect -22672 -23172 -22652 -23108
rect -22588 -23172 -22568 -23108
rect -22672 -23188 -22568 -23172
rect -22672 -23252 -22652 -23188
rect -22588 -23252 -22568 -23188
rect -22672 -23268 -22568 -23252
rect -22672 -23332 -22652 -23268
rect -22588 -23332 -22568 -23268
rect -22672 -23348 -22568 -23332
rect -22672 -23412 -22652 -23348
rect -22588 -23412 -22568 -23348
rect -22672 -23428 -22568 -23412
rect -22672 -23492 -22652 -23428
rect -22588 -23492 -22568 -23428
rect -22672 -23508 -22568 -23492
rect -22672 -23572 -22652 -23508
rect -22588 -23572 -22568 -23508
rect -22672 -23588 -22568 -23572
rect -22672 -23652 -22652 -23588
rect -22588 -23652 -22568 -23588
rect -22672 -23668 -22568 -23652
rect -22672 -23732 -22652 -23668
rect -22588 -23732 -22568 -23668
rect -22672 -23748 -22568 -23732
rect -22672 -23812 -22652 -23748
rect -22588 -23812 -22568 -23748
rect -22672 -23828 -22568 -23812
rect -22672 -23892 -22652 -23828
rect -22588 -23892 -22568 -23828
rect -22672 -23908 -22568 -23892
rect -22672 -23972 -22652 -23908
rect -22588 -23972 -22568 -23908
rect -22672 -23988 -22568 -23972
rect -22672 -24052 -22652 -23988
rect -22588 -24052 -22568 -23988
rect -22672 -24068 -22568 -24052
rect -22672 -24132 -22652 -24068
rect -22588 -24132 -22568 -24068
rect -22672 -24148 -22568 -24132
rect -22672 -24212 -22652 -24148
rect -22588 -24212 -22568 -24148
rect -22672 -24228 -22568 -24212
rect -22672 -24292 -22652 -24228
rect -22588 -24292 -22568 -24228
rect -22672 -24308 -22568 -24292
rect -22672 -24372 -22652 -24308
rect -22588 -24372 -22568 -24308
rect -22672 -24388 -22568 -24372
rect -22672 -24452 -22652 -24388
rect -22588 -24452 -22568 -24388
rect -22672 -24468 -22568 -24452
rect -22672 -24532 -22652 -24468
rect -22588 -24532 -22568 -24468
rect -22672 -24548 -22568 -24532
rect -22672 -24612 -22652 -24548
rect -22588 -24612 -22568 -24548
rect -22672 -24628 -22568 -24612
rect -22672 -24692 -22652 -24628
rect -22588 -24692 -22568 -24628
rect -22672 -24708 -22568 -24692
rect -22672 -24772 -22652 -24708
rect -22588 -24772 -22568 -24708
rect -22672 -24788 -22568 -24772
rect -22672 -24852 -22652 -24788
rect -22588 -24852 -22568 -24788
rect -22672 -24868 -22568 -24852
rect -22672 -24932 -22652 -24868
rect -22588 -24932 -22568 -24868
rect -22672 -24948 -22568 -24932
rect -22672 -25012 -22652 -24948
rect -22588 -25012 -22568 -24948
rect -22672 -25028 -22568 -25012
rect -22672 -25092 -22652 -25028
rect -22588 -25092 -22568 -25028
rect -22672 -25108 -22568 -25092
rect -22672 -25172 -22652 -25108
rect -22588 -25172 -22568 -25108
rect -22672 -25188 -22568 -25172
rect -22672 -25252 -22652 -25188
rect -22588 -25252 -22568 -25188
rect -22672 -25268 -22568 -25252
rect -22672 -25332 -22652 -25268
rect -22588 -25332 -22568 -25268
rect -22672 -25348 -22568 -25332
rect -22672 -25412 -22652 -25348
rect -22588 -25412 -22568 -25348
rect -22672 -25428 -22568 -25412
rect -22672 -25492 -22652 -25428
rect -22588 -25492 -22568 -25428
rect -22672 -25508 -22568 -25492
rect -22672 -25572 -22652 -25508
rect -22588 -25572 -22568 -25508
rect -22672 -25588 -22568 -25572
rect -22672 -25652 -22652 -25588
rect -22588 -25652 -22568 -25588
rect -22672 -25668 -22568 -25652
rect -22672 -25732 -22652 -25668
rect -22588 -25732 -22568 -25668
rect -22672 -25748 -22568 -25732
rect -22672 -25812 -22652 -25748
rect -22588 -25812 -22568 -25748
rect -22672 -25828 -22568 -25812
rect -22672 -25892 -22652 -25828
rect -22588 -25892 -22568 -25828
rect -22672 -25908 -22568 -25892
rect -22672 -25972 -22652 -25908
rect -22588 -25972 -22568 -25908
rect -22672 -25988 -22568 -25972
rect -22672 -26052 -22652 -25988
rect -22588 -26052 -22568 -25988
rect -22672 -26068 -22568 -26052
rect -22672 -26132 -22652 -26068
rect -22588 -26132 -22568 -26068
rect -22672 -26148 -22568 -26132
rect -22672 -26212 -22652 -26148
rect -22588 -26212 -22568 -26148
rect -22672 -26228 -22568 -26212
rect -22672 -26292 -22652 -26228
rect -22588 -26292 -22568 -26228
rect -22672 -26308 -22568 -26292
rect -22672 -26372 -22652 -26308
rect -22588 -26372 -22568 -26308
rect -22672 -26388 -22568 -26372
rect -28284 -26748 -28180 -26452
rect -33896 -26828 -33792 -26812
rect -33896 -26892 -33876 -26828
rect -33812 -26892 -33792 -26828
rect -33896 -26908 -33792 -26892
rect -33896 -26972 -33876 -26908
rect -33812 -26972 -33792 -26908
rect -33896 -26988 -33792 -26972
rect -33896 -27052 -33876 -26988
rect -33812 -27052 -33792 -26988
rect -33896 -27068 -33792 -27052
rect -33896 -27132 -33876 -27068
rect -33812 -27132 -33792 -27068
rect -33896 -27148 -33792 -27132
rect -33896 -27212 -33876 -27148
rect -33812 -27212 -33792 -27148
rect -33896 -27228 -33792 -27212
rect -33896 -27292 -33876 -27228
rect -33812 -27292 -33792 -27228
rect -33896 -27308 -33792 -27292
rect -33896 -27372 -33876 -27308
rect -33812 -27372 -33792 -27308
rect -33896 -27388 -33792 -27372
rect -33896 -27452 -33876 -27388
rect -33812 -27452 -33792 -27388
rect -33896 -27468 -33792 -27452
rect -33896 -27532 -33876 -27468
rect -33812 -27532 -33792 -27468
rect -33896 -27548 -33792 -27532
rect -33896 -27612 -33876 -27548
rect -33812 -27612 -33792 -27548
rect -33896 -27628 -33792 -27612
rect -33896 -27692 -33876 -27628
rect -33812 -27692 -33792 -27628
rect -33896 -27708 -33792 -27692
rect -33896 -27772 -33876 -27708
rect -33812 -27772 -33792 -27708
rect -33896 -27788 -33792 -27772
rect -33896 -27852 -33876 -27788
rect -33812 -27852 -33792 -27788
rect -33896 -27868 -33792 -27852
rect -33896 -27932 -33876 -27868
rect -33812 -27932 -33792 -27868
rect -33896 -27948 -33792 -27932
rect -33896 -28012 -33876 -27948
rect -33812 -28012 -33792 -27948
rect -33896 -28028 -33792 -28012
rect -33896 -28092 -33876 -28028
rect -33812 -28092 -33792 -28028
rect -33896 -28108 -33792 -28092
rect -33896 -28172 -33876 -28108
rect -33812 -28172 -33792 -28108
rect -33896 -28188 -33792 -28172
rect -33896 -28252 -33876 -28188
rect -33812 -28252 -33792 -28188
rect -33896 -28268 -33792 -28252
rect -33896 -28332 -33876 -28268
rect -33812 -28332 -33792 -28268
rect -33896 -28348 -33792 -28332
rect -33896 -28412 -33876 -28348
rect -33812 -28412 -33792 -28348
rect -33896 -28428 -33792 -28412
rect -33896 -28492 -33876 -28428
rect -33812 -28492 -33792 -28428
rect -33896 -28508 -33792 -28492
rect -33896 -28572 -33876 -28508
rect -33812 -28572 -33792 -28508
rect -33896 -28588 -33792 -28572
rect -33896 -28652 -33876 -28588
rect -33812 -28652 -33792 -28588
rect -33896 -28668 -33792 -28652
rect -33896 -28732 -33876 -28668
rect -33812 -28732 -33792 -28668
rect -33896 -28748 -33792 -28732
rect -33896 -28812 -33876 -28748
rect -33812 -28812 -33792 -28748
rect -33896 -28828 -33792 -28812
rect -33896 -28892 -33876 -28828
rect -33812 -28892 -33792 -28828
rect -33896 -28908 -33792 -28892
rect -33896 -28972 -33876 -28908
rect -33812 -28972 -33792 -28908
rect -33896 -28988 -33792 -28972
rect -33896 -29052 -33876 -28988
rect -33812 -29052 -33792 -28988
rect -33896 -29068 -33792 -29052
rect -33896 -29132 -33876 -29068
rect -33812 -29132 -33792 -29068
rect -33896 -29148 -33792 -29132
rect -33896 -29212 -33876 -29148
rect -33812 -29212 -33792 -29148
rect -33896 -29228 -33792 -29212
rect -33896 -29292 -33876 -29228
rect -33812 -29292 -33792 -29228
rect -33896 -29308 -33792 -29292
rect -33896 -29372 -33876 -29308
rect -33812 -29372 -33792 -29308
rect -33896 -29388 -33792 -29372
rect -33896 -29452 -33876 -29388
rect -33812 -29452 -33792 -29388
rect -33896 -29468 -33792 -29452
rect -33896 -29532 -33876 -29468
rect -33812 -29532 -33792 -29468
rect -33896 -29548 -33792 -29532
rect -33896 -29612 -33876 -29548
rect -33812 -29612 -33792 -29548
rect -33896 -29628 -33792 -29612
rect -33896 -29692 -33876 -29628
rect -33812 -29692 -33792 -29628
rect -33896 -29708 -33792 -29692
rect -33896 -29772 -33876 -29708
rect -33812 -29772 -33792 -29708
rect -33896 -29788 -33792 -29772
rect -33896 -29852 -33876 -29788
rect -33812 -29852 -33792 -29788
rect -33896 -29868 -33792 -29852
rect -33896 -29932 -33876 -29868
rect -33812 -29932 -33792 -29868
rect -33896 -29948 -33792 -29932
rect -33896 -30012 -33876 -29948
rect -33812 -30012 -33792 -29948
rect -33896 -30028 -33792 -30012
rect -33896 -30092 -33876 -30028
rect -33812 -30092 -33792 -30028
rect -33896 -30108 -33792 -30092
rect -33896 -30172 -33876 -30108
rect -33812 -30172 -33792 -30108
rect -33896 -30188 -33792 -30172
rect -33896 -30252 -33876 -30188
rect -33812 -30252 -33792 -30188
rect -33896 -30268 -33792 -30252
rect -33896 -30332 -33876 -30268
rect -33812 -30332 -33792 -30268
rect -33896 -30348 -33792 -30332
rect -33896 -30412 -33876 -30348
rect -33812 -30412 -33792 -30348
rect -33896 -30428 -33792 -30412
rect -33896 -30492 -33876 -30428
rect -33812 -30492 -33792 -30428
rect -33896 -30508 -33792 -30492
rect -33896 -30572 -33876 -30508
rect -33812 -30572 -33792 -30508
rect -33896 -30588 -33792 -30572
rect -33896 -30652 -33876 -30588
rect -33812 -30652 -33792 -30588
rect -33896 -30668 -33792 -30652
rect -33896 -30732 -33876 -30668
rect -33812 -30732 -33792 -30668
rect -33896 -30748 -33792 -30732
rect -33896 -30812 -33876 -30748
rect -33812 -30812 -33792 -30748
rect -33896 -30828 -33792 -30812
rect -33896 -30892 -33876 -30828
rect -33812 -30892 -33792 -30828
rect -33896 -30908 -33792 -30892
rect -33896 -30972 -33876 -30908
rect -33812 -30972 -33792 -30908
rect -33896 -30988 -33792 -30972
rect -33896 -31052 -33876 -30988
rect -33812 -31052 -33792 -30988
rect -33896 -31068 -33792 -31052
rect -33896 -31132 -33876 -31068
rect -33812 -31132 -33792 -31068
rect -33896 -31148 -33792 -31132
rect -33896 -31212 -33876 -31148
rect -33812 -31212 -33792 -31148
rect -33896 -31228 -33792 -31212
rect -33896 -31292 -33876 -31228
rect -33812 -31292 -33792 -31228
rect -33896 -31308 -33792 -31292
rect -33896 -31372 -33876 -31308
rect -33812 -31372 -33792 -31308
rect -33896 -31388 -33792 -31372
rect -33896 -31452 -33876 -31388
rect -33812 -31452 -33792 -31388
rect -33896 -31468 -33792 -31452
rect -33896 -31532 -33876 -31468
rect -33812 -31532 -33792 -31468
rect -33896 -31548 -33792 -31532
rect -33896 -31612 -33876 -31548
rect -33812 -31612 -33792 -31548
rect -33896 -31628 -33792 -31612
rect -33896 -31692 -33876 -31628
rect -33812 -31692 -33792 -31628
rect -33896 -31708 -33792 -31692
rect -36676 -32119 -36572 -31721
rect -33896 -31772 -33876 -31708
rect -33812 -31772 -33792 -31708
rect -33473 -26828 -28551 -26799
rect -33473 -31692 -33444 -26828
rect -28580 -31692 -28551 -26828
rect -33473 -31721 -28551 -31692
rect -28284 -26812 -28264 -26748
rect -28200 -26812 -28180 -26748
rect -25452 -26799 -25348 -26401
rect -22672 -26452 -22652 -26388
rect -22588 -26452 -22568 -26388
rect -22249 -21508 -17327 -21479
rect -22249 -26372 -22220 -21508
rect -17356 -26372 -17327 -21508
rect -22249 -26401 -17327 -26372
rect -17060 -21492 -17040 -21428
rect -16976 -21492 -16956 -21428
rect -14228 -21479 -14124 -21081
rect -11448 -21132 -11428 -21068
rect -11364 -21132 -11344 -21068
rect -11025 -16188 -6103 -16159
rect -11025 -21052 -10996 -16188
rect -6132 -21052 -6103 -16188
rect -11025 -21081 -6103 -21052
rect -5836 -16172 -5816 -16108
rect -5752 -16172 -5732 -16108
rect -3004 -16159 -2900 -15761
rect -224 -15812 -204 -15748
rect -140 -15812 -120 -15748
rect 199 -10868 5121 -10839
rect 199 -15732 228 -10868
rect 5092 -15732 5121 -10868
rect 199 -15761 5121 -15732
rect 5388 -10852 5408 -10788
rect 5472 -10852 5492 -10788
rect 8220 -10839 8324 -10441
rect 11000 -10492 11020 -10428
rect 11084 -10492 11104 -10428
rect 11423 -5548 16345 -5519
rect 11423 -10412 11452 -5548
rect 16316 -10412 16345 -5548
rect 11423 -10441 16345 -10412
rect 16612 -5532 16632 -5468
rect 16696 -5532 16716 -5468
rect 19444 -5519 19548 -5121
rect 22224 -5172 22244 -5108
rect 22308 -5172 22328 -5108
rect 22647 -228 27569 -199
rect 22647 -5092 22676 -228
rect 27540 -5092 27569 -228
rect 22647 -5121 27569 -5092
rect 27836 -212 27856 -148
rect 27920 -212 27940 -148
rect 30668 -199 30772 199
rect 33448 148 33468 212
rect 33532 148 33552 212
rect 33871 5092 38793 5121
rect 33871 228 33900 5092
rect 38764 228 38793 5092
rect 33871 199 38793 228
rect 39060 5108 39080 5172
rect 39144 5108 39164 5172
rect 39060 5092 39164 5108
rect 39060 5028 39080 5092
rect 39144 5028 39164 5092
rect 39060 5012 39164 5028
rect 39060 4948 39080 5012
rect 39144 4948 39164 5012
rect 39060 4932 39164 4948
rect 39060 4868 39080 4932
rect 39144 4868 39164 4932
rect 39060 4852 39164 4868
rect 39060 4788 39080 4852
rect 39144 4788 39164 4852
rect 39060 4772 39164 4788
rect 39060 4708 39080 4772
rect 39144 4708 39164 4772
rect 39060 4692 39164 4708
rect 39060 4628 39080 4692
rect 39144 4628 39164 4692
rect 39060 4612 39164 4628
rect 39060 4548 39080 4612
rect 39144 4548 39164 4612
rect 39060 4532 39164 4548
rect 39060 4468 39080 4532
rect 39144 4468 39164 4532
rect 39060 4452 39164 4468
rect 39060 4388 39080 4452
rect 39144 4388 39164 4452
rect 39060 4372 39164 4388
rect 39060 4308 39080 4372
rect 39144 4308 39164 4372
rect 39060 4292 39164 4308
rect 39060 4228 39080 4292
rect 39144 4228 39164 4292
rect 39060 4212 39164 4228
rect 39060 4148 39080 4212
rect 39144 4148 39164 4212
rect 39060 4132 39164 4148
rect 39060 4068 39080 4132
rect 39144 4068 39164 4132
rect 39060 4052 39164 4068
rect 39060 3988 39080 4052
rect 39144 3988 39164 4052
rect 39060 3972 39164 3988
rect 39060 3908 39080 3972
rect 39144 3908 39164 3972
rect 39060 3892 39164 3908
rect 39060 3828 39080 3892
rect 39144 3828 39164 3892
rect 39060 3812 39164 3828
rect 39060 3748 39080 3812
rect 39144 3748 39164 3812
rect 39060 3732 39164 3748
rect 39060 3668 39080 3732
rect 39144 3668 39164 3732
rect 39060 3652 39164 3668
rect 39060 3588 39080 3652
rect 39144 3588 39164 3652
rect 39060 3572 39164 3588
rect 39060 3508 39080 3572
rect 39144 3508 39164 3572
rect 39060 3492 39164 3508
rect 39060 3428 39080 3492
rect 39144 3428 39164 3492
rect 39060 3412 39164 3428
rect 39060 3348 39080 3412
rect 39144 3348 39164 3412
rect 39060 3332 39164 3348
rect 39060 3268 39080 3332
rect 39144 3268 39164 3332
rect 39060 3252 39164 3268
rect 39060 3188 39080 3252
rect 39144 3188 39164 3252
rect 39060 3172 39164 3188
rect 39060 3108 39080 3172
rect 39144 3108 39164 3172
rect 39060 3092 39164 3108
rect 39060 3028 39080 3092
rect 39144 3028 39164 3092
rect 39060 3012 39164 3028
rect 39060 2948 39080 3012
rect 39144 2948 39164 3012
rect 39060 2932 39164 2948
rect 39060 2868 39080 2932
rect 39144 2868 39164 2932
rect 39060 2852 39164 2868
rect 39060 2788 39080 2852
rect 39144 2788 39164 2852
rect 39060 2772 39164 2788
rect 39060 2708 39080 2772
rect 39144 2708 39164 2772
rect 39060 2692 39164 2708
rect 39060 2628 39080 2692
rect 39144 2628 39164 2692
rect 39060 2612 39164 2628
rect 39060 2548 39080 2612
rect 39144 2548 39164 2612
rect 39060 2532 39164 2548
rect 39060 2468 39080 2532
rect 39144 2468 39164 2532
rect 39060 2452 39164 2468
rect 39060 2388 39080 2452
rect 39144 2388 39164 2452
rect 39060 2372 39164 2388
rect 39060 2308 39080 2372
rect 39144 2308 39164 2372
rect 39060 2292 39164 2308
rect 39060 2228 39080 2292
rect 39144 2228 39164 2292
rect 39060 2212 39164 2228
rect 39060 2148 39080 2212
rect 39144 2148 39164 2212
rect 39060 2132 39164 2148
rect 39060 2068 39080 2132
rect 39144 2068 39164 2132
rect 39060 2052 39164 2068
rect 39060 1988 39080 2052
rect 39144 1988 39164 2052
rect 39060 1972 39164 1988
rect 39060 1908 39080 1972
rect 39144 1908 39164 1972
rect 39060 1892 39164 1908
rect 39060 1828 39080 1892
rect 39144 1828 39164 1892
rect 39060 1812 39164 1828
rect 39060 1748 39080 1812
rect 39144 1748 39164 1812
rect 39060 1732 39164 1748
rect 39060 1668 39080 1732
rect 39144 1668 39164 1732
rect 39060 1652 39164 1668
rect 39060 1588 39080 1652
rect 39144 1588 39164 1652
rect 39060 1572 39164 1588
rect 39060 1508 39080 1572
rect 39144 1508 39164 1572
rect 39060 1492 39164 1508
rect 39060 1428 39080 1492
rect 39144 1428 39164 1492
rect 39060 1412 39164 1428
rect 39060 1348 39080 1412
rect 39144 1348 39164 1412
rect 39060 1332 39164 1348
rect 39060 1268 39080 1332
rect 39144 1268 39164 1332
rect 39060 1252 39164 1268
rect 39060 1188 39080 1252
rect 39144 1188 39164 1252
rect 39060 1172 39164 1188
rect 39060 1108 39080 1172
rect 39144 1108 39164 1172
rect 39060 1092 39164 1108
rect 39060 1028 39080 1092
rect 39144 1028 39164 1092
rect 39060 1012 39164 1028
rect 39060 948 39080 1012
rect 39144 948 39164 1012
rect 39060 932 39164 948
rect 39060 868 39080 932
rect 39144 868 39164 932
rect 39060 852 39164 868
rect 39060 788 39080 852
rect 39144 788 39164 852
rect 39060 772 39164 788
rect 39060 708 39080 772
rect 39144 708 39164 772
rect 39060 692 39164 708
rect 39060 628 39080 692
rect 39144 628 39164 692
rect 39060 612 39164 628
rect 39060 548 39080 612
rect 39144 548 39164 612
rect 39060 532 39164 548
rect 39060 468 39080 532
rect 39144 468 39164 532
rect 39060 452 39164 468
rect 39060 388 39080 452
rect 39144 388 39164 452
rect 39060 372 39164 388
rect 39060 308 39080 372
rect 39144 308 39164 372
rect 39060 292 39164 308
rect 39060 228 39080 292
rect 39144 228 39164 292
rect 39060 212 39164 228
rect 33448 -148 33552 148
rect 27836 -228 27940 -212
rect 27836 -292 27856 -228
rect 27920 -292 27940 -228
rect 27836 -308 27940 -292
rect 27836 -372 27856 -308
rect 27920 -372 27940 -308
rect 27836 -388 27940 -372
rect 27836 -452 27856 -388
rect 27920 -452 27940 -388
rect 27836 -468 27940 -452
rect 27836 -532 27856 -468
rect 27920 -532 27940 -468
rect 27836 -548 27940 -532
rect 27836 -612 27856 -548
rect 27920 -612 27940 -548
rect 27836 -628 27940 -612
rect 27836 -692 27856 -628
rect 27920 -692 27940 -628
rect 27836 -708 27940 -692
rect 27836 -772 27856 -708
rect 27920 -772 27940 -708
rect 27836 -788 27940 -772
rect 27836 -852 27856 -788
rect 27920 -852 27940 -788
rect 27836 -868 27940 -852
rect 27836 -932 27856 -868
rect 27920 -932 27940 -868
rect 27836 -948 27940 -932
rect 27836 -1012 27856 -948
rect 27920 -1012 27940 -948
rect 27836 -1028 27940 -1012
rect 27836 -1092 27856 -1028
rect 27920 -1092 27940 -1028
rect 27836 -1108 27940 -1092
rect 27836 -1172 27856 -1108
rect 27920 -1172 27940 -1108
rect 27836 -1188 27940 -1172
rect 27836 -1252 27856 -1188
rect 27920 -1252 27940 -1188
rect 27836 -1268 27940 -1252
rect 27836 -1332 27856 -1268
rect 27920 -1332 27940 -1268
rect 27836 -1348 27940 -1332
rect 27836 -1412 27856 -1348
rect 27920 -1412 27940 -1348
rect 27836 -1428 27940 -1412
rect 27836 -1492 27856 -1428
rect 27920 -1492 27940 -1428
rect 27836 -1508 27940 -1492
rect 27836 -1572 27856 -1508
rect 27920 -1572 27940 -1508
rect 27836 -1588 27940 -1572
rect 27836 -1652 27856 -1588
rect 27920 -1652 27940 -1588
rect 27836 -1668 27940 -1652
rect 27836 -1732 27856 -1668
rect 27920 -1732 27940 -1668
rect 27836 -1748 27940 -1732
rect 27836 -1812 27856 -1748
rect 27920 -1812 27940 -1748
rect 27836 -1828 27940 -1812
rect 27836 -1892 27856 -1828
rect 27920 -1892 27940 -1828
rect 27836 -1908 27940 -1892
rect 27836 -1972 27856 -1908
rect 27920 -1972 27940 -1908
rect 27836 -1988 27940 -1972
rect 27836 -2052 27856 -1988
rect 27920 -2052 27940 -1988
rect 27836 -2068 27940 -2052
rect 27836 -2132 27856 -2068
rect 27920 -2132 27940 -2068
rect 27836 -2148 27940 -2132
rect 27836 -2212 27856 -2148
rect 27920 -2212 27940 -2148
rect 27836 -2228 27940 -2212
rect 27836 -2292 27856 -2228
rect 27920 -2292 27940 -2228
rect 27836 -2308 27940 -2292
rect 27836 -2372 27856 -2308
rect 27920 -2372 27940 -2308
rect 27836 -2388 27940 -2372
rect 27836 -2452 27856 -2388
rect 27920 -2452 27940 -2388
rect 27836 -2468 27940 -2452
rect 27836 -2532 27856 -2468
rect 27920 -2532 27940 -2468
rect 27836 -2548 27940 -2532
rect 27836 -2612 27856 -2548
rect 27920 -2612 27940 -2548
rect 27836 -2628 27940 -2612
rect 27836 -2692 27856 -2628
rect 27920 -2692 27940 -2628
rect 27836 -2708 27940 -2692
rect 27836 -2772 27856 -2708
rect 27920 -2772 27940 -2708
rect 27836 -2788 27940 -2772
rect 27836 -2852 27856 -2788
rect 27920 -2852 27940 -2788
rect 27836 -2868 27940 -2852
rect 27836 -2932 27856 -2868
rect 27920 -2932 27940 -2868
rect 27836 -2948 27940 -2932
rect 27836 -3012 27856 -2948
rect 27920 -3012 27940 -2948
rect 27836 -3028 27940 -3012
rect 27836 -3092 27856 -3028
rect 27920 -3092 27940 -3028
rect 27836 -3108 27940 -3092
rect 27836 -3172 27856 -3108
rect 27920 -3172 27940 -3108
rect 27836 -3188 27940 -3172
rect 27836 -3252 27856 -3188
rect 27920 -3252 27940 -3188
rect 27836 -3268 27940 -3252
rect 27836 -3332 27856 -3268
rect 27920 -3332 27940 -3268
rect 27836 -3348 27940 -3332
rect 27836 -3412 27856 -3348
rect 27920 -3412 27940 -3348
rect 27836 -3428 27940 -3412
rect 27836 -3492 27856 -3428
rect 27920 -3492 27940 -3428
rect 27836 -3508 27940 -3492
rect 27836 -3572 27856 -3508
rect 27920 -3572 27940 -3508
rect 27836 -3588 27940 -3572
rect 27836 -3652 27856 -3588
rect 27920 -3652 27940 -3588
rect 27836 -3668 27940 -3652
rect 27836 -3732 27856 -3668
rect 27920 -3732 27940 -3668
rect 27836 -3748 27940 -3732
rect 27836 -3812 27856 -3748
rect 27920 -3812 27940 -3748
rect 27836 -3828 27940 -3812
rect 27836 -3892 27856 -3828
rect 27920 -3892 27940 -3828
rect 27836 -3908 27940 -3892
rect 27836 -3972 27856 -3908
rect 27920 -3972 27940 -3908
rect 27836 -3988 27940 -3972
rect 27836 -4052 27856 -3988
rect 27920 -4052 27940 -3988
rect 27836 -4068 27940 -4052
rect 27836 -4132 27856 -4068
rect 27920 -4132 27940 -4068
rect 27836 -4148 27940 -4132
rect 27836 -4212 27856 -4148
rect 27920 -4212 27940 -4148
rect 27836 -4228 27940 -4212
rect 27836 -4292 27856 -4228
rect 27920 -4292 27940 -4228
rect 27836 -4308 27940 -4292
rect 27836 -4372 27856 -4308
rect 27920 -4372 27940 -4308
rect 27836 -4388 27940 -4372
rect 27836 -4452 27856 -4388
rect 27920 -4452 27940 -4388
rect 27836 -4468 27940 -4452
rect 27836 -4532 27856 -4468
rect 27920 -4532 27940 -4468
rect 27836 -4548 27940 -4532
rect 27836 -4612 27856 -4548
rect 27920 -4612 27940 -4548
rect 27836 -4628 27940 -4612
rect 27836 -4692 27856 -4628
rect 27920 -4692 27940 -4628
rect 27836 -4708 27940 -4692
rect 27836 -4772 27856 -4708
rect 27920 -4772 27940 -4708
rect 27836 -4788 27940 -4772
rect 27836 -4852 27856 -4788
rect 27920 -4852 27940 -4788
rect 27836 -4868 27940 -4852
rect 27836 -4932 27856 -4868
rect 27920 -4932 27940 -4868
rect 27836 -4948 27940 -4932
rect 27836 -5012 27856 -4948
rect 27920 -5012 27940 -4948
rect 27836 -5028 27940 -5012
rect 27836 -5092 27856 -5028
rect 27920 -5092 27940 -5028
rect 27836 -5108 27940 -5092
rect 22224 -5468 22328 -5172
rect 16612 -5548 16716 -5532
rect 16612 -5612 16632 -5548
rect 16696 -5612 16716 -5548
rect 16612 -5628 16716 -5612
rect 16612 -5692 16632 -5628
rect 16696 -5692 16716 -5628
rect 16612 -5708 16716 -5692
rect 16612 -5772 16632 -5708
rect 16696 -5772 16716 -5708
rect 16612 -5788 16716 -5772
rect 16612 -5852 16632 -5788
rect 16696 -5852 16716 -5788
rect 16612 -5868 16716 -5852
rect 16612 -5932 16632 -5868
rect 16696 -5932 16716 -5868
rect 16612 -5948 16716 -5932
rect 16612 -6012 16632 -5948
rect 16696 -6012 16716 -5948
rect 16612 -6028 16716 -6012
rect 16612 -6092 16632 -6028
rect 16696 -6092 16716 -6028
rect 16612 -6108 16716 -6092
rect 16612 -6172 16632 -6108
rect 16696 -6172 16716 -6108
rect 16612 -6188 16716 -6172
rect 16612 -6252 16632 -6188
rect 16696 -6252 16716 -6188
rect 16612 -6268 16716 -6252
rect 16612 -6332 16632 -6268
rect 16696 -6332 16716 -6268
rect 16612 -6348 16716 -6332
rect 16612 -6412 16632 -6348
rect 16696 -6412 16716 -6348
rect 16612 -6428 16716 -6412
rect 16612 -6492 16632 -6428
rect 16696 -6492 16716 -6428
rect 16612 -6508 16716 -6492
rect 16612 -6572 16632 -6508
rect 16696 -6572 16716 -6508
rect 16612 -6588 16716 -6572
rect 16612 -6652 16632 -6588
rect 16696 -6652 16716 -6588
rect 16612 -6668 16716 -6652
rect 16612 -6732 16632 -6668
rect 16696 -6732 16716 -6668
rect 16612 -6748 16716 -6732
rect 16612 -6812 16632 -6748
rect 16696 -6812 16716 -6748
rect 16612 -6828 16716 -6812
rect 16612 -6892 16632 -6828
rect 16696 -6892 16716 -6828
rect 16612 -6908 16716 -6892
rect 16612 -6972 16632 -6908
rect 16696 -6972 16716 -6908
rect 16612 -6988 16716 -6972
rect 16612 -7052 16632 -6988
rect 16696 -7052 16716 -6988
rect 16612 -7068 16716 -7052
rect 16612 -7132 16632 -7068
rect 16696 -7132 16716 -7068
rect 16612 -7148 16716 -7132
rect 16612 -7212 16632 -7148
rect 16696 -7212 16716 -7148
rect 16612 -7228 16716 -7212
rect 16612 -7292 16632 -7228
rect 16696 -7292 16716 -7228
rect 16612 -7308 16716 -7292
rect 16612 -7372 16632 -7308
rect 16696 -7372 16716 -7308
rect 16612 -7388 16716 -7372
rect 16612 -7452 16632 -7388
rect 16696 -7452 16716 -7388
rect 16612 -7468 16716 -7452
rect 16612 -7532 16632 -7468
rect 16696 -7532 16716 -7468
rect 16612 -7548 16716 -7532
rect 16612 -7612 16632 -7548
rect 16696 -7612 16716 -7548
rect 16612 -7628 16716 -7612
rect 16612 -7692 16632 -7628
rect 16696 -7692 16716 -7628
rect 16612 -7708 16716 -7692
rect 16612 -7772 16632 -7708
rect 16696 -7772 16716 -7708
rect 16612 -7788 16716 -7772
rect 16612 -7852 16632 -7788
rect 16696 -7852 16716 -7788
rect 16612 -7868 16716 -7852
rect 16612 -7932 16632 -7868
rect 16696 -7932 16716 -7868
rect 16612 -7948 16716 -7932
rect 16612 -8012 16632 -7948
rect 16696 -8012 16716 -7948
rect 16612 -8028 16716 -8012
rect 16612 -8092 16632 -8028
rect 16696 -8092 16716 -8028
rect 16612 -8108 16716 -8092
rect 16612 -8172 16632 -8108
rect 16696 -8172 16716 -8108
rect 16612 -8188 16716 -8172
rect 16612 -8252 16632 -8188
rect 16696 -8252 16716 -8188
rect 16612 -8268 16716 -8252
rect 16612 -8332 16632 -8268
rect 16696 -8332 16716 -8268
rect 16612 -8348 16716 -8332
rect 16612 -8412 16632 -8348
rect 16696 -8412 16716 -8348
rect 16612 -8428 16716 -8412
rect 16612 -8492 16632 -8428
rect 16696 -8492 16716 -8428
rect 16612 -8508 16716 -8492
rect 16612 -8572 16632 -8508
rect 16696 -8572 16716 -8508
rect 16612 -8588 16716 -8572
rect 16612 -8652 16632 -8588
rect 16696 -8652 16716 -8588
rect 16612 -8668 16716 -8652
rect 16612 -8732 16632 -8668
rect 16696 -8732 16716 -8668
rect 16612 -8748 16716 -8732
rect 16612 -8812 16632 -8748
rect 16696 -8812 16716 -8748
rect 16612 -8828 16716 -8812
rect 16612 -8892 16632 -8828
rect 16696 -8892 16716 -8828
rect 16612 -8908 16716 -8892
rect 16612 -8972 16632 -8908
rect 16696 -8972 16716 -8908
rect 16612 -8988 16716 -8972
rect 16612 -9052 16632 -8988
rect 16696 -9052 16716 -8988
rect 16612 -9068 16716 -9052
rect 16612 -9132 16632 -9068
rect 16696 -9132 16716 -9068
rect 16612 -9148 16716 -9132
rect 16612 -9212 16632 -9148
rect 16696 -9212 16716 -9148
rect 16612 -9228 16716 -9212
rect 16612 -9292 16632 -9228
rect 16696 -9292 16716 -9228
rect 16612 -9308 16716 -9292
rect 16612 -9372 16632 -9308
rect 16696 -9372 16716 -9308
rect 16612 -9388 16716 -9372
rect 16612 -9452 16632 -9388
rect 16696 -9452 16716 -9388
rect 16612 -9468 16716 -9452
rect 16612 -9532 16632 -9468
rect 16696 -9532 16716 -9468
rect 16612 -9548 16716 -9532
rect 16612 -9612 16632 -9548
rect 16696 -9612 16716 -9548
rect 16612 -9628 16716 -9612
rect 16612 -9692 16632 -9628
rect 16696 -9692 16716 -9628
rect 16612 -9708 16716 -9692
rect 16612 -9772 16632 -9708
rect 16696 -9772 16716 -9708
rect 16612 -9788 16716 -9772
rect 16612 -9852 16632 -9788
rect 16696 -9852 16716 -9788
rect 16612 -9868 16716 -9852
rect 16612 -9932 16632 -9868
rect 16696 -9932 16716 -9868
rect 16612 -9948 16716 -9932
rect 16612 -10012 16632 -9948
rect 16696 -10012 16716 -9948
rect 16612 -10028 16716 -10012
rect 16612 -10092 16632 -10028
rect 16696 -10092 16716 -10028
rect 16612 -10108 16716 -10092
rect 16612 -10172 16632 -10108
rect 16696 -10172 16716 -10108
rect 16612 -10188 16716 -10172
rect 16612 -10252 16632 -10188
rect 16696 -10252 16716 -10188
rect 16612 -10268 16716 -10252
rect 16612 -10332 16632 -10268
rect 16696 -10332 16716 -10268
rect 16612 -10348 16716 -10332
rect 16612 -10412 16632 -10348
rect 16696 -10412 16716 -10348
rect 16612 -10428 16716 -10412
rect 11000 -10788 11104 -10492
rect 5388 -10868 5492 -10852
rect 5388 -10932 5408 -10868
rect 5472 -10932 5492 -10868
rect 5388 -10948 5492 -10932
rect 5388 -11012 5408 -10948
rect 5472 -11012 5492 -10948
rect 5388 -11028 5492 -11012
rect 5388 -11092 5408 -11028
rect 5472 -11092 5492 -11028
rect 5388 -11108 5492 -11092
rect 5388 -11172 5408 -11108
rect 5472 -11172 5492 -11108
rect 5388 -11188 5492 -11172
rect 5388 -11252 5408 -11188
rect 5472 -11252 5492 -11188
rect 5388 -11268 5492 -11252
rect 5388 -11332 5408 -11268
rect 5472 -11332 5492 -11268
rect 5388 -11348 5492 -11332
rect 5388 -11412 5408 -11348
rect 5472 -11412 5492 -11348
rect 5388 -11428 5492 -11412
rect 5388 -11492 5408 -11428
rect 5472 -11492 5492 -11428
rect 5388 -11508 5492 -11492
rect 5388 -11572 5408 -11508
rect 5472 -11572 5492 -11508
rect 5388 -11588 5492 -11572
rect 5388 -11652 5408 -11588
rect 5472 -11652 5492 -11588
rect 5388 -11668 5492 -11652
rect 5388 -11732 5408 -11668
rect 5472 -11732 5492 -11668
rect 5388 -11748 5492 -11732
rect 5388 -11812 5408 -11748
rect 5472 -11812 5492 -11748
rect 5388 -11828 5492 -11812
rect 5388 -11892 5408 -11828
rect 5472 -11892 5492 -11828
rect 5388 -11908 5492 -11892
rect 5388 -11972 5408 -11908
rect 5472 -11972 5492 -11908
rect 5388 -11988 5492 -11972
rect 5388 -12052 5408 -11988
rect 5472 -12052 5492 -11988
rect 5388 -12068 5492 -12052
rect 5388 -12132 5408 -12068
rect 5472 -12132 5492 -12068
rect 5388 -12148 5492 -12132
rect 5388 -12212 5408 -12148
rect 5472 -12212 5492 -12148
rect 5388 -12228 5492 -12212
rect 5388 -12292 5408 -12228
rect 5472 -12292 5492 -12228
rect 5388 -12308 5492 -12292
rect 5388 -12372 5408 -12308
rect 5472 -12372 5492 -12308
rect 5388 -12388 5492 -12372
rect 5388 -12452 5408 -12388
rect 5472 -12452 5492 -12388
rect 5388 -12468 5492 -12452
rect 5388 -12532 5408 -12468
rect 5472 -12532 5492 -12468
rect 5388 -12548 5492 -12532
rect 5388 -12612 5408 -12548
rect 5472 -12612 5492 -12548
rect 5388 -12628 5492 -12612
rect 5388 -12692 5408 -12628
rect 5472 -12692 5492 -12628
rect 5388 -12708 5492 -12692
rect 5388 -12772 5408 -12708
rect 5472 -12772 5492 -12708
rect 5388 -12788 5492 -12772
rect 5388 -12852 5408 -12788
rect 5472 -12852 5492 -12788
rect 5388 -12868 5492 -12852
rect 5388 -12932 5408 -12868
rect 5472 -12932 5492 -12868
rect 5388 -12948 5492 -12932
rect 5388 -13012 5408 -12948
rect 5472 -13012 5492 -12948
rect 5388 -13028 5492 -13012
rect 5388 -13092 5408 -13028
rect 5472 -13092 5492 -13028
rect 5388 -13108 5492 -13092
rect 5388 -13172 5408 -13108
rect 5472 -13172 5492 -13108
rect 5388 -13188 5492 -13172
rect 5388 -13252 5408 -13188
rect 5472 -13252 5492 -13188
rect 5388 -13268 5492 -13252
rect 5388 -13332 5408 -13268
rect 5472 -13332 5492 -13268
rect 5388 -13348 5492 -13332
rect 5388 -13412 5408 -13348
rect 5472 -13412 5492 -13348
rect 5388 -13428 5492 -13412
rect 5388 -13492 5408 -13428
rect 5472 -13492 5492 -13428
rect 5388 -13508 5492 -13492
rect 5388 -13572 5408 -13508
rect 5472 -13572 5492 -13508
rect 5388 -13588 5492 -13572
rect 5388 -13652 5408 -13588
rect 5472 -13652 5492 -13588
rect 5388 -13668 5492 -13652
rect 5388 -13732 5408 -13668
rect 5472 -13732 5492 -13668
rect 5388 -13748 5492 -13732
rect 5388 -13812 5408 -13748
rect 5472 -13812 5492 -13748
rect 5388 -13828 5492 -13812
rect 5388 -13892 5408 -13828
rect 5472 -13892 5492 -13828
rect 5388 -13908 5492 -13892
rect 5388 -13972 5408 -13908
rect 5472 -13972 5492 -13908
rect 5388 -13988 5492 -13972
rect 5388 -14052 5408 -13988
rect 5472 -14052 5492 -13988
rect 5388 -14068 5492 -14052
rect 5388 -14132 5408 -14068
rect 5472 -14132 5492 -14068
rect 5388 -14148 5492 -14132
rect 5388 -14212 5408 -14148
rect 5472 -14212 5492 -14148
rect 5388 -14228 5492 -14212
rect 5388 -14292 5408 -14228
rect 5472 -14292 5492 -14228
rect 5388 -14308 5492 -14292
rect 5388 -14372 5408 -14308
rect 5472 -14372 5492 -14308
rect 5388 -14388 5492 -14372
rect 5388 -14452 5408 -14388
rect 5472 -14452 5492 -14388
rect 5388 -14468 5492 -14452
rect 5388 -14532 5408 -14468
rect 5472 -14532 5492 -14468
rect 5388 -14548 5492 -14532
rect 5388 -14612 5408 -14548
rect 5472 -14612 5492 -14548
rect 5388 -14628 5492 -14612
rect 5388 -14692 5408 -14628
rect 5472 -14692 5492 -14628
rect 5388 -14708 5492 -14692
rect 5388 -14772 5408 -14708
rect 5472 -14772 5492 -14708
rect 5388 -14788 5492 -14772
rect 5388 -14852 5408 -14788
rect 5472 -14852 5492 -14788
rect 5388 -14868 5492 -14852
rect 5388 -14932 5408 -14868
rect 5472 -14932 5492 -14868
rect 5388 -14948 5492 -14932
rect 5388 -15012 5408 -14948
rect 5472 -15012 5492 -14948
rect 5388 -15028 5492 -15012
rect 5388 -15092 5408 -15028
rect 5472 -15092 5492 -15028
rect 5388 -15108 5492 -15092
rect 5388 -15172 5408 -15108
rect 5472 -15172 5492 -15108
rect 5388 -15188 5492 -15172
rect 5388 -15252 5408 -15188
rect 5472 -15252 5492 -15188
rect 5388 -15268 5492 -15252
rect 5388 -15332 5408 -15268
rect 5472 -15332 5492 -15268
rect 5388 -15348 5492 -15332
rect 5388 -15412 5408 -15348
rect 5472 -15412 5492 -15348
rect 5388 -15428 5492 -15412
rect 5388 -15492 5408 -15428
rect 5472 -15492 5492 -15428
rect 5388 -15508 5492 -15492
rect 5388 -15572 5408 -15508
rect 5472 -15572 5492 -15508
rect 5388 -15588 5492 -15572
rect 5388 -15652 5408 -15588
rect 5472 -15652 5492 -15588
rect 5388 -15668 5492 -15652
rect 5388 -15732 5408 -15668
rect 5472 -15732 5492 -15668
rect 5388 -15748 5492 -15732
rect -224 -16108 -120 -15812
rect -5836 -16188 -5732 -16172
rect -5836 -16252 -5816 -16188
rect -5752 -16252 -5732 -16188
rect -5836 -16268 -5732 -16252
rect -5836 -16332 -5816 -16268
rect -5752 -16332 -5732 -16268
rect -5836 -16348 -5732 -16332
rect -5836 -16412 -5816 -16348
rect -5752 -16412 -5732 -16348
rect -5836 -16428 -5732 -16412
rect -5836 -16492 -5816 -16428
rect -5752 -16492 -5732 -16428
rect -5836 -16508 -5732 -16492
rect -5836 -16572 -5816 -16508
rect -5752 -16572 -5732 -16508
rect -5836 -16588 -5732 -16572
rect -5836 -16652 -5816 -16588
rect -5752 -16652 -5732 -16588
rect -5836 -16668 -5732 -16652
rect -5836 -16732 -5816 -16668
rect -5752 -16732 -5732 -16668
rect -5836 -16748 -5732 -16732
rect -5836 -16812 -5816 -16748
rect -5752 -16812 -5732 -16748
rect -5836 -16828 -5732 -16812
rect -5836 -16892 -5816 -16828
rect -5752 -16892 -5732 -16828
rect -5836 -16908 -5732 -16892
rect -5836 -16972 -5816 -16908
rect -5752 -16972 -5732 -16908
rect -5836 -16988 -5732 -16972
rect -5836 -17052 -5816 -16988
rect -5752 -17052 -5732 -16988
rect -5836 -17068 -5732 -17052
rect -5836 -17132 -5816 -17068
rect -5752 -17132 -5732 -17068
rect -5836 -17148 -5732 -17132
rect -5836 -17212 -5816 -17148
rect -5752 -17212 -5732 -17148
rect -5836 -17228 -5732 -17212
rect -5836 -17292 -5816 -17228
rect -5752 -17292 -5732 -17228
rect -5836 -17308 -5732 -17292
rect -5836 -17372 -5816 -17308
rect -5752 -17372 -5732 -17308
rect -5836 -17388 -5732 -17372
rect -5836 -17452 -5816 -17388
rect -5752 -17452 -5732 -17388
rect -5836 -17468 -5732 -17452
rect -5836 -17532 -5816 -17468
rect -5752 -17532 -5732 -17468
rect -5836 -17548 -5732 -17532
rect -5836 -17612 -5816 -17548
rect -5752 -17612 -5732 -17548
rect -5836 -17628 -5732 -17612
rect -5836 -17692 -5816 -17628
rect -5752 -17692 -5732 -17628
rect -5836 -17708 -5732 -17692
rect -5836 -17772 -5816 -17708
rect -5752 -17772 -5732 -17708
rect -5836 -17788 -5732 -17772
rect -5836 -17852 -5816 -17788
rect -5752 -17852 -5732 -17788
rect -5836 -17868 -5732 -17852
rect -5836 -17932 -5816 -17868
rect -5752 -17932 -5732 -17868
rect -5836 -17948 -5732 -17932
rect -5836 -18012 -5816 -17948
rect -5752 -18012 -5732 -17948
rect -5836 -18028 -5732 -18012
rect -5836 -18092 -5816 -18028
rect -5752 -18092 -5732 -18028
rect -5836 -18108 -5732 -18092
rect -5836 -18172 -5816 -18108
rect -5752 -18172 -5732 -18108
rect -5836 -18188 -5732 -18172
rect -5836 -18252 -5816 -18188
rect -5752 -18252 -5732 -18188
rect -5836 -18268 -5732 -18252
rect -5836 -18332 -5816 -18268
rect -5752 -18332 -5732 -18268
rect -5836 -18348 -5732 -18332
rect -5836 -18412 -5816 -18348
rect -5752 -18412 -5732 -18348
rect -5836 -18428 -5732 -18412
rect -5836 -18492 -5816 -18428
rect -5752 -18492 -5732 -18428
rect -5836 -18508 -5732 -18492
rect -5836 -18572 -5816 -18508
rect -5752 -18572 -5732 -18508
rect -5836 -18588 -5732 -18572
rect -5836 -18652 -5816 -18588
rect -5752 -18652 -5732 -18588
rect -5836 -18668 -5732 -18652
rect -5836 -18732 -5816 -18668
rect -5752 -18732 -5732 -18668
rect -5836 -18748 -5732 -18732
rect -5836 -18812 -5816 -18748
rect -5752 -18812 -5732 -18748
rect -5836 -18828 -5732 -18812
rect -5836 -18892 -5816 -18828
rect -5752 -18892 -5732 -18828
rect -5836 -18908 -5732 -18892
rect -5836 -18972 -5816 -18908
rect -5752 -18972 -5732 -18908
rect -5836 -18988 -5732 -18972
rect -5836 -19052 -5816 -18988
rect -5752 -19052 -5732 -18988
rect -5836 -19068 -5732 -19052
rect -5836 -19132 -5816 -19068
rect -5752 -19132 -5732 -19068
rect -5836 -19148 -5732 -19132
rect -5836 -19212 -5816 -19148
rect -5752 -19212 -5732 -19148
rect -5836 -19228 -5732 -19212
rect -5836 -19292 -5816 -19228
rect -5752 -19292 -5732 -19228
rect -5836 -19308 -5732 -19292
rect -5836 -19372 -5816 -19308
rect -5752 -19372 -5732 -19308
rect -5836 -19388 -5732 -19372
rect -5836 -19452 -5816 -19388
rect -5752 -19452 -5732 -19388
rect -5836 -19468 -5732 -19452
rect -5836 -19532 -5816 -19468
rect -5752 -19532 -5732 -19468
rect -5836 -19548 -5732 -19532
rect -5836 -19612 -5816 -19548
rect -5752 -19612 -5732 -19548
rect -5836 -19628 -5732 -19612
rect -5836 -19692 -5816 -19628
rect -5752 -19692 -5732 -19628
rect -5836 -19708 -5732 -19692
rect -5836 -19772 -5816 -19708
rect -5752 -19772 -5732 -19708
rect -5836 -19788 -5732 -19772
rect -5836 -19852 -5816 -19788
rect -5752 -19852 -5732 -19788
rect -5836 -19868 -5732 -19852
rect -5836 -19932 -5816 -19868
rect -5752 -19932 -5732 -19868
rect -5836 -19948 -5732 -19932
rect -5836 -20012 -5816 -19948
rect -5752 -20012 -5732 -19948
rect -5836 -20028 -5732 -20012
rect -5836 -20092 -5816 -20028
rect -5752 -20092 -5732 -20028
rect -5836 -20108 -5732 -20092
rect -5836 -20172 -5816 -20108
rect -5752 -20172 -5732 -20108
rect -5836 -20188 -5732 -20172
rect -5836 -20252 -5816 -20188
rect -5752 -20252 -5732 -20188
rect -5836 -20268 -5732 -20252
rect -5836 -20332 -5816 -20268
rect -5752 -20332 -5732 -20268
rect -5836 -20348 -5732 -20332
rect -5836 -20412 -5816 -20348
rect -5752 -20412 -5732 -20348
rect -5836 -20428 -5732 -20412
rect -5836 -20492 -5816 -20428
rect -5752 -20492 -5732 -20428
rect -5836 -20508 -5732 -20492
rect -5836 -20572 -5816 -20508
rect -5752 -20572 -5732 -20508
rect -5836 -20588 -5732 -20572
rect -5836 -20652 -5816 -20588
rect -5752 -20652 -5732 -20588
rect -5836 -20668 -5732 -20652
rect -5836 -20732 -5816 -20668
rect -5752 -20732 -5732 -20668
rect -5836 -20748 -5732 -20732
rect -5836 -20812 -5816 -20748
rect -5752 -20812 -5732 -20748
rect -5836 -20828 -5732 -20812
rect -5836 -20892 -5816 -20828
rect -5752 -20892 -5732 -20828
rect -5836 -20908 -5732 -20892
rect -5836 -20972 -5816 -20908
rect -5752 -20972 -5732 -20908
rect -5836 -20988 -5732 -20972
rect -5836 -21052 -5816 -20988
rect -5752 -21052 -5732 -20988
rect -5836 -21068 -5732 -21052
rect -11448 -21428 -11344 -21132
rect -17060 -21508 -16956 -21492
rect -17060 -21572 -17040 -21508
rect -16976 -21572 -16956 -21508
rect -17060 -21588 -16956 -21572
rect -17060 -21652 -17040 -21588
rect -16976 -21652 -16956 -21588
rect -17060 -21668 -16956 -21652
rect -17060 -21732 -17040 -21668
rect -16976 -21732 -16956 -21668
rect -17060 -21748 -16956 -21732
rect -17060 -21812 -17040 -21748
rect -16976 -21812 -16956 -21748
rect -17060 -21828 -16956 -21812
rect -17060 -21892 -17040 -21828
rect -16976 -21892 -16956 -21828
rect -17060 -21908 -16956 -21892
rect -17060 -21972 -17040 -21908
rect -16976 -21972 -16956 -21908
rect -17060 -21988 -16956 -21972
rect -17060 -22052 -17040 -21988
rect -16976 -22052 -16956 -21988
rect -17060 -22068 -16956 -22052
rect -17060 -22132 -17040 -22068
rect -16976 -22132 -16956 -22068
rect -17060 -22148 -16956 -22132
rect -17060 -22212 -17040 -22148
rect -16976 -22212 -16956 -22148
rect -17060 -22228 -16956 -22212
rect -17060 -22292 -17040 -22228
rect -16976 -22292 -16956 -22228
rect -17060 -22308 -16956 -22292
rect -17060 -22372 -17040 -22308
rect -16976 -22372 -16956 -22308
rect -17060 -22388 -16956 -22372
rect -17060 -22452 -17040 -22388
rect -16976 -22452 -16956 -22388
rect -17060 -22468 -16956 -22452
rect -17060 -22532 -17040 -22468
rect -16976 -22532 -16956 -22468
rect -17060 -22548 -16956 -22532
rect -17060 -22612 -17040 -22548
rect -16976 -22612 -16956 -22548
rect -17060 -22628 -16956 -22612
rect -17060 -22692 -17040 -22628
rect -16976 -22692 -16956 -22628
rect -17060 -22708 -16956 -22692
rect -17060 -22772 -17040 -22708
rect -16976 -22772 -16956 -22708
rect -17060 -22788 -16956 -22772
rect -17060 -22852 -17040 -22788
rect -16976 -22852 -16956 -22788
rect -17060 -22868 -16956 -22852
rect -17060 -22932 -17040 -22868
rect -16976 -22932 -16956 -22868
rect -17060 -22948 -16956 -22932
rect -17060 -23012 -17040 -22948
rect -16976 -23012 -16956 -22948
rect -17060 -23028 -16956 -23012
rect -17060 -23092 -17040 -23028
rect -16976 -23092 -16956 -23028
rect -17060 -23108 -16956 -23092
rect -17060 -23172 -17040 -23108
rect -16976 -23172 -16956 -23108
rect -17060 -23188 -16956 -23172
rect -17060 -23252 -17040 -23188
rect -16976 -23252 -16956 -23188
rect -17060 -23268 -16956 -23252
rect -17060 -23332 -17040 -23268
rect -16976 -23332 -16956 -23268
rect -17060 -23348 -16956 -23332
rect -17060 -23412 -17040 -23348
rect -16976 -23412 -16956 -23348
rect -17060 -23428 -16956 -23412
rect -17060 -23492 -17040 -23428
rect -16976 -23492 -16956 -23428
rect -17060 -23508 -16956 -23492
rect -17060 -23572 -17040 -23508
rect -16976 -23572 -16956 -23508
rect -17060 -23588 -16956 -23572
rect -17060 -23652 -17040 -23588
rect -16976 -23652 -16956 -23588
rect -17060 -23668 -16956 -23652
rect -17060 -23732 -17040 -23668
rect -16976 -23732 -16956 -23668
rect -17060 -23748 -16956 -23732
rect -17060 -23812 -17040 -23748
rect -16976 -23812 -16956 -23748
rect -17060 -23828 -16956 -23812
rect -17060 -23892 -17040 -23828
rect -16976 -23892 -16956 -23828
rect -17060 -23908 -16956 -23892
rect -17060 -23972 -17040 -23908
rect -16976 -23972 -16956 -23908
rect -17060 -23988 -16956 -23972
rect -17060 -24052 -17040 -23988
rect -16976 -24052 -16956 -23988
rect -17060 -24068 -16956 -24052
rect -17060 -24132 -17040 -24068
rect -16976 -24132 -16956 -24068
rect -17060 -24148 -16956 -24132
rect -17060 -24212 -17040 -24148
rect -16976 -24212 -16956 -24148
rect -17060 -24228 -16956 -24212
rect -17060 -24292 -17040 -24228
rect -16976 -24292 -16956 -24228
rect -17060 -24308 -16956 -24292
rect -17060 -24372 -17040 -24308
rect -16976 -24372 -16956 -24308
rect -17060 -24388 -16956 -24372
rect -17060 -24452 -17040 -24388
rect -16976 -24452 -16956 -24388
rect -17060 -24468 -16956 -24452
rect -17060 -24532 -17040 -24468
rect -16976 -24532 -16956 -24468
rect -17060 -24548 -16956 -24532
rect -17060 -24612 -17040 -24548
rect -16976 -24612 -16956 -24548
rect -17060 -24628 -16956 -24612
rect -17060 -24692 -17040 -24628
rect -16976 -24692 -16956 -24628
rect -17060 -24708 -16956 -24692
rect -17060 -24772 -17040 -24708
rect -16976 -24772 -16956 -24708
rect -17060 -24788 -16956 -24772
rect -17060 -24852 -17040 -24788
rect -16976 -24852 -16956 -24788
rect -17060 -24868 -16956 -24852
rect -17060 -24932 -17040 -24868
rect -16976 -24932 -16956 -24868
rect -17060 -24948 -16956 -24932
rect -17060 -25012 -17040 -24948
rect -16976 -25012 -16956 -24948
rect -17060 -25028 -16956 -25012
rect -17060 -25092 -17040 -25028
rect -16976 -25092 -16956 -25028
rect -17060 -25108 -16956 -25092
rect -17060 -25172 -17040 -25108
rect -16976 -25172 -16956 -25108
rect -17060 -25188 -16956 -25172
rect -17060 -25252 -17040 -25188
rect -16976 -25252 -16956 -25188
rect -17060 -25268 -16956 -25252
rect -17060 -25332 -17040 -25268
rect -16976 -25332 -16956 -25268
rect -17060 -25348 -16956 -25332
rect -17060 -25412 -17040 -25348
rect -16976 -25412 -16956 -25348
rect -17060 -25428 -16956 -25412
rect -17060 -25492 -17040 -25428
rect -16976 -25492 -16956 -25428
rect -17060 -25508 -16956 -25492
rect -17060 -25572 -17040 -25508
rect -16976 -25572 -16956 -25508
rect -17060 -25588 -16956 -25572
rect -17060 -25652 -17040 -25588
rect -16976 -25652 -16956 -25588
rect -17060 -25668 -16956 -25652
rect -17060 -25732 -17040 -25668
rect -16976 -25732 -16956 -25668
rect -17060 -25748 -16956 -25732
rect -17060 -25812 -17040 -25748
rect -16976 -25812 -16956 -25748
rect -17060 -25828 -16956 -25812
rect -17060 -25892 -17040 -25828
rect -16976 -25892 -16956 -25828
rect -17060 -25908 -16956 -25892
rect -17060 -25972 -17040 -25908
rect -16976 -25972 -16956 -25908
rect -17060 -25988 -16956 -25972
rect -17060 -26052 -17040 -25988
rect -16976 -26052 -16956 -25988
rect -17060 -26068 -16956 -26052
rect -17060 -26132 -17040 -26068
rect -16976 -26132 -16956 -26068
rect -17060 -26148 -16956 -26132
rect -17060 -26212 -17040 -26148
rect -16976 -26212 -16956 -26148
rect -17060 -26228 -16956 -26212
rect -17060 -26292 -17040 -26228
rect -16976 -26292 -16956 -26228
rect -17060 -26308 -16956 -26292
rect -17060 -26372 -17040 -26308
rect -16976 -26372 -16956 -26308
rect -17060 -26388 -16956 -26372
rect -22672 -26748 -22568 -26452
rect -28284 -26828 -28180 -26812
rect -28284 -26892 -28264 -26828
rect -28200 -26892 -28180 -26828
rect -28284 -26908 -28180 -26892
rect -28284 -26972 -28264 -26908
rect -28200 -26972 -28180 -26908
rect -28284 -26988 -28180 -26972
rect -28284 -27052 -28264 -26988
rect -28200 -27052 -28180 -26988
rect -28284 -27068 -28180 -27052
rect -28284 -27132 -28264 -27068
rect -28200 -27132 -28180 -27068
rect -28284 -27148 -28180 -27132
rect -28284 -27212 -28264 -27148
rect -28200 -27212 -28180 -27148
rect -28284 -27228 -28180 -27212
rect -28284 -27292 -28264 -27228
rect -28200 -27292 -28180 -27228
rect -28284 -27308 -28180 -27292
rect -28284 -27372 -28264 -27308
rect -28200 -27372 -28180 -27308
rect -28284 -27388 -28180 -27372
rect -28284 -27452 -28264 -27388
rect -28200 -27452 -28180 -27388
rect -28284 -27468 -28180 -27452
rect -28284 -27532 -28264 -27468
rect -28200 -27532 -28180 -27468
rect -28284 -27548 -28180 -27532
rect -28284 -27612 -28264 -27548
rect -28200 -27612 -28180 -27548
rect -28284 -27628 -28180 -27612
rect -28284 -27692 -28264 -27628
rect -28200 -27692 -28180 -27628
rect -28284 -27708 -28180 -27692
rect -28284 -27772 -28264 -27708
rect -28200 -27772 -28180 -27708
rect -28284 -27788 -28180 -27772
rect -28284 -27852 -28264 -27788
rect -28200 -27852 -28180 -27788
rect -28284 -27868 -28180 -27852
rect -28284 -27932 -28264 -27868
rect -28200 -27932 -28180 -27868
rect -28284 -27948 -28180 -27932
rect -28284 -28012 -28264 -27948
rect -28200 -28012 -28180 -27948
rect -28284 -28028 -28180 -28012
rect -28284 -28092 -28264 -28028
rect -28200 -28092 -28180 -28028
rect -28284 -28108 -28180 -28092
rect -28284 -28172 -28264 -28108
rect -28200 -28172 -28180 -28108
rect -28284 -28188 -28180 -28172
rect -28284 -28252 -28264 -28188
rect -28200 -28252 -28180 -28188
rect -28284 -28268 -28180 -28252
rect -28284 -28332 -28264 -28268
rect -28200 -28332 -28180 -28268
rect -28284 -28348 -28180 -28332
rect -28284 -28412 -28264 -28348
rect -28200 -28412 -28180 -28348
rect -28284 -28428 -28180 -28412
rect -28284 -28492 -28264 -28428
rect -28200 -28492 -28180 -28428
rect -28284 -28508 -28180 -28492
rect -28284 -28572 -28264 -28508
rect -28200 -28572 -28180 -28508
rect -28284 -28588 -28180 -28572
rect -28284 -28652 -28264 -28588
rect -28200 -28652 -28180 -28588
rect -28284 -28668 -28180 -28652
rect -28284 -28732 -28264 -28668
rect -28200 -28732 -28180 -28668
rect -28284 -28748 -28180 -28732
rect -28284 -28812 -28264 -28748
rect -28200 -28812 -28180 -28748
rect -28284 -28828 -28180 -28812
rect -28284 -28892 -28264 -28828
rect -28200 -28892 -28180 -28828
rect -28284 -28908 -28180 -28892
rect -28284 -28972 -28264 -28908
rect -28200 -28972 -28180 -28908
rect -28284 -28988 -28180 -28972
rect -28284 -29052 -28264 -28988
rect -28200 -29052 -28180 -28988
rect -28284 -29068 -28180 -29052
rect -28284 -29132 -28264 -29068
rect -28200 -29132 -28180 -29068
rect -28284 -29148 -28180 -29132
rect -28284 -29212 -28264 -29148
rect -28200 -29212 -28180 -29148
rect -28284 -29228 -28180 -29212
rect -28284 -29292 -28264 -29228
rect -28200 -29292 -28180 -29228
rect -28284 -29308 -28180 -29292
rect -28284 -29372 -28264 -29308
rect -28200 -29372 -28180 -29308
rect -28284 -29388 -28180 -29372
rect -28284 -29452 -28264 -29388
rect -28200 -29452 -28180 -29388
rect -28284 -29468 -28180 -29452
rect -28284 -29532 -28264 -29468
rect -28200 -29532 -28180 -29468
rect -28284 -29548 -28180 -29532
rect -28284 -29612 -28264 -29548
rect -28200 -29612 -28180 -29548
rect -28284 -29628 -28180 -29612
rect -28284 -29692 -28264 -29628
rect -28200 -29692 -28180 -29628
rect -28284 -29708 -28180 -29692
rect -28284 -29772 -28264 -29708
rect -28200 -29772 -28180 -29708
rect -28284 -29788 -28180 -29772
rect -28284 -29852 -28264 -29788
rect -28200 -29852 -28180 -29788
rect -28284 -29868 -28180 -29852
rect -28284 -29932 -28264 -29868
rect -28200 -29932 -28180 -29868
rect -28284 -29948 -28180 -29932
rect -28284 -30012 -28264 -29948
rect -28200 -30012 -28180 -29948
rect -28284 -30028 -28180 -30012
rect -28284 -30092 -28264 -30028
rect -28200 -30092 -28180 -30028
rect -28284 -30108 -28180 -30092
rect -28284 -30172 -28264 -30108
rect -28200 -30172 -28180 -30108
rect -28284 -30188 -28180 -30172
rect -28284 -30252 -28264 -30188
rect -28200 -30252 -28180 -30188
rect -28284 -30268 -28180 -30252
rect -28284 -30332 -28264 -30268
rect -28200 -30332 -28180 -30268
rect -28284 -30348 -28180 -30332
rect -28284 -30412 -28264 -30348
rect -28200 -30412 -28180 -30348
rect -28284 -30428 -28180 -30412
rect -28284 -30492 -28264 -30428
rect -28200 -30492 -28180 -30428
rect -28284 -30508 -28180 -30492
rect -28284 -30572 -28264 -30508
rect -28200 -30572 -28180 -30508
rect -28284 -30588 -28180 -30572
rect -28284 -30652 -28264 -30588
rect -28200 -30652 -28180 -30588
rect -28284 -30668 -28180 -30652
rect -28284 -30732 -28264 -30668
rect -28200 -30732 -28180 -30668
rect -28284 -30748 -28180 -30732
rect -28284 -30812 -28264 -30748
rect -28200 -30812 -28180 -30748
rect -28284 -30828 -28180 -30812
rect -28284 -30892 -28264 -30828
rect -28200 -30892 -28180 -30828
rect -28284 -30908 -28180 -30892
rect -28284 -30972 -28264 -30908
rect -28200 -30972 -28180 -30908
rect -28284 -30988 -28180 -30972
rect -28284 -31052 -28264 -30988
rect -28200 -31052 -28180 -30988
rect -28284 -31068 -28180 -31052
rect -28284 -31132 -28264 -31068
rect -28200 -31132 -28180 -31068
rect -28284 -31148 -28180 -31132
rect -28284 -31212 -28264 -31148
rect -28200 -31212 -28180 -31148
rect -28284 -31228 -28180 -31212
rect -28284 -31292 -28264 -31228
rect -28200 -31292 -28180 -31228
rect -28284 -31308 -28180 -31292
rect -28284 -31372 -28264 -31308
rect -28200 -31372 -28180 -31308
rect -28284 -31388 -28180 -31372
rect -28284 -31452 -28264 -31388
rect -28200 -31452 -28180 -31388
rect -28284 -31468 -28180 -31452
rect -28284 -31532 -28264 -31468
rect -28200 -31532 -28180 -31468
rect -28284 -31548 -28180 -31532
rect -28284 -31612 -28264 -31548
rect -28200 -31612 -28180 -31548
rect -28284 -31628 -28180 -31612
rect -28284 -31692 -28264 -31628
rect -28200 -31692 -28180 -31628
rect -28284 -31708 -28180 -31692
rect -33896 -32068 -33792 -31772
rect -39085 -32148 -34163 -32119
rect -39085 -37012 -39056 -32148
rect -34192 -37012 -34163 -32148
rect -39085 -37041 -34163 -37012
rect -33896 -32132 -33876 -32068
rect -33812 -32132 -33792 -32068
rect -31064 -32119 -30960 -31721
rect -28284 -31772 -28264 -31708
rect -28200 -31772 -28180 -31708
rect -27861 -26828 -22939 -26799
rect -27861 -31692 -27832 -26828
rect -22968 -31692 -22939 -26828
rect -27861 -31721 -22939 -31692
rect -22672 -26812 -22652 -26748
rect -22588 -26812 -22568 -26748
rect -19840 -26799 -19736 -26401
rect -17060 -26452 -17040 -26388
rect -16976 -26452 -16956 -26388
rect -16637 -21508 -11715 -21479
rect -16637 -26372 -16608 -21508
rect -11744 -26372 -11715 -21508
rect -16637 -26401 -11715 -26372
rect -11448 -21492 -11428 -21428
rect -11364 -21492 -11344 -21428
rect -8616 -21479 -8512 -21081
rect -5836 -21132 -5816 -21068
rect -5752 -21132 -5732 -21068
rect -5413 -16188 -491 -16159
rect -5413 -21052 -5384 -16188
rect -520 -21052 -491 -16188
rect -5413 -21081 -491 -21052
rect -224 -16172 -204 -16108
rect -140 -16172 -120 -16108
rect 2608 -16159 2712 -15761
rect 5388 -15812 5408 -15748
rect 5472 -15812 5492 -15748
rect 5811 -10868 10733 -10839
rect 5811 -15732 5840 -10868
rect 10704 -15732 10733 -10868
rect 5811 -15761 10733 -15732
rect 11000 -10852 11020 -10788
rect 11084 -10852 11104 -10788
rect 13832 -10839 13936 -10441
rect 16612 -10492 16632 -10428
rect 16696 -10492 16716 -10428
rect 17035 -5548 21957 -5519
rect 17035 -10412 17064 -5548
rect 21928 -10412 21957 -5548
rect 17035 -10441 21957 -10412
rect 22224 -5532 22244 -5468
rect 22308 -5532 22328 -5468
rect 25056 -5519 25160 -5121
rect 27836 -5172 27856 -5108
rect 27920 -5172 27940 -5108
rect 28259 -228 33181 -199
rect 28259 -5092 28288 -228
rect 33152 -5092 33181 -228
rect 28259 -5121 33181 -5092
rect 33448 -212 33468 -148
rect 33532 -212 33552 -148
rect 36280 -199 36384 199
rect 39060 148 39080 212
rect 39144 148 39164 212
rect 39060 -148 39164 148
rect 33448 -228 33552 -212
rect 33448 -292 33468 -228
rect 33532 -292 33552 -228
rect 33448 -308 33552 -292
rect 33448 -372 33468 -308
rect 33532 -372 33552 -308
rect 33448 -388 33552 -372
rect 33448 -452 33468 -388
rect 33532 -452 33552 -388
rect 33448 -468 33552 -452
rect 33448 -532 33468 -468
rect 33532 -532 33552 -468
rect 33448 -548 33552 -532
rect 33448 -612 33468 -548
rect 33532 -612 33552 -548
rect 33448 -628 33552 -612
rect 33448 -692 33468 -628
rect 33532 -692 33552 -628
rect 33448 -708 33552 -692
rect 33448 -772 33468 -708
rect 33532 -772 33552 -708
rect 33448 -788 33552 -772
rect 33448 -852 33468 -788
rect 33532 -852 33552 -788
rect 33448 -868 33552 -852
rect 33448 -932 33468 -868
rect 33532 -932 33552 -868
rect 33448 -948 33552 -932
rect 33448 -1012 33468 -948
rect 33532 -1012 33552 -948
rect 33448 -1028 33552 -1012
rect 33448 -1092 33468 -1028
rect 33532 -1092 33552 -1028
rect 33448 -1108 33552 -1092
rect 33448 -1172 33468 -1108
rect 33532 -1172 33552 -1108
rect 33448 -1188 33552 -1172
rect 33448 -1252 33468 -1188
rect 33532 -1252 33552 -1188
rect 33448 -1268 33552 -1252
rect 33448 -1332 33468 -1268
rect 33532 -1332 33552 -1268
rect 33448 -1348 33552 -1332
rect 33448 -1412 33468 -1348
rect 33532 -1412 33552 -1348
rect 33448 -1428 33552 -1412
rect 33448 -1492 33468 -1428
rect 33532 -1492 33552 -1428
rect 33448 -1508 33552 -1492
rect 33448 -1572 33468 -1508
rect 33532 -1572 33552 -1508
rect 33448 -1588 33552 -1572
rect 33448 -1652 33468 -1588
rect 33532 -1652 33552 -1588
rect 33448 -1668 33552 -1652
rect 33448 -1732 33468 -1668
rect 33532 -1732 33552 -1668
rect 33448 -1748 33552 -1732
rect 33448 -1812 33468 -1748
rect 33532 -1812 33552 -1748
rect 33448 -1828 33552 -1812
rect 33448 -1892 33468 -1828
rect 33532 -1892 33552 -1828
rect 33448 -1908 33552 -1892
rect 33448 -1972 33468 -1908
rect 33532 -1972 33552 -1908
rect 33448 -1988 33552 -1972
rect 33448 -2052 33468 -1988
rect 33532 -2052 33552 -1988
rect 33448 -2068 33552 -2052
rect 33448 -2132 33468 -2068
rect 33532 -2132 33552 -2068
rect 33448 -2148 33552 -2132
rect 33448 -2212 33468 -2148
rect 33532 -2212 33552 -2148
rect 33448 -2228 33552 -2212
rect 33448 -2292 33468 -2228
rect 33532 -2292 33552 -2228
rect 33448 -2308 33552 -2292
rect 33448 -2372 33468 -2308
rect 33532 -2372 33552 -2308
rect 33448 -2388 33552 -2372
rect 33448 -2452 33468 -2388
rect 33532 -2452 33552 -2388
rect 33448 -2468 33552 -2452
rect 33448 -2532 33468 -2468
rect 33532 -2532 33552 -2468
rect 33448 -2548 33552 -2532
rect 33448 -2612 33468 -2548
rect 33532 -2612 33552 -2548
rect 33448 -2628 33552 -2612
rect 33448 -2692 33468 -2628
rect 33532 -2692 33552 -2628
rect 33448 -2708 33552 -2692
rect 33448 -2772 33468 -2708
rect 33532 -2772 33552 -2708
rect 33448 -2788 33552 -2772
rect 33448 -2852 33468 -2788
rect 33532 -2852 33552 -2788
rect 33448 -2868 33552 -2852
rect 33448 -2932 33468 -2868
rect 33532 -2932 33552 -2868
rect 33448 -2948 33552 -2932
rect 33448 -3012 33468 -2948
rect 33532 -3012 33552 -2948
rect 33448 -3028 33552 -3012
rect 33448 -3092 33468 -3028
rect 33532 -3092 33552 -3028
rect 33448 -3108 33552 -3092
rect 33448 -3172 33468 -3108
rect 33532 -3172 33552 -3108
rect 33448 -3188 33552 -3172
rect 33448 -3252 33468 -3188
rect 33532 -3252 33552 -3188
rect 33448 -3268 33552 -3252
rect 33448 -3332 33468 -3268
rect 33532 -3332 33552 -3268
rect 33448 -3348 33552 -3332
rect 33448 -3412 33468 -3348
rect 33532 -3412 33552 -3348
rect 33448 -3428 33552 -3412
rect 33448 -3492 33468 -3428
rect 33532 -3492 33552 -3428
rect 33448 -3508 33552 -3492
rect 33448 -3572 33468 -3508
rect 33532 -3572 33552 -3508
rect 33448 -3588 33552 -3572
rect 33448 -3652 33468 -3588
rect 33532 -3652 33552 -3588
rect 33448 -3668 33552 -3652
rect 33448 -3732 33468 -3668
rect 33532 -3732 33552 -3668
rect 33448 -3748 33552 -3732
rect 33448 -3812 33468 -3748
rect 33532 -3812 33552 -3748
rect 33448 -3828 33552 -3812
rect 33448 -3892 33468 -3828
rect 33532 -3892 33552 -3828
rect 33448 -3908 33552 -3892
rect 33448 -3972 33468 -3908
rect 33532 -3972 33552 -3908
rect 33448 -3988 33552 -3972
rect 33448 -4052 33468 -3988
rect 33532 -4052 33552 -3988
rect 33448 -4068 33552 -4052
rect 33448 -4132 33468 -4068
rect 33532 -4132 33552 -4068
rect 33448 -4148 33552 -4132
rect 33448 -4212 33468 -4148
rect 33532 -4212 33552 -4148
rect 33448 -4228 33552 -4212
rect 33448 -4292 33468 -4228
rect 33532 -4292 33552 -4228
rect 33448 -4308 33552 -4292
rect 33448 -4372 33468 -4308
rect 33532 -4372 33552 -4308
rect 33448 -4388 33552 -4372
rect 33448 -4452 33468 -4388
rect 33532 -4452 33552 -4388
rect 33448 -4468 33552 -4452
rect 33448 -4532 33468 -4468
rect 33532 -4532 33552 -4468
rect 33448 -4548 33552 -4532
rect 33448 -4612 33468 -4548
rect 33532 -4612 33552 -4548
rect 33448 -4628 33552 -4612
rect 33448 -4692 33468 -4628
rect 33532 -4692 33552 -4628
rect 33448 -4708 33552 -4692
rect 33448 -4772 33468 -4708
rect 33532 -4772 33552 -4708
rect 33448 -4788 33552 -4772
rect 33448 -4852 33468 -4788
rect 33532 -4852 33552 -4788
rect 33448 -4868 33552 -4852
rect 33448 -4932 33468 -4868
rect 33532 -4932 33552 -4868
rect 33448 -4948 33552 -4932
rect 33448 -5012 33468 -4948
rect 33532 -5012 33552 -4948
rect 33448 -5028 33552 -5012
rect 33448 -5092 33468 -5028
rect 33532 -5092 33552 -5028
rect 33448 -5108 33552 -5092
rect 27836 -5468 27940 -5172
rect 22224 -5548 22328 -5532
rect 22224 -5612 22244 -5548
rect 22308 -5612 22328 -5548
rect 22224 -5628 22328 -5612
rect 22224 -5692 22244 -5628
rect 22308 -5692 22328 -5628
rect 22224 -5708 22328 -5692
rect 22224 -5772 22244 -5708
rect 22308 -5772 22328 -5708
rect 22224 -5788 22328 -5772
rect 22224 -5852 22244 -5788
rect 22308 -5852 22328 -5788
rect 22224 -5868 22328 -5852
rect 22224 -5932 22244 -5868
rect 22308 -5932 22328 -5868
rect 22224 -5948 22328 -5932
rect 22224 -6012 22244 -5948
rect 22308 -6012 22328 -5948
rect 22224 -6028 22328 -6012
rect 22224 -6092 22244 -6028
rect 22308 -6092 22328 -6028
rect 22224 -6108 22328 -6092
rect 22224 -6172 22244 -6108
rect 22308 -6172 22328 -6108
rect 22224 -6188 22328 -6172
rect 22224 -6252 22244 -6188
rect 22308 -6252 22328 -6188
rect 22224 -6268 22328 -6252
rect 22224 -6332 22244 -6268
rect 22308 -6332 22328 -6268
rect 22224 -6348 22328 -6332
rect 22224 -6412 22244 -6348
rect 22308 -6412 22328 -6348
rect 22224 -6428 22328 -6412
rect 22224 -6492 22244 -6428
rect 22308 -6492 22328 -6428
rect 22224 -6508 22328 -6492
rect 22224 -6572 22244 -6508
rect 22308 -6572 22328 -6508
rect 22224 -6588 22328 -6572
rect 22224 -6652 22244 -6588
rect 22308 -6652 22328 -6588
rect 22224 -6668 22328 -6652
rect 22224 -6732 22244 -6668
rect 22308 -6732 22328 -6668
rect 22224 -6748 22328 -6732
rect 22224 -6812 22244 -6748
rect 22308 -6812 22328 -6748
rect 22224 -6828 22328 -6812
rect 22224 -6892 22244 -6828
rect 22308 -6892 22328 -6828
rect 22224 -6908 22328 -6892
rect 22224 -6972 22244 -6908
rect 22308 -6972 22328 -6908
rect 22224 -6988 22328 -6972
rect 22224 -7052 22244 -6988
rect 22308 -7052 22328 -6988
rect 22224 -7068 22328 -7052
rect 22224 -7132 22244 -7068
rect 22308 -7132 22328 -7068
rect 22224 -7148 22328 -7132
rect 22224 -7212 22244 -7148
rect 22308 -7212 22328 -7148
rect 22224 -7228 22328 -7212
rect 22224 -7292 22244 -7228
rect 22308 -7292 22328 -7228
rect 22224 -7308 22328 -7292
rect 22224 -7372 22244 -7308
rect 22308 -7372 22328 -7308
rect 22224 -7388 22328 -7372
rect 22224 -7452 22244 -7388
rect 22308 -7452 22328 -7388
rect 22224 -7468 22328 -7452
rect 22224 -7532 22244 -7468
rect 22308 -7532 22328 -7468
rect 22224 -7548 22328 -7532
rect 22224 -7612 22244 -7548
rect 22308 -7612 22328 -7548
rect 22224 -7628 22328 -7612
rect 22224 -7692 22244 -7628
rect 22308 -7692 22328 -7628
rect 22224 -7708 22328 -7692
rect 22224 -7772 22244 -7708
rect 22308 -7772 22328 -7708
rect 22224 -7788 22328 -7772
rect 22224 -7852 22244 -7788
rect 22308 -7852 22328 -7788
rect 22224 -7868 22328 -7852
rect 22224 -7932 22244 -7868
rect 22308 -7932 22328 -7868
rect 22224 -7948 22328 -7932
rect 22224 -8012 22244 -7948
rect 22308 -8012 22328 -7948
rect 22224 -8028 22328 -8012
rect 22224 -8092 22244 -8028
rect 22308 -8092 22328 -8028
rect 22224 -8108 22328 -8092
rect 22224 -8172 22244 -8108
rect 22308 -8172 22328 -8108
rect 22224 -8188 22328 -8172
rect 22224 -8252 22244 -8188
rect 22308 -8252 22328 -8188
rect 22224 -8268 22328 -8252
rect 22224 -8332 22244 -8268
rect 22308 -8332 22328 -8268
rect 22224 -8348 22328 -8332
rect 22224 -8412 22244 -8348
rect 22308 -8412 22328 -8348
rect 22224 -8428 22328 -8412
rect 22224 -8492 22244 -8428
rect 22308 -8492 22328 -8428
rect 22224 -8508 22328 -8492
rect 22224 -8572 22244 -8508
rect 22308 -8572 22328 -8508
rect 22224 -8588 22328 -8572
rect 22224 -8652 22244 -8588
rect 22308 -8652 22328 -8588
rect 22224 -8668 22328 -8652
rect 22224 -8732 22244 -8668
rect 22308 -8732 22328 -8668
rect 22224 -8748 22328 -8732
rect 22224 -8812 22244 -8748
rect 22308 -8812 22328 -8748
rect 22224 -8828 22328 -8812
rect 22224 -8892 22244 -8828
rect 22308 -8892 22328 -8828
rect 22224 -8908 22328 -8892
rect 22224 -8972 22244 -8908
rect 22308 -8972 22328 -8908
rect 22224 -8988 22328 -8972
rect 22224 -9052 22244 -8988
rect 22308 -9052 22328 -8988
rect 22224 -9068 22328 -9052
rect 22224 -9132 22244 -9068
rect 22308 -9132 22328 -9068
rect 22224 -9148 22328 -9132
rect 22224 -9212 22244 -9148
rect 22308 -9212 22328 -9148
rect 22224 -9228 22328 -9212
rect 22224 -9292 22244 -9228
rect 22308 -9292 22328 -9228
rect 22224 -9308 22328 -9292
rect 22224 -9372 22244 -9308
rect 22308 -9372 22328 -9308
rect 22224 -9388 22328 -9372
rect 22224 -9452 22244 -9388
rect 22308 -9452 22328 -9388
rect 22224 -9468 22328 -9452
rect 22224 -9532 22244 -9468
rect 22308 -9532 22328 -9468
rect 22224 -9548 22328 -9532
rect 22224 -9612 22244 -9548
rect 22308 -9612 22328 -9548
rect 22224 -9628 22328 -9612
rect 22224 -9692 22244 -9628
rect 22308 -9692 22328 -9628
rect 22224 -9708 22328 -9692
rect 22224 -9772 22244 -9708
rect 22308 -9772 22328 -9708
rect 22224 -9788 22328 -9772
rect 22224 -9852 22244 -9788
rect 22308 -9852 22328 -9788
rect 22224 -9868 22328 -9852
rect 22224 -9932 22244 -9868
rect 22308 -9932 22328 -9868
rect 22224 -9948 22328 -9932
rect 22224 -10012 22244 -9948
rect 22308 -10012 22328 -9948
rect 22224 -10028 22328 -10012
rect 22224 -10092 22244 -10028
rect 22308 -10092 22328 -10028
rect 22224 -10108 22328 -10092
rect 22224 -10172 22244 -10108
rect 22308 -10172 22328 -10108
rect 22224 -10188 22328 -10172
rect 22224 -10252 22244 -10188
rect 22308 -10252 22328 -10188
rect 22224 -10268 22328 -10252
rect 22224 -10332 22244 -10268
rect 22308 -10332 22328 -10268
rect 22224 -10348 22328 -10332
rect 22224 -10412 22244 -10348
rect 22308 -10412 22328 -10348
rect 22224 -10428 22328 -10412
rect 16612 -10788 16716 -10492
rect 11000 -10868 11104 -10852
rect 11000 -10932 11020 -10868
rect 11084 -10932 11104 -10868
rect 11000 -10948 11104 -10932
rect 11000 -11012 11020 -10948
rect 11084 -11012 11104 -10948
rect 11000 -11028 11104 -11012
rect 11000 -11092 11020 -11028
rect 11084 -11092 11104 -11028
rect 11000 -11108 11104 -11092
rect 11000 -11172 11020 -11108
rect 11084 -11172 11104 -11108
rect 11000 -11188 11104 -11172
rect 11000 -11252 11020 -11188
rect 11084 -11252 11104 -11188
rect 11000 -11268 11104 -11252
rect 11000 -11332 11020 -11268
rect 11084 -11332 11104 -11268
rect 11000 -11348 11104 -11332
rect 11000 -11412 11020 -11348
rect 11084 -11412 11104 -11348
rect 11000 -11428 11104 -11412
rect 11000 -11492 11020 -11428
rect 11084 -11492 11104 -11428
rect 11000 -11508 11104 -11492
rect 11000 -11572 11020 -11508
rect 11084 -11572 11104 -11508
rect 11000 -11588 11104 -11572
rect 11000 -11652 11020 -11588
rect 11084 -11652 11104 -11588
rect 11000 -11668 11104 -11652
rect 11000 -11732 11020 -11668
rect 11084 -11732 11104 -11668
rect 11000 -11748 11104 -11732
rect 11000 -11812 11020 -11748
rect 11084 -11812 11104 -11748
rect 11000 -11828 11104 -11812
rect 11000 -11892 11020 -11828
rect 11084 -11892 11104 -11828
rect 11000 -11908 11104 -11892
rect 11000 -11972 11020 -11908
rect 11084 -11972 11104 -11908
rect 11000 -11988 11104 -11972
rect 11000 -12052 11020 -11988
rect 11084 -12052 11104 -11988
rect 11000 -12068 11104 -12052
rect 11000 -12132 11020 -12068
rect 11084 -12132 11104 -12068
rect 11000 -12148 11104 -12132
rect 11000 -12212 11020 -12148
rect 11084 -12212 11104 -12148
rect 11000 -12228 11104 -12212
rect 11000 -12292 11020 -12228
rect 11084 -12292 11104 -12228
rect 11000 -12308 11104 -12292
rect 11000 -12372 11020 -12308
rect 11084 -12372 11104 -12308
rect 11000 -12388 11104 -12372
rect 11000 -12452 11020 -12388
rect 11084 -12452 11104 -12388
rect 11000 -12468 11104 -12452
rect 11000 -12532 11020 -12468
rect 11084 -12532 11104 -12468
rect 11000 -12548 11104 -12532
rect 11000 -12612 11020 -12548
rect 11084 -12612 11104 -12548
rect 11000 -12628 11104 -12612
rect 11000 -12692 11020 -12628
rect 11084 -12692 11104 -12628
rect 11000 -12708 11104 -12692
rect 11000 -12772 11020 -12708
rect 11084 -12772 11104 -12708
rect 11000 -12788 11104 -12772
rect 11000 -12852 11020 -12788
rect 11084 -12852 11104 -12788
rect 11000 -12868 11104 -12852
rect 11000 -12932 11020 -12868
rect 11084 -12932 11104 -12868
rect 11000 -12948 11104 -12932
rect 11000 -13012 11020 -12948
rect 11084 -13012 11104 -12948
rect 11000 -13028 11104 -13012
rect 11000 -13092 11020 -13028
rect 11084 -13092 11104 -13028
rect 11000 -13108 11104 -13092
rect 11000 -13172 11020 -13108
rect 11084 -13172 11104 -13108
rect 11000 -13188 11104 -13172
rect 11000 -13252 11020 -13188
rect 11084 -13252 11104 -13188
rect 11000 -13268 11104 -13252
rect 11000 -13332 11020 -13268
rect 11084 -13332 11104 -13268
rect 11000 -13348 11104 -13332
rect 11000 -13412 11020 -13348
rect 11084 -13412 11104 -13348
rect 11000 -13428 11104 -13412
rect 11000 -13492 11020 -13428
rect 11084 -13492 11104 -13428
rect 11000 -13508 11104 -13492
rect 11000 -13572 11020 -13508
rect 11084 -13572 11104 -13508
rect 11000 -13588 11104 -13572
rect 11000 -13652 11020 -13588
rect 11084 -13652 11104 -13588
rect 11000 -13668 11104 -13652
rect 11000 -13732 11020 -13668
rect 11084 -13732 11104 -13668
rect 11000 -13748 11104 -13732
rect 11000 -13812 11020 -13748
rect 11084 -13812 11104 -13748
rect 11000 -13828 11104 -13812
rect 11000 -13892 11020 -13828
rect 11084 -13892 11104 -13828
rect 11000 -13908 11104 -13892
rect 11000 -13972 11020 -13908
rect 11084 -13972 11104 -13908
rect 11000 -13988 11104 -13972
rect 11000 -14052 11020 -13988
rect 11084 -14052 11104 -13988
rect 11000 -14068 11104 -14052
rect 11000 -14132 11020 -14068
rect 11084 -14132 11104 -14068
rect 11000 -14148 11104 -14132
rect 11000 -14212 11020 -14148
rect 11084 -14212 11104 -14148
rect 11000 -14228 11104 -14212
rect 11000 -14292 11020 -14228
rect 11084 -14292 11104 -14228
rect 11000 -14308 11104 -14292
rect 11000 -14372 11020 -14308
rect 11084 -14372 11104 -14308
rect 11000 -14388 11104 -14372
rect 11000 -14452 11020 -14388
rect 11084 -14452 11104 -14388
rect 11000 -14468 11104 -14452
rect 11000 -14532 11020 -14468
rect 11084 -14532 11104 -14468
rect 11000 -14548 11104 -14532
rect 11000 -14612 11020 -14548
rect 11084 -14612 11104 -14548
rect 11000 -14628 11104 -14612
rect 11000 -14692 11020 -14628
rect 11084 -14692 11104 -14628
rect 11000 -14708 11104 -14692
rect 11000 -14772 11020 -14708
rect 11084 -14772 11104 -14708
rect 11000 -14788 11104 -14772
rect 11000 -14852 11020 -14788
rect 11084 -14852 11104 -14788
rect 11000 -14868 11104 -14852
rect 11000 -14932 11020 -14868
rect 11084 -14932 11104 -14868
rect 11000 -14948 11104 -14932
rect 11000 -15012 11020 -14948
rect 11084 -15012 11104 -14948
rect 11000 -15028 11104 -15012
rect 11000 -15092 11020 -15028
rect 11084 -15092 11104 -15028
rect 11000 -15108 11104 -15092
rect 11000 -15172 11020 -15108
rect 11084 -15172 11104 -15108
rect 11000 -15188 11104 -15172
rect 11000 -15252 11020 -15188
rect 11084 -15252 11104 -15188
rect 11000 -15268 11104 -15252
rect 11000 -15332 11020 -15268
rect 11084 -15332 11104 -15268
rect 11000 -15348 11104 -15332
rect 11000 -15412 11020 -15348
rect 11084 -15412 11104 -15348
rect 11000 -15428 11104 -15412
rect 11000 -15492 11020 -15428
rect 11084 -15492 11104 -15428
rect 11000 -15508 11104 -15492
rect 11000 -15572 11020 -15508
rect 11084 -15572 11104 -15508
rect 11000 -15588 11104 -15572
rect 11000 -15652 11020 -15588
rect 11084 -15652 11104 -15588
rect 11000 -15668 11104 -15652
rect 11000 -15732 11020 -15668
rect 11084 -15732 11104 -15668
rect 11000 -15748 11104 -15732
rect 5388 -16108 5492 -15812
rect -224 -16188 -120 -16172
rect -224 -16252 -204 -16188
rect -140 -16252 -120 -16188
rect -224 -16268 -120 -16252
rect -224 -16332 -204 -16268
rect -140 -16332 -120 -16268
rect -224 -16348 -120 -16332
rect -224 -16412 -204 -16348
rect -140 -16412 -120 -16348
rect -224 -16428 -120 -16412
rect -224 -16492 -204 -16428
rect -140 -16492 -120 -16428
rect -224 -16508 -120 -16492
rect -224 -16572 -204 -16508
rect -140 -16572 -120 -16508
rect -224 -16588 -120 -16572
rect -224 -16652 -204 -16588
rect -140 -16652 -120 -16588
rect -224 -16668 -120 -16652
rect -224 -16732 -204 -16668
rect -140 -16732 -120 -16668
rect -224 -16748 -120 -16732
rect -224 -16812 -204 -16748
rect -140 -16812 -120 -16748
rect -224 -16828 -120 -16812
rect -224 -16892 -204 -16828
rect -140 -16892 -120 -16828
rect -224 -16908 -120 -16892
rect -224 -16972 -204 -16908
rect -140 -16972 -120 -16908
rect -224 -16988 -120 -16972
rect -224 -17052 -204 -16988
rect -140 -17052 -120 -16988
rect -224 -17068 -120 -17052
rect -224 -17132 -204 -17068
rect -140 -17132 -120 -17068
rect -224 -17148 -120 -17132
rect -224 -17212 -204 -17148
rect -140 -17212 -120 -17148
rect -224 -17228 -120 -17212
rect -224 -17292 -204 -17228
rect -140 -17292 -120 -17228
rect -224 -17308 -120 -17292
rect -224 -17372 -204 -17308
rect -140 -17372 -120 -17308
rect -224 -17388 -120 -17372
rect -224 -17452 -204 -17388
rect -140 -17452 -120 -17388
rect -224 -17468 -120 -17452
rect -224 -17532 -204 -17468
rect -140 -17532 -120 -17468
rect -224 -17548 -120 -17532
rect -224 -17612 -204 -17548
rect -140 -17612 -120 -17548
rect -224 -17628 -120 -17612
rect -224 -17692 -204 -17628
rect -140 -17692 -120 -17628
rect -224 -17708 -120 -17692
rect -224 -17772 -204 -17708
rect -140 -17772 -120 -17708
rect -224 -17788 -120 -17772
rect -224 -17852 -204 -17788
rect -140 -17852 -120 -17788
rect -224 -17868 -120 -17852
rect -224 -17932 -204 -17868
rect -140 -17932 -120 -17868
rect -224 -17948 -120 -17932
rect -224 -18012 -204 -17948
rect -140 -18012 -120 -17948
rect -224 -18028 -120 -18012
rect -224 -18092 -204 -18028
rect -140 -18092 -120 -18028
rect -224 -18108 -120 -18092
rect -224 -18172 -204 -18108
rect -140 -18172 -120 -18108
rect -224 -18188 -120 -18172
rect -224 -18252 -204 -18188
rect -140 -18252 -120 -18188
rect -224 -18268 -120 -18252
rect -224 -18332 -204 -18268
rect -140 -18332 -120 -18268
rect -224 -18348 -120 -18332
rect -224 -18412 -204 -18348
rect -140 -18412 -120 -18348
rect -224 -18428 -120 -18412
rect -224 -18492 -204 -18428
rect -140 -18492 -120 -18428
rect -224 -18508 -120 -18492
rect -224 -18572 -204 -18508
rect -140 -18572 -120 -18508
rect -224 -18588 -120 -18572
rect -224 -18652 -204 -18588
rect -140 -18652 -120 -18588
rect -224 -18668 -120 -18652
rect -224 -18732 -204 -18668
rect -140 -18732 -120 -18668
rect -224 -18748 -120 -18732
rect -224 -18812 -204 -18748
rect -140 -18812 -120 -18748
rect -224 -18828 -120 -18812
rect -224 -18892 -204 -18828
rect -140 -18892 -120 -18828
rect -224 -18908 -120 -18892
rect -224 -18972 -204 -18908
rect -140 -18972 -120 -18908
rect -224 -18988 -120 -18972
rect -224 -19052 -204 -18988
rect -140 -19052 -120 -18988
rect -224 -19068 -120 -19052
rect -224 -19132 -204 -19068
rect -140 -19132 -120 -19068
rect -224 -19148 -120 -19132
rect -224 -19212 -204 -19148
rect -140 -19212 -120 -19148
rect -224 -19228 -120 -19212
rect -224 -19292 -204 -19228
rect -140 -19292 -120 -19228
rect -224 -19308 -120 -19292
rect -224 -19372 -204 -19308
rect -140 -19372 -120 -19308
rect -224 -19388 -120 -19372
rect -224 -19452 -204 -19388
rect -140 -19452 -120 -19388
rect -224 -19468 -120 -19452
rect -224 -19532 -204 -19468
rect -140 -19532 -120 -19468
rect -224 -19548 -120 -19532
rect -224 -19612 -204 -19548
rect -140 -19612 -120 -19548
rect -224 -19628 -120 -19612
rect -224 -19692 -204 -19628
rect -140 -19692 -120 -19628
rect -224 -19708 -120 -19692
rect -224 -19772 -204 -19708
rect -140 -19772 -120 -19708
rect -224 -19788 -120 -19772
rect -224 -19852 -204 -19788
rect -140 -19852 -120 -19788
rect -224 -19868 -120 -19852
rect -224 -19932 -204 -19868
rect -140 -19932 -120 -19868
rect -224 -19948 -120 -19932
rect -224 -20012 -204 -19948
rect -140 -20012 -120 -19948
rect -224 -20028 -120 -20012
rect -224 -20092 -204 -20028
rect -140 -20092 -120 -20028
rect -224 -20108 -120 -20092
rect -224 -20172 -204 -20108
rect -140 -20172 -120 -20108
rect -224 -20188 -120 -20172
rect -224 -20252 -204 -20188
rect -140 -20252 -120 -20188
rect -224 -20268 -120 -20252
rect -224 -20332 -204 -20268
rect -140 -20332 -120 -20268
rect -224 -20348 -120 -20332
rect -224 -20412 -204 -20348
rect -140 -20412 -120 -20348
rect -224 -20428 -120 -20412
rect -224 -20492 -204 -20428
rect -140 -20492 -120 -20428
rect -224 -20508 -120 -20492
rect -224 -20572 -204 -20508
rect -140 -20572 -120 -20508
rect -224 -20588 -120 -20572
rect -224 -20652 -204 -20588
rect -140 -20652 -120 -20588
rect -224 -20668 -120 -20652
rect -224 -20732 -204 -20668
rect -140 -20732 -120 -20668
rect -224 -20748 -120 -20732
rect -224 -20812 -204 -20748
rect -140 -20812 -120 -20748
rect -224 -20828 -120 -20812
rect -224 -20892 -204 -20828
rect -140 -20892 -120 -20828
rect -224 -20908 -120 -20892
rect -224 -20972 -204 -20908
rect -140 -20972 -120 -20908
rect -224 -20988 -120 -20972
rect -224 -21052 -204 -20988
rect -140 -21052 -120 -20988
rect -224 -21068 -120 -21052
rect -5836 -21428 -5732 -21132
rect -11448 -21508 -11344 -21492
rect -11448 -21572 -11428 -21508
rect -11364 -21572 -11344 -21508
rect -11448 -21588 -11344 -21572
rect -11448 -21652 -11428 -21588
rect -11364 -21652 -11344 -21588
rect -11448 -21668 -11344 -21652
rect -11448 -21732 -11428 -21668
rect -11364 -21732 -11344 -21668
rect -11448 -21748 -11344 -21732
rect -11448 -21812 -11428 -21748
rect -11364 -21812 -11344 -21748
rect -11448 -21828 -11344 -21812
rect -11448 -21892 -11428 -21828
rect -11364 -21892 -11344 -21828
rect -11448 -21908 -11344 -21892
rect -11448 -21972 -11428 -21908
rect -11364 -21972 -11344 -21908
rect -11448 -21988 -11344 -21972
rect -11448 -22052 -11428 -21988
rect -11364 -22052 -11344 -21988
rect -11448 -22068 -11344 -22052
rect -11448 -22132 -11428 -22068
rect -11364 -22132 -11344 -22068
rect -11448 -22148 -11344 -22132
rect -11448 -22212 -11428 -22148
rect -11364 -22212 -11344 -22148
rect -11448 -22228 -11344 -22212
rect -11448 -22292 -11428 -22228
rect -11364 -22292 -11344 -22228
rect -11448 -22308 -11344 -22292
rect -11448 -22372 -11428 -22308
rect -11364 -22372 -11344 -22308
rect -11448 -22388 -11344 -22372
rect -11448 -22452 -11428 -22388
rect -11364 -22452 -11344 -22388
rect -11448 -22468 -11344 -22452
rect -11448 -22532 -11428 -22468
rect -11364 -22532 -11344 -22468
rect -11448 -22548 -11344 -22532
rect -11448 -22612 -11428 -22548
rect -11364 -22612 -11344 -22548
rect -11448 -22628 -11344 -22612
rect -11448 -22692 -11428 -22628
rect -11364 -22692 -11344 -22628
rect -11448 -22708 -11344 -22692
rect -11448 -22772 -11428 -22708
rect -11364 -22772 -11344 -22708
rect -11448 -22788 -11344 -22772
rect -11448 -22852 -11428 -22788
rect -11364 -22852 -11344 -22788
rect -11448 -22868 -11344 -22852
rect -11448 -22932 -11428 -22868
rect -11364 -22932 -11344 -22868
rect -11448 -22948 -11344 -22932
rect -11448 -23012 -11428 -22948
rect -11364 -23012 -11344 -22948
rect -11448 -23028 -11344 -23012
rect -11448 -23092 -11428 -23028
rect -11364 -23092 -11344 -23028
rect -11448 -23108 -11344 -23092
rect -11448 -23172 -11428 -23108
rect -11364 -23172 -11344 -23108
rect -11448 -23188 -11344 -23172
rect -11448 -23252 -11428 -23188
rect -11364 -23252 -11344 -23188
rect -11448 -23268 -11344 -23252
rect -11448 -23332 -11428 -23268
rect -11364 -23332 -11344 -23268
rect -11448 -23348 -11344 -23332
rect -11448 -23412 -11428 -23348
rect -11364 -23412 -11344 -23348
rect -11448 -23428 -11344 -23412
rect -11448 -23492 -11428 -23428
rect -11364 -23492 -11344 -23428
rect -11448 -23508 -11344 -23492
rect -11448 -23572 -11428 -23508
rect -11364 -23572 -11344 -23508
rect -11448 -23588 -11344 -23572
rect -11448 -23652 -11428 -23588
rect -11364 -23652 -11344 -23588
rect -11448 -23668 -11344 -23652
rect -11448 -23732 -11428 -23668
rect -11364 -23732 -11344 -23668
rect -11448 -23748 -11344 -23732
rect -11448 -23812 -11428 -23748
rect -11364 -23812 -11344 -23748
rect -11448 -23828 -11344 -23812
rect -11448 -23892 -11428 -23828
rect -11364 -23892 -11344 -23828
rect -11448 -23908 -11344 -23892
rect -11448 -23972 -11428 -23908
rect -11364 -23972 -11344 -23908
rect -11448 -23988 -11344 -23972
rect -11448 -24052 -11428 -23988
rect -11364 -24052 -11344 -23988
rect -11448 -24068 -11344 -24052
rect -11448 -24132 -11428 -24068
rect -11364 -24132 -11344 -24068
rect -11448 -24148 -11344 -24132
rect -11448 -24212 -11428 -24148
rect -11364 -24212 -11344 -24148
rect -11448 -24228 -11344 -24212
rect -11448 -24292 -11428 -24228
rect -11364 -24292 -11344 -24228
rect -11448 -24308 -11344 -24292
rect -11448 -24372 -11428 -24308
rect -11364 -24372 -11344 -24308
rect -11448 -24388 -11344 -24372
rect -11448 -24452 -11428 -24388
rect -11364 -24452 -11344 -24388
rect -11448 -24468 -11344 -24452
rect -11448 -24532 -11428 -24468
rect -11364 -24532 -11344 -24468
rect -11448 -24548 -11344 -24532
rect -11448 -24612 -11428 -24548
rect -11364 -24612 -11344 -24548
rect -11448 -24628 -11344 -24612
rect -11448 -24692 -11428 -24628
rect -11364 -24692 -11344 -24628
rect -11448 -24708 -11344 -24692
rect -11448 -24772 -11428 -24708
rect -11364 -24772 -11344 -24708
rect -11448 -24788 -11344 -24772
rect -11448 -24852 -11428 -24788
rect -11364 -24852 -11344 -24788
rect -11448 -24868 -11344 -24852
rect -11448 -24932 -11428 -24868
rect -11364 -24932 -11344 -24868
rect -11448 -24948 -11344 -24932
rect -11448 -25012 -11428 -24948
rect -11364 -25012 -11344 -24948
rect -11448 -25028 -11344 -25012
rect -11448 -25092 -11428 -25028
rect -11364 -25092 -11344 -25028
rect -11448 -25108 -11344 -25092
rect -11448 -25172 -11428 -25108
rect -11364 -25172 -11344 -25108
rect -11448 -25188 -11344 -25172
rect -11448 -25252 -11428 -25188
rect -11364 -25252 -11344 -25188
rect -11448 -25268 -11344 -25252
rect -11448 -25332 -11428 -25268
rect -11364 -25332 -11344 -25268
rect -11448 -25348 -11344 -25332
rect -11448 -25412 -11428 -25348
rect -11364 -25412 -11344 -25348
rect -11448 -25428 -11344 -25412
rect -11448 -25492 -11428 -25428
rect -11364 -25492 -11344 -25428
rect -11448 -25508 -11344 -25492
rect -11448 -25572 -11428 -25508
rect -11364 -25572 -11344 -25508
rect -11448 -25588 -11344 -25572
rect -11448 -25652 -11428 -25588
rect -11364 -25652 -11344 -25588
rect -11448 -25668 -11344 -25652
rect -11448 -25732 -11428 -25668
rect -11364 -25732 -11344 -25668
rect -11448 -25748 -11344 -25732
rect -11448 -25812 -11428 -25748
rect -11364 -25812 -11344 -25748
rect -11448 -25828 -11344 -25812
rect -11448 -25892 -11428 -25828
rect -11364 -25892 -11344 -25828
rect -11448 -25908 -11344 -25892
rect -11448 -25972 -11428 -25908
rect -11364 -25972 -11344 -25908
rect -11448 -25988 -11344 -25972
rect -11448 -26052 -11428 -25988
rect -11364 -26052 -11344 -25988
rect -11448 -26068 -11344 -26052
rect -11448 -26132 -11428 -26068
rect -11364 -26132 -11344 -26068
rect -11448 -26148 -11344 -26132
rect -11448 -26212 -11428 -26148
rect -11364 -26212 -11344 -26148
rect -11448 -26228 -11344 -26212
rect -11448 -26292 -11428 -26228
rect -11364 -26292 -11344 -26228
rect -11448 -26308 -11344 -26292
rect -11448 -26372 -11428 -26308
rect -11364 -26372 -11344 -26308
rect -11448 -26388 -11344 -26372
rect -17060 -26748 -16956 -26452
rect -22672 -26828 -22568 -26812
rect -22672 -26892 -22652 -26828
rect -22588 -26892 -22568 -26828
rect -22672 -26908 -22568 -26892
rect -22672 -26972 -22652 -26908
rect -22588 -26972 -22568 -26908
rect -22672 -26988 -22568 -26972
rect -22672 -27052 -22652 -26988
rect -22588 -27052 -22568 -26988
rect -22672 -27068 -22568 -27052
rect -22672 -27132 -22652 -27068
rect -22588 -27132 -22568 -27068
rect -22672 -27148 -22568 -27132
rect -22672 -27212 -22652 -27148
rect -22588 -27212 -22568 -27148
rect -22672 -27228 -22568 -27212
rect -22672 -27292 -22652 -27228
rect -22588 -27292 -22568 -27228
rect -22672 -27308 -22568 -27292
rect -22672 -27372 -22652 -27308
rect -22588 -27372 -22568 -27308
rect -22672 -27388 -22568 -27372
rect -22672 -27452 -22652 -27388
rect -22588 -27452 -22568 -27388
rect -22672 -27468 -22568 -27452
rect -22672 -27532 -22652 -27468
rect -22588 -27532 -22568 -27468
rect -22672 -27548 -22568 -27532
rect -22672 -27612 -22652 -27548
rect -22588 -27612 -22568 -27548
rect -22672 -27628 -22568 -27612
rect -22672 -27692 -22652 -27628
rect -22588 -27692 -22568 -27628
rect -22672 -27708 -22568 -27692
rect -22672 -27772 -22652 -27708
rect -22588 -27772 -22568 -27708
rect -22672 -27788 -22568 -27772
rect -22672 -27852 -22652 -27788
rect -22588 -27852 -22568 -27788
rect -22672 -27868 -22568 -27852
rect -22672 -27932 -22652 -27868
rect -22588 -27932 -22568 -27868
rect -22672 -27948 -22568 -27932
rect -22672 -28012 -22652 -27948
rect -22588 -28012 -22568 -27948
rect -22672 -28028 -22568 -28012
rect -22672 -28092 -22652 -28028
rect -22588 -28092 -22568 -28028
rect -22672 -28108 -22568 -28092
rect -22672 -28172 -22652 -28108
rect -22588 -28172 -22568 -28108
rect -22672 -28188 -22568 -28172
rect -22672 -28252 -22652 -28188
rect -22588 -28252 -22568 -28188
rect -22672 -28268 -22568 -28252
rect -22672 -28332 -22652 -28268
rect -22588 -28332 -22568 -28268
rect -22672 -28348 -22568 -28332
rect -22672 -28412 -22652 -28348
rect -22588 -28412 -22568 -28348
rect -22672 -28428 -22568 -28412
rect -22672 -28492 -22652 -28428
rect -22588 -28492 -22568 -28428
rect -22672 -28508 -22568 -28492
rect -22672 -28572 -22652 -28508
rect -22588 -28572 -22568 -28508
rect -22672 -28588 -22568 -28572
rect -22672 -28652 -22652 -28588
rect -22588 -28652 -22568 -28588
rect -22672 -28668 -22568 -28652
rect -22672 -28732 -22652 -28668
rect -22588 -28732 -22568 -28668
rect -22672 -28748 -22568 -28732
rect -22672 -28812 -22652 -28748
rect -22588 -28812 -22568 -28748
rect -22672 -28828 -22568 -28812
rect -22672 -28892 -22652 -28828
rect -22588 -28892 -22568 -28828
rect -22672 -28908 -22568 -28892
rect -22672 -28972 -22652 -28908
rect -22588 -28972 -22568 -28908
rect -22672 -28988 -22568 -28972
rect -22672 -29052 -22652 -28988
rect -22588 -29052 -22568 -28988
rect -22672 -29068 -22568 -29052
rect -22672 -29132 -22652 -29068
rect -22588 -29132 -22568 -29068
rect -22672 -29148 -22568 -29132
rect -22672 -29212 -22652 -29148
rect -22588 -29212 -22568 -29148
rect -22672 -29228 -22568 -29212
rect -22672 -29292 -22652 -29228
rect -22588 -29292 -22568 -29228
rect -22672 -29308 -22568 -29292
rect -22672 -29372 -22652 -29308
rect -22588 -29372 -22568 -29308
rect -22672 -29388 -22568 -29372
rect -22672 -29452 -22652 -29388
rect -22588 -29452 -22568 -29388
rect -22672 -29468 -22568 -29452
rect -22672 -29532 -22652 -29468
rect -22588 -29532 -22568 -29468
rect -22672 -29548 -22568 -29532
rect -22672 -29612 -22652 -29548
rect -22588 -29612 -22568 -29548
rect -22672 -29628 -22568 -29612
rect -22672 -29692 -22652 -29628
rect -22588 -29692 -22568 -29628
rect -22672 -29708 -22568 -29692
rect -22672 -29772 -22652 -29708
rect -22588 -29772 -22568 -29708
rect -22672 -29788 -22568 -29772
rect -22672 -29852 -22652 -29788
rect -22588 -29852 -22568 -29788
rect -22672 -29868 -22568 -29852
rect -22672 -29932 -22652 -29868
rect -22588 -29932 -22568 -29868
rect -22672 -29948 -22568 -29932
rect -22672 -30012 -22652 -29948
rect -22588 -30012 -22568 -29948
rect -22672 -30028 -22568 -30012
rect -22672 -30092 -22652 -30028
rect -22588 -30092 -22568 -30028
rect -22672 -30108 -22568 -30092
rect -22672 -30172 -22652 -30108
rect -22588 -30172 -22568 -30108
rect -22672 -30188 -22568 -30172
rect -22672 -30252 -22652 -30188
rect -22588 -30252 -22568 -30188
rect -22672 -30268 -22568 -30252
rect -22672 -30332 -22652 -30268
rect -22588 -30332 -22568 -30268
rect -22672 -30348 -22568 -30332
rect -22672 -30412 -22652 -30348
rect -22588 -30412 -22568 -30348
rect -22672 -30428 -22568 -30412
rect -22672 -30492 -22652 -30428
rect -22588 -30492 -22568 -30428
rect -22672 -30508 -22568 -30492
rect -22672 -30572 -22652 -30508
rect -22588 -30572 -22568 -30508
rect -22672 -30588 -22568 -30572
rect -22672 -30652 -22652 -30588
rect -22588 -30652 -22568 -30588
rect -22672 -30668 -22568 -30652
rect -22672 -30732 -22652 -30668
rect -22588 -30732 -22568 -30668
rect -22672 -30748 -22568 -30732
rect -22672 -30812 -22652 -30748
rect -22588 -30812 -22568 -30748
rect -22672 -30828 -22568 -30812
rect -22672 -30892 -22652 -30828
rect -22588 -30892 -22568 -30828
rect -22672 -30908 -22568 -30892
rect -22672 -30972 -22652 -30908
rect -22588 -30972 -22568 -30908
rect -22672 -30988 -22568 -30972
rect -22672 -31052 -22652 -30988
rect -22588 -31052 -22568 -30988
rect -22672 -31068 -22568 -31052
rect -22672 -31132 -22652 -31068
rect -22588 -31132 -22568 -31068
rect -22672 -31148 -22568 -31132
rect -22672 -31212 -22652 -31148
rect -22588 -31212 -22568 -31148
rect -22672 -31228 -22568 -31212
rect -22672 -31292 -22652 -31228
rect -22588 -31292 -22568 -31228
rect -22672 -31308 -22568 -31292
rect -22672 -31372 -22652 -31308
rect -22588 -31372 -22568 -31308
rect -22672 -31388 -22568 -31372
rect -22672 -31452 -22652 -31388
rect -22588 -31452 -22568 -31388
rect -22672 -31468 -22568 -31452
rect -22672 -31532 -22652 -31468
rect -22588 -31532 -22568 -31468
rect -22672 -31548 -22568 -31532
rect -22672 -31612 -22652 -31548
rect -22588 -31612 -22568 -31548
rect -22672 -31628 -22568 -31612
rect -22672 -31692 -22652 -31628
rect -22588 -31692 -22568 -31628
rect -22672 -31708 -22568 -31692
rect -28284 -32068 -28180 -31772
rect -33896 -32148 -33792 -32132
rect -33896 -32212 -33876 -32148
rect -33812 -32212 -33792 -32148
rect -33896 -32228 -33792 -32212
rect -33896 -32292 -33876 -32228
rect -33812 -32292 -33792 -32228
rect -33896 -32308 -33792 -32292
rect -33896 -32372 -33876 -32308
rect -33812 -32372 -33792 -32308
rect -33896 -32388 -33792 -32372
rect -33896 -32452 -33876 -32388
rect -33812 -32452 -33792 -32388
rect -33896 -32468 -33792 -32452
rect -33896 -32532 -33876 -32468
rect -33812 -32532 -33792 -32468
rect -33896 -32548 -33792 -32532
rect -33896 -32612 -33876 -32548
rect -33812 -32612 -33792 -32548
rect -33896 -32628 -33792 -32612
rect -33896 -32692 -33876 -32628
rect -33812 -32692 -33792 -32628
rect -33896 -32708 -33792 -32692
rect -33896 -32772 -33876 -32708
rect -33812 -32772 -33792 -32708
rect -33896 -32788 -33792 -32772
rect -33896 -32852 -33876 -32788
rect -33812 -32852 -33792 -32788
rect -33896 -32868 -33792 -32852
rect -33896 -32932 -33876 -32868
rect -33812 -32932 -33792 -32868
rect -33896 -32948 -33792 -32932
rect -33896 -33012 -33876 -32948
rect -33812 -33012 -33792 -32948
rect -33896 -33028 -33792 -33012
rect -33896 -33092 -33876 -33028
rect -33812 -33092 -33792 -33028
rect -33896 -33108 -33792 -33092
rect -33896 -33172 -33876 -33108
rect -33812 -33172 -33792 -33108
rect -33896 -33188 -33792 -33172
rect -33896 -33252 -33876 -33188
rect -33812 -33252 -33792 -33188
rect -33896 -33268 -33792 -33252
rect -33896 -33332 -33876 -33268
rect -33812 -33332 -33792 -33268
rect -33896 -33348 -33792 -33332
rect -33896 -33412 -33876 -33348
rect -33812 -33412 -33792 -33348
rect -33896 -33428 -33792 -33412
rect -33896 -33492 -33876 -33428
rect -33812 -33492 -33792 -33428
rect -33896 -33508 -33792 -33492
rect -33896 -33572 -33876 -33508
rect -33812 -33572 -33792 -33508
rect -33896 -33588 -33792 -33572
rect -33896 -33652 -33876 -33588
rect -33812 -33652 -33792 -33588
rect -33896 -33668 -33792 -33652
rect -33896 -33732 -33876 -33668
rect -33812 -33732 -33792 -33668
rect -33896 -33748 -33792 -33732
rect -33896 -33812 -33876 -33748
rect -33812 -33812 -33792 -33748
rect -33896 -33828 -33792 -33812
rect -33896 -33892 -33876 -33828
rect -33812 -33892 -33792 -33828
rect -33896 -33908 -33792 -33892
rect -33896 -33972 -33876 -33908
rect -33812 -33972 -33792 -33908
rect -33896 -33988 -33792 -33972
rect -33896 -34052 -33876 -33988
rect -33812 -34052 -33792 -33988
rect -33896 -34068 -33792 -34052
rect -33896 -34132 -33876 -34068
rect -33812 -34132 -33792 -34068
rect -33896 -34148 -33792 -34132
rect -33896 -34212 -33876 -34148
rect -33812 -34212 -33792 -34148
rect -33896 -34228 -33792 -34212
rect -33896 -34292 -33876 -34228
rect -33812 -34292 -33792 -34228
rect -33896 -34308 -33792 -34292
rect -33896 -34372 -33876 -34308
rect -33812 -34372 -33792 -34308
rect -33896 -34388 -33792 -34372
rect -33896 -34452 -33876 -34388
rect -33812 -34452 -33792 -34388
rect -33896 -34468 -33792 -34452
rect -33896 -34532 -33876 -34468
rect -33812 -34532 -33792 -34468
rect -33896 -34548 -33792 -34532
rect -33896 -34612 -33876 -34548
rect -33812 -34612 -33792 -34548
rect -33896 -34628 -33792 -34612
rect -33896 -34692 -33876 -34628
rect -33812 -34692 -33792 -34628
rect -33896 -34708 -33792 -34692
rect -33896 -34772 -33876 -34708
rect -33812 -34772 -33792 -34708
rect -33896 -34788 -33792 -34772
rect -33896 -34852 -33876 -34788
rect -33812 -34852 -33792 -34788
rect -33896 -34868 -33792 -34852
rect -33896 -34932 -33876 -34868
rect -33812 -34932 -33792 -34868
rect -33896 -34948 -33792 -34932
rect -33896 -35012 -33876 -34948
rect -33812 -35012 -33792 -34948
rect -33896 -35028 -33792 -35012
rect -33896 -35092 -33876 -35028
rect -33812 -35092 -33792 -35028
rect -33896 -35108 -33792 -35092
rect -33896 -35172 -33876 -35108
rect -33812 -35172 -33792 -35108
rect -33896 -35188 -33792 -35172
rect -33896 -35252 -33876 -35188
rect -33812 -35252 -33792 -35188
rect -33896 -35268 -33792 -35252
rect -33896 -35332 -33876 -35268
rect -33812 -35332 -33792 -35268
rect -33896 -35348 -33792 -35332
rect -33896 -35412 -33876 -35348
rect -33812 -35412 -33792 -35348
rect -33896 -35428 -33792 -35412
rect -33896 -35492 -33876 -35428
rect -33812 -35492 -33792 -35428
rect -33896 -35508 -33792 -35492
rect -33896 -35572 -33876 -35508
rect -33812 -35572 -33792 -35508
rect -33896 -35588 -33792 -35572
rect -33896 -35652 -33876 -35588
rect -33812 -35652 -33792 -35588
rect -33896 -35668 -33792 -35652
rect -33896 -35732 -33876 -35668
rect -33812 -35732 -33792 -35668
rect -33896 -35748 -33792 -35732
rect -33896 -35812 -33876 -35748
rect -33812 -35812 -33792 -35748
rect -33896 -35828 -33792 -35812
rect -33896 -35892 -33876 -35828
rect -33812 -35892 -33792 -35828
rect -33896 -35908 -33792 -35892
rect -33896 -35972 -33876 -35908
rect -33812 -35972 -33792 -35908
rect -33896 -35988 -33792 -35972
rect -33896 -36052 -33876 -35988
rect -33812 -36052 -33792 -35988
rect -33896 -36068 -33792 -36052
rect -33896 -36132 -33876 -36068
rect -33812 -36132 -33792 -36068
rect -33896 -36148 -33792 -36132
rect -33896 -36212 -33876 -36148
rect -33812 -36212 -33792 -36148
rect -33896 -36228 -33792 -36212
rect -33896 -36292 -33876 -36228
rect -33812 -36292 -33792 -36228
rect -33896 -36308 -33792 -36292
rect -33896 -36372 -33876 -36308
rect -33812 -36372 -33792 -36308
rect -33896 -36388 -33792 -36372
rect -33896 -36452 -33876 -36388
rect -33812 -36452 -33792 -36388
rect -33896 -36468 -33792 -36452
rect -33896 -36532 -33876 -36468
rect -33812 -36532 -33792 -36468
rect -33896 -36548 -33792 -36532
rect -33896 -36612 -33876 -36548
rect -33812 -36612 -33792 -36548
rect -33896 -36628 -33792 -36612
rect -33896 -36692 -33876 -36628
rect -33812 -36692 -33792 -36628
rect -33896 -36708 -33792 -36692
rect -33896 -36772 -33876 -36708
rect -33812 -36772 -33792 -36708
rect -33896 -36788 -33792 -36772
rect -33896 -36852 -33876 -36788
rect -33812 -36852 -33792 -36788
rect -33896 -36868 -33792 -36852
rect -33896 -36932 -33876 -36868
rect -33812 -36932 -33792 -36868
rect -33896 -36948 -33792 -36932
rect -33896 -37012 -33876 -36948
rect -33812 -37012 -33792 -36948
rect -33896 -37028 -33792 -37012
rect -36676 -37240 -36572 -37041
rect -33896 -37092 -33876 -37028
rect -33812 -37092 -33792 -37028
rect -33473 -32148 -28551 -32119
rect -33473 -37012 -33444 -32148
rect -28580 -37012 -28551 -32148
rect -33473 -37041 -28551 -37012
rect -28284 -32132 -28264 -32068
rect -28200 -32132 -28180 -32068
rect -25452 -32119 -25348 -31721
rect -22672 -31772 -22652 -31708
rect -22588 -31772 -22568 -31708
rect -22249 -26828 -17327 -26799
rect -22249 -31692 -22220 -26828
rect -17356 -31692 -17327 -26828
rect -22249 -31721 -17327 -31692
rect -17060 -26812 -17040 -26748
rect -16976 -26812 -16956 -26748
rect -14228 -26799 -14124 -26401
rect -11448 -26452 -11428 -26388
rect -11364 -26452 -11344 -26388
rect -11025 -21508 -6103 -21479
rect -11025 -26372 -10996 -21508
rect -6132 -26372 -6103 -21508
rect -11025 -26401 -6103 -26372
rect -5836 -21492 -5816 -21428
rect -5752 -21492 -5732 -21428
rect -3004 -21479 -2900 -21081
rect -224 -21132 -204 -21068
rect -140 -21132 -120 -21068
rect 199 -16188 5121 -16159
rect 199 -21052 228 -16188
rect 5092 -21052 5121 -16188
rect 199 -21081 5121 -21052
rect 5388 -16172 5408 -16108
rect 5472 -16172 5492 -16108
rect 8220 -16159 8324 -15761
rect 11000 -15812 11020 -15748
rect 11084 -15812 11104 -15748
rect 11423 -10868 16345 -10839
rect 11423 -15732 11452 -10868
rect 16316 -15732 16345 -10868
rect 11423 -15761 16345 -15732
rect 16612 -10852 16632 -10788
rect 16696 -10852 16716 -10788
rect 19444 -10839 19548 -10441
rect 22224 -10492 22244 -10428
rect 22308 -10492 22328 -10428
rect 22647 -5548 27569 -5519
rect 22647 -10412 22676 -5548
rect 27540 -10412 27569 -5548
rect 22647 -10441 27569 -10412
rect 27836 -5532 27856 -5468
rect 27920 -5532 27940 -5468
rect 30668 -5519 30772 -5121
rect 33448 -5172 33468 -5108
rect 33532 -5172 33552 -5108
rect 33871 -228 38793 -199
rect 33871 -5092 33900 -228
rect 38764 -5092 38793 -228
rect 33871 -5121 38793 -5092
rect 39060 -212 39080 -148
rect 39144 -212 39164 -148
rect 39060 -228 39164 -212
rect 39060 -292 39080 -228
rect 39144 -292 39164 -228
rect 39060 -308 39164 -292
rect 39060 -372 39080 -308
rect 39144 -372 39164 -308
rect 39060 -388 39164 -372
rect 39060 -452 39080 -388
rect 39144 -452 39164 -388
rect 39060 -468 39164 -452
rect 39060 -532 39080 -468
rect 39144 -532 39164 -468
rect 39060 -548 39164 -532
rect 39060 -612 39080 -548
rect 39144 -612 39164 -548
rect 39060 -628 39164 -612
rect 39060 -692 39080 -628
rect 39144 -692 39164 -628
rect 39060 -708 39164 -692
rect 39060 -772 39080 -708
rect 39144 -772 39164 -708
rect 39060 -788 39164 -772
rect 39060 -852 39080 -788
rect 39144 -852 39164 -788
rect 39060 -868 39164 -852
rect 39060 -932 39080 -868
rect 39144 -932 39164 -868
rect 39060 -948 39164 -932
rect 39060 -1012 39080 -948
rect 39144 -1012 39164 -948
rect 39060 -1028 39164 -1012
rect 39060 -1092 39080 -1028
rect 39144 -1092 39164 -1028
rect 39060 -1108 39164 -1092
rect 39060 -1172 39080 -1108
rect 39144 -1172 39164 -1108
rect 39060 -1188 39164 -1172
rect 39060 -1252 39080 -1188
rect 39144 -1252 39164 -1188
rect 39060 -1268 39164 -1252
rect 39060 -1332 39080 -1268
rect 39144 -1332 39164 -1268
rect 39060 -1348 39164 -1332
rect 39060 -1412 39080 -1348
rect 39144 -1412 39164 -1348
rect 39060 -1428 39164 -1412
rect 39060 -1492 39080 -1428
rect 39144 -1492 39164 -1428
rect 39060 -1508 39164 -1492
rect 39060 -1572 39080 -1508
rect 39144 -1572 39164 -1508
rect 39060 -1588 39164 -1572
rect 39060 -1652 39080 -1588
rect 39144 -1652 39164 -1588
rect 39060 -1668 39164 -1652
rect 39060 -1732 39080 -1668
rect 39144 -1732 39164 -1668
rect 39060 -1748 39164 -1732
rect 39060 -1812 39080 -1748
rect 39144 -1812 39164 -1748
rect 39060 -1828 39164 -1812
rect 39060 -1892 39080 -1828
rect 39144 -1892 39164 -1828
rect 39060 -1908 39164 -1892
rect 39060 -1972 39080 -1908
rect 39144 -1972 39164 -1908
rect 39060 -1988 39164 -1972
rect 39060 -2052 39080 -1988
rect 39144 -2052 39164 -1988
rect 39060 -2068 39164 -2052
rect 39060 -2132 39080 -2068
rect 39144 -2132 39164 -2068
rect 39060 -2148 39164 -2132
rect 39060 -2212 39080 -2148
rect 39144 -2212 39164 -2148
rect 39060 -2228 39164 -2212
rect 39060 -2292 39080 -2228
rect 39144 -2292 39164 -2228
rect 39060 -2308 39164 -2292
rect 39060 -2372 39080 -2308
rect 39144 -2372 39164 -2308
rect 39060 -2388 39164 -2372
rect 39060 -2452 39080 -2388
rect 39144 -2452 39164 -2388
rect 39060 -2468 39164 -2452
rect 39060 -2532 39080 -2468
rect 39144 -2532 39164 -2468
rect 39060 -2548 39164 -2532
rect 39060 -2612 39080 -2548
rect 39144 -2612 39164 -2548
rect 39060 -2628 39164 -2612
rect 39060 -2692 39080 -2628
rect 39144 -2692 39164 -2628
rect 39060 -2708 39164 -2692
rect 39060 -2772 39080 -2708
rect 39144 -2772 39164 -2708
rect 39060 -2788 39164 -2772
rect 39060 -2852 39080 -2788
rect 39144 -2852 39164 -2788
rect 39060 -2868 39164 -2852
rect 39060 -2932 39080 -2868
rect 39144 -2932 39164 -2868
rect 39060 -2948 39164 -2932
rect 39060 -3012 39080 -2948
rect 39144 -3012 39164 -2948
rect 39060 -3028 39164 -3012
rect 39060 -3092 39080 -3028
rect 39144 -3092 39164 -3028
rect 39060 -3108 39164 -3092
rect 39060 -3172 39080 -3108
rect 39144 -3172 39164 -3108
rect 39060 -3188 39164 -3172
rect 39060 -3252 39080 -3188
rect 39144 -3252 39164 -3188
rect 39060 -3268 39164 -3252
rect 39060 -3332 39080 -3268
rect 39144 -3332 39164 -3268
rect 39060 -3348 39164 -3332
rect 39060 -3412 39080 -3348
rect 39144 -3412 39164 -3348
rect 39060 -3428 39164 -3412
rect 39060 -3492 39080 -3428
rect 39144 -3492 39164 -3428
rect 39060 -3508 39164 -3492
rect 39060 -3572 39080 -3508
rect 39144 -3572 39164 -3508
rect 39060 -3588 39164 -3572
rect 39060 -3652 39080 -3588
rect 39144 -3652 39164 -3588
rect 39060 -3668 39164 -3652
rect 39060 -3732 39080 -3668
rect 39144 -3732 39164 -3668
rect 39060 -3748 39164 -3732
rect 39060 -3812 39080 -3748
rect 39144 -3812 39164 -3748
rect 39060 -3828 39164 -3812
rect 39060 -3892 39080 -3828
rect 39144 -3892 39164 -3828
rect 39060 -3908 39164 -3892
rect 39060 -3972 39080 -3908
rect 39144 -3972 39164 -3908
rect 39060 -3988 39164 -3972
rect 39060 -4052 39080 -3988
rect 39144 -4052 39164 -3988
rect 39060 -4068 39164 -4052
rect 39060 -4132 39080 -4068
rect 39144 -4132 39164 -4068
rect 39060 -4148 39164 -4132
rect 39060 -4212 39080 -4148
rect 39144 -4212 39164 -4148
rect 39060 -4228 39164 -4212
rect 39060 -4292 39080 -4228
rect 39144 -4292 39164 -4228
rect 39060 -4308 39164 -4292
rect 39060 -4372 39080 -4308
rect 39144 -4372 39164 -4308
rect 39060 -4388 39164 -4372
rect 39060 -4452 39080 -4388
rect 39144 -4452 39164 -4388
rect 39060 -4468 39164 -4452
rect 39060 -4532 39080 -4468
rect 39144 -4532 39164 -4468
rect 39060 -4548 39164 -4532
rect 39060 -4612 39080 -4548
rect 39144 -4612 39164 -4548
rect 39060 -4628 39164 -4612
rect 39060 -4692 39080 -4628
rect 39144 -4692 39164 -4628
rect 39060 -4708 39164 -4692
rect 39060 -4772 39080 -4708
rect 39144 -4772 39164 -4708
rect 39060 -4788 39164 -4772
rect 39060 -4852 39080 -4788
rect 39144 -4852 39164 -4788
rect 39060 -4868 39164 -4852
rect 39060 -4932 39080 -4868
rect 39144 -4932 39164 -4868
rect 39060 -4948 39164 -4932
rect 39060 -5012 39080 -4948
rect 39144 -5012 39164 -4948
rect 39060 -5028 39164 -5012
rect 39060 -5092 39080 -5028
rect 39144 -5092 39164 -5028
rect 39060 -5108 39164 -5092
rect 33448 -5468 33552 -5172
rect 27836 -5548 27940 -5532
rect 27836 -5612 27856 -5548
rect 27920 -5612 27940 -5548
rect 27836 -5628 27940 -5612
rect 27836 -5692 27856 -5628
rect 27920 -5692 27940 -5628
rect 27836 -5708 27940 -5692
rect 27836 -5772 27856 -5708
rect 27920 -5772 27940 -5708
rect 27836 -5788 27940 -5772
rect 27836 -5852 27856 -5788
rect 27920 -5852 27940 -5788
rect 27836 -5868 27940 -5852
rect 27836 -5932 27856 -5868
rect 27920 -5932 27940 -5868
rect 27836 -5948 27940 -5932
rect 27836 -6012 27856 -5948
rect 27920 -6012 27940 -5948
rect 27836 -6028 27940 -6012
rect 27836 -6092 27856 -6028
rect 27920 -6092 27940 -6028
rect 27836 -6108 27940 -6092
rect 27836 -6172 27856 -6108
rect 27920 -6172 27940 -6108
rect 27836 -6188 27940 -6172
rect 27836 -6252 27856 -6188
rect 27920 -6252 27940 -6188
rect 27836 -6268 27940 -6252
rect 27836 -6332 27856 -6268
rect 27920 -6332 27940 -6268
rect 27836 -6348 27940 -6332
rect 27836 -6412 27856 -6348
rect 27920 -6412 27940 -6348
rect 27836 -6428 27940 -6412
rect 27836 -6492 27856 -6428
rect 27920 -6492 27940 -6428
rect 27836 -6508 27940 -6492
rect 27836 -6572 27856 -6508
rect 27920 -6572 27940 -6508
rect 27836 -6588 27940 -6572
rect 27836 -6652 27856 -6588
rect 27920 -6652 27940 -6588
rect 27836 -6668 27940 -6652
rect 27836 -6732 27856 -6668
rect 27920 -6732 27940 -6668
rect 27836 -6748 27940 -6732
rect 27836 -6812 27856 -6748
rect 27920 -6812 27940 -6748
rect 27836 -6828 27940 -6812
rect 27836 -6892 27856 -6828
rect 27920 -6892 27940 -6828
rect 27836 -6908 27940 -6892
rect 27836 -6972 27856 -6908
rect 27920 -6972 27940 -6908
rect 27836 -6988 27940 -6972
rect 27836 -7052 27856 -6988
rect 27920 -7052 27940 -6988
rect 27836 -7068 27940 -7052
rect 27836 -7132 27856 -7068
rect 27920 -7132 27940 -7068
rect 27836 -7148 27940 -7132
rect 27836 -7212 27856 -7148
rect 27920 -7212 27940 -7148
rect 27836 -7228 27940 -7212
rect 27836 -7292 27856 -7228
rect 27920 -7292 27940 -7228
rect 27836 -7308 27940 -7292
rect 27836 -7372 27856 -7308
rect 27920 -7372 27940 -7308
rect 27836 -7388 27940 -7372
rect 27836 -7452 27856 -7388
rect 27920 -7452 27940 -7388
rect 27836 -7468 27940 -7452
rect 27836 -7532 27856 -7468
rect 27920 -7532 27940 -7468
rect 27836 -7548 27940 -7532
rect 27836 -7612 27856 -7548
rect 27920 -7612 27940 -7548
rect 27836 -7628 27940 -7612
rect 27836 -7692 27856 -7628
rect 27920 -7692 27940 -7628
rect 27836 -7708 27940 -7692
rect 27836 -7772 27856 -7708
rect 27920 -7772 27940 -7708
rect 27836 -7788 27940 -7772
rect 27836 -7852 27856 -7788
rect 27920 -7852 27940 -7788
rect 27836 -7868 27940 -7852
rect 27836 -7932 27856 -7868
rect 27920 -7932 27940 -7868
rect 27836 -7948 27940 -7932
rect 27836 -8012 27856 -7948
rect 27920 -8012 27940 -7948
rect 27836 -8028 27940 -8012
rect 27836 -8092 27856 -8028
rect 27920 -8092 27940 -8028
rect 27836 -8108 27940 -8092
rect 27836 -8172 27856 -8108
rect 27920 -8172 27940 -8108
rect 27836 -8188 27940 -8172
rect 27836 -8252 27856 -8188
rect 27920 -8252 27940 -8188
rect 27836 -8268 27940 -8252
rect 27836 -8332 27856 -8268
rect 27920 -8332 27940 -8268
rect 27836 -8348 27940 -8332
rect 27836 -8412 27856 -8348
rect 27920 -8412 27940 -8348
rect 27836 -8428 27940 -8412
rect 27836 -8492 27856 -8428
rect 27920 -8492 27940 -8428
rect 27836 -8508 27940 -8492
rect 27836 -8572 27856 -8508
rect 27920 -8572 27940 -8508
rect 27836 -8588 27940 -8572
rect 27836 -8652 27856 -8588
rect 27920 -8652 27940 -8588
rect 27836 -8668 27940 -8652
rect 27836 -8732 27856 -8668
rect 27920 -8732 27940 -8668
rect 27836 -8748 27940 -8732
rect 27836 -8812 27856 -8748
rect 27920 -8812 27940 -8748
rect 27836 -8828 27940 -8812
rect 27836 -8892 27856 -8828
rect 27920 -8892 27940 -8828
rect 27836 -8908 27940 -8892
rect 27836 -8972 27856 -8908
rect 27920 -8972 27940 -8908
rect 27836 -8988 27940 -8972
rect 27836 -9052 27856 -8988
rect 27920 -9052 27940 -8988
rect 27836 -9068 27940 -9052
rect 27836 -9132 27856 -9068
rect 27920 -9132 27940 -9068
rect 27836 -9148 27940 -9132
rect 27836 -9212 27856 -9148
rect 27920 -9212 27940 -9148
rect 27836 -9228 27940 -9212
rect 27836 -9292 27856 -9228
rect 27920 -9292 27940 -9228
rect 27836 -9308 27940 -9292
rect 27836 -9372 27856 -9308
rect 27920 -9372 27940 -9308
rect 27836 -9388 27940 -9372
rect 27836 -9452 27856 -9388
rect 27920 -9452 27940 -9388
rect 27836 -9468 27940 -9452
rect 27836 -9532 27856 -9468
rect 27920 -9532 27940 -9468
rect 27836 -9548 27940 -9532
rect 27836 -9612 27856 -9548
rect 27920 -9612 27940 -9548
rect 27836 -9628 27940 -9612
rect 27836 -9692 27856 -9628
rect 27920 -9692 27940 -9628
rect 27836 -9708 27940 -9692
rect 27836 -9772 27856 -9708
rect 27920 -9772 27940 -9708
rect 27836 -9788 27940 -9772
rect 27836 -9852 27856 -9788
rect 27920 -9852 27940 -9788
rect 27836 -9868 27940 -9852
rect 27836 -9932 27856 -9868
rect 27920 -9932 27940 -9868
rect 27836 -9948 27940 -9932
rect 27836 -10012 27856 -9948
rect 27920 -10012 27940 -9948
rect 27836 -10028 27940 -10012
rect 27836 -10092 27856 -10028
rect 27920 -10092 27940 -10028
rect 27836 -10108 27940 -10092
rect 27836 -10172 27856 -10108
rect 27920 -10172 27940 -10108
rect 27836 -10188 27940 -10172
rect 27836 -10252 27856 -10188
rect 27920 -10252 27940 -10188
rect 27836 -10268 27940 -10252
rect 27836 -10332 27856 -10268
rect 27920 -10332 27940 -10268
rect 27836 -10348 27940 -10332
rect 27836 -10412 27856 -10348
rect 27920 -10412 27940 -10348
rect 27836 -10428 27940 -10412
rect 22224 -10788 22328 -10492
rect 16612 -10868 16716 -10852
rect 16612 -10932 16632 -10868
rect 16696 -10932 16716 -10868
rect 16612 -10948 16716 -10932
rect 16612 -11012 16632 -10948
rect 16696 -11012 16716 -10948
rect 16612 -11028 16716 -11012
rect 16612 -11092 16632 -11028
rect 16696 -11092 16716 -11028
rect 16612 -11108 16716 -11092
rect 16612 -11172 16632 -11108
rect 16696 -11172 16716 -11108
rect 16612 -11188 16716 -11172
rect 16612 -11252 16632 -11188
rect 16696 -11252 16716 -11188
rect 16612 -11268 16716 -11252
rect 16612 -11332 16632 -11268
rect 16696 -11332 16716 -11268
rect 16612 -11348 16716 -11332
rect 16612 -11412 16632 -11348
rect 16696 -11412 16716 -11348
rect 16612 -11428 16716 -11412
rect 16612 -11492 16632 -11428
rect 16696 -11492 16716 -11428
rect 16612 -11508 16716 -11492
rect 16612 -11572 16632 -11508
rect 16696 -11572 16716 -11508
rect 16612 -11588 16716 -11572
rect 16612 -11652 16632 -11588
rect 16696 -11652 16716 -11588
rect 16612 -11668 16716 -11652
rect 16612 -11732 16632 -11668
rect 16696 -11732 16716 -11668
rect 16612 -11748 16716 -11732
rect 16612 -11812 16632 -11748
rect 16696 -11812 16716 -11748
rect 16612 -11828 16716 -11812
rect 16612 -11892 16632 -11828
rect 16696 -11892 16716 -11828
rect 16612 -11908 16716 -11892
rect 16612 -11972 16632 -11908
rect 16696 -11972 16716 -11908
rect 16612 -11988 16716 -11972
rect 16612 -12052 16632 -11988
rect 16696 -12052 16716 -11988
rect 16612 -12068 16716 -12052
rect 16612 -12132 16632 -12068
rect 16696 -12132 16716 -12068
rect 16612 -12148 16716 -12132
rect 16612 -12212 16632 -12148
rect 16696 -12212 16716 -12148
rect 16612 -12228 16716 -12212
rect 16612 -12292 16632 -12228
rect 16696 -12292 16716 -12228
rect 16612 -12308 16716 -12292
rect 16612 -12372 16632 -12308
rect 16696 -12372 16716 -12308
rect 16612 -12388 16716 -12372
rect 16612 -12452 16632 -12388
rect 16696 -12452 16716 -12388
rect 16612 -12468 16716 -12452
rect 16612 -12532 16632 -12468
rect 16696 -12532 16716 -12468
rect 16612 -12548 16716 -12532
rect 16612 -12612 16632 -12548
rect 16696 -12612 16716 -12548
rect 16612 -12628 16716 -12612
rect 16612 -12692 16632 -12628
rect 16696 -12692 16716 -12628
rect 16612 -12708 16716 -12692
rect 16612 -12772 16632 -12708
rect 16696 -12772 16716 -12708
rect 16612 -12788 16716 -12772
rect 16612 -12852 16632 -12788
rect 16696 -12852 16716 -12788
rect 16612 -12868 16716 -12852
rect 16612 -12932 16632 -12868
rect 16696 -12932 16716 -12868
rect 16612 -12948 16716 -12932
rect 16612 -13012 16632 -12948
rect 16696 -13012 16716 -12948
rect 16612 -13028 16716 -13012
rect 16612 -13092 16632 -13028
rect 16696 -13092 16716 -13028
rect 16612 -13108 16716 -13092
rect 16612 -13172 16632 -13108
rect 16696 -13172 16716 -13108
rect 16612 -13188 16716 -13172
rect 16612 -13252 16632 -13188
rect 16696 -13252 16716 -13188
rect 16612 -13268 16716 -13252
rect 16612 -13332 16632 -13268
rect 16696 -13332 16716 -13268
rect 16612 -13348 16716 -13332
rect 16612 -13412 16632 -13348
rect 16696 -13412 16716 -13348
rect 16612 -13428 16716 -13412
rect 16612 -13492 16632 -13428
rect 16696 -13492 16716 -13428
rect 16612 -13508 16716 -13492
rect 16612 -13572 16632 -13508
rect 16696 -13572 16716 -13508
rect 16612 -13588 16716 -13572
rect 16612 -13652 16632 -13588
rect 16696 -13652 16716 -13588
rect 16612 -13668 16716 -13652
rect 16612 -13732 16632 -13668
rect 16696 -13732 16716 -13668
rect 16612 -13748 16716 -13732
rect 16612 -13812 16632 -13748
rect 16696 -13812 16716 -13748
rect 16612 -13828 16716 -13812
rect 16612 -13892 16632 -13828
rect 16696 -13892 16716 -13828
rect 16612 -13908 16716 -13892
rect 16612 -13972 16632 -13908
rect 16696 -13972 16716 -13908
rect 16612 -13988 16716 -13972
rect 16612 -14052 16632 -13988
rect 16696 -14052 16716 -13988
rect 16612 -14068 16716 -14052
rect 16612 -14132 16632 -14068
rect 16696 -14132 16716 -14068
rect 16612 -14148 16716 -14132
rect 16612 -14212 16632 -14148
rect 16696 -14212 16716 -14148
rect 16612 -14228 16716 -14212
rect 16612 -14292 16632 -14228
rect 16696 -14292 16716 -14228
rect 16612 -14308 16716 -14292
rect 16612 -14372 16632 -14308
rect 16696 -14372 16716 -14308
rect 16612 -14388 16716 -14372
rect 16612 -14452 16632 -14388
rect 16696 -14452 16716 -14388
rect 16612 -14468 16716 -14452
rect 16612 -14532 16632 -14468
rect 16696 -14532 16716 -14468
rect 16612 -14548 16716 -14532
rect 16612 -14612 16632 -14548
rect 16696 -14612 16716 -14548
rect 16612 -14628 16716 -14612
rect 16612 -14692 16632 -14628
rect 16696 -14692 16716 -14628
rect 16612 -14708 16716 -14692
rect 16612 -14772 16632 -14708
rect 16696 -14772 16716 -14708
rect 16612 -14788 16716 -14772
rect 16612 -14852 16632 -14788
rect 16696 -14852 16716 -14788
rect 16612 -14868 16716 -14852
rect 16612 -14932 16632 -14868
rect 16696 -14932 16716 -14868
rect 16612 -14948 16716 -14932
rect 16612 -15012 16632 -14948
rect 16696 -15012 16716 -14948
rect 16612 -15028 16716 -15012
rect 16612 -15092 16632 -15028
rect 16696 -15092 16716 -15028
rect 16612 -15108 16716 -15092
rect 16612 -15172 16632 -15108
rect 16696 -15172 16716 -15108
rect 16612 -15188 16716 -15172
rect 16612 -15252 16632 -15188
rect 16696 -15252 16716 -15188
rect 16612 -15268 16716 -15252
rect 16612 -15332 16632 -15268
rect 16696 -15332 16716 -15268
rect 16612 -15348 16716 -15332
rect 16612 -15412 16632 -15348
rect 16696 -15412 16716 -15348
rect 16612 -15428 16716 -15412
rect 16612 -15492 16632 -15428
rect 16696 -15492 16716 -15428
rect 16612 -15508 16716 -15492
rect 16612 -15572 16632 -15508
rect 16696 -15572 16716 -15508
rect 16612 -15588 16716 -15572
rect 16612 -15652 16632 -15588
rect 16696 -15652 16716 -15588
rect 16612 -15668 16716 -15652
rect 16612 -15732 16632 -15668
rect 16696 -15732 16716 -15668
rect 16612 -15748 16716 -15732
rect 11000 -16108 11104 -15812
rect 5388 -16188 5492 -16172
rect 5388 -16252 5408 -16188
rect 5472 -16252 5492 -16188
rect 5388 -16268 5492 -16252
rect 5388 -16332 5408 -16268
rect 5472 -16332 5492 -16268
rect 5388 -16348 5492 -16332
rect 5388 -16412 5408 -16348
rect 5472 -16412 5492 -16348
rect 5388 -16428 5492 -16412
rect 5388 -16492 5408 -16428
rect 5472 -16492 5492 -16428
rect 5388 -16508 5492 -16492
rect 5388 -16572 5408 -16508
rect 5472 -16572 5492 -16508
rect 5388 -16588 5492 -16572
rect 5388 -16652 5408 -16588
rect 5472 -16652 5492 -16588
rect 5388 -16668 5492 -16652
rect 5388 -16732 5408 -16668
rect 5472 -16732 5492 -16668
rect 5388 -16748 5492 -16732
rect 5388 -16812 5408 -16748
rect 5472 -16812 5492 -16748
rect 5388 -16828 5492 -16812
rect 5388 -16892 5408 -16828
rect 5472 -16892 5492 -16828
rect 5388 -16908 5492 -16892
rect 5388 -16972 5408 -16908
rect 5472 -16972 5492 -16908
rect 5388 -16988 5492 -16972
rect 5388 -17052 5408 -16988
rect 5472 -17052 5492 -16988
rect 5388 -17068 5492 -17052
rect 5388 -17132 5408 -17068
rect 5472 -17132 5492 -17068
rect 5388 -17148 5492 -17132
rect 5388 -17212 5408 -17148
rect 5472 -17212 5492 -17148
rect 5388 -17228 5492 -17212
rect 5388 -17292 5408 -17228
rect 5472 -17292 5492 -17228
rect 5388 -17308 5492 -17292
rect 5388 -17372 5408 -17308
rect 5472 -17372 5492 -17308
rect 5388 -17388 5492 -17372
rect 5388 -17452 5408 -17388
rect 5472 -17452 5492 -17388
rect 5388 -17468 5492 -17452
rect 5388 -17532 5408 -17468
rect 5472 -17532 5492 -17468
rect 5388 -17548 5492 -17532
rect 5388 -17612 5408 -17548
rect 5472 -17612 5492 -17548
rect 5388 -17628 5492 -17612
rect 5388 -17692 5408 -17628
rect 5472 -17692 5492 -17628
rect 5388 -17708 5492 -17692
rect 5388 -17772 5408 -17708
rect 5472 -17772 5492 -17708
rect 5388 -17788 5492 -17772
rect 5388 -17852 5408 -17788
rect 5472 -17852 5492 -17788
rect 5388 -17868 5492 -17852
rect 5388 -17932 5408 -17868
rect 5472 -17932 5492 -17868
rect 5388 -17948 5492 -17932
rect 5388 -18012 5408 -17948
rect 5472 -18012 5492 -17948
rect 5388 -18028 5492 -18012
rect 5388 -18092 5408 -18028
rect 5472 -18092 5492 -18028
rect 5388 -18108 5492 -18092
rect 5388 -18172 5408 -18108
rect 5472 -18172 5492 -18108
rect 5388 -18188 5492 -18172
rect 5388 -18252 5408 -18188
rect 5472 -18252 5492 -18188
rect 5388 -18268 5492 -18252
rect 5388 -18332 5408 -18268
rect 5472 -18332 5492 -18268
rect 5388 -18348 5492 -18332
rect 5388 -18412 5408 -18348
rect 5472 -18412 5492 -18348
rect 5388 -18428 5492 -18412
rect 5388 -18492 5408 -18428
rect 5472 -18492 5492 -18428
rect 5388 -18508 5492 -18492
rect 5388 -18572 5408 -18508
rect 5472 -18572 5492 -18508
rect 5388 -18588 5492 -18572
rect 5388 -18652 5408 -18588
rect 5472 -18652 5492 -18588
rect 5388 -18668 5492 -18652
rect 5388 -18732 5408 -18668
rect 5472 -18732 5492 -18668
rect 5388 -18748 5492 -18732
rect 5388 -18812 5408 -18748
rect 5472 -18812 5492 -18748
rect 5388 -18828 5492 -18812
rect 5388 -18892 5408 -18828
rect 5472 -18892 5492 -18828
rect 5388 -18908 5492 -18892
rect 5388 -18972 5408 -18908
rect 5472 -18972 5492 -18908
rect 5388 -18988 5492 -18972
rect 5388 -19052 5408 -18988
rect 5472 -19052 5492 -18988
rect 5388 -19068 5492 -19052
rect 5388 -19132 5408 -19068
rect 5472 -19132 5492 -19068
rect 5388 -19148 5492 -19132
rect 5388 -19212 5408 -19148
rect 5472 -19212 5492 -19148
rect 5388 -19228 5492 -19212
rect 5388 -19292 5408 -19228
rect 5472 -19292 5492 -19228
rect 5388 -19308 5492 -19292
rect 5388 -19372 5408 -19308
rect 5472 -19372 5492 -19308
rect 5388 -19388 5492 -19372
rect 5388 -19452 5408 -19388
rect 5472 -19452 5492 -19388
rect 5388 -19468 5492 -19452
rect 5388 -19532 5408 -19468
rect 5472 -19532 5492 -19468
rect 5388 -19548 5492 -19532
rect 5388 -19612 5408 -19548
rect 5472 -19612 5492 -19548
rect 5388 -19628 5492 -19612
rect 5388 -19692 5408 -19628
rect 5472 -19692 5492 -19628
rect 5388 -19708 5492 -19692
rect 5388 -19772 5408 -19708
rect 5472 -19772 5492 -19708
rect 5388 -19788 5492 -19772
rect 5388 -19852 5408 -19788
rect 5472 -19852 5492 -19788
rect 5388 -19868 5492 -19852
rect 5388 -19932 5408 -19868
rect 5472 -19932 5492 -19868
rect 5388 -19948 5492 -19932
rect 5388 -20012 5408 -19948
rect 5472 -20012 5492 -19948
rect 5388 -20028 5492 -20012
rect 5388 -20092 5408 -20028
rect 5472 -20092 5492 -20028
rect 5388 -20108 5492 -20092
rect 5388 -20172 5408 -20108
rect 5472 -20172 5492 -20108
rect 5388 -20188 5492 -20172
rect 5388 -20252 5408 -20188
rect 5472 -20252 5492 -20188
rect 5388 -20268 5492 -20252
rect 5388 -20332 5408 -20268
rect 5472 -20332 5492 -20268
rect 5388 -20348 5492 -20332
rect 5388 -20412 5408 -20348
rect 5472 -20412 5492 -20348
rect 5388 -20428 5492 -20412
rect 5388 -20492 5408 -20428
rect 5472 -20492 5492 -20428
rect 5388 -20508 5492 -20492
rect 5388 -20572 5408 -20508
rect 5472 -20572 5492 -20508
rect 5388 -20588 5492 -20572
rect 5388 -20652 5408 -20588
rect 5472 -20652 5492 -20588
rect 5388 -20668 5492 -20652
rect 5388 -20732 5408 -20668
rect 5472 -20732 5492 -20668
rect 5388 -20748 5492 -20732
rect 5388 -20812 5408 -20748
rect 5472 -20812 5492 -20748
rect 5388 -20828 5492 -20812
rect 5388 -20892 5408 -20828
rect 5472 -20892 5492 -20828
rect 5388 -20908 5492 -20892
rect 5388 -20972 5408 -20908
rect 5472 -20972 5492 -20908
rect 5388 -20988 5492 -20972
rect 5388 -21052 5408 -20988
rect 5472 -21052 5492 -20988
rect 5388 -21068 5492 -21052
rect -224 -21428 -120 -21132
rect -5836 -21508 -5732 -21492
rect -5836 -21572 -5816 -21508
rect -5752 -21572 -5732 -21508
rect -5836 -21588 -5732 -21572
rect -5836 -21652 -5816 -21588
rect -5752 -21652 -5732 -21588
rect -5836 -21668 -5732 -21652
rect -5836 -21732 -5816 -21668
rect -5752 -21732 -5732 -21668
rect -5836 -21748 -5732 -21732
rect -5836 -21812 -5816 -21748
rect -5752 -21812 -5732 -21748
rect -5836 -21828 -5732 -21812
rect -5836 -21892 -5816 -21828
rect -5752 -21892 -5732 -21828
rect -5836 -21908 -5732 -21892
rect -5836 -21972 -5816 -21908
rect -5752 -21972 -5732 -21908
rect -5836 -21988 -5732 -21972
rect -5836 -22052 -5816 -21988
rect -5752 -22052 -5732 -21988
rect -5836 -22068 -5732 -22052
rect -5836 -22132 -5816 -22068
rect -5752 -22132 -5732 -22068
rect -5836 -22148 -5732 -22132
rect -5836 -22212 -5816 -22148
rect -5752 -22212 -5732 -22148
rect -5836 -22228 -5732 -22212
rect -5836 -22292 -5816 -22228
rect -5752 -22292 -5732 -22228
rect -5836 -22308 -5732 -22292
rect -5836 -22372 -5816 -22308
rect -5752 -22372 -5732 -22308
rect -5836 -22388 -5732 -22372
rect -5836 -22452 -5816 -22388
rect -5752 -22452 -5732 -22388
rect -5836 -22468 -5732 -22452
rect -5836 -22532 -5816 -22468
rect -5752 -22532 -5732 -22468
rect -5836 -22548 -5732 -22532
rect -5836 -22612 -5816 -22548
rect -5752 -22612 -5732 -22548
rect -5836 -22628 -5732 -22612
rect -5836 -22692 -5816 -22628
rect -5752 -22692 -5732 -22628
rect -5836 -22708 -5732 -22692
rect -5836 -22772 -5816 -22708
rect -5752 -22772 -5732 -22708
rect -5836 -22788 -5732 -22772
rect -5836 -22852 -5816 -22788
rect -5752 -22852 -5732 -22788
rect -5836 -22868 -5732 -22852
rect -5836 -22932 -5816 -22868
rect -5752 -22932 -5732 -22868
rect -5836 -22948 -5732 -22932
rect -5836 -23012 -5816 -22948
rect -5752 -23012 -5732 -22948
rect -5836 -23028 -5732 -23012
rect -5836 -23092 -5816 -23028
rect -5752 -23092 -5732 -23028
rect -5836 -23108 -5732 -23092
rect -5836 -23172 -5816 -23108
rect -5752 -23172 -5732 -23108
rect -5836 -23188 -5732 -23172
rect -5836 -23252 -5816 -23188
rect -5752 -23252 -5732 -23188
rect -5836 -23268 -5732 -23252
rect -5836 -23332 -5816 -23268
rect -5752 -23332 -5732 -23268
rect -5836 -23348 -5732 -23332
rect -5836 -23412 -5816 -23348
rect -5752 -23412 -5732 -23348
rect -5836 -23428 -5732 -23412
rect -5836 -23492 -5816 -23428
rect -5752 -23492 -5732 -23428
rect -5836 -23508 -5732 -23492
rect -5836 -23572 -5816 -23508
rect -5752 -23572 -5732 -23508
rect -5836 -23588 -5732 -23572
rect -5836 -23652 -5816 -23588
rect -5752 -23652 -5732 -23588
rect -5836 -23668 -5732 -23652
rect -5836 -23732 -5816 -23668
rect -5752 -23732 -5732 -23668
rect -5836 -23748 -5732 -23732
rect -5836 -23812 -5816 -23748
rect -5752 -23812 -5732 -23748
rect -5836 -23828 -5732 -23812
rect -5836 -23892 -5816 -23828
rect -5752 -23892 -5732 -23828
rect -5836 -23908 -5732 -23892
rect -5836 -23972 -5816 -23908
rect -5752 -23972 -5732 -23908
rect -5836 -23988 -5732 -23972
rect -5836 -24052 -5816 -23988
rect -5752 -24052 -5732 -23988
rect -5836 -24068 -5732 -24052
rect -5836 -24132 -5816 -24068
rect -5752 -24132 -5732 -24068
rect -5836 -24148 -5732 -24132
rect -5836 -24212 -5816 -24148
rect -5752 -24212 -5732 -24148
rect -5836 -24228 -5732 -24212
rect -5836 -24292 -5816 -24228
rect -5752 -24292 -5732 -24228
rect -5836 -24308 -5732 -24292
rect -5836 -24372 -5816 -24308
rect -5752 -24372 -5732 -24308
rect -5836 -24388 -5732 -24372
rect -5836 -24452 -5816 -24388
rect -5752 -24452 -5732 -24388
rect -5836 -24468 -5732 -24452
rect -5836 -24532 -5816 -24468
rect -5752 -24532 -5732 -24468
rect -5836 -24548 -5732 -24532
rect -5836 -24612 -5816 -24548
rect -5752 -24612 -5732 -24548
rect -5836 -24628 -5732 -24612
rect -5836 -24692 -5816 -24628
rect -5752 -24692 -5732 -24628
rect -5836 -24708 -5732 -24692
rect -5836 -24772 -5816 -24708
rect -5752 -24772 -5732 -24708
rect -5836 -24788 -5732 -24772
rect -5836 -24852 -5816 -24788
rect -5752 -24852 -5732 -24788
rect -5836 -24868 -5732 -24852
rect -5836 -24932 -5816 -24868
rect -5752 -24932 -5732 -24868
rect -5836 -24948 -5732 -24932
rect -5836 -25012 -5816 -24948
rect -5752 -25012 -5732 -24948
rect -5836 -25028 -5732 -25012
rect -5836 -25092 -5816 -25028
rect -5752 -25092 -5732 -25028
rect -5836 -25108 -5732 -25092
rect -5836 -25172 -5816 -25108
rect -5752 -25172 -5732 -25108
rect -5836 -25188 -5732 -25172
rect -5836 -25252 -5816 -25188
rect -5752 -25252 -5732 -25188
rect -5836 -25268 -5732 -25252
rect -5836 -25332 -5816 -25268
rect -5752 -25332 -5732 -25268
rect -5836 -25348 -5732 -25332
rect -5836 -25412 -5816 -25348
rect -5752 -25412 -5732 -25348
rect -5836 -25428 -5732 -25412
rect -5836 -25492 -5816 -25428
rect -5752 -25492 -5732 -25428
rect -5836 -25508 -5732 -25492
rect -5836 -25572 -5816 -25508
rect -5752 -25572 -5732 -25508
rect -5836 -25588 -5732 -25572
rect -5836 -25652 -5816 -25588
rect -5752 -25652 -5732 -25588
rect -5836 -25668 -5732 -25652
rect -5836 -25732 -5816 -25668
rect -5752 -25732 -5732 -25668
rect -5836 -25748 -5732 -25732
rect -5836 -25812 -5816 -25748
rect -5752 -25812 -5732 -25748
rect -5836 -25828 -5732 -25812
rect -5836 -25892 -5816 -25828
rect -5752 -25892 -5732 -25828
rect -5836 -25908 -5732 -25892
rect -5836 -25972 -5816 -25908
rect -5752 -25972 -5732 -25908
rect -5836 -25988 -5732 -25972
rect -5836 -26052 -5816 -25988
rect -5752 -26052 -5732 -25988
rect -5836 -26068 -5732 -26052
rect -5836 -26132 -5816 -26068
rect -5752 -26132 -5732 -26068
rect -5836 -26148 -5732 -26132
rect -5836 -26212 -5816 -26148
rect -5752 -26212 -5732 -26148
rect -5836 -26228 -5732 -26212
rect -5836 -26292 -5816 -26228
rect -5752 -26292 -5732 -26228
rect -5836 -26308 -5732 -26292
rect -5836 -26372 -5816 -26308
rect -5752 -26372 -5732 -26308
rect -5836 -26388 -5732 -26372
rect -11448 -26748 -11344 -26452
rect -17060 -26828 -16956 -26812
rect -17060 -26892 -17040 -26828
rect -16976 -26892 -16956 -26828
rect -17060 -26908 -16956 -26892
rect -17060 -26972 -17040 -26908
rect -16976 -26972 -16956 -26908
rect -17060 -26988 -16956 -26972
rect -17060 -27052 -17040 -26988
rect -16976 -27052 -16956 -26988
rect -17060 -27068 -16956 -27052
rect -17060 -27132 -17040 -27068
rect -16976 -27132 -16956 -27068
rect -17060 -27148 -16956 -27132
rect -17060 -27212 -17040 -27148
rect -16976 -27212 -16956 -27148
rect -17060 -27228 -16956 -27212
rect -17060 -27292 -17040 -27228
rect -16976 -27292 -16956 -27228
rect -17060 -27308 -16956 -27292
rect -17060 -27372 -17040 -27308
rect -16976 -27372 -16956 -27308
rect -17060 -27388 -16956 -27372
rect -17060 -27452 -17040 -27388
rect -16976 -27452 -16956 -27388
rect -17060 -27468 -16956 -27452
rect -17060 -27532 -17040 -27468
rect -16976 -27532 -16956 -27468
rect -17060 -27548 -16956 -27532
rect -17060 -27612 -17040 -27548
rect -16976 -27612 -16956 -27548
rect -17060 -27628 -16956 -27612
rect -17060 -27692 -17040 -27628
rect -16976 -27692 -16956 -27628
rect -17060 -27708 -16956 -27692
rect -17060 -27772 -17040 -27708
rect -16976 -27772 -16956 -27708
rect -17060 -27788 -16956 -27772
rect -17060 -27852 -17040 -27788
rect -16976 -27852 -16956 -27788
rect -17060 -27868 -16956 -27852
rect -17060 -27932 -17040 -27868
rect -16976 -27932 -16956 -27868
rect -17060 -27948 -16956 -27932
rect -17060 -28012 -17040 -27948
rect -16976 -28012 -16956 -27948
rect -17060 -28028 -16956 -28012
rect -17060 -28092 -17040 -28028
rect -16976 -28092 -16956 -28028
rect -17060 -28108 -16956 -28092
rect -17060 -28172 -17040 -28108
rect -16976 -28172 -16956 -28108
rect -17060 -28188 -16956 -28172
rect -17060 -28252 -17040 -28188
rect -16976 -28252 -16956 -28188
rect -17060 -28268 -16956 -28252
rect -17060 -28332 -17040 -28268
rect -16976 -28332 -16956 -28268
rect -17060 -28348 -16956 -28332
rect -17060 -28412 -17040 -28348
rect -16976 -28412 -16956 -28348
rect -17060 -28428 -16956 -28412
rect -17060 -28492 -17040 -28428
rect -16976 -28492 -16956 -28428
rect -17060 -28508 -16956 -28492
rect -17060 -28572 -17040 -28508
rect -16976 -28572 -16956 -28508
rect -17060 -28588 -16956 -28572
rect -17060 -28652 -17040 -28588
rect -16976 -28652 -16956 -28588
rect -17060 -28668 -16956 -28652
rect -17060 -28732 -17040 -28668
rect -16976 -28732 -16956 -28668
rect -17060 -28748 -16956 -28732
rect -17060 -28812 -17040 -28748
rect -16976 -28812 -16956 -28748
rect -17060 -28828 -16956 -28812
rect -17060 -28892 -17040 -28828
rect -16976 -28892 -16956 -28828
rect -17060 -28908 -16956 -28892
rect -17060 -28972 -17040 -28908
rect -16976 -28972 -16956 -28908
rect -17060 -28988 -16956 -28972
rect -17060 -29052 -17040 -28988
rect -16976 -29052 -16956 -28988
rect -17060 -29068 -16956 -29052
rect -17060 -29132 -17040 -29068
rect -16976 -29132 -16956 -29068
rect -17060 -29148 -16956 -29132
rect -17060 -29212 -17040 -29148
rect -16976 -29212 -16956 -29148
rect -17060 -29228 -16956 -29212
rect -17060 -29292 -17040 -29228
rect -16976 -29292 -16956 -29228
rect -17060 -29308 -16956 -29292
rect -17060 -29372 -17040 -29308
rect -16976 -29372 -16956 -29308
rect -17060 -29388 -16956 -29372
rect -17060 -29452 -17040 -29388
rect -16976 -29452 -16956 -29388
rect -17060 -29468 -16956 -29452
rect -17060 -29532 -17040 -29468
rect -16976 -29532 -16956 -29468
rect -17060 -29548 -16956 -29532
rect -17060 -29612 -17040 -29548
rect -16976 -29612 -16956 -29548
rect -17060 -29628 -16956 -29612
rect -17060 -29692 -17040 -29628
rect -16976 -29692 -16956 -29628
rect -17060 -29708 -16956 -29692
rect -17060 -29772 -17040 -29708
rect -16976 -29772 -16956 -29708
rect -17060 -29788 -16956 -29772
rect -17060 -29852 -17040 -29788
rect -16976 -29852 -16956 -29788
rect -17060 -29868 -16956 -29852
rect -17060 -29932 -17040 -29868
rect -16976 -29932 -16956 -29868
rect -17060 -29948 -16956 -29932
rect -17060 -30012 -17040 -29948
rect -16976 -30012 -16956 -29948
rect -17060 -30028 -16956 -30012
rect -17060 -30092 -17040 -30028
rect -16976 -30092 -16956 -30028
rect -17060 -30108 -16956 -30092
rect -17060 -30172 -17040 -30108
rect -16976 -30172 -16956 -30108
rect -17060 -30188 -16956 -30172
rect -17060 -30252 -17040 -30188
rect -16976 -30252 -16956 -30188
rect -17060 -30268 -16956 -30252
rect -17060 -30332 -17040 -30268
rect -16976 -30332 -16956 -30268
rect -17060 -30348 -16956 -30332
rect -17060 -30412 -17040 -30348
rect -16976 -30412 -16956 -30348
rect -17060 -30428 -16956 -30412
rect -17060 -30492 -17040 -30428
rect -16976 -30492 -16956 -30428
rect -17060 -30508 -16956 -30492
rect -17060 -30572 -17040 -30508
rect -16976 -30572 -16956 -30508
rect -17060 -30588 -16956 -30572
rect -17060 -30652 -17040 -30588
rect -16976 -30652 -16956 -30588
rect -17060 -30668 -16956 -30652
rect -17060 -30732 -17040 -30668
rect -16976 -30732 -16956 -30668
rect -17060 -30748 -16956 -30732
rect -17060 -30812 -17040 -30748
rect -16976 -30812 -16956 -30748
rect -17060 -30828 -16956 -30812
rect -17060 -30892 -17040 -30828
rect -16976 -30892 -16956 -30828
rect -17060 -30908 -16956 -30892
rect -17060 -30972 -17040 -30908
rect -16976 -30972 -16956 -30908
rect -17060 -30988 -16956 -30972
rect -17060 -31052 -17040 -30988
rect -16976 -31052 -16956 -30988
rect -17060 -31068 -16956 -31052
rect -17060 -31132 -17040 -31068
rect -16976 -31132 -16956 -31068
rect -17060 -31148 -16956 -31132
rect -17060 -31212 -17040 -31148
rect -16976 -31212 -16956 -31148
rect -17060 -31228 -16956 -31212
rect -17060 -31292 -17040 -31228
rect -16976 -31292 -16956 -31228
rect -17060 -31308 -16956 -31292
rect -17060 -31372 -17040 -31308
rect -16976 -31372 -16956 -31308
rect -17060 -31388 -16956 -31372
rect -17060 -31452 -17040 -31388
rect -16976 -31452 -16956 -31388
rect -17060 -31468 -16956 -31452
rect -17060 -31532 -17040 -31468
rect -16976 -31532 -16956 -31468
rect -17060 -31548 -16956 -31532
rect -17060 -31612 -17040 -31548
rect -16976 -31612 -16956 -31548
rect -17060 -31628 -16956 -31612
rect -17060 -31692 -17040 -31628
rect -16976 -31692 -16956 -31628
rect -17060 -31708 -16956 -31692
rect -22672 -32068 -22568 -31772
rect -28284 -32148 -28180 -32132
rect -28284 -32212 -28264 -32148
rect -28200 -32212 -28180 -32148
rect -28284 -32228 -28180 -32212
rect -28284 -32292 -28264 -32228
rect -28200 -32292 -28180 -32228
rect -28284 -32308 -28180 -32292
rect -28284 -32372 -28264 -32308
rect -28200 -32372 -28180 -32308
rect -28284 -32388 -28180 -32372
rect -28284 -32452 -28264 -32388
rect -28200 -32452 -28180 -32388
rect -28284 -32468 -28180 -32452
rect -28284 -32532 -28264 -32468
rect -28200 -32532 -28180 -32468
rect -28284 -32548 -28180 -32532
rect -28284 -32612 -28264 -32548
rect -28200 -32612 -28180 -32548
rect -28284 -32628 -28180 -32612
rect -28284 -32692 -28264 -32628
rect -28200 -32692 -28180 -32628
rect -28284 -32708 -28180 -32692
rect -28284 -32772 -28264 -32708
rect -28200 -32772 -28180 -32708
rect -28284 -32788 -28180 -32772
rect -28284 -32852 -28264 -32788
rect -28200 -32852 -28180 -32788
rect -28284 -32868 -28180 -32852
rect -28284 -32932 -28264 -32868
rect -28200 -32932 -28180 -32868
rect -28284 -32948 -28180 -32932
rect -28284 -33012 -28264 -32948
rect -28200 -33012 -28180 -32948
rect -28284 -33028 -28180 -33012
rect -28284 -33092 -28264 -33028
rect -28200 -33092 -28180 -33028
rect -28284 -33108 -28180 -33092
rect -28284 -33172 -28264 -33108
rect -28200 -33172 -28180 -33108
rect -28284 -33188 -28180 -33172
rect -28284 -33252 -28264 -33188
rect -28200 -33252 -28180 -33188
rect -28284 -33268 -28180 -33252
rect -28284 -33332 -28264 -33268
rect -28200 -33332 -28180 -33268
rect -28284 -33348 -28180 -33332
rect -28284 -33412 -28264 -33348
rect -28200 -33412 -28180 -33348
rect -28284 -33428 -28180 -33412
rect -28284 -33492 -28264 -33428
rect -28200 -33492 -28180 -33428
rect -28284 -33508 -28180 -33492
rect -28284 -33572 -28264 -33508
rect -28200 -33572 -28180 -33508
rect -28284 -33588 -28180 -33572
rect -28284 -33652 -28264 -33588
rect -28200 -33652 -28180 -33588
rect -28284 -33668 -28180 -33652
rect -28284 -33732 -28264 -33668
rect -28200 -33732 -28180 -33668
rect -28284 -33748 -28180 -33732
rect -28284 -33812 -28264 -33748
rect -28200 -33812 -28180 -33748
rect -28284 -33828 -28180 -33812
rect -28284 -33892 -28264 -33828
rect -28200 -33892 -28180 -33828
rect -28284 -33908 -28180 -33892
rect -28284 -33972 -28264 -33908
rect -28200 -33972 -28180 -33908
rect -28284 -33988 -28180 -33972
rect -28284 -34052 -28264 -33988
rect -28200 -34052 -28180 -33988
rect -28284 -34068 -28180 -34052
rect -28284 -34132 -28264 -34068
rect -28200 -34132 -28180 -34068
rect -28284 -34148 -28180 -34132
rect -28284 -34212 -28264 -34148
rect -28200 -34212 -28180 -34148
rect -28284 -34228 -28180 -34212
rect -28284 -34292 -28264 -34228
rect -28200 -34292 -28180 -34228
rect -28284 -34308 -28180 -34292
rect -28284 -34372 -28264 -34308
rect -28200 -34372 -28180 -34308
rect -28284 -34388 -28180 -34372
rect -28284 -34452 -28264 -34388
rect -28200 -34452 -28180 -34388
rect -28284 -34468 -28180 -34452
rect -28284 -34532 -28264 -34468
rect -28200 -34532 -28180 -34468
rect -28284 -34548 -28180 -34532
rect -28284 -34612 -28264 -34548
rect -28200 -34612 -28180 -34548
rect -28284 -34628 -28180 -34612
rect -28284 -34692 -28264 -34628
rect -28200 -34692 -28180 -34628
rect -28284 -34708 -28180 -34692
rect -28284 -34772 -28264 -34708
rect -28200 -34772 -28180 -34708
rect -28284 -34788 -28180 -34772
rect -28284 -34852 -28264 -34788
rect -28200 -34852 -28180 -34788
rect -28284 -34868 -28180 -34852
rect -28284 -34932 -28264 -34868
rect -28200 -34932 -28180 -34868
rect -28284 -34948 -28180 -34932
rect -28284 -35012 -28264 -34948
rect -28200 -35012 -28180 -34948
rect -28284 -35028 -28180 -35012
rect -28284 -35092 -28264 -35028
rect -28200 -35092 -28180 -35028
rect -28284 -35108 -28180 -35092
rect -28284 -35172 -28264 -35108
rect -28200 -35172 -28180 -35108
rect -28284 -35188 -28180 -35172
rect -28284 -35252 -28264 -35188
rect -28200 -35252 -28180 -35188
rect -28284 -35268 -28180 -35252
rect -28284 -35332 -28264 -35268
rect -28200 -35332 -28180 -35268
rect -28284 -35348 -28180 -35332
rect -28284 -35412 -28264 -35348
rect -28200 -35412 -28180 -35348
rect -28284 -35428 -28180 -35412
rect -28284 -35492 -28264 -35428
rect -28200 -35492 -28180 -35428
rect -28284 -35508 -28180 -35492
rect -28284 -35572 -28264 -35508
rect -28200 -35572 -28180 -35508
rect -28284 -35588 -28180 -35572
rect -28284 -35652 -28264 -35588
rect -28200 -35652 -28180 -35588
rect -28284 -35668 -28180 -35652
rect -28284 -35732 -28264 -35668
rect -28200 -35732 -28180 -35668
rect -28284 -35748 -28180 -35732
rect -28284 -35812 -28264 -35748
rect -28200 -35812 -28180 -35748
rect -28284 -35828 -28180 -35812
rect -28284 -35892 -28264 -35828
rect -28200 -35892 -28180 -35828
rect -28284 -35908 -28180 -35892
rect -28284 -35972 -28264 -35908
rect -28200 -35972 -28180 -35908
rect -28284 -35988 -28180 -35972
rect -28284 -36052 -28264 -35988
rect -28200 -36052 -28180 -35988
rect -28284 -36068 -28180 -36052
rect -28284 -36132 -28264 -36068
rect -28200 -36132 -28180 -36068
rect -28284 -36148 -28180 -36132
rect -28284 -36212 -28264 -36148
rect -28200 -36212 -28180 -36148
rect -28284 -36228 -28180 -36212
rect -28284 -36292 -28264 -36228
rect -28200 -36292 -28180 -36228
rect -28284 -36308 -28180 -36292
rect -28284 -36372 -28264 -36308
rect -28200 -36372 -28180 -36308
rect -28284 -36388 -28180 -36372
rect -28284 -36452 -28264 -36388
rect -28200 -36452 -28180 -36388
rect -28284 -36468 -28180 -36452
rect -28284 -36532 -28264 -36468
rect -28200 -36532 -28180 -36468
rect -28284 -36548 -28180 -36532
rect -28284 -36612 -28264 -36548
rect -28200 -36612 -28180 -36548
rect -28284 -36628 -28180 -36612
rect -28284 -36692 -28264 -36628
rect -28200 -36692 -28180 -36628
rect -28284 -36708 -28180 -36692
rect -28284 -36772 -28264 -36708
rect -28200 -36772 -28180 -36708
rect -28284 -36788 -28180 -36772
rect -28284 -36852 -28264 -36788
rect -28200 -36852 -28180 -36788
rect -28284 -36868 -28180 -36852
rect -28284 -36932 -28264 -36868
rect -28200 -36932 -28180 -36868
rect -28284 -36948 -28180 -36932
rect -28284 -37012 -28264 -36948
rect -28200 -37012 -28180 -36948
rect -28284 -37028 -28180 -37012
rect -33896 -37240 -33792 -37092
rect -31064 -37240 -30960 -37041
rect -28284 -37092 -28264 -37028
rect -28200 -37092 -28180 -37028
rect -27861 -32148 -22939 -32119
rect -27861 -37012 -27832 -32148
rect -22968 -37012 -22939 -32148
rect -27861 -37041 -22939 -37012
rect -22672 -32132 -22652 -32068
rect -22588 -32132 -22568 -32068
rect -19840 -32119 -19736 -31721
rect -17060 -31772 -17040 -31708
rect -16976 -31772 -16956 -31708
rect -16637 -26828 -11715 -26799
rect -16637 -31692 -16608 -26828
rect -11744 -31692 -11715 -26828
rect -16637 -31721 -11715 -31692
rect -11448 -26812 -11428 -26748
rect -11364 -26812 -11344 -26748
rect -8616 -26799 -8512 -26401
rect -5836 -26452 -5816 -26388
rect -5752 -26452 -5732 -26388
rect -5413 -21508 -491 -21479
rect -5413 -26372 -5384 -21508
rect -520 -26372 -491 -21508
rect -5413 -26401 -491 -26372
rect -224 -21492 -204 -21428
rect -140 -21492 -120 -21428
rect 2608 -21479 2712 -21081
rect 5388 -21132 5408 -21068
rect 5472 -21132 5492 -21068
rect 5811 -16188 10733 -16159
rect 5811 -21052 5840 -16188
rect 10704 -21052 10733 -16188
rect 5811 -21081 10733 -21052
rect 11000 -16172 11020 -16108
rect 11084 -16172 11104 -16108
rect 13832 -16159 13936 -15761
rect 16612 -15812 16632 -15748
rect 16696 -15812 16716 -15748
rect 17035 -10868 21957 -10839
rect 17035 -15732 17064 -10868
rect 21928 -15732 21957 -10868
rect 17035 -15761 21957 -15732
rect 22224 -10852 22244 -10788
rect 22308 -10852 22328 -10788
rect 25056 -10839 25160 -10441
rect 27836 -10492 27856 -10428
rect 27920 -10492 27940 -10428
rect 28259 -5548 33181 -5519
rect 28259 -10412 28288 -5548
rect 33152 -10412 33181 -5548
rect 28259 -10441 33181 -10412
rect 33448 -5532 33468 -5468
rect 33532 -5532 33552 -5468
rect 36280 -5519 36384 -5121
rect 39060 -5172 39080 -5108
rect 39144 -5172 39164 -5108
rect 39060 -5468 39164 -5172
rect 33448 -5548 33552 -5532
rect 33448 -5612 33468 -5548
rect 33532 -5612 33552 -5548
rect 33448 -5628 33552 -5612
rect 33448 -5692 33468 -5628
rect 33532 -5692 33552 -5628
rect 33448 -5708 33552 -5692
rect 33448 -5772 33468 -5708
rect 33532 -5772 33552 -5708
rect 33448 -5788 33552 -5772
rect 33448 -5852 33468 -5788
rect 33532 -5852 33552 -5788
rect 33448 -5868 33552 -5852
rect 33448 -5932 33468 -5868
rect 33532 -5932 33552 -5868
rect 33448 -5948 33552 -5932
rect 33448 -6012 33468 -5948
rect 33532 -6012 33552 -5948
rect 33448 -6028 33552 -6012
rect 33448 -6092 33468 -6028
rect 33532 -6092 33552 -6028
rect 33448 -6108 33552 -6092
rect 33448 -6172 33468 -6108
rect 33532 -6172 33552 -6108
rect 33448 -6188 33552 -6172
rect 33448 -6252 33468 -6188
rect 33532 -6252 33552 -6188
rect 33448 -6268 33552 -6252
rect 33448 -6332 33468 -6268
rect 33532 -6332 33552 -6268
rect 33448 -6348 33552 -6332
rect 33448 -6412 33468 -6348
rect 33532 -6412 33552 -6348
rect 33448 -6428 33552 -6412
rect 33448 -6492 33468 -6428
rect 33532 -6492 33552 -6428
rect 33448 -6508 33552 -6492
rect 33448 -6572 33468 -6508
rect 33532 -6572 33552 -6508
rect 33448 -6588 33552 -6572
rect 33448 -6652 33468 -6588
rect 33532 -6652 33552 -6588
rect 33448 -6668 33552 -6652
rect 33448 -6732 33468 -6668
rect 33532 -6732 33552 -6668
rect 33448 -6748 33552 -6732
rect 33448 -6812 33468 -6748
rect 33532 -6812 33552 -6748
rect 33448 -6828 33552 -6812
rect 33448 -6892 33468 -6828
rect 33532 -6892 33552 -6828
rect 33448 -6908 33552 -6892
rect 33448 -6972 33468 -6908
rect 33532 -6972 33552 -6908
rect 33448 -6988 33552 -6972
rect 33448 -7052 33468 -6988
rect 33532 -7052 33552 -6988
rect 33448 -7068 33552 -7052
rect 33448 -7132 33468 -7068
rect 33532 -7132 33552 -7068
rect 33448 -7148 33552 -7132
rect 33448 -7212 33468 -7148
rect 33532 -7212 33552 -7148
rect 33448 -7228 33552 -7212
rect 33448 -7292 33468 -7228
rect 33532 -7292 33552 -7228
rect 33448 -7308 33552 -7292
rect 33448 -7372 33468 -7308
rect 33532 -7372 33552 -7308
rect 33448 -7388 33552 -7372
rect 33448 -7452 33468 -7388
rect 33532 -7452 33552 -7388
rect 33448 -7468 33552 -7452
rect 33448 -7532 33468 -7468
rect 33532 -7532 33552 -7468
rect 33448 -7548 33552 -7532
rect 33448 -7612 33468 -7548
rect 33532 -7612 33552 -7548
rect 33448 -7628 33552 -7612
rect 33448 -7692 33468 -7628
rect 33532 -7692 33552 -7628
rect 33448 -7708 33552 -7692
rect 33448 -7772 33468 -7708
rect 33532 -7772 33552 -7708
rect 33448 -7788 33552 -7772
rect 33448 -7852 33468 -7788
rect 33532 -7852 33552 -7788
rect 33448 -7868 33552 -7852
rect 33448 -7932 33468 -7868
rect 33532 -7932 33552 -7868
rect 33448 -7948 33552 -7932
rect 33448 -8012 33468 -7948
rect 33532 -8012 33552 -7948
rect 33448 -8028 33552 -8012
rect 33448 -8092 33468 -8028
rect 33532 -8092 33552 -8028
rect 33448 -8108 33552 -8092
rect 33448 -8172 33468 -8108
rect 33532 -8172 33552 -8108
rect 33448 -8188 33552 -8172
rect 33448 -8252 33468 -8188
rect 33532 -8252 33552 -8188
rect 33448 -8268 33552 -8252
rect 33448 -8332 33468 -8268
rect 33532 -8332 33552 -8268
rect 33448 -8348 33552 -8332
rect 33448 -8412 33468 -8348
rect 33532 -8412 33552 -8348
rect 33448 -8428 33552 -8412
rect 33448 -8492 33468 -8428
rect 33532 -8492 33552 -8428
rect 33448 -8508 33552 -8492
rect 33448 -8572 33468 -8508
rect 33532 -8572 33552 -8508
rect 33448 -8588 33552 -8572
rect 33448 -8652 33468 -8588
rect 33532 -8652 33552 -8588
rect 33448 -8668 33552 -8652
rect 33448 -8732 33468 -8668
rect 33532 -8732 33552 -8668
rect 33448 -8748 33552 -8732
rect 33448 -8812 33468 -8748
rect 33532 -8812 33552 -8748
rect 33448 -8828 33552 -8812
rect 33448 -8892 33468 -8828
rect 33532 -8892 33552 -8828
rect 33448 -8908 33552 -8892
rect 33448 -8972 33468 -8908
rect 33532 -8972 33552 -8908
rect 33448 -8988 33552 -8972
rect 33448 -9052 33468 -8988
rect 33532 -9052 33552 -8988
rect 33448 -9068 33552 -9052
rect 33448 -9132 33468 -9068
rect 33532 -9132 33552 -9068
rect 33448 -9148 33552 -9132
rect 33448 -9212 33468 -9148
rect 33532 -9212 33552 -9148
rect 33448 -9228 33552 -9212
rect 33448 -9292 33468 -9228
rect 33532 -9292 33552 -9228
rect 33448 -9308 33552 -9292
rect 33448 -9372 33468 -9308
rect 33532 -9372 33552 -9308
rect 33448 -9388 33552 -9372
rect 33448 -9452 33468 -9388
rect 33532 -9452 33552 -9388
rect 33448 -9468 33552 -9452
rect 33448 -9532 33468 -9468
rect 33532 -9532 33552 -9468
rect 33448 -9548 33552 -9532
rect 33448 -9612 33468 -9548
rect 33532 -9612 33552 -9548
rect 33448 -9628 33552 -9612
rect 33448 -9692 33468 -9628
rect 33532 -9692 33552 -9628
rect 33448 -9708 33552 -9692
rect 33448 -9772 33468 -9708
rect 33532 -9772 33552 -9708
rect 33448 -9788 33552 -9772
rect 33448 -9852 33468 -9788
rect 33532 -9852 33552 -9788
rect 33448 -9868 33552 -9852
rect 33448 -9932 33468 -9868
rect 33532 -9932 33552 -9868
rect 33448 -9948 33552 -9932
rect 33448 -10012 33468 -9948
rect 33532 -10012 33552 -9948
rect 33448 -10028 33552 -10012
rect 33448 -10092 33468 -10028
rect 33532 -10092 33552 -10028
rect 33448 -10108 33552 -10092
rect 33448 -10172 33468 -10108
rect 33532 -10172 33552 -10108
rect 33448 -10188 33552 -10172
rect 33448 -10252 33468 -10188
rect 33532 -10252 33552 -10188
rect 33448 -10268 33552 -10252
rect 33448 -10332 33468 -10268
rect 33532 -10332 33552 -10268
rect 33448 -10348 33552 -10332
rect 33448 -10412 33468 -10348
rect 33532 -10412 33552 -10348
rect 33448 -10428 33552 -10412
rect 27836 -10788 27940 -10492
rect 22224 -10868 22328 -10852
rect 22224 -10932 22244 -10868
rect 22308 -10932 22328 -10868
rect 22224 -10948 22328 -10932
rect 22224 -11012 22244 -10948
rect 22308 -11012 22328 -10948
rect 22224 -11028 22328 -11012
rect 22224 -11092 22244 -11028
rect 22308 -11092 22328 -11028
rect 22224 -11108 22328 -11092
rect 22224 -11172 22244 -11108
rect 22308 -11172 22328 -11108
rect 22224 -11188 22328 -11172
rect 22224 -11252 22244 -11188
rect 22308 -11252 22328 -11188
rect 22224 -11268 22328 -11252
rect 22224 -11332 22244 -11268
rect 22308 -11332 22328 -11268
rect 22224 -11348 22328 -11332
rect 22224 -11412 22244 -11348
rect 22308 -11412 22328 -11348
rect 22224 -11428 22328 -11412
rect 22224 -11492 22244 -11428
rect 22308 -11492 22328 -11428
rect 22224 -11508 22328 -11492
rect 22224 -11572 22244 -11508
rect 22308 -11572 22328 -11508
rect 22224 -11588 22328 -11572
rect 22224 -11652 22244 -11588
rect 22308 -11652 22328 -11588
rect 22224 -11668 22328 -11652
rect 22224 -11732 22244 -11668
rect 22308 -11732 22328 -11668
rect 22224 -11748 22328 -11732
rect 22224 -11812 22244 -11748
rect 22308 -11812 22328 -11748
rect 22224 -11828 22328 -11812
rect 22224 -11892 22244 -11828
rect 22308 -11892 22328 -11828
rect 22224 -11908 22328 -11892
rect 22224 -11972 22244 -11908
rect 22308 -11972 22328 -11908
rect 22224 -11988 22328 -11972
rect 22224 -12052 22244 -11988
rect 22308 -12052 22328 -11988
rect 22224 -12068 22328 -12052
rect 22224 -12132 22244 -12068
rect 22308 -12132 22328 -12068
rect 22224 -12148 22328 -12132
rect 22224 -12212 22244 -12148
rect 22308 -12212 22328 -12148
rect 22224 -12228 22328 -12212
rect 22224 -12292 22244 -12228
rect 22308 -12292 22328 -12228
rect 22224 -12308 22328 -12292
rect 22224 -12372 22244 -12308
rect 22308 -12372 22328 -12308
rect 22224 -12388 22328 -12372
rect 22224 -12452 22244 -12388
rect 22308 -12452 22328 -12388
rect 22224 -12468 22328 -12452
rect 22224 -12532 22244 -12468
rect 22308 -12532 22328 -12468
rect 22224 -12548 22328 -12532
rect 22224 -12612 22244 -12548
rect 22308 -12612 22328 -12548
rect 22224 -12628 22328 -12612
rect 22224 -12692 22244 -12628
rect 22308 -12692 22328 -12628
rect 22224 -12708 22328 -12692
rect 22224 -12772 22244 -12708
rect 22308 -12772 22328 -12708
rect 22224 -12788 22328 -12772
rect 22224 -12852 22244 -12788
rect 22308 -12852 22328 -12788
rect 22224 -12868 22328 -12852
rect 22224 -12932 22244 -12868
rect 22308 -12932 22328 -12868
rect 22224 -12948 22328 -12932
rect 22224 -13012 22244 -12948
rect 22308 -13012 22328 -12948
rect 22224 -13028 22328 -13012
rect 22224 -13092 22244 -13028
rect 22308 -13092 22328 -13028
rect 22224 -13108 22328 -13092
rect 22224 -13172 22244 -13108
rect 22308 -13172 22328 -13108
rect 22224 -13188 22328 -13172
rect 22224 -13252 22244 -13188
rect 22308 -13252 22328 -13188
rect 22224 -13268 22328 -13252
rect 22224 -13332 22244 -13268
rect 22308 -13332 22328 -13268
rect 22224 -13348 22328 -13332
rect 22224 -13412 22244 -13348
rect 22308 -13412 22328 -13348
rect 22224 -13428 22328 -13412
rect 22224 -13492 22244 -13428
rect 22308 -13492 22328 -13428
rect 22224 -13508 22328 -13492
rect 22224 -13572 22244 -13508
rect 22308 -13572 22328 -13508
rect 22224 -13588 22328 -13572
rect 22224 -13652 22244 -13588
rect 22308 -13652 22328 -13588
rect 22224 -13668 22328 -13652
rect 22224 -13732 22244 -13668
rect 22308 -13732 22328 -13668
rect 22224 -13748 22328 -13732
rect 22224 -13812 22244 -13748
rect 22308 -13812 22328 -13748
rect 22224 -13828 22328 -13812
rect 22224 -13892 22244 -13828
rect 22308 -13892 22328 -13828
rect 22224 -13908 22328 -13892
rect 22224 -13972 22244 -13908
rect 22308 -13972 22328 -13908
rect 22224 -13988 22328 -13972
rect 22224 -14052 22244 -13988
rect 22308 -14052 22328 -13988
rect 22224 -14068 22328 -14052
rect 22224 -14132 22244 -14068
rect 22308 -14132 22328 -14068
rect 22224 -14148 22328 -14132
rect 22224 -14212 22244 -14148
rect 22308 -14212 22328 -14148
rect 22224 -14228 22328 -14212
rect 22224 -14292 22244 -14228
rect 22308 -14292 22328 -14228
rect 22224 -14308 22328 -14292
rect 22224 -14372 22244 -14308
rect 22308 -14372 22328 -14308
rect 22224 -14388 22328 -14372
rect 22224 -14452 22244 -14388
rect 22308 -14452 22328 -14388
rect 22224 -14468 22328 -14452
rect 22224 -14532 22244 -14468
rect 22308 -14532 22328 -14468
rect 22224 -14548 22328 -14532
rect 22224 -14612 22244 -14548
rect 22308 -14612 22328 -14548
rect 22224 -14628 22328 -14612
rect 22224 -14692 22244 -14628
rect 22308 -14692 22328 -14628
rect 22224 -14708 22328 -14692
rect 22224 -14772 22244 -14708
rect 22308 -14772 22328 -14708
rect 22224 -14788 22328 -14772
rect 22224 -14852 22244 -14788
rect 22308 -14852 22328 -14788
rect 22224 -14868 22328 -14852
rect 22224 -14932 22244 -14868
rect 22308 -14932 22328 -14868
rect 22224 -14948 22328 -14932
rect 22224 -15012 22244 -14948
rect 22308 -15012 22328 -14948
rect 22224 -15028 22328 -15012
rect 22224 -15092 22244 -15028
rect 22308 -15092 22328 -15028
rect 22224 -15108 22328 -15092
rect 22224 -15172 22244 -15108
rect 22308 -15172 22328 -15108
rect 22224 -15188 22328 -15172
rect 22224 -15252 22244 -15188
rect 22308 -15252 22328 -15188
rect 22224 -15268 22328 -15252
rect 22224 -15332 22244 -15268
rect 22308 -15332 22328 -15268
rect 22224 -15348 22328 -15332
rect 22224 -15412 22244 -15348
rect 22308 -15412 22328 -15348
rect 22224 -15428 22328 -15412
rect 22224 -15492 22244 -15428
rect 22308 -15492 22328 -15428
rect 22224 -15508 22328 -15492
rect 22224 -15572 22244 -15508
rect 22308 -15572 22328 -15508
rect 22224 -15588 22328 -15572
rect 22224 -15652 22244 -15588
rect 22308 -15652 22328 -15588
rect 22224 -15668 22328 -15652
rect 22224 -15732 22244 -15668
rect 22308 -15732 22328 -15668
rect 22224 -15748 22328 -15732
rect 16612 -16108 16716 -15812
rect 11000 -16188 11104 -16172
rect 11000 -16252 11020 -16188
rect 11084 -16252 11104 -16188
rect 11000 -16268 11104 -16252
rect 11000 -16332 11020 -16268
rect 11084 -16332 11104 -16268
rect 11000 -16348 11104 -16332
rect 11000 -16412 11020 -16348
rect 11084 -16412 11104 -16348
rect 11000 -16428 11104 -16412
rect 11000 -16492 11020 -16428
rect 11084 -16492 11104 -16428
rect 11000 -16508 11104 -16492
rect 11000 -16572 11020 -16508
rect 11084 -16572 11104 -16508
rect 11000 -16588 11104 -16572
rect 11000 -16652 11020 -16588
rect 11084 -16652 11104 -16588
rect 11000 -16668 11104 -16652
rect 11000 -16732 11020 -16668
rect 11084 -16732 11104 -16668
rect 11000 -16748 11104 -16732
rect 11000 -16812 11020 -16748
rect 11084 -16812 11104 -16748
rect 11000 -16828 11104 -16812
rect 11000 -16892 11020 -16828
rect 11084 -16892 11104 -16828
rect 11000 -16908 11104 -16892
rect 11000 -16972 11020 -16908
rect 11084 -16972 11104 -16908
rect 11000 -16988 11104 -16972
rect 11000 -17052 11020 -16988
rect 11084 -17052 11104 -16988
rect 11000 -17068 11104 -17052
rect 11000 -17132 11020 -17068
rect 11084 -17132 11104 -17068
rect 11000 -17148 11104 -17132
rect 11000 -17212 11020 -17148
rect 11084 -17212 11104 -17148
rect 11000 -17228 11104 -17212
rect 11000 -17292 11020 -17228
rect 11084 -17292 11104 -17228
rect 11000 -17308 11104 -17292
rect 11000 -17372 11020 -17308
rect 11084 -17372 11104 -17308
rect 11000 -17388 11104 -17372
rect 11000 -17452 11020 -17388
rect 11084 -17452 11104 -17388
rect 11000 -17468 11104 -17452
rect 11000 -17532 11020 -17468
rect 11084 -17532 11104 -17468
rect 11000 -17548 11104 -17532
rect 11000 -17612 11020 -17548
rect 11084 -17612 11104 -17548
rect 11000 -17628 11104 -17612
rect 11000 -17692 11020 -17628
rect 11084 -17692 11104 -17628
rect 11000 -17708 11104 -17692
rect 11000 -17772 11020 -17708
rect 11084 -17772 11104 -17708
rect 11000 -17788 11104 -17772
rect 11000 -17852 11020 -17788
rect 11084 -17852 11104 -17788
rect 11000 -17868 11104 -17852
rect 11000 -17932 11020 -17868
rect 11084 -17932 11104 -17868
rect 11000 -17948 11104 -17932
rect 11000 -18012 11020 -17948
rect 11084 -18012 11104 -17948
rect 11000 -18028 11104 -18012
rect 11000 -18092 11020 -18028
rect 11084 -18092 11104 -18028
rect 11000 -18108 11104 -18092
rect 11000 -18172 11020 -18108
rect 11084 -18172 11104 -18108
rect 11000 -18188 11104 -18172
rect 11000 -18252 11020 -18188
rect 11084 -18252 11104 -18188
rect 11000 -18268 11104 -18252
rect 11000 -18332 11020 -18268
rect 11084 -18332 11104 -18268
rect 11000 -18348 11104 -18332
rect 11000 -18412 11020 -18348
rect 11084 -18412 11104 -18348
rect 11000 -18428 11104 -18412
rect 11000 -18492 11020 -18428
rect 11084 -18492 11104 -18428
rect 11000 -18508 11104 -18492
rect 11000 -18572 11020 -18508
rect 11084 -18572 11104 -18508
rect 11000 -18588 11104 -18572
rect 11000 -18652 11020 -18588
rect 11084 -18652 11104 -18588
rect 11000 -18668 11104 -18652
rect 11000 -18732 11020 -18668
rect 11084 -18732 11104 -18668
rect 11000 -18748 11104 -18732
rect 11000 -18812 11020 -18748
rect 11084 -18812 11104 -18748
rect 11000 -18828 11104 -18812
rect 11000 -18892 11020 -18828
rect 11084 -18892 11104 -18828
rect 11000 -18908 11104 -18892
rect 11000 -18972 11020 -18908
rect 11084 -18972 11104 -18908
rect 11000 -18988 11104 -18972
rect 11000 -19052 11020 -18988
rect 11084 -19052 11104 -18988
rect 11000 -19068 11104 -19052
rect 11000 -19132 11020 -19068
rect 11084 -19132 11104 -19068
rect 11000 -19148 11104 -19132
rect 11000 -19212 11020 -19148
rect 11084 -19212 11104 -19148
rect 11000 -19228 11104 -19212
rect 11000 -19292 11020 -19228
rect 11084 -19292 11104 -19228
rect 11000 -19308 11104 -19292
rect 11000 -19372 11020 -19308
rect 11084 -19372 11104 -19308
rect 11000 -19388 11104 -19372
rect 11000 -19452 11020 -19388
rect 11084 -19452 11104 -19388
rect 11000 -19468 11104 -19452
rect 11000 -19532 11020 -19468
rect 11084 -19532 11104 -19468
rect 11000 -19548 11104 -19532
rect 11000 -19612 11020 -19548
rect 11084 -19612 11104 -19548
rect 11000 -19628 11104 -19612
rect 11000 -19692 11020 -19628
rect 11084 -19692 11104 -19628
rect 11000 -19708 11104 -19692
rect 11000 -19772 11020 -19708
rect 11084 -19772 11104 -19708
rect 11000 -19788 11104 -19772
rect 11000 -19852 11020 -19788
rect 11084 -19852 11104 -19788
rect 11000 -19868 11104 -19852
rect 11000 -19932 11020 -19868
rect 11084 -19932 11104 -19868
rect 11000 -19948 11104 -19932
rect 11000 -20012 11020 -19948
rect 11084 -20012 11104 -19948
rect 11000 -20028 11104 -20012
rect 11000 -20092 11020 -20028
rect 11084 -20092 11104 -20028
rect 11000 -20108 11104 -20092
rect 11000 -20172 11020 -20108
rect 11084 -20172 11104 -20108
rect 11000 -20188 11104 -20172
rect 11000 -20252 11020 -20188
rect 11084 -20252 11104 -20188
rect 11000 -20268 11104 -20252
rect 11000 -20332 11020 -20268
rect 11084 -20332 11104 -20268
rect 11000 -20348 11104 -20332
rect 11000 -20412 11020 -20348
rect 11084 -20412 11104 -20348
rect 11000 -20428 11104 -20412
rect 11000 -20492 11020 -20428
rect 11084 -20492 11104 -20428
rect 11000 -20508 11104 -20492
rect 11000 -20572 11020 -20508
rect 11084 -20572 11104 -20508
rect 11000 -20588 11104 -20572
rect 11000 -20652 11020 -20588
rect 11084 -20652 11104 -20588
rect 11000 -20668 11104 -20652
rect 11000 -20732 11020 -20668
rect 11084 -20732 11104 -20668
rect 11000 -20748 11104 -20732
rect 11000 -20812 11020 -20748
rect 11084 -20812 11104 -20748
rect 11000 -20828 11104 -20812
rect 11000 -20892 11020 -20828
rect 11084 -20892 11104 -20828
rect 11000 -20908 11104 -20892
rect 11000 -20972 11020 -20908
rect 11084 -20972 11104 -20908
rect 11000 -20988 11104 -20972
rect 11000 -21052 11020 -20988
rect 11084 -21052 11104 -20988
rect 11000 -21068 11104 -21052
rect 5388 -21428 5492 -21132
rect -224 -21508 -120 -21492
rect -224 -21572 -204 -21508
rect -140 -21572 -120 -21508
rect -224 -21588 -120 -21572
rect -224 -21652 -204 -21588
rect -140 -21652 -120 -21588
rect -224 -21668 -120 -21652
rect -224 -21732 -204 -21668
rect -140 -21732 -120 -21668
rect -224 -21748 -120 -21732
rect -224 -21812 -204 -21748
rect -140 -21812 -120 -21748
rect -224 -21828 -120 -21812
rect -224 -21892 -204 -21828
rect -140 -21892 -120 -21828
rect -224 -21908 -120 -21892
rect -224 -21972 -204 -21908
rect -140 -21972 -120 -21908
rect -224 -21988 -120 -21972
rect -224 -22052 -204 -21988
rect -140 -22052 -120 -21988
rect -224 -22068 -120 -22052
rect -224 -22132 -204 -22068
rect -140 -22132 -120 -22068
rect -224 -22148 -120 -22132
rect -224 -22212 -204 -22148
rect -140 -22212 -120 -22148
rect -224 -22228 -120 -22212
rect -224 -22292 -204 -22228
rect -140 -22292 -120 -22228
rect -224 -22308 -120 -22292
rect -224 -22372 -204 -22308
rect -140 -22372 -120 -22308
rect -224 -22388 -120 -22372
rect -224 -22452 -204 -22388
rect -140 -22452 -120 -22388
rect -224 -22468 -120 -22452
rect -224 -22532 -204 -22468
rect -140 -22532 -120 -22468
rect -224 -22548 -120 -22532
rect -224 -22612 -204 -22548
rect -140 -22612 -120 -22548
rect -224 -22628 -120 -22612
rect -224 -22692 -204 -22628
rect -140 -22692 -120 -22628
rect -224 -22708 -120 -22692
rect -224 -22772 -204 -22708
rect -140 -22772 -120 -22708
rect -224 -22788 -120 -22772
rect -224 -22852 -204 -22788
rect -140 -22852 -120 -22788
rect -224 -22868 -120 -22852
rect -224 -22932 -204 -22868
rect -140 -22932 -120 -22868
rect -224 -22948 -120 -22932
rect -224 -23012 -204 -22948
rect -140 -23012 -120 -22948
rect -224 -23028 -120 -23012
rect -224 -23092 -204 -23028
rect -140 -23092 -120 -23028
rect -224 -23108 -120 -23092
rect -224 -23172 -204 -23108
rect -140 -23172 -120 -23108
rect -224 -23188 -120 -23172
rect -224 -23252 -204 -23188
rect -140 -23252 -120 -23188
rect -224 -23268 -120 -23252
rect -224 -23332 -204 -23268
rect -140 -23332 -120 -23268
rect -224 -23348 -120 -23332
rect -224 -23412 -204 -23348
rect -140 -23412 -120 -23348
rect -224 -23428 -120 -23412
rect -224 -23492 -204 -23428
rect -140 -23492 -120 -23428
rect -224 -23508 -120 -23492
rect -224 -23572 -204 -23508
rect -140 -23572 -120 -23508
rect -224 -23588 -120 -23572
rect -224 -23652 -204 -23588
rect -140 -23652 -120 -23588
rect -224 -23668 -120 -23652
rect -224 -23732 -204 -23668
rect -140 -23732 -120 -23668
rect -224 -23748 -120 -23732
rect -224 -23812 -204 -23748
rect -140 -23812 -120 -23748
rect -224 -23828 -120 -23812
rect -224 -23892 -204 -23828
rect -140 -23892 -120 -23828
rect -224 -23908 -120 -23892
rect -224 -23972 -204 -23908
rect -140 -23972 -120 -23908
rect -224 -23988 -120 -23972
rect -224 -24052 -204 -23988
rect -140 -24052 -120 -23988
rect -224 -24068 -120 -24052
rect -224 -24132 -204 -24068
rect -140 -24132 -120 -24068
rect -224 -24148 -120 -24132
rect -224 -24212 -204 -24148
rect -140 -24212 -120 -24148
rect -224 -24228 -120 -24212
rect -224 -24292 -204 -24228
rect -140 -24292 -120 -24228
rect -224 -24308 -120 -24292
rect -224 -24372 -204 -24308
rect -140 -24372 -120 -24308
rect -224 -24388 -120 -24372
rect -224 -24452 -204 -24388
rect -140 -24452 -120 -24388
rect -224 -24468 -120 -24452
rect -224 -24532 -204 -24468
rect -140 -24532 -120 -24468
rect -224 -24548 -120 -24532
rect -224 -24612 -204 -24548
rect -140 -24612 -120 -24548
rect -224 -24628 -120 -24612
rect -224 -24692 -204 -24628
rect -140 -24692 -120 -24628
rect -224 -24708 -120 -24692
rect -224 -24772 -204 -24708
rect -140 -24772 -120 -24708
rect -224 -24788 -120 -24772
rect -224 -24852 -204 -24788
rect -140 -24852 -120 -24788
rect -224 -24868 -120 -24852
rect -224 -24932 -204 -24868
rect -140 -24932 -120 -24868
rect -224 -24948 -120 -24932
rect -224 -25012 -204 -24948
rect -140 -25012 -120 -24948
rect -224 -25028 -120 -25012
rect -224 -25092 -204 -25028
rect -140 -25092 -120 -25028
rect -224 -25108 -120 -25092
rect -224 -25172 -204 -25108
rect -140 -25172 -120 -25108
rect -224 -25188 -120 -25172
rect -224 -25252 -204 -25188
rect -140 -25252 -120 -25188
rect -224 -25268 -120 -25252
rect -224 -25332 -204 -25268
rect -140 -25332 -120 -25268
rect -224 -25348 -120 -25332
rect -224 -25412 -204 -25348
rect -140 -25412 -120 -25348
rect -224 -25428 -120 -25412
rect -224 -25492 -204 -25428
rect -140 -25492 -120 -25428
rect -224 -25508 -120 -25492
rect -224 -25572 -204 -25508
rect -140 -25572 -120 -25508
rect -224 -25588 -120 -25572
rect -224 -25652 -204 -25588
rect -140 -25652 -120 -25588
rect -224 -25668 -120 -25652
rect -224 -25732 -204 -25668
rect -140 -25732 -120 -25668
rect -224 -25748 -120 -25732
rect -224 -25812 -204 -25748
rect -140 -25812 -120 -25748
rect -224 -25828 -120 -25812
rect -224 -25892 -204 -25828
rect -140 -25892 -120 -25828
rect -224 -25908 -120 -25892
rect -224 -25972 -204 -25908
rect -140 -25972 -120 -25908
rect -224 -25988 -120 -25972
rect -224 -26052 -204 -25988
rect -140 -26052 -120 -25988
rect -224 -26068 -120 -26052
rect -224 -26132 -204 -26068
rect -140 -26132 -120 -26068
rect -224 -26148 -120 -26132
rect -224 -26212 -204 -26148
rect -140 -26212 -120 -26148
rect -224 -26228 -120 -26212
rect -224 -26292 -204 -26228
rect -140 -26292 -120 -26228
rect -224 -26308 -120 -26292
rect -224 -26372 -204 -26308
rect -140 -26372 -120 -26308
rect -224 -26388 -120 -26372
rect -5836 -26748 -5732 -26452
rect -11448 -26828 -11344 -26812
rect -11448 -26892 -11428 -26828
rect -11364 -26892 -11344 -26828
rect -11448 -26908 -11344 -26892
rect -11448 -26972 -11428 -26908
rect -11364 -26972 -11344 -26908
rect -11448 -26988 -11344 -26972
rect -11448 -27052 -11428 -26988
rect -11364 -27052 -11344 -26988
rect -11448 -27068 -11344 -27052
rect -11448 -27132 -11428 -27068
rect -11364 -27132 -11344 -27068
rect -11448 -27148 -11344 -27132
rect -11448 -27212 -11428 -27148
rect -11364 -27212 -11344 -27148
rect -11448 -27228 -11344 -27212
rect -11448 -27292 -11428 -27228
rect -11364 -27292 -11344 -27228
rect -11448 -27308 -11344 -27292
rect -11448 -27372 -11428 -27308
rect -11364 -27372 -11344 -27308
rect -11448 -27388 -11344 -27372
rect -11448 -27452 -11428 -27388
rect -11364 -27452 -11344 -27388
rect -11448 -27468 -11344 -27452
rect -11448 -27532 -11428 -27468
rect -11364 -27532 -11344 -27468
rect -11448 -27548 -11344 -27532
rect -11448 -27612 -11428 -27548
rect -11364 -27612 -11344 -27548
rect -11448 -27628 -11344 -27612
rect -11448 -27692 -11428 -27628
rect -11364 -27692 -11344 -27628
rect -11448 -27708 -11344 -27692
rect -11448 -27772 -11428 -27708
rect -11364 -27772 -11344 -27708
rect -11448 -27788 -11344 -27772
rect -11448 -27852 -11428 -27788
rect -11364 -27852 -11344 -27788
rect -11448 -27868 -11344 -27852
rect -11448 -27932 -11428 -27868
rect -11364 -27932 -11344 -27868
rect -11448 -27948 -11344 -27932
rect -11448 -28012 -11428 -27948
rect -11364 -28012 -11344 -27948
rect -11448 -28028 -11344 -28012
rect -11448 -28092 -11428 -28028
rect -11364 -28092 -11344 -28028
rect -11448 -28108 -11344 -28092
rect -11448 -28172 -11428 -28108
rect -11364 -28172 -11344 -28108
rect -11448 -28188 -11344 -28172
rect -11448 -28252 -11428 -28188
rect -11364 -28252 -11344 -28188
rect -11448 -28268 -11344 -28252
rect -11448 -28332 -11428 -28268
rect -11364 -28332 -11344 -28268
rect -11448 -28348 -11344 -28332
rect -11448 -28412 -11428 -28348
rect -11364 -28412 -11344 -28348
rect -11448 -28428 -11344 -28412
rect -11448 -28492 -11428 -28428
rect -11364 -28492 -11344 -28428
rect -11448 -28508 -11344 -28492
rect -11448 -28572 -11428 -28508
rect -11364 -28572 -11344 -28508
rect -11448 -28588 -11344 -28572
rect -11448 -28652 -11428 -28588
rect -11364 -28652 -11344 -28588
rect -11448 -28668 -11344 -28652
rect -11448 -28732 -11428 -28668
rect -11364 -28732 -11344 -28668
rect -11448 -28748 -11344 -28732
rect -11448 -28812 -11428 -28748
rect -11364 -28812 -11344 -28748
rect -11448 -28828 -11344 -28812
rect -11448 -28892 -11428 -28828
rect -11364 -28892 -11344 -28828
rect -11448 -28908 -11344 -28892
rect -11448 -28972 -11428 -28908
rect -11364 -28972 -11344 -28908
rect -11448 -28988 -11344 -28972
rect -11448 -29052 -11428 -28988
rect -11364 -29052 -11344 -28988
rect -11448 -29068 -11344 -29052
rect -11448 -29132 -11428 -29068
rect -11364 -29132 -11344 -29068
rect -11448 -29148 -11344 -29132
rect -11448 -29212 -11428 -29148
rect -11364 -29212 -11344 -29148
rect -11448 -29228 -11344 -29212
rect -11448 -29292 -11428 -29228
rect -11364 -29292 -11344 -29228
rect -11448 -29308 -11344 -29292
rect -11448 -29372 -11428 -29308
rect -11364 -29372 -11344 -29308
rect -11448 -29388 -11344 -29372
rect -11448 -29452 -11428 -29388
rect -11364 -29452 -11344 -29388
rect -11448 -29468 -11344 -29452
rect -11448 -29532 -11428 -29468
rect -11364 -29532 -11344 -29468
rect -11448 -29548 -11344 -29532
rect -11448 -29612 -11428 -29548
rect -11364 -29612 -11344 -29548
rect -11448 -29628 -11344 -29612
rect -11448 -29692 -11428 -29628
rect -11364 -29692 -11344 -29628
rect -11448 -29708 -11344 -29692
rect -11448 -29772 -11428 -29708
rect -11364 -29772 -11344 -29708
rect -11448 -29788 -11344 -29772
rect -11448 -29852 -11428 -29788
rect -11364 -29852 -11344 -29788
rect -11448 -29868 -11344 -29852
rect -11448 -29932 -11428 -29868
rect -11364 -29932 -11344 -29868
rect -11448 -29948 -11344 -29932
rect -11448 -30012 -11428 -29948
rect -11364 -30012 -11344 -29948
rect -11448 -30028 -11344 -30012
rect -11448 -30092 -11428 -30028
rect -11364 -30092 -11344 -30028
rect -11448 -30108 -11344 -30092
rect -11448 -30172 -11428 -30108
rect -11364 -30172 -11344 -30108
rect -11448 -30188 -11344 -30172
rect -11448 -30252 -11428 -30188
rect -11364 -30252 -11344 -30188
rect -11448 -30268 -11344 -30252
rect -11448 -30332 -11428 -30268
rect -11364 -30332 -11344 -30268
rect -11448 -30348 -11344 -30332
rect -11448 -30412 -11428 -30348
rect -11364 -30412 -11344 -30348
rect -11448 -30428 -11344 -30412
rect -11448 -30492 -11428 -30428
rect -11364 -30492 -11344 -30428
rect -11448 -30508 -11344 -30492
rect -11448 -30572 -11428 -30508
rect -11364 -30572 -11344 -30508
rect -11448 -30588 -11344 -30572
rect -11448 -30652 -11428 -30588
rect -11364 -30652 -11344 -30588
rect -11448 -30668 -11344 -30652
rect -11448 -30732 -11428 -30668
rect -11364 -30732 -11344 -30668
rect -11448 -30748 -11344 -30732
rect -11448 -30812 -11428 -30748
rect -11364 -30812 -11344 -30748
rect -11448 -30828 -11344 -30812
rect -11448 -30892 -11428 -30828
rect -11364 -30892 -11344 -30828
rect -11448 -30908 -11344 -30892
rect -11448 -30972 -11428 -30908
rect -11364 -30972 -11344 -30908
rect -11448 -30988 -11344 -30972
rect -11448 -31052 -11428 -30988
rect -11364 -31052 -11344 -30988
rect -11448 -31068 -11344 -31052
rect -11448 -31132 -11428 -31068
rect -11364 -31132 -11344 -31068
rect -11448 -31148 -11344 -31132
rect -11448 -31212 -11428 -31148
rect -11364 -31212 -11344 -31148
rect -11448 -31228 -11344 -31212
rect -11448 -31292 -11428 -31228
rect -11364 -31292 -11344 -31228
rect -11448 -31308 -11344 -31292
rect -11448 -31372 -11428 -31308
rect -11364 -31372 -11344 -31308
rect -11448 -31388 -11344 -31372
rect -11448 -31452 -11428 -31388
rect -11364 -31452 -11344 -31388
rect -11448 -31468 -11344 -31452
rect -11448 -31532 -11428 -31468
rect -11364 -31532 -11344 -31468
rect -11448 -31548 -11344 -31532
rect -11448 -31612 -11428 -31548
rect -11364 -31612 -11344 -31548
rect -11448 -31628 -11344 -31612
rect -11448 -31692 -11428 -31628
rect -11364 -31692 -11344 -31628
rect -11448 -31708 -11344 -31692
rect -17060 -32068 -16956 -31772
rect -22672 -32148 -22568 -32132
rect -22672 -32212 -22652 -32148
rect -22588 -32212 -22568 -32148
rect -22672 -32228 -22568 -32212
rect -22672 -32292 -22652 -32228
rect -22588 -32292 -22568 -32228
rect -22672 -32308 -22568 -32292
rect -22672 -32372 -22652 -32308
rect -22588 -32372 -22568 -32308
rect -22672 -32388 -22568 -32372
rect -22672 -32452 -22652 -32388
rect -22588 -32452 -22568 -32388
rect -22672 -32468 -22568 -32452
rect -22672 -32532 -22652 -32468
rect -22588 -32532 -22568 -32468
rect -22672 -32548 -22568 -32532
rect -22672 -32612 -22652 -32548
rect -22588 -32612 -22568 -32548
rect -22672 -32628 -22568 -32612
rect -22672 -32692 -22652 -32628
rect -22588 -32692 -22568 -32628
rect -22672 -32708 -22568 -32692
rect -22672 -32772 -22652 -32708
rect -22588 -32772 -22568 -32708
rect -22672 -32788 -22568 -32772
rect -22672 -32852 -22652 -32788
rect -22588 -32852 -22568 -32788
rect -22672 -32868 -22568 -32852
rect -22672 -32932 -22652 -32868
rect -22588 -32932 -22568 -32868
rect -22672 -32948 -22568 -32932
rect -22672 -33012 -22652 -32948
rect -22588 -33012 -22568 -32948
rect -22672 -33028 -22568 -33012
rect -22672 -33092 -22652 -33028
rect -22588 -33092 -22568 -33028
rect -22672 -33108 -22568 -33092
rect -22672 -33172 -22652 -33108
rect -22588 -33172 -22568 -33108
rect -22672 -33188 -22568 -33172
rect -22672 -33252 -22652 -33188
rect -22588 -33252 -22568 -33188
rect -22672 -33268 -22568 -33252
rect -22672 -33332 -22652 -33268
rect -22588 -33332 -22568 -33268
rect -22672 -33348 -22568 -33332
rect -22672 -33412 -22652 -33348
rect -22588 -33412 -22568 -33348
rect -22672 -33428 -22568 -33412
rect -22672 -33492 -22652 -33428
rect -22588 -33492 -22568 -33428
rect -22672 -33508 -22568 -33492
rect -22672 -33572 -22652 -33508
rect -22588 -33572 -22568 -33508
rect -22672 -33588 -22568 -33572
rect -22672 -33652 -22652 -33588
rect -22588 -33652 -22568 -33588
rect -22672 -33668 -22568 -33652
rect -22672 -33732 -22652 -33668
rect -22588 -33732 -22568 -33668
rect -22672 -33748 -22568 -33732
rect -22672 -33812 -22652 -33748
rect -22588 -33812 -22568 -33748
rect -22672 -33828 -22568 -33812
rect -22672 -33892 -22652 -33828
rect -22588 -33892 -22568 -33828
rect -22672 -33908 -22568 -33892
rect -22672 -33972 -22652 -33908
rect -22588 -33972 -22568 -33908
rect -22672 -33988 -22568 -33972
rect -22672 -34052 -22652 -33988
rect -22588 -34052 -22568 -33988
rect -22672 -34068 -22568 -34052
rect -22672 -34132 -22652 -34068
rect -22588 -34132 -22568 -34068
rect -22672 -34148 -22568 -34132
rect -22672 -34212 -22652 -34148
rect -22588 -34212 -22568 -34148
rect -22672 -34228 -22568 -34212
rect -22672 -34292 -22652 -34228
rect -22588 -34292 -22568 -34228
rect -22672 -34308 -22568 -34292
rect -22672 -34372 -22652 -34308
rect -22588 -34372 -22568 -34308
rect -22672 -34388 -22568 -34372
rect -22672 -34452 -22652 -34388
rect -22588 -34452 -22568 -34388
rect -22672 -34468 -22568 -34452
rect -22672 -34532 -22652 -34468
rect -22588 -34532 -22568 -34468
rect -22672 -34548 -22568 -34532
rect -22672 -34612 -22652 -34548
rect -22588 -34612 -22568 -34548
rect -22672 -34628 -22568 -34612
rect -22672 -34692 -22652 -34628
rect -22588 -34692 -22568 -34628
rect -22672 -34708 -22568 -34692
rect -22672 -34772 -22652 -34708
rect -22588 -34772 -22568 -34708
rect -22672 -34788 -22568 -34772
rect -22672 -34852 -22652 -34788
rect -22588 -34852 -22568 -34788
rect -22672 -34868 -22568 -34852
rect -22672 -34932 -22652 -34868
rect -22588 -34932 -22568 -34868
rect -22672 -34948 -22568 -34932
rect -22672 -35012 -22652 -34948
rect -22588 -35012 -22568 -34948
rect -22672 -35028 -22568 -35012
rect -22672 -35092 -22652 -35028
rect -22588 -35092 -22568 -35028
rect -22672 -35108 -22568 -35092
rect -22672 -35172 -22652 -35108
rect -22588 -35172 -22568 -35108
rect -22672 -35188 -22568 -35172
rect -22672 -35252 -22652 -35188
rect -22588 -35252 -22568 -35188
rect -22672 -35268 -22568 -35252
rect -22672 -35332 -22652 -35268
rect -22588 -35332 -22568 -35268
rect -22672 -35348 -22568 -35332
rect -22672 -35412 -22652 -35348
rect -22588 -35412 -22568 -35348
rect -22672 -35428 -22568 -35412
rect -22672 -35492 -22652 -35428
rect -22588 -35492 -22568 -35428
rect -22672 -35508 -22568 -35492
rect -22672 -35572 -22652 -35508
rect -22588 -35572 -22568 -35508
rect -22672 -35588 -22568 -35572
rect -22672 -35652 -22652 -35588
rect -22588 -35652 -22568 -35588
rect -22672 -35668 -22568 -35652
rect -22672 -35732 -22652 -35668
rect -22588 -35732 -22568 -35668
rect -22672 -35748 -22568 -35732
rect -22672 -35812 -22652 -35748
rect -22588 -35812 -22568 -35748
rect -22672 -35828 -22568 -35812
rect -22672 -35892 -22652 -35828
rect -22588 -35892 -22568 -35828
rect -22672 -35908 -22568 -35892
rect -22672 -35972 -22652 -35908
rect -22588 -35972 -22568 -35908
rect -22672 -35988 -22568 -35972
rect -22672 -36052 -22652 -35988
rect -22588 -36052 -22568 -35988
rect -22672 -36068 -22568 -36052
rect -22672 -36132 -22652 -36068
rect -22588 -36132 -22568 -36068
rect -22672 -36148 -22568 -36132
rect -22672 -36212 -22652 -36148
rect -22588 -36212 -22568 -36148
rect -22672 -36228 -22568 -36212
rect -22672 -36292 -22652 -36228
rect -22588 -36292 -22568 -36228
rect -22672 -36308 -22568 -36292
rect -22672 -36372 -22652 -36308
rect -22588 -36372 -22568 -36308
rect -22672 -36388 -22568 -36372
rect -22672 -36452 -22652 -36388
rect -22588 -36452 -22568 -36388
rect -22672 -36468 -22568 -36452
rect -22672 -36532 -22652 -36468
rect -22588 -36532 -22568 -36468
rect -22672 -36548 -22568 -36532
rect -22672 -36612 -22652 -36548
rect -22588 -36612 -22568 -36548
rect -22672 -36628 -22568 -36612
rect -22672 -36692 -22652 -36628
rect -22588 -36692 -22568 -36628
rect -22672 -36708 -22568 -36692
rect -22672 -36772 -22652 -36708
rect -22588 -36772 -22568 -36708
rect -22672 -36788 -22568 -36772
rect -22672 -36852 -22652 -36788
rect -22588 -36852 -22568 -36788
rect -22672 -36868 -22568 -36852
rect -22672 -36932 -22652 -36868
rect -22588 -36932 -22568 -36868
rect -22672 -36948 -22568 -36932
rect -22672 -37012 -22652 -36948
rect -22588 -37012 -22568 -36948
rect -22672 -37028 -22568 -37012
rect -28284 -37240 -28180 -37092
rect -25452 -37240 -25348 -37041
rect -22672 -37092 -22652 -37028
rect -22588 -37092 -22568 -37028
rect -22249 -32148 -17327 -32119
rect -22249 -37012 -22220 -32148
rect -17356 -37012 -17327 -32148
rect -22249 -37041 -17327 -37012
rect -17060 -32132 -17040 -32068
rect -16976 -32132 -16956 -32068
rect -14228 -32119 -14124 -31721
rect -11448 -31772 -11428 -31708
rect -11364 -31772 -11344 -31708
rect -11025 -26828 -6103 -26799
rect -11025 -31692 -10996 -26828
rect -6132 -31692 -6103 -26828
rect -11025 -31721 -6103 -31692
rect -5836 -26812 -5816 -26748
rect -5752 -26812 -5732 -26748
rect -3004 -26799 -2900 -26401
rect -224 -26452 -204 -26388
rect -140 -26452 -120 -26388
rect 199 -21508 5121 -21479
rect 199 -26372 228 -21508
rect 5092 -26372 5121 -21508
rect 199 -26401 5121 -26372
rect 5388 -21492 5408 -21428
rect 5472 -21492 5492 -21428
rect 8220 -21479 8324 -21081
rect 11000 -21132 11020 -21068
rect 11084 -21132 11104 -21068
rect 11423 -16188 16345 -16159
rect 11423 -21052 11452 -16188
rect 16316 -21052 16345 -16188
rect 11423 -21081 16345 -21052
rect 16612 -16172 16632 -16108
rect 16696 -16172 16716 -16108
rect 19444 -16159 19548 -15761
rect 22224 -15812 22244 -15748
rect 22308 -15812 22328 -15748
rect 22647 -10868 27569 -10839
rect 22647 -15732 22676 -10868
rect 27540 -15732 27569 -10868
rect 22647 -15761 27569 -15732
rect 27836 -10852 27856 -10788
rect 27920 -10852 27940 -10788
rect 30668 -10839 30772 -10441
rect 33448 -10492 33468 -10428
rect 33532 -10492 33552 -10428
rect 33871 -5548 38793 -5519
rect 33871 -10412 33900 -5548
rect 38764 -10412 38793 -5548
rect 33871 -10441 38793 -10412
rect 39060 -5532 39080 -5468
rect 39144 -5532 39164 -5468
rect 39060 -5548 39164 -5532
rect 39060 -5612 39080 -5548
rect 39144 -5612 39164 -5548
rect 39060 -5628 39164 -5612
rect 39060 -5692 39080 -5628
rect 39144 -5692 39164 -5628
rect 39060 -5708 39164 -5692
rect 39060 -5772 39080 -5708
rect 39144 -5772 39164 -5708
rect 39060 -5788 39164 -5772
rect 39060 -5852 39080 -5788
rect 39144 -5852 39164 -5788
rect 39060 -5868 39164 -5852
rect 39060 -5932 39080 -5868
rect 39144 -5932 39164 -5868
rect 39060 -5948 39164 -5932
rect 39060 -6012 39080 -5948
rect 39144 -6012 39164 -5948
rect 39060 -6028 39164 -6012
rect 39060 -6092 39080 -6028
rect 39144 -6092 39164 -6028
rect 39060 -6108 39164 -6092
rect 39060 -6172 39080 -6108
rect 39144 -6172 39164 -6108
rect 39060 -6188 39164 -6172
rect 39060 -6252 39080 -6188
rect 39144 -6252 39164 -6188
rect 39060 -6268 39164 -6252
rect 39060 -6332 39080 -6268
rect 39144 -6332 39164 -6268
rect 39060 -6348 39164 -6332
rect 39060 -6412 39080 -6348
rect 39144 -6412 39164 -6348
rect 39060 -6428 39164 -6412
rect 39060 -6492 39080 -6428
rect 39144 -6492 39164 -6428
rect 39060 -6508 39164 -6492
rect 39060 -6572 39080 -6508
rect 39144 -6572 39164 -6508
rect 39060 -6588 39164 -6572
rect 39060 -6652 39080 -6588
rect 39144 -6652 39164 -6588
rect 39060 -6668 39164 -6652
rect 39060 -6732 39080 -6668
rect 39144 -6732 39164 -6668
rect 39060 -6748 39164 -6732
rect 39060 -6812 39080 -6748
rect 39144 -6812 39164 -6748
rect 39060 -6828 39164 -6812
rect 39060 -6892 39080 -6828
rect 39144 -6892 39164 -6828
rect 39060 -6908 39164 -6892
rect 39060 -6972 39080 -6908
rect 39144 -6972 39164 -6908
rect 39060 -6988 39164 -6972
rect 39060 -7052 39080 -6988
rect 39144 -7052 39164 -6988
rect 39060 -7068 39164 -7052
rect 39060 -7132 39080 -7068
rect 39144 -7132 39164 -7068
rect 39060 -7148 39164 -7132
rect 39060 -7212 39080 -7148
rect 39144 -7212 39164 -7148
rect 39060 -7228 39164 -7212
rect 39060 -7292 39080 -7228
rect 39144 -7292 39164 -7228
rect 39060 -7308 39164 -7292
rect 39060 -7372 39080 -7308
rect 39144 -7372 39164 -7308
rect 39060 -7388 39164 -7372
rect 39060 -7452 39080 -7388
rect 39144 -7452 39164 -7388
rect 39060 -7468 39164 -7452
rect 39060 -7532 39080 -7468
rect 39144 -7532 39164 -7468
rect 39060 -7548 39164 -7532
rect 39060 -7612 39080 -7548
rect 39144 -7612 39164 -7548
rect 39060 -7628 39164 -7612
rect 39060 -7692 39080 -7628
rect 39144 -7692 39164 -7628
rect 39060 -7708 39164 -7692
rect 39060 -7772 39080 -7708
rect 39144 -7772 39164 -7708
rect 39060 -7788 39164 -7772
rect 39060 -7852 39080 -7788
rect 39144 -7852 39164 -7788
rect 39060 -7868 39164 -7852
rect 39060 -7932 39080 -7868
rect 39144 -7932 39164 -7868
rect 39060 -7948 39164 -7932
rect 39060 -8012 39080 -7948
rect 39144 -8012 39164 -7948
rect 39060 -8028 39164 -8012
rect 39060 -8092 39080 -8028
rect 39144 -8092 39164 -8028
rect 39060 -8108 39164 -8092
rect 39060 -8172 39080 -8108
rect 39144 -8172 39164 -8108
rect 39060 -8188 39164 -8172
rect 39060 -8252 39080 -8188
rect 39144 -8252 39164 -8188
rect 39060 -8268 39164 -8252
rect 39060 -8332 39080 -8268
rect 39144 -8332 39164 -8268
rect 39060 -8348 39164 -8332
rect 39060 -8412 39080 -8348
rect 39144 -8412 39164 -8348
rect 39060 -8428 39164 -8412
rect 39060 -8492 39080 -8428
rect 39144 -8492 39164 -8428
rect 39060 -8508 39164 -8492
rect 39060 -8572 39080 -8508
rect 39144 -8572 39164 -8508
rect 39060 -8588 39164 -8572
rect 39060 -8652 39080 -8588
rect 39144 -8652 39164 -8588
rect 39060 -8668 39164 -8652
rect 39060 -8732 39080 -8668
rect 39144 -8732 39164 -8668
rect 39060 -8748 39164 -8732
rect 39060 -8812 39080 -8748
rect 39144 -8812 39164 -8748
rect 39060 -8828 39164 -8812
rect 39060 -8892 39080 -8828
rect 39144 -8892 39164 -8828
rect 39060 -8908 39164 -8892
rect 39060 -8972 39080 -8908
rect 39144 -8972 39164 -8908
rect 39060 -8988 39164 -8972
rect 39060 -9052 39080 -8988
rect 39144 -9052 39164 -8988
rect 39060 -9068 39164 -9052
rect 39060 -9132 39080 -9068
rect 39144 -9132 39164 -9068
rect 39060 -9148 39164 -9132
rect 39060 -9212 39080 -9148
rect 39144 -9212 39164 -9148
rect 39060 -9228 39164 -9212
rect 39060 -9292 39080 -9228
rect 39144 -9292 39164 -9228
rect 39060 -9308 39164 -9292
rect 39060 -9372 39080 -9308
rect 39144 -9372 39164 -9308
rect 39060 -9388 39164 -9372
rect 39060 -9452 39080 -9388
rect 39144 -9452 39164 -9388
rect 39060 -9468 39164 -9452
rect 39060 -9532 39080 -9468
rect 39144 -9532 39164 -9468
rect 39060 -9548 39164 -9532
rect 39060 -9612 39080 -9548
rect 39144 -9612 39164 -9548
rect 39060 -9628 39164 -9612
rect 39060 -9692 39080 -9628
rect 39144 -9692 39164 -9628
rect 39060 -9708 39164 -9692
rect 39060 -9772 39080 -9708
rect 39144 -9772 39164 -9708
rect 39060 -9788 39164 -9772
rect 39060 -9852 39080 -9788
rect 39144 -9852 39164 -9788
rect 39060 -9868 39164 -9852
rect 39060 -9932 39080 -9868
rect 39144 -9932 39164 -9868
rect 39060 -9948 39164 -9932
rect 39060 -10012 39080 -9948
rect 39144 -10012 39164 -9948
rect 39060 -10028 39164 -10012
rect 39060 -10092 39080 -10028
rect 39144 -10092 39164 -10028
rect 39060 -10108 39164 -10092
rect 39060 -10172 39080 -10108
rect 39144 -10172 39164 -10108
rect 39060 -10188 39164 -10172
rect 39060 -10252 39080 -10188
rect 39144 -10252 39164 -10188
rect 39060 -10268 39164 -10252
rect 39060 -10332 39080 -10268
rect 39144 -10332 39164 -10268
rect 39060 -10348 39164 -10332
rect 39060 -10412 39080 -10348
rect 39144 -10412 39164 -10348
rect 39060 -10428 39164 -10412
rect 33448 -10788 33552 -10492
rect 27836 -10868 27940 -10852
rect 27836 -10932 27856 -10868
rect 27920 -10932 27940 -10868
rect 27836 -10948 27940 -10932
rect 27836 -11012 27856 -10948
rect 27920 -11012 27940 -10948
rect 27836 -11028 27940 -11012
rect 27836 -11092 27856 -11028
rect 27920 -11092 27940 -11028
rect 27836 -11108 27940 -11092
rect 27836 -11172 27856 -11108
rect 27920 -11172 27940 -11108
rect 27836 -11188 27940 -11172
rect 27836 -11252 27856 -11188
rect 27920 -11252 27940 -11188
rect 27836 -11268 27940 -11252
rect 27836 -11332 27856 -11268
rect 27920 -11332 27940 -11268
rect 27836 -11348 27940 -11332
rect 27836 -11412 27856 -11348
rect 27920 -11412 27940 -11348
rect 27836 -11428 27940 -11412
rect 27836 -11492 27856 -11428
rect 27920 -11492 27940 -11428
rect 27836 -11508 27940 -11492
rect 27836 -11572 27856 -11508
rect 27920 -11572 27940 -11508
rect 27836 -11588 27940 -11572
rect 27836 -11652 27856 -11588
rect 27920 -11652 27940 -11588
rect 27836 -11668 27940 -11652
rect 27836 -11732 27856 -11668
rect 27920 -11732 27940 -11668
rect 27836 -11748 27940 -11732
rect 27836 -11812 27856 -11748
rect 27920 -11812 27940 -11748
rect 27836 -11828 27940 -11812
rect 27836 -11892 27856 -11828
rect 27920 -11892 27940 -11828
rect 27836 -11908 27940 -11892
rect 27836 -11972 27856 -11908
rect 27920 -11972 27940 -11908
rect 27836 -11988 27940 -11972
rect 27836 -12052 27856 -11988
rect 27920 -12052 27940 -11988
rect 27836 -12068 27940 -12052
rect 27836 -12132 27856 -12068
rect 27920 -12132 27940 -12068
rect 27836 -12148 27940 -12132
rect 27836 -12212 27856 -12148
rect 27920 -12212 27940 -12148
rect 27836 -12228 27940 -12212
rect 27836 -12292 27856 -12228
rect 27920 -12292 27940 -12228
rect 27836 -12308 27940 -12292
rect 27836 -12372 27856 -12308
rect 27920 -12372 27940 -12308
rect 27836 -12388 27940 -12372
rect 27836 -12452 27856 -12388
rect 27920 -12452 27940 -12388
rect 27836 -12468 27940 -12452
rect 27836 -12532 27856 -12468
rect 27920 -12532 27940 -12468
rect 27836 -12548 27940 -12532
rect 27836 -12612 27856 -12548
rect 27920 -12612 27940 -12548
rect 27836 -12628 27940 -12612
rect 27836 -12692 27856 -12628
rect 27920 -12692 27940 -12628
rect 27836 -12708 27940 -12692
rect 27836 -12772 27856 -12708
rect 27920 -12772 27940 -12708
rect 27836 -12788 27940 -12772
rect 27836 -12852 27856 -12788
rect 27920 -12852 27940 -12788
rect 27836 -12868 27940 -12852
rect 27836 -12932 27856 -12868
rect 27920 -12932 27940 -12868
rect 27836 -12948 27940 -12932
rect 27836 -13012 27856 -12948
rect 27920 -13012 27940 -12948
rect 27836 -13028 27940 -13012
rect 27836 -13092 27856 -13028
rect 27920 -13092 27940 -13028
rect 27836 -13108 27940 -13092
rect 27836 -13172 27856 -13108
rect 27920 -13172 27940 -13108
rect 27836 -13188 27940 -13172
rect 27836 -13252 27856 -13188
rect 27920 -13252 27940 -13188
rect 27836 -13268 27940 -13252
rect 27836 -13332 27856 -13268
rect 27920 -13332 27940 -13268
rect 27836 -13348 27940 -13332
rect 27836 -13412 27856 -13348
rect 27920 -13412 27940 -13348
rect 27836 -13428 27940 -13412
rect 27836 -13492 27856 -13428
rect 27920 -13492 27940 -13428
rect 27836 -13508 27940 -13492
rect 27836 -13572 27856 -13508
rect 27920 -13572 27940 -13508
rect 27836 -13588 27940 -13572
rect 27836 -13652 27856 -13588
rect 27920 -13652 27940 -13588
rect 27836 -13668 27940 -13652
rect 27836 -13732 27856 -13668
rect 27920 -13732 27940 -13668
rect 27836 -13748 27940 -13732
rect 27836 -13812 27856 -13748
rect 27920 -13812 27940 -13748
rect 27836 -13828 27940 -13812
rect 27836 -13892 27856 -13828
rect 27920 -13892 27940 -13828
rect 27836 -13908 27940 -13892
rect 27836 -13972 27856 -13908
rect 27920 -13972 27940 -13908
rect 27836 -13988 27940 -13972
rect 27836 -14052 27856 -13988
rect 27920 -14052 27940 -13988
rect 27836 -14068 27940 -14052
rect 27836 -14132 27856 -14068
rect 27920 -14132 27940 -14068
rect 27836 -14148 27940 -14132
rect 27836 -14212 27856 -14148
rect 27920 -14212 27940 -14148
rect 27836 -14228 27940 -14212
rect 27836 -14292 27856 -14228
rect 27920 -14292 27940 -14228
rect 27836 -14308 27940 -14292
rect 27836 -14372 27856 -14308
rect 27920 -14372 27940 -14308
rect 27836 -14388 27940 -14372
rect 27836 -14452 27856 -14388
rect 27920 -14452 27940 -14388
rect 27836 -14468 27940 -14452
rect 27836 -14532 27856 -14468
rect 27920 -14532 27940 -14468
rect 27836 -14548 27940 -14532
rect 27836 -14612 27856 -14548
rect 27920 -14612 27940 -14548
rect 27836 -14628 27940 -14612
rect 27836 -14692 27856 -14628
rect 27920 -14692 27940 -14628
rect 27836 -14708 27940 -14692
rect 27836 -14772 27856 -14708
rect 27920 -14772 27940 -14708
rect 27836 -14788 27940 -14772
rect 27836 -14852 27856 -14788
rect 27920 -14852 27940 -14788
rect 27836 -14868 27940 -14852
rect 27836 -14932 27856 -14868
rect 27920 -14932 27940 -14868
rect 27836 -14948 27940 -14932
rect 27836 -15012 27856 -14948
rect 27920 -15012 27940 -14948
rect 27836 -15028 27940 -15012
rect 27836 -15092 27856 -15028
rect 27920 -15092 27940 -15028
rect 27836 -15108 27940 -15092
rect 27836 -15172 27856 -15108
rect 27920 -15172 27940 -15108
rect 27836 -15188 27940 -15172
rect 27836 -15252 27856 -15188
rect 27920 -15252 27940 -15188
rect 27836 -15268 27940 -15252
rect 27836 -15332 27856 -15268
rect 27920 -15332 27940 -15268
rect 27836 -15348 27940 -15332
rect 27836 -15412 27856 -15348
rect 27920 -15412 27940 -15348
rect 27836 -15428 27940 -15412
rect 27836 -15492 27856 -15428
rect 27920 -15492 27940 -15428
rect 27836 -15508 27940 -15492
rect 27836 -15572 27856 -15508
rect 27920 -15572 27940 -15508
rect 27836 -15588 27940 -15572
rect 27836 -15652 27856 -15588
rect 27920 -15652 27940 -15588
rect 27836 -15668 27940 -15652
rect 27836 -15732 27856 -15668
rect 27920 -15732 27940 -15668
rect 27836 -15748 27940 -15732
rect 22224 -16108 22328 -15812
rect 16612 -16188 16716 -16172
rect 16612 -16252 16632 -16188
rect 16696 -16252 16716 -16188
rect 16612 -16268 16716 -16252
rect 16612 -16332 16632 -16268
rect 16696 -16332 16716 -16268
rect 16612 -16348 16716 -16332
rect 16612 -16412 16632 -16348
rect 16696 -16412 16716 -16348
rect 16612 -16428 16716 -16412
rect 16612 -16492 16632 -16428
rect 16696 -16492 16716 -16428
rect 16612 -16508 16716 -16492
rect 16612 -16572 16632 -16508
rect 16696 -16572 16716 -16508
rect 16612 -16588 16716 -16572
rect 16612 -16652 16632 -16588
rect 16696 -16652 16716 -16588
rect 16612 -16668 16716 -16652
rect 16612 -16732 16632 -16668
rect 16696 -16732 16716 -16668
rect 16612 -16748 16716 -16732
rect 16612 -16812 16632 -16748
rect 16696 -16812 16716 -16748
rect 16612 -16828 16716 -16812
rect 16612 -16892 16632 -16828
rect 16696 -16892 16716 -16828
rect 16612 -16908 16716 -16892
rect 16612 -16972 16632 -16908
rect 16696 -16972 16716 -16908
rect 16612 -16988 16716 -16972
rect 16612 -17052 16632 -16988
rect 16696 -17052 16716 -16988
rect 16612 -17068 16716 -17052
rect 16612 -17132 16632 -17068
rect 16696 -17132 16716 -17068
rect 16612 -17148 16716 -17132
rect 16612 -17212 16632 -17148
rect 16696 -17212 16716 -17148
rect 16612 -17228 16716 -17212
rect 16612 -17292 16632 -17228
rect 16696 -17292 16716 -17228
rect 16612 -17308 16716 -17292
rect 16612 -17372 16632 -17308
rect 16696 -17372 16716 -17308
rect 16612 -17388 16716 -17372
rect 16612 -17452 16632 -17388
rect 16696 -17452 16716 -17388
rect 16612 -17468 16716 -17452
rect 16612 -17532 16632 -17468
rect 16696 -17532 16716 -17468
rect 16612 -17548 16716 -17532
rect 16612 -17612 16632 -17548
rect 16696 -17612 16716 -17548
rect 16612 -17628 16716 -17612
rect 16612 -17692 16632 -17628
rect 16696 -17692 16716 -17628
rect 16612 -17708 16716 -17692
rect 16612 -17772 16632 -17708
rect 16696 -17772 16716 -17708
rect 16612 -17788 16716 -17772
rect 16612 -17852 16632 -17788
rect 16696 -17852 16716 -17788
rect 16612 -17868 16716 -17852
rect 16612 -17932 16632 -17868
rect 16696 -17932 16716 -17868
rect 16612 -17948 16716 -17932
rect 16612 -18012 16632 -17948
rect 16696 -18012 16716 -17948
rect 16612 -18028 16716 -18012
rect 16612 -18092 16632 -18028
rect 16696 -18092 16716 -18028
rect 16612 -18108 16716 -18092
rect 16612 -18172 16632 -18108
rect 16696 -18172 16716 -18108
rect 16612 -18188 16716 -18172
rect 16612 -18252 16632 -18188
rect 16696 -18252 16716 -18188
rect 16612 -18268 16716 -18252
rect 16612 -18332 16632 -18268
rect 16696 -18332 16716 -18268
rect 16612 -18348 16716 -18332
rect 16612 -18412 16632 -18348
rect 16696 -18412 16716 -18348
rect 16612 -18428 16716 -18412
rect 16612 -18492 16632 -18428
rect 16696 -18492 16716 -18428
rect 16612 -18508 16716 -18492
rect 16612 -18572 16632 -18508
rect 16696 -18572 16716 -18508
rect 16612 -18588 16716 -18572
rect 16612 -18652 16632 -18588
rect 16696 -18652 16716 -18588
rect 16612 -18668 16716 -18652
rect 16612 -18732 16632 -18668
rect 16696 -18732 16716 -18668
rect 16612 -18748 16716 -18732
rect 16612 -18812 16632 -18748
rect 16696 -18812 16716 -18748
rect 16612 -18828 16716 -18812
rect 16612 -18892 16632 -18828
rect 16696 -18892 16716 -18828
rect 16612 -18908 16716 -18892
rect 16612 -18972 16632 -18908
rect 16696 -18972 16716 -18908
rect 16612 -18988 16716 -18972
rect 16612 -19052 16632 -18988
rect 16696 -19052 16716 -18988
rect 16612 -19068 16716 -19052
rect 16612 -19132 16632 -19068
rect 16696 -19132 16716 -19068
rect 16612 -19148 16716 -19132
rect 16612 -19212 16632 -19148
rect 16696 -19212 16716 -19148
rect 16612 -19228 16716 -19212
rect 16612 -19292 16632 -19228
rect 16696 -19292 16716 -19228
rect 16612 -19308 16716 -19292
rect 16612 -19372 16632 -19308
rect 16696 -19372 16716 -19308
rect 16612 -19388 16716 -19372
rect 16612 -19452 16632 -19388
rect 16696 -19452 16716 -19388
rect 16612 -19468 16716 -19452
rect 16612 -19532 16632 -19468
rect 16696 -19532 16716 -19468
rect 16612 -19548 16716 -19532
rect 16612 -19612 16632 -19548
rect 16696 -19612 16716 -19548
rect 16612 -19628 16716 -19612
rect 16612 -19692 16632 -19628
rect 16696 -19692 16716 -19628
rect 16612 -19708 16716 -19692
rect 16612 -19772 16632 -19708
rect 16696 -19772 16716 -19708
rect 16612 -19788 16716 -19772
rect 16612 -19852 16632 -19788
rect 16696 -19852 16716 -19788
rect 16612 -19868 16716 -19852
rect 16612 -19932 16632 -19868
rect 16696 -19932 16716 -19868
rect 16612 -19948 16716 -19932
rect 16612 -20012 16632 -19948
rect 16696 -20012 16716 -19948
rect 16612 -20028 16716 -20012
rect 16612 -20092 16632 -20028
rect 16696 -20092 16716 -20028
rect 16612 -20108 16716 -20092
rect 16612 -20172 16632 -20108
rect 16696 -20172 16716 -20108
rect 16612 -20188 16716 -20172
rect 16612 -20252 16632 -20188
rect 16696 -20252 16716 -20188
rect 16612 -20268 16716 -20252
rect 16612 -20332 16632 -20268
rect 16696 -20332 16716 -20268
rect 16612 -20348 16716 -20332
rect 16612 -20412 16632 -20348
rect 16696 -20412 16716 -20348
rect 16612 -20428 16716 -20412
rect 16612 -20492 16632 -20428
rect 16696 -20492 16716 -20428
rect 16612 -20508 16716 -20492
rect 16612 -20572 16632 -20508
rect 16696 -20572 16716 -20508
rect 16612 -20588 16716 -20572
rect 16612 -20652 16632 -20588
rect 16696 -20652 16716 -20588
rect 16612 -20668 16716 -20652
rect 16612 -20732 16632 -20668
rect 16696 -20732 16716 -20668
rect 16612 -20748 16716 -20732
rect 16612 -20812 16632 -20748
rect 16696 -20812 16716 -20748
rect 16612 -20828 16716 -20812
rect 16612 -20892 16632 -20828
rect 16696 -20892 16716 -20828
rect 16612 -20908 16716 -20892
rect 16612 -20972 16632 -20908
rect 16696 -20972 16716 -20908
rect 16612 -20988 16716 -20972
rect 16612 -21052 16632 -20988
rect 16696 -21052 16716 -20988
rect 16612 -21068 16716 -21052
rect 11000 -21428 11104 -21132
rect 5388 -21508 5492 -21492
rect 5388 -21572 5408 -21508
rect 5472 -21572 5492 -21508
rect 5388 -21588 5492 -21572
rect 5388 -21652 5408 -21588
rect 5472 -21652 5492 -21588
rect 5388 -21668 5492 -21652
rect 5388 -21732 5408 -21668
rect 5472 -21732 5492 -21668
rect 5388 -21748 5492 -21732
rect 5388 -21812 5408 -21748
rect 5472 -21812 5492 -21748
rect 5388 -21828 5492 -21812
rect 5388 -21892 5408 -21828
rect 5472 -21892 5492 -21828
rect 5388 -21908 5492 -21892
rect 5388 -21972 5408 -21908
rect 5472 -21972 5492 -21908
rect 5388 -21988 5492 -21972
rect 5388 -22052 5408 -21988
rect 5472 -22052 5492 -21988
rect 5388 -22068 5492 -22052
rect 5388 -22132 5408 -22068
rect 5472 -22132 5492 -22068
rect 5388 -22148 5492 -22132
rect 5388 -22212 5408 -22148
rect 5472 -22212 5492 -22148
rect 5388 -22228 5492 -22212
rect 5388 -22292 5408 -22228
rect 5472 -22292 5492 -22228
rect 5388 -22308 5492 -22292
rect 5388 -22372 5408 -22308
rect 5472 -22372 5492 -22308
rect 5388 -22388 5492 -22372
rect 5388 -22452 5408 -22388
rect 5472 -22452 5492 -22388
rect 5388 -22468 5492 -22452
rect 5388 -22532 5408 -22468
rect 5472 -22532 5492 -22468
rect 5388 -22548 5492 -22532
rect 5388 -22612 5408 -22548
rect 5472 -22612 5492 -22548
rect 5388 -22628 5492 -22612
rect 5388 -22692 5408 -22628
rect 5472 -22692 5492 -22628
rect 5388 -22708 5492 -22692
rect 5388 -22772 5408 -22708
rect 5472 -22772 5492 -22708
rect 5388 -22788 5492 -22772
rect 5388 -22852 5408 -22788
rect 5472 -22852 5492 -22788
rect 5388 -22868 5492 -22852
rect 5388 -22932 5408 -22868
rect 5472 -22932 5492 -22868
rect 5388 -22948 5492 -22932
rect 5388 -23012 5408 -22948
rect 5472 -23012 5492 -22948
rect 5388 -23028 5492 -23012
rect 5388 -23092 5408 -23028
rect 5472 -23092 5492 -23028
rect 5388 -23108 5492 -23092
rect 5388 -23172 5408 -23108
rect 5472 -23172 5492 -23108
rect 5388 -23188 5492 -23172
rect 5388 -23252 5408 -23188
rect 5472 -23252 5492 -23188
rect 5388 -23268 5492 -23252
rect 5388 -23332 5408 -23268
rect 5472 -23332 5492 -23268
rect 5388 -23348 5492 -23332
rect 5388 -23412 5408 -23348
rect 5472 -23412 5492 -23348
rect 5388 -23428 5492 -23412
rect 5388 -23492 5408 -23428
rect 5472 -23492 5492 -23428
rect 5388 -23508 5492 -23492
rect 5388 -23572 5408 -23508
rect 5472 -23572 5492 -23508
rect 5388 -23588 5492 -23572
rect 5388 -23652 5408 -23588
rect 5472 -23652 5492 -23588
rect 5388 -23668 5492 -23652
rect 5388 -23732 5408 -23668
rect 5472 -23732 5492 -23668
rect 5388 -23748 5492 -23732
rect 5388 -23812 5408 -23748
rect 5472 -23812 5492 -23748
rect 5388 -23828 5492 -23812
rect 5388 -23892 5408 -23828
rect 5472 -23892 5492 -23828
rect 5388 -23908 5492 -23892
rect 5388 -23972 5408 -23908
rect 5472 -23972 5492 -23908
rect 5388 -23988 5492 -23972
rect 5388 -24052 5408 -23988
rect 5472 -24052 5492 -23988
rect 5388 -24068 5492 -24052
rect 5388 -24132 5408 -24068
rect 5472 -24132 5492 -24068
rect 5388 -24148 5492 -24132
rect 5388 -24212 5408 -24148
rect 5472 -24212 5492 -24148
rect 5388 -24228 5492 -24212
rect 5388 -24292 5408 -24228
rect 5472 -24292 5492 -24228
rect 5388 -24308 5492 -24292
rect 5388 -24372 5408 -24308
rect 5472 -24372 5492 -24308
rect 5388 -24388 5492 -24372
rect 5388 -24452 5408 -24388
rect 5472 -24452 5492 -24388
rect 5388 -24468 5492 -24452
rect 5388 -24532 5408 -24468
rect 5472 -24532 5492 -24468
rect 5388 -24548 5492 -24532
rect 5388 -24612 5408 -24548
rect 5472 -24612 5492 -24548
rect 5388 -24628 5492 -24612
rect 5388 -24692 5408 -24628
rect 5472 -24692 5492 -24628
rect 5388 -24708 5492 -24692
rect 5388 -24772 5408 -24708
rect 5472 -24772 5492 -24708
rect 5388 -24788 5492 -24772
rect 5388 -24852 5408 -24788
rect 5472 -24852 5492 -24788
rect 5388 -24868 5492 -24852
rect 5388 -24932 5408 -24868
rect 5472 -24932 5492 -24868
rect 5388 -24948 5492 -24932
rect 5388 -25012 5408 -24948
rect 5472 -25012 5492 -24948
rect 5388 -25028 5492 -25012
rect 5388 -25092 5408 -25028
rect 5472 -25092 5492 -25028
rect 5388 -25108 5492 -25092
rect 5388 -25172 5408 -25108
rect 5472 -25172 5492 -25108
rect 5388 -25188 5492 -25172
rect 5388 -25252 5408 -25188
rect 5472 -25252 5492 -25188
rect 5388 -25268 5492 -25252
rect 5388 -25332 5408 -25268
rect 5472 -25332 5492 -25268
rect 5388 -25348 5492 -25332
rect 5388 -25412 5408 -25348
rect 5472 -25412 5492 -25348
rect 5388 -25428 5492 -25412
rect 5388 -25492 5408 -25428
rect 5472 -25492 5492 -25428
rect 5388 -25508 5492 -25492
rect 5388 -25572 5408 -25508
rect 5472 -25572 5492 -25508
rect 5388 -25588 5492 -25572
rect 5388 -25652 5408 -25588
rect 5472 -25652 5492 -25588
rect 5388 -25668 5492 -25652
rect 5388 -25732 5408 -25668
rect 5472 -25732 5492 -25668
rect 5388 -25748 5492 -25732
rect 5388 -25812 5408 -25748
rect 5472 -25812 5492 -25748
rect 5388 -25828 5492 -25812
rect 5388 -25892 5408 -25828
rect 5472 -25892 5492 -25828
rect 5388 -25908 5492 -25892
rect 5388 -25972 5408 -25908
rect 5472 -25972 5492 -25908
rect 5388 -25988 5492 -25972
rect 5388 -26052 5408 -25988
rect 5472 -26052 5492 -25988
rect 5388 -26068 5492 -26052
rect 5388 -26132 5408 -26068
rect 5472 -26132 5492 -26068
rect 5388 -26148 5492 -26132
rect 5388 -26212 5408 -26148
rect 5472 -26212 5492 -26148
rect 5388 -26228 5492 -26212
rect 5388 -26292 5408 -26228
rect 5472 -26292 5492 -26228
rect 5388 -26308 5492 -26292
rect 5388 -26372 5408 -26308
rect 5472 -26372 5492 -26308
rect 5388 -26388 5492 -26372
rect -224 -26748 -120 -26452
rect -5836 -26828 -5732 -26812
rect -5836 -26892 -5816 -26828
rect -5752 -26892 -5732 -26828
rect -5836 -26908 -5732 -26892
rect -5836 -26972 -5816 -26908
rect -5752 -26972 -5732 -26908
rect -5836 -26988 -5732 -26972
rect -5836 -27052 -5816 -26988
rect -5752 -27052 -5732 -26988
rect -5836 -27068 -5732 -27052
rect -5836 -27132 -5816 -27068
rect -5752 -27132 -5732 -27068
rect -5836 -27148 -5732 -27132
rect -5836 -27212 -5816 -27148
rect -5752 -27212 -5732 -27148
rect -5836 -27228 -5732 -27212
rect -5836 -27292 -5816 -27228
rect -5752 -27292 -5732 -27228
rect -5836 -27308 -5732 -27292
rect -5836 -27372 -5816 -27308
rect -5752 -27372 -5732 -27308
rect -5836 -27388 -5732 -27372
rect -5836 -27452 -5816 -27388
rect -5752 -27452 -5732 -27388
rect -5836 -27468 -5732 -27452
rect -5836 -27532 -5816 -27468
rect -5752 -27532 -5732 -27468
rect -5836 -27548 -5732 -27532
rect -5836 -27612 -5816 -27548
rect -5752 -27612 -5732 -27548
rect -5836 -27628 -5732 -27612
rect -5836 -27692 -5816 -27628
rect -5752 -27692 -5732 -27628
rect -5836 -27708 -5732 -27692
rect -5836 -27772 -5816 -27708
rect -5752 -27772 -5732 -27708
rect -5836 -27788 -5732 -27772
rect -5836 -27852 -5816 -27788
rect -5752 -27852 -5732 -27788
rect -5836 -27868 -5732 -27852
rect -5836 -27932 -5816 -27868
rect -5752 -27932 -5732 -27868
rect -5836 -27948 -5732 -27932
rect -5836 -28012 -5816 -27948
rect -5752 -28012 -5732 -27948
rect -5836 -28028 -5732 -28012
rect -5836 -28092 -5816 -28028
rect -5752 -28092 -5732 -28028
rect -5836 -28108 -5732 -28092
rect -5836 -28172 -5816 -28108
rect -5752 -28172 -5732 -28108
rect -5836 -28188 -5732 -28172
rect -5836 -28252 -5816 -28188
rect -5752 -28252 -5732 -28188
rect -5836 -28268 -5732 -28252
rect -5836 -28332 -5816 -28268
rect -5752 -28332 -5732 -28268
rect -5836 -28348 -5732 -28332
rect -5836 -28412 -5816 -28348
rect -5752 -28412 -5732 -28348
rect -5836 -28428 -5732 -28412
rect -5836 -28492 -5816 -28428
rect -5752 -28492 -5732 -28428
rect -5836 -28508 -5732 -28492
rect -5836 -28572 -5816 -28508
rect -5752 -28572 -5732 -28508
rect -5836 -28588 -5732 -28572
rect -5836 -28652 -5816 -28588
rect -5752 -28652 -5732 -28588
rect -5836 -28668 -5732 -28652
rect -5836 -28732 -5816 -28668
rect -5752 -28732 -5732 -28668
rect -5836 -28748 -5732 -28732
rect -5836 -28812 -5816 -28748
rect -5752 -28812 -5732 -28748
rect -5836 -28828 -5732 -28812
rect -5836 -28892 -5816 -28828
rect -5752 -28892 -5732 -28828
rect -5836 -28908 -5732 -28892
rect -5836 -28972 -5816 -28908
rect -5752 -28972 -5732 -28908
rect -5836 -28988 -5732 -28972
rect -5836 -29052 -5816 -28988
rect -5752 -29052 -5732 -28988
rect -5836 -29068 -5732 -29052
rect -5836 -29132 -5816 -29068
rect -5752 -29132 -5732 -29068
rect -5836 -29148 -5732 -29132
rect -5836 -29212 -5816 -29148
rect -5752 -29212 -5732 -29148
rect -5836 -29228 -5732 -29212
rect -5836 -29292 -5816 -29228
rect -5752 -29292 -5732 -29228
rect -5836 -29308 -5732 -29292
rect -5836 -29372 -5816 -29308
rect -5752 -29372 -5732 -29308
rect -5836 -29388 -5732 -29372
rect -5836 -29452 -5816 -29388
rect -5752 -29452 -5732 -29388
rect -5836 -29468 -5732 -29452
rect -5836 -29532 -5816 -29468
rect -5752 -29532 -5732 -29468
rect -5836 -29548 -5732 -29532
rect -5836 -29612 -5816 -29548
rect -5752 -29612 -5732 -29548
rect -5836 -29628 -5732 -29612
rect -5836 -29692 -5816 -29628
rect -5752 -29692 -5732 -29628
rect -5836 -29708 -5732 -29692
rect -5836 -29772 -5816 -29708
rect -5752 -29772 -5732 -29708
rect -5836 -29788 -5732 -29772
rect -5836 -29852 -5816 -29788
rect -5752 -29852 -5732 -29788
rect -5836 -29868 -5732 -29852
rect -5836 -29932 -5816 -29868
rect -5752 -29932 -5732 -29868
rect -5836 -29948 -5732 -29932
rect -5836 -30012 -5816 -29948
rect -5752 -30012 -5732 -29948
rect -5836 -30028 -5732 -30012
rect -5836 -30092 -5816 -30028
rect -5752 -30092 -5732 -30028
rect -5836 -30108 -5732 -30092
rect -5836 -30172 -5816 -30108
rect -5752 -30172 -5732 -30108
rect -5836 -30188 -5732 -30172
rect -5836 -30252 -5816 -30188
rect -5752 -30252 -5732 -30188
rect -5836 -30268 -5732 -30252
rect -5836 -30332 -5816 -30268
rect -5752 -30332 -5732 -30268
rect -5836 -30348 -5732 -30332
rect -5836 -30412 -5816 -30348
rect -5752 -30412 -5732 -30348
rect -5836 -30428 -5732 -30412
rect -5836 -30492 -5816 -30428
rect -5752 -30492 -5732 -30428
rect -5836 -30508 -5732 -30492
rect -5836 -30572 -5816 -30508
rect -5752 -30572 -5732 -30508
rect -5836 -30588 -5732 -30572
rect -5836 -30652 -5816 -30588
rect -5752 -30652 -5732 -30588
rect -5836 -30668 -5732 -30652
rect -5836 -30732 -5816 -30668
rect -5752 -30732 -5732 -30668
rect -5836 -30748 -5732 -30732
rect -5836 -30812 -5816 -30748
rect -5752 -30812 -5732 -30748
rect -5836 -30828 -5732 -30812
rect -5836 -30892 -5816 -30828
rect -5752 -30892 -5732 -30828
rect -5836 -30908 -5732 -30892
rect -5836 -30972 -5816 -30908
rect -5752 -30972 -5732 -30908
rect -5836 -30988 -5732 -30972
rect -5836 -31052 -5816 -30988
rect -5752 -31052 -5732 -30988
rect -5836 -31068 -5732 -31052
rect -5836 -31132 -5816 -31068
rect -5752 -31132 -5732 -31068
rect -5836 -31148 -5732 -31132
rect -5836 -31212 -5816 -31148
rect -5752 -31212 -5732 -31148
rect -5836 -31228 -5732 -31212
rect -5836 -31292 -5816 -31228
rect -5752 -31292 -5732 -31228
rect -5836 -31308 -5732 -31292
rect -5836 -31372 -5816 -31308
rect -5752 -31372 -5732 -31308
rect -5836 -31388 -5732 -31372
rect -5836 -31452 -5816 -31388
rect -5752 -31452 -5732 -31388
rect -5836 -31468 -5732 -31452
rect -5836 -31532 -5816 -31468
rect -5752 -31532 -5732 -31468
rect -5836 -31548 -5732 -31532
rect -5836 -31612 -5816 -31548
rect -5752 -31612 -5732 -31548
rect -5836 -31628 -5732 -31612
rect -5836 -31692 -5816 -31628
rect -5752 -31692 -5732 -31628
rect -5836 -31708 -5732 -31692
rect -11448 -32068 -11344 -31772
rect -17060 -32148 -16956 -32132
rect -17060 -32212 -17040 -32148
rect -16976 -32212 -16956 -32148
rect -17060 -32228 -16956 -32212
rect -17060 -32292 -17040 -32228
rect -16976 -32292 -16956 -32228
rect -17060 -32308 -16956 -32292
rect -17060 -32372 -17040 -32308
rect -16976 -32372 -16956 -32308
rect -17060 -32388 -16956 -32372
rect -17060 -32452 -17040 -32388
rect -16976 -32452 -16956 -32388
rect -17060 -32468 -16956 -32452
rect -17060 -32532 -17040 -32468
rect -16976 -32532 -16956 -32468
rect -17060 -32548 -16956 -32532
rect -17060 -32612 -17040 -32548
rect -16976 -32612 -16956 -32548
rect -17060 -32628 -16956 -32612
rect -17060 -32692 -17040 -32628
rect -16976 -32692 -16956 -32628
rect -17060 -32708 -16956 -32692
rect -17060 -32772 -17040 -32708
rect -16976 -32772 -16956 -32708
rect -17060 -32788 -16956 -32772
rect -17060 -32852 -17040 -32788
rect -16976 -32852 -16956 -32788
rect -17060 -32868 -16956 -32852
rect -17060 -32932 -17040 -32868
rect -16976 -32932 -16956 -32868
rect -17060 -32948 -16956 -32932
rect -17060 -33012 -17040 -32948
rect -16976 -33012 -16956 -32948
rect -17060 -33028 -16956 -33012
rect -17060 -33092 -17040 -33028
rect -16976 -33092 -16956 -33028
rect -17060 -33108 -16956 -33092
rect -17060 -33172 -17040 -33108
rect -16976 -33172 -16956 -33108
rect -17060 -33188 -16956 -33172
rect -17060 -33252 -17040 -33188
rect -16976 -33252 -16956 -33188
rect -17060 -33268 -16956 -33252
rect -17060 -33332 -17040 -33268
rect -16976 -33332 -16956 -33268
rect -17060 -33348 -16956 -33332
rect -17060 -33412 -17040 -33348
rect -16976 -33412 -16956 -33348
rect -17060 -33428 -16956 -33412
rect -17060 -33492 -17040 -33428
rect -16976 -33492 -16956 -33428
rect -17060 -33508 -16956 -33492
rect -17060 -33572 -17040 -33508
rect -16976 -33572 -16956 -33508
rect -17060 -33588 -16956 -33572
rect -17060 -33652 -17040 -33588
rect -16976 -33652 -16956 -33588
rect -17060 -33668 -16956 -33652
rect -17060 -33732 -17040 -33668
rect -16976 -33732 -16956 -33668
rect -17060 -33748 -16956 -33732
rect -17060 -33812 -17040 -33748
rect -16976 -33812 -16956 -33748
rect -17060 -33828 -16956 -33812
rect -17060 -33892 -17040 -33828
rect -16976 -33892 -16956 -33828
rect -17060 -33908 -16956 -33892
rect -17060 -33972 -17040 -33908
rect -16976 -33972 -16956 -33908
rect -17060 -33988 -16956 -33972
rect -17060 -34052 -17040 -33988
rect -16976 -34052 -16956 -33988
rect -17060 -34068 -16956 -34052
rect -17060 -34132 -17040 -34068
rect -16976 -34132 -16956 -34068
rect -17060 -34148 -16956 -34132
rect -17060 -34212 -17040 -34148
rect -16976 -34212 -16956 -34148
rect -17060 -34228 -16956 -34212
rect -17060 -34292 -17040 -34228
rect -16976 -34292 -16956 -34228
rect -17060 -34308 -16956 -34292
rect -17060 -34372 -17040 -34308
rect -16976 -34372 -16956 -34308
rect -17060 -34388 -16956 -34372
rect -17060 -34452 -17040 -34388
rect -16976 -34452 -16956 -34388
rect -17060 -34468 -16956 -34452
rect -17060 -34532 -17040 -34468
rect -16976 -34532 -16956 -34468
rect -17060 -34548 -16956 -34532
rect -17060 -34612 -17040 -34548
rect -16976 -34612 -16956 -34548
rect -17060 -34628 -16956 -34612
rect -17060 -34692 -17040 -34628
rect -16976 -34692 -16956 -34628
rect -17060 -34708 -16956 -34692
rect -17060 -34772 -17040 -34708
rect -16976 -34772 -16956 -34708
rect -17060 -34788 -16956 -34772
rect -17060 -34852 -17040 -34788
rect -16976 -34852 -16956 -34788
rect -17060 -34868 -16956 -34852
rect -17060 -34932 -17040 -34868
rect -16976 -34932 -16956 -34868
rect -17060 -34948 -16956 -34932
rect -17060 -35012 -17040 -34948
rect -16976 -35012 -16956 -34948
rect -17060 -35028 -16956 -35012
rect -17060 -35092 -17040 -35028
rect -16976 -35092 -16956 -35028
rect -17060 -35108 -16956 -35092
rect -17060 -35172 -17040 -35108
rect -16976 -35172 -16956 -35108
rect -17060 -35188 -16956 -35172
rect -17060 -35252 -17040 -35188
rect -16976 -35252 -16956 -35188
rect -17060 -35268 -16956 -35252
rect -17060 -35332 -17040 -35268
rect -16976 -35332 -16956 -35268
rect -17060 -35348 -16956 -35332
rect -17060 -35412 -17040 -35348
rect -16976 -35412 -16956 -35348
rect -17060 -35428 -16956 -35412
rect -17060 -35492 -17040 -35428
rect -16976 -35492 -16956 -35428
rect -17060 -35508 -16956 -35492
rect -17060 -35572 -17040 -35508
rect -16976 -35572 -16956 -35508
rect -17060 -35588 -16956 -35572
rect -17060 -35652 -17040 -35588
rect -16976 -35652 -16956 -35588
rect -17060 -35668 -16956 -35652
rect -17060 -35732 -17040 -35668
rect -16976 -35732 -16956 -35668
rect -17060 -35748 -16956 -35732
rect -17060 -35812 -17040 -35748
rect -16976 -35812 -16956 -35748
rect -17060 -35828 -16956 -35812
rect -17060 -35892 -17040 -35828
rect -16976 -35892 -16956 -35828
rect -17060 -35908 -16956 -35892
rect -17060 -35972 -17040 -35908
rect -16976 -35972 -16956 -35908
rect -17060 -35988 -16956 -35972
rect -17060 -36052 -17040 -35988
rect -16976 -36052 -16956 -35988
rect -17060 -36068 -16956 -36052
rect -17060 -36132 -17040 -36068
rect -16976 -36132 -16956 -36068
rect -17060 -36148 -16956 -36132
rect -17060 -36212 -17040 -36148
rect -16976 -36212 -16956 -36148
rect -17060 -36228 -16956 -36212
rect -17060 -36292 -17040 -36228
rect -16976 -36292 -16956 -36228
rect -17060 -36308 -16956 -36292
rect -17060 -36372 -17040 -36308
rect -16976 -36372 -16956 -36308
rect -17060 -36388 -16956 -36372
rect -17060 -36452 -17040 -36388
rect -16976 -36452 -16956 -36388
rect -17060 -36468 -16956 -36452
rect -17060 -36532 -17040 -36468
rect -16976 -36532 -16956 -36468
rect -17060 -36548 -16956 -36532
rect -17060 -36612 -17040 -36548
rect -16976 -36612 -16956 -36548
rect -17060 -36628 -16956 -36612
rect -17060 -36692 -17040 -36628
rect -16976 -36692 -16956 -36628
rect -17060 -36708 -16956 -36692
rect -17060 -36772 -17040 -36708
rect -16976 -36772 -16956 -36708
rect -17060 -36788 -16956 -36772
rect -17060 -36852 -17040 -36788
rect -16976 -36852 -16956 -36788
rect -17060 -36868 -16956 -36852
rect -17060 -36932 -17040 -36868
rect -16976 -36932 -16956 -36868
rect -17060 -36948 -16956 -36932
rect -17060 -37012 -17040 -36948
rect -16976 -37012 -16956 -36948
rect -17060 -37028 -16956 -37012
rect -22672 -37240 -22568 -37092
rect -19840 -37240 -19736 -37041
rect -17060 -37092 -17040 -37028
rect -16976 -37092 -16956 -37028
rect -16637 -32148 -11715 -32119
rect -16637 -37012 -16608 -32148
rect -11744 -37012 -11715 -32148
rect -16637 -37041 -11715 -37012
rect -11448 -32132 -11428 -32068
rect -11364 -32132 -11344 -32068
rect -8616 -32119 -8512 -31721
rect -5836 -31772 -5816 -31708
rect -5752 -31772 -5732 -31708
rect -5413 -26828 -491 -26799
rect -5413 -31692 -5384 -26828
rect -520 -31692 -491 -26828
rect -5413 -31721 -491 -31692
rect -224 -26812 -204 -26748
rect -140 -26812 -120 -26748
rect 2608 -26799 2712 -26401
rect 5388 -26452 5408 -26388
rect 5472 -26452 5492 -26388
rect 5811 -21508 10733 -21479
rect 5811 -26372 5840 -21508
rect 10704 -26372 10733 -21508
rect 5811 -26401 10733 -26372
rect 11000 -21492 11020 -21428
rect 11084 -21492 11104 -21428
rect 13832 -21479 13936 -21081
rect 16612 -21132 16632 -21068
rect 16696 -21132 16716 -21068
rect 17035 -16188 21957 -16159
rect 17035 -21052 17064 -16188
rect 21928 -21052 21957 -16188
rect 17035 -21081 21957 -21052
rect 22224 -16172 22244 -16108
rect 22308 -16172 22328 -16108
rect 25056 -16159 25160 -15761
rect 27836 -15812 27856 -15748
rect 27920 -15812 27940 -15748
rect 28259 -10868 33181 -10839
rect 28259 -15732 28288 -10868
rect 33152 -15732 33181 -10868
rect 28259 -15761 33181 -15732
rect 33448 -10852 33468 -10788
rect 33532 -10852 33552 -10788
rect 36280 -10839 36384 -10441
rect 39060 -10492 39080 -10428
rect 39144 -10492 39164 -10428
rect 39060 -10788 39164 -10492
rect 33448 -10868 33552 -10852
rect 33448 -10932 33468 -10868
rect 33532 -10932 33552 -10868
rect 33448 -10948 33552 -10932
rect 33448 -11012 33468 -10948
rect 33532 -11012 33552 -10948
rect 33448 -11028 33552 -11012
rect 33448 -11092 33468 -11028
rect 33532 -11092 33552 -11028
rect 33448 -11108 33552 -11092
rect 33448 -11172 33468 -11108
rect 33532 -11172 33552 -11108
rect 33448 -11188 33552 -11172
rect 33448 -11252 33468 -11188
rect 33532 -11252 33552 -11188
rect 33448 -11268 33552 -11252
rect 33448 -11332 33468 -11268
rect 33532 -11332 33552 -11268
rect 33448 -11348 33552 -11332
rect 33448 -11412 33468 -11348
rect 33532 -11412 33552 -11348
rect 33448 -11428 33552 -11412
rect 33448 -11492 33468 -11428
rect 33532 -11492 33552 -11428
rect 33448 -11508 33552 -11492
rect 33448 -11572 33468 -11508
rect 33532 -11572 33552 -11508
rect 33448 -11588 33552 -11572
rect 33448 -11652 33468 -11588
rect 33532 -11652 33552 -11588
rect 33448 -11668 33552 -11652
rect 33448 -11732 33468 -11668
rect 33532 -11732 33552 -11668
rect 33448 -11748 33552 -11732
rect 33448 -11812 33468 -11748
rect 33532 -11812 33552 -11748
rect 33448 -11828 33552 -11812
rect 33448 -11892 33468 -11828
rect 33532 -11892 33552 -11828
rect 33448 -11908 33552 -11892
rect 33448 -11972 33468 -11908
rect 33532 -11972 33552 -11908
rect 33448 -11988 33552 -11972
rect 33448 -12052 33468 -11988
rect 33532 -12052 33552 -11988
rect 33448 -12068 33552 -12052
rect 33448 -12132 33468 -12068
rect 33532 -12132 33552 -12068
rect 33448 -12148 33552 -12132
rect 33448 -12212 33468 -12148
rect 33532 -12212 33552 -12148
rect 33448 -12228 33552 -12212
rect 33448 -12292 33468 -12228
rect 33532 -12292 33552 -12228
rect 33448 -12308 33552 -12292
rect 33448 -12372 33468 -12308
rect 33532 -12372 33552 -12308
rect 33448 -12388 33552 -12372
rect 33448 -12452 33468 -12388
rect 33532 -12452 33552 -12388
rect 33448 -12468 33552 -12452
rect 33448 -12532 33468 -12468
rect 33532 -12532 33552 -12468
rect 33448 -12548 33552 -12532
rect 33448 -12612 33468 -12548
rect 33532 -12612 33552 -12548
rect 33448 -12628 33552 -12612
rect 33448 -12692 33468 -12628
rect 33532 -12692 33552 -12628
rect 33448 -12708 33552 -12692
rect 33448 -12772 33468 -12708
rect 33532 -12772 33552 -12708
rect 33448 -12788 33552 -12772
rect 33448 -12852 33468 -12788
rect 33532 -12852 33552 -12788
rect 33448 -12868 33552 -12852
rect 33448 -12932 33468 -12868
rect 33532 -12932 33552 -12868
rect 33448 -12948 33552 -12932
rect 33448 -13012 33468 -12948
rect 33532 -13012 33552 -12948
rect 33448 -13028 33552 -13012
rect 33448 -13092 33468 -13028
rect 33532 -13092 33552 -13028
rect 33448 -13108 33552 -13092
rect 33448 -13172 33468 -13108
rect 33532 -13172 33552 -13108
rect 33448 -13188 33552 -13172
rect 33448 -13252 33468 -13188
rect 33532 -13252 33552 -13188
rect 33448 -13268 33552 -13252
rect 33448 -13332 33468 -13268
rect 33532 -13332 33552 -13268
rect 33448 -13348 33552 -13332
rect 33448 -13412 33468 -13348
rect 33532 -13412 33552 -13348
rect 33448 -13428 33552 -13412
rect 33448 -13492 33468 -13428
rect 33532 -13492 33552 -13428
rect 33448 -13508 33552 -13492
rect 33448 -13572 33468 -13508
rect 33532 -13572 33552 -13508
rect 33448 -13588 33552 -13572
rect 33448 -13652 33468 -13588
rect 33532 -13652 33552 -13588
rect 33448 -13668 33552 -13652
rect 33448 -13732 33468 -13668
rect 33532 -13732 33552 -13668
rect 33448 -13748 33552 -13732
rect 33448 -13812 33468 -13748
rect 33532 -13812 33552 -13748
rect 33448 -13828 33552 -13812
rect 33448 -13892 33468 -13828
rect 33532 -13892 33552 -13828
rect 33448 -13908 33552 -13892
rect 33448 -13972 33468 -13908
rect 33532 -13972 33552 -13908
rect 33448 -13988 33552 -13972
rect 33448 -14052 33468 -13988
rect 33532 -14052 33552 -13988
rect 33448 -14068 33552 -14052
rect 33448 -14132 33468 -14068
rect 33532 -14132 33552 -14068
rect 33448 -14148 33552 -14132
rect 33448 -14212 33468 -14148
rect 33532 -14212 33552 -14148
rect 33448 -14228 33552 -14212
rect 33448 -14292 33468 -14228
rect 33532 -14292 33552 -14228
rect 33448 -14308 33552 -14292
rect 33448 -14372 33468 -14308
rect 33532 -14372 33552 -14308
rect 33448 -14388 33552 -14372
rect 33448 -14452 33468 -14388
rect 33532 -14452 33552 -14388
rect 33448 -14468 33552 -14452
rect 33448 -14532 33468 -14468
rect 33532 -14532 33552 -14468
rect 33448 -14548 33552 -14532
rect 33448 -14612 33468 -14548
rect 33532 -14612 33552 -14548
rect 33448 -14628 33552 -14612
rect 33448 -14692 33468 -14628
rect 33532 -14692 33552 -14628
rect 33448 -14708 33552 -14692
rect 33448 -14772 33468 -14708
rect 33532 -14772 33552 -14708
rect 33448 -14788 33552 -14772
rect 33448 -14852 33468 -14788
rect 33532 -14852 33552 -14788
rect 33448 -14868 33552 -14852
rect 33448 -14932 33468 -14868
rect 33532 -14932 33552 -14868
rect 33448 -14948 33552 -14932
rect 33448 -15012 33468 -14948
rect 33532 -15012 33552 -14948
rect 33448 -15028 33552 -15012
rect 33448 -15092 33468 -15028
rect 33532 -15092 33552 -15028
rect 33448 -15108 33552 -15092
rect 33448 -15172 33468 -15108
rect 33532 -15172 33552 -15108
rect 33448 -15188 33552 -15172
rect 33448 -15252 33468 -15188
rect 33532 -15252 33552 -15188
rect 33448 -15268 33552 -15252
rect 33448 -15332 33468 -15268
rect 33532 -15332 33552 -15268
rect 33448 -15348 33552 -15332
rect 33448 -15412 33468 -15348
rect 33532 -15412 33552 -15348
rect 33448 -15428 33552 -15412
rect 33448 -15492 33468 -15428
rect 33532 -15492 33552 -15428
rect 33448 -15508 33552 -15492
rect 33448 -15572 33468 -15508
rect 33532 -15572 33552 -15508
rect 33448 -15588 33552 -15572
rect 33448 -15652 33468 -15588
rect 33532 -15652 33552 -15588
rect 33448 -15668 33552 -15652
rect 33448 -15732 33468 -15668
rect 33532 -15732 33552 -15668
rect 33448 -15748 33552 -15732
rect 27836 -16108 27940 -15812
rect 22224 -16188 22328 -16172
rect 22224 -16252 22244 -16188
rect 22308 -16252 22328 -16188
rect 22224 -16268 22328 -16252
rect 22224 -16332 22244 -16268
rect 22308 -16332 22328 -16268
rect 22224 -16348 22328 -16332
rect 22224 -16412 22244 -16348
rect 22308 -16412 22328 -16348
rect 22224 -16428 22328 -16412
rect 22224 -16492 22244 -16428
rect 22308 -16492 22328 -16428
rect 22224 -16508 22328 -16492
rect 22224 -16572 22244 -16508
rect 22308 -16572 22328 -16508
rect 22224 -16588 22328 -16572
rect 22224 -16652 22244 -16588
rect 22308 -16652 22328 -16588
rect 22224 -16668 22328 -16652
rect 22224 -16732 22244 -16668
rect 22308 -16732 22328 -16668
rect 22224 -16748 22328 -16732
rect 22224 -16812 22244 -16748
rect 22308 -16812 22328 -16748
rect 22224 -16828 22328 -16812
rect 22224 -16892 22244 -16828
rect 22308 -16892 22328 -16828
rect 22224 -16908 22328 -16892
rect 22224 -16972 22244 -16908
rect 22308 -16972 22328 -16908
rect 22224 -16988 22328 -16972
rect 22224 -17052 22244 -16988
rect 22308 -17052 22328 -16988
rect 22224 -17068 22328 -17052
rect 22224 -17132 22244 -17068
rect 22308 -17132 22328 -17068
rect 22224 -17148 22328 -17132
rect 22224 -17212 22244 -17148
rect 22308 -17212 22328 -17148
rect 22224 -17228 22328 -17212
rect 22224 -17292 22244 -17228
rect 22308 -17292 22328 -17228
rect 22224 -17308 22328 -17292
rect 22224 -17372 22244 -17308
rect 22308 -17372 22328 -17308
rect 22224 -17388 22328 -17372
rect 22224 -17452 22244 -17388
rect 22308 -17452 22328 -17388
rect 22224 -17468 22328 -17452
rect 22224 -17532 22244 -17468
rect 22308 -17532 22328 -17468
rect 22224 -17548 22328 -17532
rect 22224 -17612 22244 -17548
rect 22308 -17612 22328 -17548
rect 22224 -17628 22328 -17612
rect 22224 -17692 22244 -17628
rect 22308 -17692 22328 -17628
rect 22224 -17708 22328 -17692
rect 22224 -17772 22244 -17708
rect 22308 -17772 22328 -17708
rect 22224 -17788 22328 -17772
rect 22224 -17852 22244 -17788
rect 22308 -17852 22328 -17788
rect 22224 -17868 22328 -17852
rect 22224 -17932 22244 -17868
rect 22308 -17932 22328 -17868
rect 22224 -17948 22328 -17932
rect 22224 -18012 22244 -17948
rect 22308 -18012 22328 -17948
rect 22224 -18028 22328 -18012
rect 22224 -18092 22244 -18028
rect 22308 -18092 22328 -18028
rect 22224 -18108 22328 -18092
rect 22224 -18172 22244 -18108
rect 22308 -18172 22328 -18108
rect 22224 -18188 22328 -18172
rect 22224 -18252 22244 -18188
rect 22308 -18252 22328 -18188
rect 22224 -18268 22328 -18252
rect 22224 -18332 22244 -18268
rect 22308 -18332 22328 -18268
rect 22224 -18348 22328 -18332
rect 22224 -18412 22244 -18348
rect 22308 -18412 22328 -18348
rect 22224 -18428 22328 -18412
rect 22224 -18492 22244 -18428
rect 22308 -18492 22328 -18428
rect 22224 -18508 22328 -18492
rect 22224 -18572 22244 -18508
rect 22308 -18572 22328 -18508
rect 22224 -18588 22328 -18572
rect 22224 -18652 22244 -18588
rect 22308 -18652 22328 -18588
rect 22224 -18668 22328 -18652
rect 22224 -18732 22244 -18668
rect 22308 -18732 22328 -18668
rect 22224 -18748 22328 -18732
rect 22224 -18812 22244 -18748
rect 22308 -18812 22328 -18748
rect 22224 -18828 22328 -18812
rect 22224 -18892 22244 -18828
rect 22308 -18892 22328 -18828
rect 22224 -18908 22328 -18892
rect 22224 -18972 22244 -18908
rect 22308 -18972 22328 -18908
rect 22224 -18988 22328 -18972
rect 22224 -19052 22244 -18988
rect 22308 -19052 22328 -18988
rect 22224 -19068 22328 -19052
rect 22224 -19132 22244 -19068
rect 22308 -19132 22328 -19068
rect 22224 -19148 22328 -19132
rect 22224 -19212 22244 -19148
rect 22308 -19212 22328 -19148
rect 22224 -19228 22328 -19212
rect 22224 -19292 22244 -19228
rect 22308 -19292 22328 -19228
rect 22224 -19308 22328 -19292
rect 22224 -19372 22244 -19308
rect 22308 -19372 22328 -19308
rect 22224 -19388 22328 -19372
rect 22224 -19452 22244 -19388
rect 22308 -19452 22328 -19388
rect 22224 -19468 22328 -19452
rect 22224 -19532 22244 -19468
rect 22308 -19532 22328 -19468
rect 22224 -19548 22328 -19532
rect 22224 -19612 22244 -19548
rect 22308 -19612 22328 -19548
rect 22224 -19628 22328 -19612
rect 22224 -19692 22244 -19628
rect 22308 -19692 22328 -19628
rect 22224 -19708 22328 -19692
rect 22224 -19772 22244 -19708
rect 22308 -19772 22328 -19708
rect 22224 -19788 22328 -19772
rect 22224 -19852 22244 -19788
rect 22308 -19852 22328 -19788
rect 22224 -19868 22328 -19852
rect 22224 -19932 22244 -19868
rect 22308 -19932 22328 -19868
rect 22224 -19948 22328 -19932
rect 22224 -20012 22244 -19948
rect 22308 -20012 22328 -19948
rect 22224 -20028 22328 -20012
rect 22224 -20092 22244 -20028
rect 22308 -20092 22328 -20028
rect 22224 -20108 22328 -20092
rect 22224 -20172 22244 -20108
rect 22308 -20172 22328 -20108
rect 22224 -20188 22328 -20172
rect 22224 -20252 22244 -20188
rect 22308 -20252 22328 -20188
rect 22224 -20268 22328 -20252
rect 22224 -20332 22244 -20268
rect 22308 -20332 22328 -20268
rect 22224 -20348 22328 -20332
rect 22224 -20412 22244 -20348
rect 22308 -20412 22328 -20348
rect 22224 -20428 22328 -20412
rect 22224 -20492 22244 -20428
rect 22308 -20492 22328 -20428
rect 22224 -20508 22328 -20492
rect 22224 -20572 22244 -20508
rect 22308 -20572 22328 -20508
rect 22224 -20588 22328 -20572
rect 22224 -20652 22244 -20588
rect 22308 -20652 22328 -20588
rect 22224 -20668 22328 -20652
rect 22224 -20732 22244 -20668
rect 22308 -20732 22328 -20668
rect 22224 -20748 22328 -20732
rect 22224 -20812 22244 -20748
rect 22308 -20812 22328 -20748
rect 22224 -20828 22328 -20812
rect 22224 -20892 22244 -20828
rect 22308 -20892 22328 -20828
rect 22224 -20908 22328 -20892
rect 22224 -20972 22244 -20908
rect 22308 -20972 22328 -20908
rect 22224 -20988 22328 -20972
rect 22224 -21052 22244 -20988
rect 22308 -21052 22328 -20988
rect 22224 -21068 22328 -21052
rect 16612 -21428 16716 -21132
rect 11000 -21508 11104 -21492
rect 11000 -21572 11020 -21508
rect 11084 -21572 11104 -21508
rect 11000 -21588 11104 -21572
rect 11000 -21652 11020 -21588
rect 11084 -21652 11104 -21588
rect 11000 -21668 11104 -21652
rect 11000 -21732 11020 -21668
rect 11084 -21732 11104 -21668
rect 11000 -21748 11104 -21732
rect 11000 -21812 11020 -21748
rect 11084 -21812 11104 -21748
rect 11000 -21828 11104 -21812
rect 11000 -21892 11020 -21828
rect 11084 -21892 11104 -21828
rect 11000 -21908 11104 -21892
rect 11000 -21972 11020 -21908
rect 11084 -21972 11104 -21908
rect 11000 -21988 11104 -21972
rect 11000 -22052 11020 -21988
rect 11084 -22052 11104 -21988
rect 11000 -22068 11104 -22052
rect 11000 -22132 11020 -22068
rect 11084 -22132 11104 -22068
rect 11000 -22148 11104 -22132
rect 11000 -22212 11020 -22148
rect 11084 -22212 11104 -22148
rect 11000 -22228 11104 -22212
rect 11000 -22292 11020 -22228
rect 11084 -22292 11104 -22228
rect 11000 -22308 11104 -22292
rect 11000 -22372 11020 -22308
rect 11084 -22372 11104 -22308
rect 11000 -22388 11104 -22372
rect 11000 -22452 11020 -22388
rect 11084 -22452 11104 -22388
rect 11000 -22468 11104 -22452
rect 11000 -22532 11020 -22468
rect 11084 -22532 11104 -22468
rect 11000 -22548 11104 -22532
rect 11000 -22612 11020 -22548
rect 11084 -22612 11104 -22548
rect 11000 -22628 11104 -22612
rect 11000 -22692 11020 -22628
rect 11084 -22692 11104 -22628
rect 11000 -22708 11104 -22692
rect 11000 -22772 11020 -22708
rect 11084 -22772 11104 -22708
rect 11000 -22788 11104 -22772
rect 11000 -22852 11020 -22788
rect 11084 -22852 11104 -22788
rect 11000 -22868 11104 -22852
rect 11000 -22932 11020 -22868
rect 11084 -22932 11104 -22868
rect 11000 -22948 11104 -22932
rect 11000 -23012 11020 -22948
rect 11084 -23012 11104 -22948
rect 11000 -23028 11104 -23012
rect 11000 -23092 11020 -23028
rect 11084 -23092 11104 -23028
rect 11000 -23108 11104 -23092
rect 11000 -23172 11020 -23108
rect 11084 -23172 11104 -23108
rect 11000 -23188 11104 -23172
rect 11000 -23252 11020 -23188
rect 11084 -23252 11104 -23188
rect 11000 -23268 11104 -23252
rect 11000 -23332 11020 -23268
rect 11084 -23332 11104 -23268
rect 11000 -23348 11104 -23332
rect 11000 -23412 11020 -23348
rect 11084 -23412 11104 -23348
rect 11000 -23428 11104 -23412
rect 11000 -23492 11020 -23428
rect 11084 -23492 11104 -23428
rect 11000 -23508 11104 -23492
rect 11000 -23572 11020 -23508
rect 11084 -23572 11104 -23508
rect 11000 -23588 11104 -23572
rect 11000 -23652 11020 -23588
rect 11084 -23652 11104 -23588
rect 11000 -23668 11104 -23652
rect 11000 -23732 11020 -23668
rect 11084 -23732 11104 -23668
rect 11000 -23748 11104 -23732
rect 11000 -23812 11020 -23748
rect 11084 -23812 11104 -23748
rect 11000 -23828 11104 -23812
rect 11000 -23892 11020 -23828
rect 11084 -23892 11104 -23828
rect 11000 -23908 11104 -23892
rect 11000 -23972 11020 -23908
rect 11084 -23972 11104 -23908
rect 11000 -23988 11104 -23972
rect 11000 -24052 11020 -23988
rect 11084 -24052 11104 -23988
rect 11000 -24068 11104 -24052
rect 11000 -24132 11020 -24068
rect 11084 -24132 11104 -24068
rect 11000 -24148 11104 -24132
rect 11000 -24212 11020 -24148
rect 11084 -24212 11104 -24148
rect 11000 -24228 11104 -24212
rect 11000 -24292 11020 -24228
rect 11084 -24292 11104 -24228
rect 11000 -24308 11104 -24292
rect 11000 -24372 11020 -24308
rect 11084 -24372 11104 -24308
rect 11000 -24388 11104 -24372
rect 11000 -24452 11020 -24388
rect 11084 -24452 11104 -24388
rect 11000 -24468 11104 -24452
rect 11000 -24532 11020 -24468
rect 11084 -24532 11104 -24468
rect 11000 -24548 11104 -24532
rect 11000 -24612 11020 -24548
rect 11084 -24612 11104 -24548
rect 11000 -24628 11104 -24612
rect 11000 -24692 11020 -24628
rect 11084 -24692 11104 -24628
rect 11000 -24708 11104 -24692
rect 11000 -24772 11020 -24708
rect 11084 -24772 11104 -24708
rect 11000 -24788 11104 -24772
rect 11000 -24852 11020 -24788
rect 11084 -24852 11104 -24788
rect 11000 -24868 11104 -24852
rect 11000 -24932 11020 -24868
rect 11084 -24932 11104 -24868
rect 11000 -24948 11104 -24932
rect 11000 -25012 11020 -24948
rect 11084 -25012 11104 -24948
rect 11000 -25028 11104 -25012
rect 11000 -25092 11020 -25028
rect 11084 -25092 11104 -25028
rect 11000 -25108 11104 -25092
rect 11000 -25172 11020 -25108
rect 11084 -25172 11104 -25108
rect 11000 -25188 11104 -25172
rect 11000 -25252 11020 -25188
rect 11084 -25252 11104 -25188
rect 11000 -25268 11104 -25252
rect 11000 -25332 11020 -25268
rect 11084 -25332 11104 -25268
rect 11000 -25348 11104 -25332
rect 11000 -25412 11020 -25348
rect 11084 -25412 11104 -25348
rect 11000 -25428 11104 -25412
rect 11000 -25492 11020 -25428
rect 11084 -25492 11104 -25428
rect 11000 -25508 11104 -25492
rect 11000 -25572 11020 -25508
rect 11084 -25572 11104 -25508
rect 11000 -25588 11104 -25572
rect 11000 -25652 11020 -25588
rect 11084 -25652 11104 -25588
rect 11000 -25668 11104 -25652
rect 11000 -25732 11020 -25668
rect 11084 -25732 11104 -25668
rect 11000 -25748 11104 -25732
rect 11000 -25812 11020 -25748
rect 11084 -25812 11104 -25748
rect 11000 -25828 11104 -25812
rect 11000 -25892 11020 -25828
rect 11084 -25892 11104 -25828
rect 11000 -25908 11104 -25892
rect 11000 -25972 11020 -25908
rect 11084 -25972 11104 -25908
rect 11000 -25988 11104 -25972
rect 11000 -26052 11020 -25988
rect 11084 -26052 11104 -25988
rect 11000 -26068 11104 -26052
rect 11000 -26132 11020 -26068
rect 11084 -26132 11104 -26068
rect 11000 -26148 11104 -26132
rect 11000 -26212 11020 -26148
rect 11084 -26212 11104 -26148
rect 11000 -26228 11104 -26212
rect 11000 -26292 11020 -26228
rect 11084 -26292 11104 -26228
rect 11000 -26308 11104 -26292
rect 11000 -26372 11020 -26308
rect 11084 -26372 11104 -26308
rect 11000 -26388 11104 -26372
rect 5388 -26748 5492 -26452
rect -224 -26828 -120 -26812
rect -224 -26892 -204 -26828
rect -140 -26892 -120 -26828
rect -224 -26908 -120 -26892
rect -224 -26972 -204 -26908
rect -140 -26972 -120 -26908
rect -224 -26988 -120 -26972
rect -224 -27052 -204 -26988
rect -140 -27052 -120 -26988
rect -224 -27068 -120 -27052
rect -224 -27132 -204 -27068
rect -140 -27132 -120 -27068
rect -224 -27148 -120 -27132
rect -224 -27212 -204 -27148
rect -140 -27212 -120 -27148
rect -224 -27228 -120 -27212
rect -224 -27292 -204 -27228
rect -140 -27292 -120 -27228
rect -224 -27308 -120 -27292
rect -224 -27372 -204 -27308
rect -140 -27372 -120 -27308
rect -224 -27388 -120 -27372
rect -224 -27452 -204 -27388
rect -140 -27452 -120 -27388
rect -224 -27468 -120 -27452
rect -224 -27532 -204 -27468
rect -140 -27532 -120 -27468
rect -224 -27548 -120 -27532
rect -224 -27612 -204 -27548
rect -140 -27612 -120 -27548
rect -224 -27628 -120 -27612
rect -224 -27692 -204 -27628
rect -140 -27692 -120 -27628
rect -224 -27708 -120 -27692
rect -224 -27772 -204 -27708
rect -140 -27772 -120 -27708
rect -224 -27788 -120 -27772
rect -224 -27852 -204 -27788
rect -140 -27852 -120 -27788
rect -224 -27868 -120 -27852
rect -224 -27932 -204 -27868
rect -140 -27932 -120 -27868
rect -224 -27948 -120 -27932
rect -224 -28012 -204 -27948
rect -140 -28012 -120 -27948
rect -224 -28028 -120 -28012
rect -224 -28092 -204 -28028
rect -140 -28092 -120 -28028
rect -224 -28108 -120 -28092
rect -224 -28172 -204 -28108
rect -140 -28172 -120 -28108
rect -224 -28188 -120 -28172
rect -224 -28252 -204 -28188
rect -140 -28252 -120 -28188
rect -224 -28268 -120 -28252
rect -224 -28332 -204 -28268
rect -140 -28332 -120 -28268
rect -224 -28348 -120 -28332
rect -224 -28412 -204 -28348
rect -140 -28412 -120 -28348
rect -224 -28428 -120 -28412
rect -224 -28492 -204 -28428
rect -140 -28492 -120 -28428
rect -224 -28508 -120 -28492
rect -224 -28572 -204 -28508
rect -140 -28572 -120 -28508
rect -224 -28588 -120 -28572
rect -224 -28652 -204 -28588
rect -140 -28652 -120 -28588
rect -224 -28668 -120 -28652
rect -224 -28732 -204 -28668
rect -140 -28732 -120 -28668
rect -224 -28748 -120 -28732
rect -224 -28812 -204 -28748
rect -140 -28812 -120 -28748
rect -224 -28828 -120 -28812
rect -224 -28892 -204 -28828
rect -140 -28892 -120 -28828
rect -224 -28908 -120 -28892
rect -224 -28972 -204 -28908
rect -140 -28972 -120 -28908
rect -224 -28988 -120 -28972
rect -224 -29052 -204 -28988
rect -140 -29052 -120 -28988
rect -224 -29068 -120 -29052
rect -224 -29132 -204 -29068
rect -140 -29132 -120 -29068
rect -224 -29148 -120 -29132
rect -224 -29212 -204 -29148
rect -140 -29212 -120 -29148
rect -224 -29228 -120 -29212
rect -224 -29292 -204 -29228
rect -140 -29292 -120 -29228
rect -224 -29308 -120 -29292
rect -224 -29372 -204 -29308
rect -140 -29372 -120 -29308
rect -224 -29388 -120 -29372
rect -224 -29452 -204 -29388
rect -140 -29452 -120 -29388
rect -224 -29468 -120 -29452
rect -224 -29532 -204 -29468
rect -140 -29532 -120 -29468
rect -224 -29548 -120 -29532
rect -224 -29612 -204 -29548
rect -140 -29612 -120 -29548
rect -224 -29628 -120 -29612
rect -224 -29692 -204 -29628
rect -140 -29692 -120 -29628
rect -224 -29708 -120 -29692
rect -224 -29772 -204 -29708
rect -140 -29772 -120 -29708
rect -224 -29788 -120 -29772
rect -224 -29852 -204 -29788
rect -140 -29852 -120 -29788
rect -224 -29868 -120 -29852
rect -224 -29932 -204 -29868
rect -140 -29932 -120 -29868
rect -224 -29948 -120 -29932
rect -224 -30012 -204 -29948
rect -140 -30012 -120 -29948
rect -224 -30028 -120 -30012
rect -224 -30092 -204 -30028
rect -140 -30092 -120 -30028
rect -224 -30108 -120 -30092
rect -224 -30172 -204 -30108
rect -140 -30172 -120 -30108
rect -224 -30188 -120 -30172
rect -224 -30252 -204 -30188
rect -140 -30252 -120 -30188
rect -224 -30268 -120 -30252
rect -224 -30332 -204 -30268
rect -140 -30332 -120 -30268
rect -224 -30348 -120 -30332
rect -224 -30412 -204 -30348
rect -140 -30412 -120 -30348
rect -224 -30428 -120 -30412
rect -224 -30492 -204 -30428
rect -140 -30492 -120 -30428
rect -224 -30508 -120 -30492
rect -224 -30572 -204 -30508
rect -140 -30572 -120 -30508
rect -224 -30588 -120 -30572
rect -224 -30652 -204 -30588
rect -140 -30652 -120 -30588
rect -224 -30668 -120 -30652
rect -224 -30732 -204 -30668
rect -140 -30732 -120 -30668
rect -224 -30748 -120 -30732
rect -224 -30812 -204 -30748
rect -140 -30812 -120 -30748
rect -224 -30828 -120 -30812
rect -224 -30892 -204 -30828
rect -140 -30892 -120 -30828
rect -224 -30908 -120 -30892
rect -224 -30972 -204 -30908
rect -140 -30972 -120 -30908
rect -224 -30988 -120 -30972
rect -224 -31052 -204 -30988
rect -140 -31052 -120 -30988
rect -224 -31068 -120 -31052
rect -224 -31132 -204 -31068
rect -140 -31132 -120 -31068
rect -224 -31148 -120 -31132
rect -224 -31212 -204 -31148
rect -140 -31212 -120 -31148
rect -224 -31228 -120 -31212
rect -224 -31292 -204 -31228
rect -140 -31292 -120 -31228
rect -224 -31308 -120 -31292
rect -224 -31372 -204 -31308
rect -140 -31372 -120 -31308
rect -224 -31388 -120 -31372
rect -224 -31452 -204 -31388
rect -140 -31452 -120 -31388
rect -224 -31468 -120 -31452
rect -224 -31532 -204 -31468
rect -140 -31532 -120 -31468
rect -224 -31548 -120 -31532
rect -224 -31612 -204 -31548
rect -140 -31612 -120 -31548
rect -224 -31628 -120 -31612
rect -224 -31692 -204 -31628
rect -140 -31692 -120 -31628
rect -224 -31708 -120 -31692
rect -5836 -32068 -5732 -31772
rect -11448 -32148 -11344 -32132
rect -11448 -32212 -11428 -32148
rect -11364 -32212 -11344 -32148
rect -11448 -32228 -11344 -32212
rect -11448 -32292 -11428 -32228
rect -11364 -32292 -11344 -32228
rect -11448 -32308 -11344 -32292
rect -11448 -32372 -11428 -32308
rect -11364 -32372 -11344 -32308
rect -11448 -32388 -11344 -32372
rect -11448 -32452 -11428 -32388
rect -11364 -32452 -11344 -32388
rect -11448 -32468 -11344 -32452
rect -11448 -32532 -11428 -32468
rect -11364 -32532 -11344 -32468
rect -11448 -32548 -11344 -32532
rect -11448 -32612 -11428 -32548
rect -11364 -32612 -11344 -32548
rect -11448 -32628 -11344 -32612
rect -11448 -32692 -11428 -32628
rect -11364 -32692 -11344 -32628
rect -11448 -32708 -11344 -32692
rect -11448 -32772 -11428 -32708
rect -11364 -32772 -11344 -32708
rect -11448 -32788 -11344 -32772
rect -11448 -32852 -11428 -32788
rect -11364 -32852 -11344 -32788
rect -11448 -32868 -11344 -32852
rect -11448 -32932 -11428 -32868
rect -11364 -32932 -11344 -32868
rect -11448 -32948 -11344 -32932
rect -11448 -33012 -11428 -32948
rect -11364 -33012 -11344 -32948
rect -11448 -33028 -11344 -33012
rect -11448 -33092 -11428 -33028
rect -11364 -33092 -11344 -33028
rect -11448 -33108 -11344 -33092
rect -11448 -33172 -11428 -33108
rect -11364 -33172 -11344 -33108
rect -11448 -33188 -11344 -33172
rect -11448 -33252 -11428 -33188
rect -11364 -33252 -11344 -33188
rect -11448 -33268 -11344 -33252
rect -11448 -33332 -11428 -33268
rect -11364 -33332 -11344 -33268
rect -11448 -33348 -11344 -33332
rect -11448 -33412 -11428 -33348
rect -11364 -33412 -11344 -33348
rect -11448 -33428 -11344 -33412
rect -11448 -33492 -11428 -33428
rect -11364 -33492 -11344 -33428
rect -11448 -33508 -11344 -33492
rect -11448 -33572 -11428 -33508
rect -11364 -33572 -11344 -33508
rect -11448 -33588 -11344 -33572
rect -11448 -33652 -11428 -33588
rect -11364 -33652 -11344 -33588
rect -11448 -33668 -11344 -33652
rect -11448 -33732 -11428 -33668
rect -11364 -33732 -11344 -33668
rect -11448 -33748 -11344 -33732
rect -11448 -33812 -11428 -33748
rect -11364 -33812 -11344 -33748
rect -11448 -33828 -11344 -33812
rect -11448 -33892 -11428 -33828
rect -11364 -33892 -11344 -33828
rect -11448 -33908 -11344 -33892
rect -11448 -33972 -11428 -33908
rect -11364 -33972 -11344 -33908
rect -11448 -33988 -11344 -33972
rect -11448 -34052 -11428 -33988
rect -11364 -34052 -11344 -33988
rect -11448 -34068 -11344 -34052
rect -11448 -34132 -11428 -34068
rect -11364 -34132 -11344 -34068
rect -11448 -34148 -11344 -34132
rect -11448 -34212 -11428 -34148
rect -11364 -34212 -11344 -34148
rect -11448 -34228 -11344 -34212
rect -11448 -34292 -11428 -34228
rect -11364 -34292 -11344 -34228
rect -11448 -34308 -11344 -34292
rect -11448 -34372 -11428 -34308
rect -11364 -34372 -11344 -34308
rect -11448 -34388 -11344 -34372
rect -11448 -34452 -11428 -34388
rect -11364 -34452 -11344 -34388
rect -11448 -34468 -11344 -34452
rect -11448 -34532 -11428 -34468
rect -11364 -34532 -11344 -34468
rect -11448 -34548 -11344 -34532
rect -11448 -34612 -11428 -34548
rect -11364 -34612 -11344 -34548
rect -11448 -34628 -11344 -34612
rect -11448 -34692 -11428 -34628
rect -11364 -34692 -11344 -34628
rect -11448 -34708 -11344 -34692
rect -11448 -34772 -11428 -34708
rect -11364 -34772 -11344 -34708
rect -11448 -34788 -11344 -34772
rect -11448 -34852 -11428 -34788
rect -11364 -34852 -11344 -34788
rect -11448 -34868 -11344 -34852
rect -11448 -34932 -11428 -34868
rect -11364 -34932 -11344 -34868
rect -11448 -34948 -11344 -34932
rect -11448 -35012 -11428 -34948
rect -11364 -35012 -11344 -34948
rect -11448 -35028 -11344 -35012
rect -11448 -35092 -11428 -35028
rect -11364 -35092 -11344 -35028
rect -11448 -35108 -11344 -35092
rect -11448 -35172 -11428 -35108
rect -11364 -35172 -11344 -35108
rect -11448 -35188 -11344 -35172
rect -11448 -35252 -11428 -35188
rect -11364 -35252 -11344 -35188
rect -11448 -35268 -11344 -35252
rect -11448 -35332 -11428 -35268
rect -11364 -35332 -11344 -35268
rect -11448 -35348 -11344 -35332
rect -11448 -35412 -11428 -35348
rect -11364 -35412 -11344 -35348
rect -11448 -35428 -11344 -35412
rect -11448 -35492 -11428 -35428
rect -11364 -35492 -11344 -35428
rect -11448 -35508 -11344 -35492
rect -11448 -35572 -11428 -35508
rect -11364 -35572 -11344 -35508
rect -11448 -35588 -11344 -35572
rect -11448 -35652 -11428 -35588
rect -11364 -35652 -11344 -35588
rect -11448 -35668 -11344 -35652
rect -11448 -35732 -11428 -35668
rect -11364 -35732 -11344 -35668
rect -11448 -35748 -11344 -35732
rect -11448 -35812 -11428 -35748
rect -11364 -35812 -11344 -35748
rect -11448 -35828 -11344 -35812
rect -11448 -35892 -11428 -35828
rect -11364 -35892 -11344 -35828
rect -11448 -35908 -11344 -35892
rect -11448 -35972 -11428 -35908
rect -11364 -35972 -11344 -35908
rect -11448 -35988 -11344 -35972
rect -11448 -36052 -11428 -35988
rect -11364 -36052 -11344 -35988
rect -11448 -36068 -11344 -36052
rect -11448 -36132 -11428 -36068
rect -11364 -36132 -11344 -36068
rect -11448 -36148 -11344 -36132
rect -11448 -36212 -11428 -36148
rect -11364 -36212 -11344 -36148
rect -11448 -36228 -11344 -36212
rect -11448 -36292 -11428 -36228
rect -11364 -36292 -11344 -36228
rect -11448 -36308 -11344 -36292
rect -11448 -36372 -11428 -36308
rect -11364 -36372 -11344 -36308
rect -11448 -36388 -11344 -36372
rect -11448 -36452 -11428 -36388
rect -11364 -36452 -11344 -36388
rect -11448 -36468 -11344 -36452
rect -11448 -36532 -11428 -36468
rect -11364 -36532 -11344 -36468
rect -11448 -36548 -11344 -36532
rect -11448 -36612 -11428 -36548
rect -11364 -36612 -11344 -36548
rect -11448 -36628 -11344 -36612
rect -11448 -36692 -11428 -36628
rect -11364 -36692 -11344 -36628
rect -11448 -36708 -11344 -36692
rect -11448 -36772 -11428 -36708
rect -11364 -36772 -11344 -36708
rect -11448 -36788 -11344 -36772
rect -11448 -36852 -11428 -36788
rect -11364 -36852 -11344 -36788
rect -11448 -36868 -11344 -36852
rect -11448 -36932 -11428 -36868
rect -11364 -36932 -11344 -36868
rect -11448 -36948 -11344 -36932
rect -11448 -37012 -11428 -36948
rect -11364 -37012 -11344 -36948
rect -11448 -37028 -11344 -37012
rect -17060 -37240 -16956 -37092
rect -14228 -37240 -14124 -37041
rect -11448 -37092 -11428 -37028
rect -11364 -37092 -11344 -37028
rect -11025 -32148 -6103 -32119
rect -11025 -37012 -10996 -32148
rect -6132 -37012 -6103 -32148
rect -11025 -37041 -6103 -37012
rect -5836 -32132 -5816 -32068
rect -5752 -32132 -5732 -32068
rect -3004 -32119 -2900 -31721
rect -224 -31772 -204 -31708
rect -140 -31772 -120 -31708
rect 199 -26828 5121 -26799
rect 199 -31692 228 -26828
rect 5092 -31692 5121 -26828
rect 199 -31721 5121 -31692
rect 5388 -26812 5408 -26748
rect 5472 -26812 5492 -26748
rect 8220 -26799 8324 -26401
rect 11000 -26452 11020 -26388
rect 11084 -26452 11104 -26388
rect 11423 -21508 16345 -21479
rect 11423 -26372 11452 -21508
rect 16316 -26372 16345 -21508
rect 11423 -26401 16345 -26372
rect 16612 -21492 16632 -21428
rect 16696 -21492 16716 -21428
rect 19444 -21479 19548 -21081
rect 22224 -21132 22244 -21068
rect 22308 -21132 22328 -21068
rect 22647 -16188 27569 -16159
rect 22647 -21052 22676 -16188
rect 27540 -21052 27569 -16188
rect 22647 -21081 27569 -21052
rect 27836 -16172 27856 -16108
rect 27920 -16172 27940 -16108
rect 30668 -16159 30772 -15761
rect 33448 -15812 33468 -15748
rect 33532 -15812 33552 -15748
rect 33871 -10868 38793 -10839
rect 33871 -15732 33900 -10868
rect 38764 -15732 38793 -10868
rect 33871 -15761 38793 -15732
rect 39060 -10852 39080 -10788
rect 39144 -10852 39164 -10788
rect 39060 -10868 39164 -10852
rect 39060 -10932 39080 -10868
rect 39144 -10932 39164 -10868
rect 39060 -10948 39164 -10932
rect 39060 -11012 39080 -10948
rect 39144 -11012 39164 -10948
rect 39060 -11028 39164 -11012
rect 39060 -11092 39080 -11028
rect 39144 -11092 39164 -11028
rect 39060 -11108 39164 -11092
rect 39060 -11172 39080 -11108
rect 39144 -11172 39164 -11108
rect 39060 -11188 39164 -11172
rect 39060 -11252 39080 -11188
rect 39144 -11252 39164 -11188
rect 39060 -11268 39164 -11252
rect 39060 -11332 39080 -11268
rect 39144 -11332 39164 -11268
rect 39060 -11348 39164 -11332
rect 39060 -11412 39080 -11348
rect 39144 -11412 39164 -11348
rect 39060 -11428 39164 -11412
rect 39060 -11492 39080 -11428
rect 39144 -11492 39164 -11428
rect 39060 -11508 39164 -11492
rect 39060 -11572 39080 -11508
rect 39144 -11572 39164 -11508
rect 39060 -11588 39164 -11572
rect 39060 -11652 39080 -11588
rect 39144 -11652 39164 -11588
rect 39060 -11668 39164 -11652
rect 39060 -11732 39080 -11668
rect 39144 -11732 39164 -11668
rect 39060 -11748 39164 -11732
rect 39060 -11812 39080 -11748
rect 39144 -11812 39164 -11748
rect 39060 -11828 39164 -11812
rect 39060 -11892 39080 -11828
rect 39144 -11892 39164 -11828
rect 39060 -11908 39164 -11892
rect 39060 -11972 39080 -11908
rect 39144 -11972 39164 -11908
rect 39060 -11988 39164 -11972
rect 39060 -12052 39080 -11988
rect 39144 -12052 39164 -11988
rect 39060 -12068 39164 -12052
rect 39060 -12132 39080 -12068
rect 39144 -12132 39164 -12068
rect 39060 -12148 39164 -12132
rect 39060 -12212 39080 -12148
rect 39144 -12212 39164 -12148
rect 39060 -12228 39164 -12212
rect 39060 -12292 39080 -12228
rect 39144 -12292 39164 -12228
rect 39060 -12308 39164 -12292
rect 39060 -12372 39080 -12308
rect 39144 -12372 39164 -12308
rect 39060 -12388 39164 -12372
rect 39060 -12452 39080 -12388
rect 39144 -12452 39164 -12388
rect 39060 -12468 39164 -12452
rect 39060 -12532 39080 -12468
rect 39144 -12532 39164 -12468
rect 39060 -12548 39164 -12532
rect 39060 -12612 39080 -12548
rect 39144 -12612 39164 -12548
rect 39060 -12628 39164 -12612
rect 39060 -12692 39080 -12628
rect 39144 -12692 39164 -12628
rect 39060 -12708 39164 -12692
rect 39060 -12772 39080 -12708
rect 39144 -12772 39164 -12708
rect 39060 -12788 39164 -12772
rect 39060 -12852 39080 -12788
rect 39144 -12852 39164 -12788
rect 39060 -12868 39164 -12852
rect 39060 -12932 39080 -12868
rect 39144 -12932 39164 -12868
rect 39060 -12948 39164 -12932
rect 39060 -13012 39080 -12948
rect 39144 -13012 39164 -12948
rect 39060 -13028 39164 -13012
rect 39060 -13092 39080 -13028
rect 39144 -13092 39164 -13028
rect 39060 -13108 39164 -13092
rect 39060 -13172 39080 -13108
rect 39144 -13172 39164 -13108
rect 39060 -13188 39164 -13172
rect 39060 -13252 39080 -13188
rect 39144 -13252 39164 -13188
rect 39060 -13268 39164 -13252
rect 39060 -13332 39080 -13268
rect 39144 -13332 39164 -13268
rect 39060 -13348 39164 -13332
rect 39060 -13412 39080 -13348
rect 39144 -13412 39164 -13348
rect 39060 -13428 39164 -13412
rect 39060 -13492 39080 -13428
rect 39144 -13492 39164 -13428
rect 39060 -13508 39164 -13492
rect 39060 -13572 39080 -13508
rect 39144 -13572 39164 -13508
rect 39060 -13588 39164 -13572
rect 39060 -13652 39080 -13588
rect 39144 -13652 39164 -13588
rect 39060 -13668 39164 -13652
rect 39060 -13732 39080 -13668
rect 39144 -13732 39164 -13668
rect 39060 -13748 39164 -13732
rect 39060 -13812 39080 -13748
rect 39144 -13812 39164 -13748
rect 39060 -13828 39164 -13812
rect 39060 -13892 39080 -13828
rect 39144 -13892 39164 -13828
rect 39060 -13908 39164 -13892
rect 39060 -13972 39080 -13908
rect 39144 -13972 39164 -13908
rect 39060 -13988 39164 -13972
rect 39060 -14052 39080 -13988
rect 39144 -14052 39164 -13988
rect 39060 -14068 39164 -14052
rect 39060 -14132 39080 -14068
rect 39144 -14132 39164 -14068
rect 39060 -14148 39164 -14132
rect 39060 -14212 39080 -14148
rect 39144 -14212 39164 -14148
rect 39060 -14228 39164 -14212
rect 39060 -14292 39080 -14228
rect 39144 -14292 39164 -14228
rect 39060 -14308 39164 -14292
rect 39060 -14372 39080 -14308
rect 39144 -14372 39164 -14308
rect 39060 -14388 39164 -14372
rect 39060 -14452 39080 -14388
rect 39144 -14452 39164 -14388
rect 39060 -14468 39164 -14452
rect 39060 -14532 39080 -14468
rect 39144 -14532 39164 -14468
rect 39060 -14548 39164 -14532
rect 39060 -14612 39080 -14548
rect 39144 -14612 39164 -14548
rect 39060 -14628 39164 -14612
rect 39060 -14692 39080 -14628
rect 39144 -14692 39164 -14628
rect 39060 -14708 39164 -14692
rect 39060 -14772 39080 -14708
rect 39144 -14772 39164 -14708
rect 39060 -14788 39164 -14772
rect 39060 -14852 39080 -14788
rect 39144 -14852 39164 -14788
rect 39060 -14868 39164 -14852
rect 39060 -14932 39080 -14868
rect 39144 -14932 39164 -14868
rect 39060 -14948 39164 -14932
rect 39060 -15012 39080 -14948
rect 39144 -15012 39164 -14948
rect 39060 -15028 39164 -15012
rect 39060 -15092 39080 -15028
rect 39144 -15092 39164 -15028
rect 39060 -15108 39164 -15092
rect 39060 -15172 39080 -15108
rect 39144 -15172 39164 -15108
rect 39060 -15188 39164 -15172
rect 39060 -15252 39080 -15188
rect 39144 -15252 39164 -15188
rect 39060 -15268 39164 -15252
rect 39060 -15332 39080 -15268
rect 39144 -15332 39164 -15268
rect 39060 -15348 39164 -15332
rect 39060 -15412 39080 -15348
rect 39144 -15412 39164 -15348
rect 39060 -15428 39164 -15412
rect 39060 -15492 39080 -15428
rect 39144 -15492 39164 -15428
rect 39060 -15508 39164 -15492
rect 39060 -15572 39080 -15508
rect 39144 -15572 39164 -15508
rect 39060 -15588 39164 -15572
rect 39060 -15652 39080 -15588
rect 39144 -15652 39164 -15588
rect 39060 -15668 39164 -15652
rect 39060 -15732 39080 -15668
rect 39144 -15732 39164 -15668
rect 39060 -15748 39164 -15732
rect 33448 -16108 33552 -15812
rect 27836 -16188 27940 -16172
rect 27836 -16252 27856 -16188
rect 27920 -16252 27940 -16188
rect 27836 -16268 27940 -16252
rect 27836 -16332 27856 -16268
rect 27920 -16332 27940 -16268
rect 27836 -16348 27940 -16332
rect 27836 -16412 27856 -16348
rect 27920 -16412 27940 -16348
rect 27836 -16428 27940 -16412
rect 27836 -16492 27856 -16428
rect 27920 -16492 27940 -16428
rect 27836 -16508 27940 -16492
rect 27836 -16572 27856 -16508
rect 27920 -16572 27940 -16508
rect 27836 -16588 27940 -16572
rect 27836 -16652 27856 -16588
rect 27920 -16652 27940 -16588
rect 27836 -16668 27940 -16652
rect 27836 -16732 27856 -16668
rect 27920 -16732 27940 -16668
rect 27836 -16748 27940 -16732
rect 27836 -16812 27856 -16748
rect 27920 -16812 27940 -16748
rect 27836 -16828 27940 -16812
rect 27836 -16892 27856 -16828
rect 27920 -16892 27940 -16828
rect 27836 -16908 27940 -16892
rect 27836 -16972 27856 -16908
rect 27920 -16972 27940 -16908
rect 27836 -16988 27940 -16972
rect 27836 -17052 27856 -16988
rect 27920 -17052 27940 -16988
rect 27836 -17068 27940 -17052
rect 27836 -17132 27856 -17068
rect 27920 -17132 27940 -17068
rect 27836 -17148 27940 -17132
rect 27836 -17212 27856 -17148
rect 27920 -17212 27940 -17148
rect 27836 -17228 27940 -17212
rect 27836 -17292 27856 -17228
rect 27920 -17292 27940 -17228
rect 27836 -17308 27940 -17292
rect 27836 -17372 27856 -17308
rect 27920 -17372 27940 -17308
rect 27836 -17388 27940 -17372
rect 27836 -17452 27856 -17388
rect 27920 -17452 27940 -17388
rect 27836 -17468 27940 -17452
rect 27836 -17532 27856 -17468
rect 27920 -17532 27940 -17468
rect 27836 -17548 27940 -17532
rect 27836 -17612 27856 -17548
rect 27920 -17612 27940 -17548
rect 27836 -17628 27940 -17612
rect 27836 -17692 27856 -17628
rect 27920 -17692 27940 -17628
rect 27836 -17708 27940 -17692
rect 27836 -17772 27856 -17708
rect 27920 -17772 27940 -17708
rect 27836 -17788 27940 -17772
rect 27836 -17852 27856 -17788
rect 27920 -17852 27940 -17788
rect 27836 -17868 27940 -17852
rect 27836 -17932 27856 -17868
rect 27920 -17932 27940 -17868
rect 27836 -17948 27940 -17932
rect 27836 -18012 27856 -17948
rect 27920 -18012 27940 -17948
rect 27836 -18028 27940 -18012
rect 27836 -18092 27856 -18028
rect 27920 -18092 27940 -18028
rect 27836 -18108 27940 -18092
rect 27836 -18172 27856 -18108
rect 27920 -18172 27940 -18108
rect 27836 -18188 27940 -18172
rect 27836 -18252 27856 -18188
rect 27920 -18252 27940 -18188
rect 27836 -18268 27940 -18252
rect 27836 -18332 27856 -18268
rect 27920 -18332 27940 -18268
rect 27836 -18348 27940 -18332
rect 27836 -18412 27856 -18348
rect 27920 -18412 27940 -18348
rect 27836 -18428 27940 -18412
rect 27836 -18492 27856 -18428
rect 27920 -18492 27940 -18428
rect 27836 -18508 27940 -18492
rect 27836 -18572 27856 -18508
rect 27920 -18572 27940 -18508
rect 27836 -18588 27940 -18572
rect 27836 -18652 27856 -18588
rect 27920 -18652 27940 -18588
rect 27836 -18668 27940 -18652
rect 27836 -18732 27856 -18668
rect 27920 -18732 27940 -18668
rect 27836 -18748 27940 -18732
rect 27836 -18812 27856 -18748
rect 27920 -18812 27940 -18748
rect 27836 -18828 27940 -18812
rect 27836 -18892 27856 -18828
rect 27920 -18892 27940 -18828
rect 27836 -18908 27940 -18892
rect 27836 -18972 27856 -18908
rect 27920 -18972 27940 -18908
rect 27836 -18988 27940 -18972
rect 27836 -19052 27856 -18988
rect 27920 -19052 27940 -18988
rect 27836 -19068 27940 -19052
rect 27836 -19132 27856 -19068
rect 27920 -19132 27940 -19068
rect 27836 -19148 27940 -19132
rect 27836 -19212 27856 -19148
rect 27920 -19212 27940 -19148
rect 27836 -19228 27940 -19212
rect 27836 -19292 27856 -19228
rect 27920 -19292 27940 -19228
rect 27836 -19308 27940 -19292
rect 27836 -19372 27856 -19308
rect 27920 -19372 27940 -19308
rect 27836 -19388 27940 -19372
rect 27836 -19452 27856 -19388
rect 27920 -19452 27940 -19388
rect 27836 -19468 27940 -19452
rect 27836 -19532 27856 -19468
rect 27920 -19532 27940 -19468
rect 27836 -19548 27940 -19532
rect 27836 -19612 27856 -19548
rect 27920 -19612 27940 -19548
rect 27836 -19628 27940 -19612
rect 27836 -19692 27856 -19628
rect 27920 -19692 27940 -19628
rect 27836 -19708 27940 -19692
rect 27836 -19772 27856 -19708
rect 27920 -19772 27940 -19708
rect 27836 -19788 27940 -19772
rect 27836 -19852 27856 -19788
rect 27920 -19852 27940 -19788
rect 27836 -19868 27940 -19852
rect 27836 -19932 27856 -19868
rect 27920 -19932 27940 -19868
rect 27836 -19948 27940 -19932
rect 27836 -20012 27856 -19948
rect 27920 -20012 27940 -19948
rect 27836 -20028 27940 -20012
rect 27836 -20092 27856 -20028
rect 27920 -20092 27940 -20028
rect 27836 -20108 27940 -20092
rect 27836 -20172 27856 -20108
rect 27920 -20172 27940 -20108
rect 27836 -20188 27940 -20172
rect 27836 -20252 27856 -20188
rect 27920 -20252 27940 -20188
rect 27836 -20268 27940 -20252
rect 27836 -20332 27856 -20268
rect 27920 -20332 27940 -20268
rect 27836 -20348 27940 -20332
rect 27836 -20412 27856 -20348
rect 27920 -20412 27940 -20348
rect 27836 -20428 27940 -20412
rect 27836 -20492 27856 -20428
rect 27920 -20492 27940 -20428
rect 27836 -20508 27940 -20492
rect 27836 -20572 27856 -20508
rect 27920 -20572 27940 -20508
rect 27836 -20588 27940 -20572
rect 27836 -20652 27856 -20588
rect 27920 -20652 27940 -20588
rect 27836 -20668 27940 -20652
rect 27836 -20732 27856 -20668
rect 27920 -20732 27940 -20668
rect 27836 -20748 27940 -20732
rect 27836 -20812 27856 -20748
rect 27920 -20812 27940 -20748
rect 27836 -20828 27940 -20812
rect 27836 -20892 27856 -20828
rect 27920 -20892 27940 -20828
rect 27836 -20908 27940 -20892
rect 27836 -20972 27856 -20908
rect 27920 -20972 27940 -20908
rect 27836 -20988 27940 -20972
rect 27836 -21052 27856 -20988
rect 27920 -21052 27940 -20988
rect 27836 -21068 27940 -21052
rect 22224 -21428 22328 -21132
rect 16612 -21508 16716 -21492
rect 16612 -21572 16632 -21508
rect 16696 -21572 16716 -21508
rect 16612 -21588 16716 -21572
rect 16612 -21652 16632 -21588
rect 16696 -21652 16716 -21588
rect 16612 -21668 16716 -21652
rect 16612 -21732 16632 -21668
rect 16696 -21732 16716 -21668
rect 16612 -21748 16716 -21732
rect 16612 -21812 16632 -21748
rect 16696 -21812 16716 -21748
rect 16612 -21828 16716 -21812
rect 16612 -21892 16632 -21828
rect 16696 -21892 16716 -21828
rect 16612 -21908 16716 -21892
rect 16612 -21972 16632 -21908
rect 16696 -21972 16716 -21908
rect 16612 -21988 16716 -21972
rect 16612 -22052 16632 -21988
rect 16696 -22052 16716 -21988
rect 16612 -22068 16716 -22052
rect 16612 -22132 16632 -22068
rect 16696 -22132 16716 -22068
rect 16612 -22148 16716 -22132
rect 16612 -22212 16632 -22148
rect 16696 -22212 16716 -22148
rect 16612 -22228 16716 -22212
rect 16612 -22292 16632 -22228
rect 16696 -22292 16716 -22228
rect 16612 -22308 16716 -22292
rect 16612 -22372 16632 -22308
rect 16696 -22372 16716 -22308
rect 16612 -22388 16716 -22372
rect 16612 -22452 16632 -22388
rect 16696 -22452 16716 -22388
rect 16612 -22468 16716 -22452
rect 16612 -22532 16632 -22468
rect 16696 -22532 16716 -22468
rect 16612 -22548 16716 -22532
rect 16612 -22612 16632 -22548
rect 16696 -22612 16716 -22548
rect 16612 -22628 16716 -22612
rect 16612 -22692 16632 -22628
rect 16696 -22692 16716 -22628
rect 16612 -22708 16716 -22692
rect 16612 -22772 16632 -22708
rect 16696 -22772 16716 -22708
rect 16612 -22788 16716 -22772
rect 16612 -22852 16632 -22788
rect 16696 -22852 16716 -22788
rect 16612 -22868 16716 -22852
rect 16612 -22932 16632 -22868
rect 16696 -22932 16716 -22868
rect 16612 -22948 16716 -22932
rect 16612 -23012 16632 -22948
rect 16696 -23012 16716 -22948
rect 16612 -23028 16716 -23012
rect 16612 -23092 16632 -23028
rect 16696 -23092 16716 -23028
rect 16612 -23108 16716 -23092
rect 16612 -23172 16632 -23108
rect 16696 -23172 16716 -23108
rect 16612 -23188 16716 -23172
rect 16612 -23252 16632 -23188
rect 16696 -23252 16716 -23188
rect 16612 -23268 16716 -23252
rect 16612 -23332 16632 -23268
rect 16696 -23332 16716 -23268
rect 16612 -23348 16716 -23332
rect 16612 -23412 16632 -23348
rect 16696 -23412 16716 -23348
rect 16612 -23428 16716 -23412
rect 16612 -23492 16632 -23428
rect 16696 -23492 16716 -23428
rect 16612 -23508 16716 -23492
rect 16612 -23572 16632 -23508
rect 16696 -23572 16716 -23508
rect 16612 -23588 16716 -23572
rect 16612 -23652 16632 -23588
rect 16696 -23652 16716 -23588
rect 16612 -23668 16716 -23652
rect 16612 -23732 16632 -23668
rect 16696 -23732 16716 -23668
rect 16612 -23748 16716 -23732
rect 16612 -23812 16632 -23748
rect 16696 -23812 16716 -23748
rect 16612 -23828 16716 -23812
rect 16612 -23892 16632 -23828
rect 16696 -23892 16716 -23828
rect 16612 -23908 16716 -23892
rect 16612 -23972 16632 -23908
rect 16696 -23972 16716 -23908
rect 16612 -23988 16716 -23972
rect 16612 -24052 16632 -23988
rect 16696 -24052 16716 -23988
rect 16612 -24068 16716 -24052
rect 16612 -24132 16632 -24068
rect 16696 -24132 16716 -24068
rect 16612 -24148 16716 -24132
rect 16612 -24212 16632 -24148
rect 16696 -24212 16716 -24148
rect 16612 -24228 16716 -24212
rect 16612 -24292 16632 -24228
rect 16696 -24292 16716 -24228
rect 16612 -24308 16716 -24292
rect 16612 -24372 16632 -24308
rect 16696 -24372 16716 -24308
rect 16612 -24388 16716 -24372
rect 16612 -24452 16632 -24388
rect 16696 -24452 16716 -24388
rect 16612 -24468 16716 -24452
rect 16612 -24532 16632 -24468
rect 16696 -24532 16716 -24468
rect 16612 -24548 16716 -24532
rect 16612 -24612 16632 -24548
rect 16696 -24612 16716 -24548
rect 16612 -24628 16716 -24612
rect 16612 -24692 16632 -24628
rect 16696 -24692 16716 -24628
rect 16612 -24708 16716 -24692
rect 16612 -24772 16632 -24708
rect 16696 -24772 16716 -24708
rect 16612 -24788 16716 -24772
rect 16612 -24852 16632 -24788
rect 16696 -24852 16716 -24788
rect 16612 -24868 16716 -24852
rect 16612 -24932 16632 -24868
rect 16696 -24932 16716 -24868
rect 16612 -24948 16716 -24932
rect 16612 -25012 16632 -24948
rect 16696 -25012 16716 -24948
rect 16612 -25028 16716 -25012
rect 16612 -25092 16632 -25028
rect 16696 -25092 16716 -25028
rect 16612 -25108 16716 -25092
rect 16612 -25172 16632 -25108
rect 16696 -25172 16716 -25108
rect 16612 -25188 16716 -25172
rect 16612 -25252 16632 -25188
rect 16696 -25252 16716 -25188
rect 16612 -25268 16716 -25252
rect 16612 -25332 16632 -25268
rect 16696 -25332 16716 -25268
rect 16612 -25348 16716 -25332
rect 16612 -25412 16632 -25348
rect 16696 -25412 16716 -25348
rect 16612 -25428 16716 -25412
rect 16612 -25492 16632 -25428
rect 16696 -25492 16716 -25428
rect 16612 -25508 16716 -25492
rect 16612 -25572 16632 -25508
rect 16696 -25572 16716 -25508
rect 16612 -25588 16716 -25572
rect 16612 -25652 16632 -25588
rect 16696 -25652 16716 -25588
rect 16612 -25668 16716 -25652
rect 16612 -25732 16632 -25668
rect 16696 -25732 16716 -25668
rect 16612 -25748 16716 -25732
rect 16612 -25812 16632 -25748
rect 16696 -25812 16716 -25748
rect 16612 -25828 16716 -25812
rect 16612 -25892 16632 -25828
rect 16696 -25892 16716 -25828
rect 16612 -25908 16716 -25892
rect 16612 -25972 16632 -25908
rect 16696 -25972 16716 -25908
rect 16612 -25988 16716 -25972
rect 16612 -26052 16632 -25988
rect 16696 -26052 16716 -25988
rect 16612 -26068 16716 -26052
rect 16612 -26132 16632 -26068
rect 16696 -26132 16716 -26068
rect 16612 -26148 16716 -26132
rect 16612 -26212 16632 -26148
rect 16696 -26212 16716 -26148
rect 16612 -26228 16716 -26212
rect 16612 -26292 16632 -26228
rect 16696 -26292 16716 -26228
rect 16612 -26308 16716 -26292
rect 16612 -26372 16632 -26308
rect 16696 -26372 16716 -26308
rect 16612 -26388 16716 -26372
rect 11000 -26748 11104 -26452
rect 5388 -26828 5492 -26812
rect 5388 -26892 5408 -26828
rect 5472 -26892 5492 -26828
rect 5388 -26908 5492 -26892
rect 5388 -26972 5408 -26908
rect 5472 -26972 5492 -26908
rect 5388 -26988 5492 -26972
rect 5388 -27052 5408 -26988
rect 5472 -27052 5492 -26988
rect 5388 -27068 5492 -27052
rect 5388 -27132 5408 -27068
rect 5472 -27132 5492 -27068
rect 5388 -27148 5492 -27132
rect 5388 -27212 5408 -27148
rect 5472 -27212 5492 -27148
rect 5388 -27228 5492 -27212
rect 5388 -27292 5408 -27228
rect 5472 -27292 5492 -27228
rect 5388 -27308 5492 -27292
rect 5388 -27372 5408 -27308
rect 5472 -27372 5492 -27308
rect 5388 -27388 5492 -27372
rect 5388 -27452 5408 -27388
rect 5472 -27452 5492 -27388
rect 5388 -27468 5492 -27452
rect 5388 -27532 5408 -27468
rect 5472 -27532 5492 -27468
rect 5388 -27548 5492 -27532
rect 5388 -27612 5408 -27548
rect 5472 -27612 5492 -27548
rect 5388 -27628 5492 -27612
rect 5388 -27692 5408 -27628
rect 5472 -27692 5492 -27628
rect 5388 -27708 5492 -27692
rect 5388 -27772 5408 -27708
rect 5472 -27772 5492 -27708
rect 5388 -27788 5492 -27772
rect 5388 -27852 5408 -27788
rect 5472 -27852 5492 -27788
rect 5388 -27868 5492 -27852
rect 5388 -27932 5408 -27868
rect 5472 -27932 5492 -27868
rect 5388 -27948 5492 -27932
rect 5388 -28012 5408 -27948
rect 5472 -28012 5492 -27948
rect 5388 -28028 5492 -28012
rect 5388 -28092 5408 -28028
rect 5472 -28092 5492 -28028
rect 5388 -28108 5492 -28092
rect 5388 -28172 5408 -28108
rect 5472 -28172 5492 -28108
rect 5388 -28188 5492 -28172
rect 5388 -28252 5408 -28188
rect 5472 -28252 5492 -28188
rect 5388 -28268 5492 -28252
rect 5388 -28332 5408 -28268
rect 5472 -28332 5492 -28268
rect 5388 -28348 5492 -28332
rect 5388 -28412 5408 -28348
rect 5472 -28412 5492 -28348
rect 5388 -28428 5492 -28412
rect 5388 -28492 5408 -28428
rect 5472 -28492 5492 -28428
rect 5388 -28508 5492 -28492
rect 5388 -28572 5408 -28508
rect 5472 -28572 5492 -28508
rect 5388 -28588 5492 -28572
rect 5388 -28652 5408 -28588
rect 5472 -28652 5492 -28588
rect 5388 -28668 5492 -28652
rect 5388 -28732 5408 -28668
rect 5472 -28732 5492 -28668
rect 5388 -28748 5492 -28732
rect 5388 -28812 5408 -28748
rect 5472 -28812 5492 -28748
rect 5388 -28828 5492 -28812
rect 5388 -28892 5408 -28828
rect 5472 -28892 5492 -28828
rect 5388 -28908 5492 -28892
rect 5388 -28972 5408 -28908
rect 5472 -28972 5492 -28908
rect 5388 -28988 5492 -28972
rect 5388 -29052 5408 -28988
rect 5472 -29052 5492 -28988
rect 5388 -29068 5492 -29052
rect 5388 -29132 5408 -29068
rect 5472 -29132 5492 -29068
rect 5388 -29148 5492 -29132
rect 5388 -29212 5408 -29148
rect 5472 -29212 5492 -29148
rect 5388 -29228 5492 -29212
rect 5388 -29292 5408 -29228
rect 5472 -29292 5492 -29228
rect 5388 -29308 5492 -29292
rect 5388 -29372 5408 -29308
rect 5472 -29372 5492 -29308
rect 5388 -29388 5492 -29372
rect 5388 -29452 5408 -29388
rect 5472 -29452 5492 -29388
rect 5388 -29468 5492 -29452
rect 5388 -29532 5408 -29468
rect 5472 -29532 5492 -29468
rect 5388 -29548 5492 -29532
rect 5388 -29612 5408 -29548
rect 5472 -29612 5492 -29548
rect 5388 -29628 5492 -29612
rect 5388 -29692 5408 -29628
rect 5472 -29692 5492 -29628
rect 5388 -29708 5492 -29692
rect 5388 -29772 5408 -29708
rect 5472 -29772 5492 -29708
rect 5388 -29788 5492 -29772
rect 5388 -29852 5408 -29788
rect 5472 -29852 5492 -29788
rect 5388 -29868 5492 -29852
rect 5388 -29932 5408 -29868
rect 5472 -29932 5492 -29868
rect 5388 -29948 5492 -29932
rect 5388 -30012 5408 -29948
rect 5472 -30012 5492 -29948
rect 5388 -30028 5492 -30012
rect 5388 -30092 5408 -30028
rect 5472 -30092 5492 -30028
rect 5388 -30108 5492 -30092
rect 5388 -30172 5408 -30108
rect 5472 -30172 5492 -30108
rect 5388 -30188 5492 -30172
rect 5388 -30252 5408 -30188
rect 5472 -30252 5492 -30188
rect 5388 -30268 5492 -30252
rect 5388 -30332 5408 -30268
rect 5472 -30332 5492 -30268
rect 5388 -30348 5492 -30332
rect 5388 -30412 5408 -30348
rect 5472 -30412 5492 -30348
rect 5388 -30428 5492 -30412
rect 5388 -30492 5408 -30428
rect 5472 -30492 5492 -30428
rect 5388 -30508 5492 -30492
rect 5388 -30572 5408 -30508
rect 5472 -30572 5492 -30508
rect 5388 -30588 5492 -30572
rect 5388 -30652 5408 -30588
rect 5472 -30652 5492 -30588
rect 5388 -30668 5492 -30652
rect 5388 -30732 5408 -30668
rect 5472 -30732 5492 -30668
rect 5388 -30748 5492 -30732
rect 5388 -30812 5408 -30748
rect 5472 -30812 5492 -30748
rect 5388 -30828 5492 -30812
rect 5388 -30892 5408 -30828
rect 5472 -30892 5492 -30828
rect 5388 -30908 5492 -30892
rect 5388 -30972 5408 -30908
rect 5472 -30972 5492 -30908
rect 5388 -30988 5492 -30972
rect 5388 -31052 5408 -30988
rect 5472 -31052 5492 -30988
rect 5388 -31068 5492 -31052
rect 5388 -31132 5408 -31068
rect 5472 -31132 5492 -31068
rect 5388 -31148 5492 -31132
rect 5388 -31212 5408 -31148
rect 5472 -31212 5492 -31148
rect 5388 -31228 5492 -31212
rect 5388 -31292 5408 -31228
rect 5472 -31292 5492 -31228
rect 5388 -31308 5492 -31292
rect 5388 -31372 5408 -31308
rect 5472 -31372 5492 -31308
rect 5388 -31388 5492 -31372
rect 5388 -31452 5408 -31388
rect 5472 -31452 5492 -31388
rect 5388 -31468 5492 -31452
rect 5388 -31532 5408 -31468
rect 5472 -31532 5492 -31468
rect 5388 -31548 5492 -31532
rect 5388 -31612 5408 -31548
rect 5472 -31612 5492 -31548
rect 5388 -31628 5492 -31612
rect 5388 -31692 5408 -31628
rect 5472 -31692 5492 -31628
rect 5388 -31708 5492 -31692
rect -224 -32068 -120 -31772
rect -5836 -32148 -5732 -32132
rect -5836 -32212 -5816 -32148
rect -5752 -32212 -5732 -32148
rect -5836 -32228 -5732 -32212
rect -5836 -32292 -5816 -32228
rect -5752 -32292 -5732 -32228
rect -5836 -32308 -5732 -32292
rect -5836 -32372 -5816 -32308
rect -5752 -32372 -5732 -32308
rect -5836 -32388 -5732 -32372
rect -5836 -32452 -5816 -32388
rect -5752 -32452 -5732 -32388
rect -5836 -32468 -5732 -32452
rect -5836 -32532 -5816 -32468
rect -5752 -32532 -5732 -32468
rect -5836 -32548 -5732 -32532
rect -5836 -32612 -5816 -32548
rect -5752 -32612 -5732 -32548
rect -5836 -32628 -5732 -32612
rect -5836 -32692 -5816 -32628
rect -5752 -32692 -5732 -32628
rect -5836 -32708 -5732 -32692
rect -5836 -32772 -5816 -32708
rect -5752 -32772 -5732 -32708
rect -5836 -32788 -5732 -32772
rect -5836 -32852 -5816 -32788
rect -5752 -32852 -5732 -32788
rect -5836 -32868 -5732 -32852
rect -5836 -32932 -5816 -32868
rect -5752 -32932 -5732 -32868
rect -5836 -32948 -5732 -32932
rect -5836 -33012 -5816 -32948
rect -5752 -33012 -5732 -32948
rect -5836 -33028 -5732 -33012
rect -5836 -33092 -5816 -33028
rect -5752 -33092 -5732 -33028
rect -5836 -33108 -5732 -33092
rect -5836 -33172 -5816 -33108
rect -5752 -33172 -5732 -33108
rect -5836 -33188 -5732 -33172
rect -5836 -33252 -5816 -33188
rect -5752 -33252 -5732 -33188
rect -5836 -33268 -5732 -33252
rect -5836 -33332 -5816 -33268
rect -5752 -33332 -5732 -33268
rect -5836 -33348 -5732 -33332
rect -5836 -33412 -5816 -33348
rect -5752 -33412 -5732 -33348
rect -5836 -33428 -5732 -33412
rect -5836 -33492 -5816 -33428
rect -5752 -33492 -5732 -33428
rect -5836 -33508 -5732 -33492
rect -5836 -33572 -5816 -33508
rect -5752 -33572 -5732 -33508
rect -5836 -33588 -5732 -33572
rect -5836 -33652 -5816 -33588
rect -5752 -33652 -5732 -33588
rect -5836 -33668 -5732 -33652
rect -5836 -33732 -5816 -33668
rect -5752 -33732 -5732 -33668
rect -5836 -33748 -5732 -33732
rect -5836 -33812 -5816 -33748
rect -5752 -33812 -5732 -33748
rect -5836 -33828 -5732 -33812
rect -5836 -33892 -5816 -33828
rect -5752 -33892 -5732 -33828
rect -5836 -33908 -5732 -33892
rect -5836 -33972 -5816 -33908
rect -5752 -33972 -5732 -33908
rect -5836 -33988 -5732 -33972
rect -5836 -34052 -5816 -33988
rect -5752 -34052 -5732 -33988
rect -5836 -34068 -5732 -34052
rect -5836 -34132 -5816 -34068
rect -5752 -34132 -5732 -34068
rect -5836 -34148 -5732 -34132
rect -5836 -34212 -5816 -34148
rect -5752 -34212 -5732 -34148
rect -5836 -34228 -5732 -34212
rect -5836 -34292 -5816 -34228
rect -5752 -34292 -5732 -34228
rect -5836 -34308 -5732 -34292
rect -5836 -34372 -5816 -34308
rect -5752 -34372 -5732 -34308
rect -5836 -34388 -5732 -34372
rect -5836 -34452 -5816 -34388
rect -5752 -34452 -5732 -34388
rect -5836 -34468 -5732 -34452
rect -5836 -34532 -5816 -34468
rect -5752 -34532 -5732 -34468
rect -5836 -34548 -5732 -34532
rect -5836 -34612 -5816 -34548
rect -5752 -34612 -5732 -34548
rect -5836 -34628 -5732 -34612
rect -5836 -34692 -5816 -34628
rect -5752 -34692 -5732 -34628
rect -5836 -34708 -5732 -34692
rect -5836 -34772 -5816 -34708
rect -5752 -34772 -5732 -34708
rect -5836 -34788 -5732 -34772
rect -5836 -34852 -5816 -34788
rect -5752 -34852 -5732 -34788
rect -5836 -34868 -5732 -34852
rect -5836 -34932 -5816 -34868
rect -5752 -34932 -5732 -34868
rect -5836 -34948 -5732 -34932
rect -5836 -35012 -5816 -34948
rect -5752 -35012 -5732 -34948
rect -5836 -35028 -5732 -35012
rect -5836 -35092 -5816 -35028
rect -5752 -35092 -5732 -35028
rect -5836 -35108 -5732 -35092
rect -5836 -35172 -5816 -35108
rect -5752 -35172 -5732 -35108
rect -5836 -35188 -5732 -35172
rect -5836 -35252 -5816 -35188
rect -5752 -35252 -5732 -35188
rect -5836 -35268 -5732 -35252
rect -5836 -35332 -5816 -35268
rect -5752 -35332 -5732 -35268
rect -5836 -35348 -5732 -35332
rect -5836 -35412 -5816 -35348
rect -5752 -35412 -5732 -35348
rect -5836 -35428 -5732 -35412
rect -5836 -35492 -5816 -35428
rect -5752 -35492 -5732 -35428
rect -5836 -35508 -5732 -35492
rect -5836 -35572 -5816 -35508
rect -5752 -35572 -5732 -35508
rect -5836 -35588 -5732 -35572
rect -5836 -35652 -5816 -35588
rect -5752 -35652 -5732 -35588
rect -5836 -35668 -5732 -35652
rect -5836 -35732 -5816 -35668
rect -5752 -35732 -5732 -35668
rect -5836 -35748 -5732 -35732
rect -5836 -35812 -5816 -35748
rect -5752 -35812 -5732 -35748
rect -5836 -35828 -5732 -35812
rect -5836 -35892 -5816 -35828
rect -5752 -35892 -5732 -35828
rect -5836 -35908 -5732 -35892
rect -5836 -35972 -5816 -35908
rect -5752 -35972 -5732 -35908
rect -5836 -35988 -5732 -35972
rect -5836 -36052 -5816 -35988
rect -5752 -36052 -5732 -35988
rect -5836 -36068 -5732 -36052
rect -5836 -36132 -5816 -36068
rect -5752 -36132 -5732 -36068
rect -5836 -36148 -5732 -36132
rect -5836 -36212 -5816 -36148
rect -5752 -36212 -5732 -36148
rect -5836 -36228 -5732 -36212
rect -5836 -36292 -5816 -36228
rect -5752 -36292 -5732 -36228
rect -5836 -36308 -5732 -36292
rect -5836 -36372 -5816 -36308
rect -5752 -36372 -5732 -36308
rect -5836 -36388 -5732 -36372
rect -5836 -36452 -5816 -36388
rect -5752 -36452 -5732 -36388
rect -5836 -36468 -5732 -36452
rect -5836 -36532 -5816 -36468
rect -5752 -36532 -5732 -36468
rect -5836 -36548 -5732 -36532
rect -5836 -36612 -5816 -36548
rect -5752 -36612 -5732 -36548
rect -5836 -36628 -5732 -36612
rect -5836 -36692 -5816 -36628
rect -5752 -36692 -5732 -36628
rect -5836 -36708 -5732 -36692
rect -5836 -36772 -5816 -36708
rect -5752 -36772 -5732 -36708
rect -5836 -36788 -5732 -36772
rect -5836 -36852 -5816 -36788
rect -5752 -36852 -5732 -36788
rect -5836 -36868 -5732 -36852
rect -5836 -36932 -5816 -36868
rect -5752 -36932 -5732 -36868
rect -5836 -36948 -5732 -36932
rect -5836 -37012 -5816 -36948
rect -5752 -37012 -5732 -36948
rect -5836 -37028 -5732 -37012
rect -11448 -37240 -11344 -37092
rect -8616 -37240 -8512 -37041
rect -5836 -37092 -5816 -37028
rect -5752 -37092 -5732 -37028
rect -5413 -32148 -491 -32119
rect -5413 -37012 -5384 -32148
rect -520 -37012 -491 -32148
rect -5413 -37041 -491 -37012
rect -224 -32132 -204 -32068
rect -140 -32132 -120 -32068
rect 2608 -32119 2712 -31721
rect 5388 -31772 5408 -31708
rect 5472 -31772 5492 -31708
rect 5811 -26828 10733 -26799
rect 5811 -31692 5840 -26828
rect 10704 -31692 10733 -26828
rect 5811 -31721 10733 -31692
rect 11000 -26812 11020 -26748
rect 11084 -26812 11104 -26748
rect 13832 -26799 13936 -26401
rect 16612 -26452 16632 -26388
rect 16696 -26452 16716 -26388
rect 17035 -21508 21957 -21479
rect 17035 -26372 17064 -21508
rect 21928 -26372 21957 -21508
rect 17035 -26401 21957 -26372
rect 22224 -21492 22244 -21428
rect 22308 -21492 22328 -21428
rect 25056 -21479 25160 -21081
rect 27836 -21132 27856 -21068
rect 27920 -21132 27940 -21068
rect 28259 -16188 33181 -16159
rect 28259 -21052 28288 -16188
rect 33152 -21052 33181 -16188
rect 28259 -21081 33181 -21052
rect 33448 -16172 33468 -16108
rect 33532 -16172 33552 -16108
rect 36280 -16159 36384 -15761
rect 39060 -15812 39080 -15748
rect 39144 -15812 39164 -15748
rect 39060 -16108 39164 -15812
rect 33448 -16188 33552 -16172
rect 33448 -16252 33468 -16188
rect 33532 -16252 33552 -16188
rect 33448 -16268 33552 -16252
rect 33448 -16332 33468 -16268
rect 33532 -16332 33552 -16268
rect 33448 -16348 33552 -16332
rect 33448 -16412 33468 -16348
rect 33532 -16412 33552 -16348
rect 33448 -16428 33552 -16412
rect 33448 -16492 33468 -16428
rect 33532 -16492 33552 -16428
rect 33448 -16508 33552 -16492
rect 33448 -16572 33468 -16508
rect 33532 -16572 33552 -16508
rect 33448 -16588 33552 -16572
rect 33448 -16652 33468 -16588
rect 33532 -16652 33552 -16588
rect 33448 -16668 33552 -16652
rect 33448 -16732 33468 -16668
rect 33532 -16732 33552 -16668
rect 33448 -16748 33552 -16732
rect 33448 -16812 33468 -16748
rect 33532 -16812 33552 -16748
rect 33448 -16828 33552 -16812
rect 33448 -16892 33468 -16828
rect 33532 -16892 33552 -16828
rect 33448 -16908 33552 -16892
rect 33448 -16972 33468 -16908
rect 33532 -16972 33552 -16908
rect 33448 -16988 33552 -16972
rect 33448 -17052 33468 -16988
rect 33532 -17052 33552 -16988
rect 33448 -17068 33552 -17052
rect 33448 -17132 33468 -17068
rect 33532 -17132 33552 -17068
rect 33448 -17148 33552 -17132
rect 33448 -17212 33468 -17148
rect 33532 -17212 33552 -17148
rect 33448 -17228 33552 -17212
rect 33448 -17292 33468 -17228
rect 33532 -17292 33552 -17228
rect 33448 -17308 33552 -17292
rect 33448 -17372 33468 -17308
rect 33532 -17372 33552 -17308
rect 33448 -17388 33552 -17372
rect 33448 -17452 33468 -17388
rect 33532 -17452 33552 -17388
rect 33448 -17468 33552 -17452
rect 33448 -17532 33468 -17468
rect 33532 -17532 33552 -17468
rect 33448 -17548 33552 -17532
rect 33448 -17612 33468 -17548
rect 33532 -17612 33552 -17548
rect 33448 -17628 33552 -17612
rect 33448 -17692 33468 -17628
rect 33532 -17692 33552 -17628
rect 33448 -17708 33552 -17692
rect 33448 -17772 33468 -17708
rect 33532 -17772 33552 -17708
rect 33448 -17788 33552 -17772
rect 33448 -17852 33468 -17788
rect 33532 -17852 33552 -17788
rect 33448 -17868 33552 -17852
rect 33448 -17932 33468 -17868
rect 33532 -17932 33552 -17868
rect 33448 -17948 33552 -17932
rect 33448 -18012 33468 -17948
rect 33532 -18012 33552 -17948
rect 33448 -18028 33552 -18012
rect 33448 -18092 33468 -18028
rect 33532 -18092 33552 -18028
rect 33448 -18108 33552 -18092
rect 33448 -18172 33468 -18108
rect 33532 -18172 33552 -18108
rect 33448 -18188 33552 -18172
rect 33448 -18252 33468 -18188
rect 33532 -18252 33552 -18188
rect 33448 -18268 33552 -18252
rect 33448 -18332 33468 -18268
rect 33532 -18332 33552 -18268
rect 33448 -18348 33552 -18332
rect 33448 -18412 33468 -18348
rect 33532 -18412 33552 -18348
rect 33448 -18428 33552 -18412
rect 33448 -18492 33468 -18428
rect 33532 -18492 33552 -18428
rect 33448 -18508 33552 -18492
rect 33448 -18572 33468 -18508
rect 33532 -18572 33552 -18508
rect 33448 -18588 33552 -18572
rect 33448 -18652 33468 -18588
rect 33532 -18652 33552 -18588
rect 33448 -18668 33552 -18652
rect 33448 -18732 33468 -18668
rect 33532 -18732 33552 -18668
rect 33448 -18748 33552 -18732
rect 33448 -18812 33468 -18748
rect 33532 -18812 33552 -18748
rect 33448 -18828 33552 -18812
rect 33448 -18892 33468 -18828
rect 33532 -18892 33552 -18828
rect 33448 -18908 33552 -18892
rect 33448 -18972 33468 -18908
rect 33532 -18972 33552 -18908
rect 33448 -18988 33552 -18972
rect 33448 -19052 33468 -18988
rect 33532 -19052 33552 -18988
rect 33448 -19068 33552 -19052
rect 33448 -19132 33468 -19068
rect 33532 -19132 33552 -19068
rect 33448 -19148 33552 -19132
rect 33448 -19212 33468 -19148
rect 33532 -19212 33552 -19148
rect 33448 -19228 33552 -19212
rect 33448 -19292 33468 -19228
rect 33532 -19292 33552 -19228
rect 33448 -19308 33552 -19292
rect 33448 -19372 33468 -19308
rect 33532 -19372 33552 -19308
rect 33448 -19388 33552 -19372
rect 33448 -19452 33468 -19388
rect 33532 -19452 33552 -19388
rect 33448 -19468 33552 -19452
rect 33448 -19532 33468 -19468
rect 33532 -19532 33552 -19468
rect 33448 -19548 33552 -19532
rect 33448 -19612 33468 -19548
rect 33532 -19612 33552 -19548
rect 33448 -19628 33552 -19612
rect 33448 -19692 33468 -19628
rect 33532 -19692 33552 -19628
rect 33448 -19708 33552 -19692
rect 33448 -19772 33468 -19708
rect 33532 -19772 33552 -19708
rect 33448 -19788 33552 -19772
rect 33448 -19852 33468 -19788
rect 33532 -19852 33552 -19788
rect 33448 -19868 33552 -19852
rect 33448 -19932 33468 -19868
rect 33532 -19932 33552 -19868
rect 33448 -19948 33552 -19932
rect 33448 -20012 33468 -19948
rect 33532 -20012 33552 -19948
rect 33448 -20028 33552 -20012
rect 33448 -20092 33468 -20028
rect 33532 -20092 33552 -20028
rect 33448 -20108 33552 -20092
rect 33448 -20172 33468 -20108
rect 33532 -20172 33552 -20108
rect 33448 -20188 33552 -20172
rect 33448 -20252 33468 -20188
rect 33532 -20252 33552 -20188
rect 33448 -20268 33552 -20252
rect 33448 -20332 33468 -20268
rect 33532 -20332 33552 -20268
rect 33448 -20348 33552 -20332
rect 33448 -20412 33468 -20348
rect 33532 -20412 33552 -20348
rect 33448 -20428 33552 -20412
rect 33448 -20492 33468 -20428
rect 33532 -20492 33552 -20428
rect 33448 -20508 33552 -20492
rect 33448 -20572 33468 -20508
rect 33532 -20572 33552 -20508
rect 33448 -20588 33552 -20572
rect 33448 -20652 33468 -20588
rect 33532 -20652 33552 -20588
rect 33448 -20668 33552 -20652
rect 33448 -20732 33468 -20668
rect 33532 -20732 33552 -20668
rect 33448 -20748 33552 -20732
rect 33448 -20812 33468 -20748
rect 33532 -20812 33552 -20748
rect 33448 -20828 33552 -20812
rect 33448 -20892 33468 -20828
rect 33532 -20892 33552 -20828
rect 33448 -20908 33552 -20892
rect 33448 -20972 33468 -20908
rect 33532 -20972 33552 -20908
rect 33448 -20988 33552 -20972
rect 33448 -21052 33468 -20988
rect 33532 -21052 33552 -20988
rect 33448 -21068 33552 -21052
rect 27836 -21428 27940 -21132
rect 22224 -21508 22328 -21492
rect 22224 -21572 22244 -21508
rect 22308 -21572 22328 -21508
rect 22224 -21588 22328 -21572
rect 22224 -21652 22244 -21588
rect 22308 -21652 22328 -21588
rect 22224 -21668 22328 -21652
rect 22224 -21732 22244 -21668
rect 22308 -21732 22328 -21668
rect 22224 -21748 22328 -21732
rect 22224 -21812 22244 -21748
rect 22308 -21812 22328 -21748
rect 22224 -21828 22328 -21812
rect 22224 -21892 22244 -21828
rect 22308 -21892 22328 -21828
rect 22224 -21908 22328 -21892
rect 22224 -21972 22244 -21908
rect 22308 -21972 22328 -21908
rect 22224 -21988 22328 -21972
rect 22224 -22052 22244 -21988
rect 22308 -22052 22328 -21988
rect 22224 -22068 22328 -22052
rect 22224 -22132 22244 -22068
rect 22308 -22132 22328 -22068
rect 22224 -22148 22328 -22132
rect 22224 -22212 22244 -22148
rect 22308 -22212 22328 -22148
rect 22224 -22228 22328 -22212
rect 22224 -22292 22244 -22228
rect 22308 -22292 22328 -22228
rect 22224 -22308 22328 -22292
rect 22224 -22372 22244 -22308
rect 22308 -22372 22328 -22308
rect 22224 -22388 22328 -22372
rect 22224 -22452 22244 -22388
rect 22308 -22452 22328 -22388
rect 22224 -22468 22328 -22452
rect 22224 -22532 22244 -22468
rect 22308 -22532 22328 -22468
rect 22224 -22548 22328 -22532
rect 22224 -22612 22244 -22548
rect 22308 -22612 22328 -22548
rect 22224 -22628 22328 -22612
rect 22224 -22692 22244 -22628
rect 22308 -22692 22328 -22628
rect 22224 -22708 22328 -22692
rect 22224 -22772 22244 -22708
rect 22308 -22772 22328 -22708
rect 22224 -22788 22328 -22772
rect 22224 -22852 22244 -22788
rect 22308 -22852 22328 -22788
rect 22224 -22868 22328 -22852
rect 22224 -22932 22244 -22868
rect 22308 -22932 22328 -22868
rect 22224 -22948 22328 -22932
rect 22224 -23012 22244 -22948
rect 22308 -23012 22328 -22948
rect 22224 -23028 22328 -23012
rect 22224 -23092 22244 -23028
rect 22308 -23092 22328 -23028
rect 22224 -23108 22328 -23092
rect 22224 -23172 22244 -23108
rect 22308 -23172 22328 -23108
rect 22224 -23188 22328 -23172
rect 22224 -23252 22244 -23188
rect 22308 -23252 22328 -23188
rect 22224 -23268 22328 -23252
rect 22224 -23332 22244 -23268
rect 22308 -23332 22328 -23268
rect 22224 -23348 22328 -23332
rect 22224 -23412 22244 -23348
rect 22308 -23412 22328 -23348
rect 22224 -23428 22328 -23412
rect 22224 -23492 22244 -23428
rect 22308 -23492 22328 -23428
rect 22224 -23508 22328 -23492
rect 22224 -23572 22244 -23508
rect 22308 -23572 22328 -23508
rect 22224 -23588 22328 -23572
rect 22224 -23652 22244 -23588
rect 22308 -23652 22328 -23588
rect 22224 -23668 22328 -23652
rect 22224 -23732 22244 -23668
rect 22308 -23732 22328 -23668
rect 22224 -23748 22328 -23732
rect 22224 -23812 22244 -23748
rect 22308 -23812 22328 -23748
rect 22224 -23828 22328 -23812
rect 22224 -23892 22244 -23828
rect 22308 -23892 22328 -23828
rect 22224 -23908 22328 -23892
rect 22224 -23972 22244 -23908
rect 22308 -23972 22328 -23908
rect 22224 -23988 22328 -23972
rect 22224 -24052 22244 -23988
rect 22308 -24052 22328 -23988
rect 22224 -24068 22328 -24052
rect 22224 -24132 22244 -24068
rect 22308 -24132 22328 -24068
rect 22224 -24148 22328 -24132
rect 22224 -24212 22244 -24148
rect 22308 -24212 22328 -24148
rect 22224 -24228 22328 -24212
rect 22224 -24292 22244 -24228
rect 22308 -24292 22328 -24228
rect 22224 -24308 22328 -24292
rect 22224 -24372 22244 -24308
rect 22308 -24372 22328 -24308
rect 22224 -24388 22328 -24372
rect 22224 -24452 22244 -24388
rect 22308 -24452 22328 -24388
rect 22224 -24468 22328 -24452
rect 22224 -24532 22244 -24468
rect 22308 -24532 22328 -24468
rect 22224 -24548 22328 -24532
rect 22224 -24612 22244 -24548
rect 22308 -24612 22328 -24548
rect 22224 -24628 22328 -24612
rect 22224 -24692 22244 -24628
rect 22308 -24692 22328 -24628
rect 22224 -24708 22328 -24692
rect 22224 -24772 22244 -24708
rect 22308 -24772 22328 -24708
rect 22224 -24788 22328 -24772
rect 22224 -24852 22244 -24788
rect 22308 -24852 22328 -24788
rect 22224 -24868 22328 -24852
rect 22224 -24932 22244 -24868
rect 22308 -24932 22328 -24868
rect 22224 -24948 22328 -24932
rect 22224 -25012 22244 -24948
rect 22308 -25012 22328 -24948
rect 22224 -25028 22328 -25012
rect 22224 -25092 22244 -25028
rect 22308 -25092 22328 -25028
rect 22224 -25108 22328 -25092
rect 22224 -25172 22244 -25108
rect 22308 -25172 22328 -25108
rect 22224 -25188 22328 -25172
rect 22224 -25252 22244 -25188
rect 22308 -25252 22328 -25188
rect 22224 -25268 22328 -25252
rect 22224 -25332 22244 -25268
rect 22308 -25332 22328 -25268
rect 22224 -25348 22328 -25332
rect 22224 -25412 22244 -25348
rect 22308 -25412 22328 -25348
rect 22224 -25428 22328 -25412
rect 22224 -25492 22244 -25428
rect 22308 -25492 22328 -25428
rect 22224 -25508 22328 -25492
rect 22224 -25572 22244 -25508
rect 22308 -25572 22328 -25508
rect 22224 -25588 22328 -25572
rect 22224 -25652 22244 -25588
rect 22308 -25652 22328 -25588
rect 22224 -25668 22328 -25652
rect 22224 -25732 22244 -25668
rect 22308 -25732 22328 -25668
rect 22224 -25748 22328 -25732
rect 22224 -25812 22244 -25748
rect 22308 -25812 22328 -25748
rect 22224 -25828 22328 -25812
rect 22224 -25892 22244 -25828
rect 22308 -25892 22328 -25828
rect 22224 -25908 22328 -25892
rect 22224 -25972 22244 -25908
rect 22308 -25972 22328 -25908
rect 22224 -25988 22328 -25972
rect 22224 -26052 22244 -25988
rect 22308 -26052 22328 -25988
rect 22224 -26068 22328 -26052
rect 22224 -26132 22244 -26068
rect 22308 -26132 22328 -26068
rect 22224 -26148 22328 -26132
rect 22224 -26212 22244 -26148
rect 22308 -26212 22328 -26148
rect 22224 -26228 22328 -26212
rect 22224 -26292 22244 -26228
rect 22308 -26292 22328 -26228
rect 22224 -26308 22328 -26292
rect 22224 -26372 22244 -26308
rect 22308 -26372 22328 -26308
rect 22224 -26388 22328 -26372
rect 16612 -26748 16716 -26452
rect 11000 -26828 11104 -26812
rect 11000 -26892 11020 -26828
rect 11084 -26892 11104 -26828
rect 11000 -26908 11104 -26892
rect 11000 -26972 11020 -26908
rect 11084 -26972 11104 -26908
rect 11000 -26988 11104 -26972
rect 11000 -27052 11020 -26988
rect 11084 -27052 11104 -26988
rect 11000 -27068 11104 -27052
rect 11000 -27132 11020 -27068
rect 11084 -27132 11104 -27068
rect 11000 -27148 11104 -27132
rect 11000 -27212 11020 -27148
rect 11084 -27212 11104 -27148
rect 11000 -27228 11104 -27212
rect 11000 -27292 11020 -27228
rect 11084 -27292 11104 -27228
rect 11000 -27308 11104 -27292
rect 11000 -27372 11020 -27308
rect 11084 -27372 11104 -27308
rect 11000 -27388 11104 -27372
rect 11000 -27452 11020 -27388
rect 11084 -27452 11104 -27388
rect 11000 -27468 11104 -27452
rect 11000 -27532 11020 -27468
rect 11084 -27532 11104 -27468
rect 11000 -27548 11104 -27532
rect 11000 -27612 11020 -27548
rect 11084 -27612 11104 -27548
rect 11000 -27628 11104 -27612
rect 11000 -27692 11020 -27628
rect 11084 -27692 11104 -27628
rect 11000 -27708 11104 -27692
rect 11000 -27772 11020 -27708
rect 11084 -27772 11104 -27708
rect 11000 -27788 11104 -27772
rect 11000 -27852 11020 -27788
rect 11084 -27852 11104 -27788
rect 11000 -27868 11104 -27852
rect 11000 -27932 11020 -27868
rect 11084 -27932 11104 -27868
rect 11000 -27948 11104 -27932
rect 11000 -28012 11020 -27948
rect 11084 -28012 11104 -27948
rect 11000 -28028 11104 -28012
rect 11000 -28092 11020 -28028
rect 11084 -28092 11104 -28028
rect 11000 -28108 11104 -28092
rect 11000 -28172 11020 -28108
rect 11084 -28172 11104 -28108
rect 11000 -28188 11104 -28172
rect 11000 -28252 11020 -28188
rect 11084 -28252 11104 -28188
rect 11000 -28268 11104 -28252
rect 11000 -28332 11020 -28268
rect 11084 -28332 11104 -28268
rect 11000 -28348 11104 -28332
rect 11000 -28412 11020 -28348
rect 11084 -28412 11104 -28348
rect 11000 -28428 11104 -28412
rect 11000 -28492 11020 -28428
rect 11084 -28492 11104 -28428
rect 11000 -28508 11104 -28492
rect 11000 -28572 11020 -28508
rect 11084 -28572 11104 -28508
rect 11000 -28588 11104 -28572
rect 11000 -28652 11020 -28588
rect 11084 -28652 11104 -28588
rect 11000 -28668 11104 -28652
rect 11000 -28732 11020 -28668
rect 11084 -28732 11104 -28668
rect 11000 -28748 11104 -28732
rect 11000 -28812 11020 -28748
rect 11084 -28812 11104 -28748
rect 11000 -28828 11104 -28812
rect 11000 -28892 11020 -28828
rect 11084 -28892 11104 -28828
rect 11000 -28908 11104 -28892
rect 11000 -28972 11020 -28908
rect 11084 -28972 11104 -28908
rect 11000 -28988 11104 -28972
rect 11000 -29052 11020 -28988
rect 11084 -29052 11104 -28988
rect 11000 -29068 11104 -29052
rect 11000 -29132 11020 -29068
rect 11084 -29132 11104 -29068
rect 11000 -29148 11104 -29132
rect 11000 -29212 11020 -29148
rect 11084 -29212 11104 -29148
rect 11000 -29228 11104 -29212
rect 11000 -29292 11020 -29228
rect 11084 -29292 11104 -29228
rect 11000 -29308 11104 -29292
rect 11000 -29372 11020 -29308
rect 11084 -29372 11104 -29308
rect 11000 -29388 11104 -29372
rect 11000 -29452 11020 -29388
rect 11084 -29452 11104 -29388
rect 11000 -29468 11104 -29452
rect 11000 -29532 11020 -29468
rect 11084 -29532 11104 -29468
rect 11000 -29548 11104 -29532
rect 11000 -29612 11020 -29548
rect 11084 -29612 11104 -29548
rect 11000 -29628 11104 -29612
rect 11000 -29692 11020 -29628
rect 11084 -29692 11104 -29628
rect 11000 -29708 11104 -29692
rect 11000 -29772 11020 -29708
rect 11084 -29772 11104 -29708
rect 11000 -29788 11104 -29772
rect 11000 -29852 11020 -29788
rect 11084 -29852 11104 -29788
rect 11000 -29868 11104 -29852
rect 11000 -29932 11020 -29868
rect 11084 -29932 11104 -29868
rect 11000 -29948 11104 -29932
rect 11000 -30012 11020 -29948
rect 11084 -30012 11104 -29948
rect 11000 -30028 11104 -30012
rect 11000 -30092 11020 -30028
rect 11084 -30092 11104 -30028
rect 11000 -30108 11104 -30092
rect 11000 -30172 11020 -30108
rect 11084 -30172 11104 -30108
rect 11000 -30188 11104 -30172
rect 11000 -30252 11020 -30188
rect 11084 -30252 11104 -30188
rect 11000 -30268 11104 -30252
rect 11000 -30332 11020 -30268
rect 11084 -30332 11104 -30268
rect 11000 -30348 11104 -30332
rect 11000 -30412 11020 -30348
rect 11084 -30412 11104 -30348
rect 11000 -30428 11104 -30412
rect 11000 -30492 11020 -30428
rect 11084 -30492 11104 -30428
rect 11000 -30508 11104 -30492
rect 11000 -30572 11020 -30508
rect 11084 -30572 11104 -30508
rect 11000 -30588 11104 -30572
rect 11000 -30652 11020 -30588
rect 11084 -30652 11104 -30588
rect 11000 -30668 11104 -30652
rect 11000 -30732 11020 -30668
rect 11084 -30732 11104 -30668
rect 11000 -30748 11104 -30732
rect 11000 -30812 11020 -30748
rect 11084 -30812 11104 -30748
rect 11000 -30828 11104 -30812
rect 11000 -30892 11020 -30828
rect 11084 -30892 11104 -30828
rect 11000 -30908 11104 -30892
rect 11000 -30972 11020 -30908
rect 11084 -30972 11104 -30908
rect 11000 -30988 11104 -30972
rect 11000 -31052 11020 -30988
rect 11084 -31052 11104 -30988
rect 11000 -31068 11104 -31052
rect 11000 -31132 11020 -31068
rect 11084 -31132 11104 -31068
rect 11000 -31148 11104 -31132
rect 11000 -31212 11020 -31148
rect 11084 -31212 11104 -31148
rect 11000 -31228 11104 -31212
rect 11000 -31292 11020 -31228
rect 11084 -31292 11104 -31228
rect 11000 -31308 11104 -31292
rect 11000 -31372 11020 -31308
rect 11084 -31372 11104 -31308
rect 11000 -31388 11104 -31372
rect 11000 -31452 11020 -31388
rect 11084 -31452 11104 -31388
rect 11000 -31468 11104 -31452
rect 11000 -31532 11020 -31468
rect 11084 -31532 11104 -31468
rect 11000 -31548 11104 -31532
rect 11000 -31612 11020 -31548
rect 11084 -31612 11104 -31548
rect 11000 -31628 11104 -31612
rect 11000 -31692 11020 -31628
rect 11084 -31692 11104 -31628
rect 11000 -31708 11104 -31692
rect 5388 -32068 5492 -31772
rect -224 -32148 -120 -32132
rect -224 -32212 -204 -32148
rect -140 -32212 -120 -32148
rect -224 -32228 -120 -32212
rect -224 -32292 -204 -32228
rect -140 -32292 -120 -32228
rect -224 -32308 -120 -32292
rect -224 -32372 -204 -32308
rect -140 -32372 -120 -32308
rect -224 -32388 -120 -32372
rect -224 -32452 -204 -32388
rect -140 -32452 -120 -32388
rect -224 -32468 -120 -32452
rect -224 -32532 -204 -32468
rect -140 -32532 -120 -32468
rect -224 -32548 -120 -32532
rect -224 -32612 -204 -32548
rect -140 -32612 -120 -32548
rect -224 -32628 -120 -32612
rect -224 -32692 -204 -32628
rect -140 -32692 -120 -32628
rect -224 -32708 -120 -32692
rect -224 -32772 -204 -32708
rect -140 -32772 -120 -32708
rect -224 -32788 -120 -32772
rect -224 -32852 -204 -32788
rect -140 -32852 -120 -32788
rect -224 -32868 -120 -32852
rect -224 -32932 -204 -32868
rect -140 -32932 -120 -32868
rect -224 -32948 -120 -32932
rect -224 -33012 -204 -32948
rect -140 -33012 -120 -32948
rect -224 -33028 -120 -33012
rect -224 -33092 -204 -33028
rect -140 -33092 -120 -33028
rect -224 -33108 -120 -33092
rect -224 -33172 -204 -33108
rect -140 -33172 -120 -33108
rect -224 -33188 -120 -33172
rect -224 -33252 -204 -33188
rect -140 -33252 -120 -33188
rect -224 -33268 -120 -33252
rect -224 -33332 -204 -33268
rect -140 -33332 -120 -33268
rect -224 -33348 -120 -33332
rect -224 -33412 -204 -33348
rect -140 -33412 -120 -33348
rect -224 -33428 -120 -33412
rect -224 -33492 -204 -33428
rect -140 -33492 -120 -33428
rect -224 -33508 -120 -33492
rect -224 -33572 -204 -33508
rect -140 -33572 -120 -33508
rect -224 -33588 -120 -33572
rect -224 -33652 -204 -33588
rect -140 -33652 -120 -33588
rect -224 -33668 -120 -33652
rect -224 -33732 -204 -33668
rect -140 -33732 -120 -33668
rect -224 -33748 -120 -33732
rect -224 -33812 -204 -33748
rect -140 -33812 -120 -33748
rect -224 -33828 -120 -33812
rect -224 -33892 -204 -33828
rect -140 -33892 -120 -33828
rect -224 -33908 -120 -33892
rect -224 -33972 -204 -33908
rect -140 -33972 -120 -33908
rect -224 -33988 -120 -33972
rect -224 -34052 -204 -33988
rect -140 -34052 -120 -33988
rect -224 -34068 -120 -34052
rect -224 -34132 -204 -34068
rect -140 -34132 -120 -34068
rect -224 -34148 -120 -34132
rect -224 -34212 -204 -34148
rect -140 -34212 -120 -34148
rect -224 -34228 -120 -34212
rect -224 -34292 -204 -34228
rect -140 -34292 -120 -34228
rect -224 -34308 -120 -34292
rect -224 -34372 -204 -34308
rect -140 -34372 -120 -34308
rect -224 -34388 -120 -34372
rect -224 -34452 -204 -34388
rect -140 -34452 -120 -34388
rect -224 -34468 -120 -34452
rect -224 -34532 -204 -34468
rect -140 -34532 -120 -34468
rect -224 -34548 -120 -34532
rect -224 -34612 -204 -34548
rect -140 -34612 -120 -34548
rect -224 -34628 -120 -34612
rect -224 -34692 -204 -34628
rect -140 -34692 -120 -34628
rect -224 -34708 -120 -34692
rect -224 -34772 -204 -34708
rect -140 -34772 -120 -34708
rect -224 -34788 -120 -34772
rect -224 -34852 -204 -34788
rect -140 -34852 -120 -34788
rect -224 -34868 -120 -34852
rect -224 -34932 -204 -34868
rect -140 -34932 -120 -34868
rect -224 -34948 -120 -34932
rect -224 -35012 -204 -34948
rect -140 -35012 -120 -34948
rect -224 -35028 -120 -35012
rect -224 -35092 -204 -35028
rect -140 -35092 -120 -35028
rect -224 -35108 -120 -35092
rect -224 -35172 -204 -35108
rect -140 -35172 -120 -35108
rect -224 -35188 -120 -35172
rect -224 -35252 -204 -35188
rect -140 -35252 -120 -35188
rect -224 -35268 -120 -35252
rect -224 -35332 -204 -35268
rect -140 -35332 -120 -35268
rect -224 -35348 -120 -35332
rect -224 -35412 -204 -35348
rect -140 -35412 -120 -35348
rect -224 -35428 -120 -35412
rect -224 -35492 -204 -35428
rect -140 -35492 -120 -35428
rect -224 -35508 -120 -35492
rect -224 -35572 -204 -35508
rect -140 -35572 -120 -35508
rect -224 -35588 -120 -35572
rect -224 -35652 -204 -35588
rect -140 -35652 -120 -35588
rect -224 -35668 -120 -35652
rect -224 -35732 -204 -35668
rect -140 -35732 -120 -35668
rect -224 -35748 -120 -35732
rect -224 -35812 -204 -35748
rect -140 -35812 -120 -35748
rect -224 -35828 -120 -35812
rect -224 -35892 -204 -35828
rect -140 -35892 -120 -35828
rect -224 -35908 -120 -35892
rect -224 -35972 -204 -35908
rect -140 -35972 -120 -35908
rect -224 -35988 -120 -35972
rect -224 -36052 -204 -35988
rect -140 -36052 -120 -35988
rect -224 -36068 -120 -36052
rect -224 -36132 -204 -36068
rect -140 -36132 -120 -36068
rect -224 -36148 -120 -36132
rect -224 -36212 -204 -36148
rect -140 -36212 -120 -36148
rect -224 -36228 -120 -36212
rect -224 -36292 -204 -36228
rect -140 -36292 -120 -36228
rect -224 -36308 -120 -36292
rect -224 -36372 -204 -36308
rect -140 -36372 -120 -36308
rect -224 -36388 -120 -36372
rect -224 -36452 -204 -36388
rect -140 -36452 -120 -36388
rect -224 -36468 -120 -36452
rect -224 -36532 -204 -36468
rect -140 -36532 -120 -36468
rect -224 -36548 -120 -36532
rect -224 -36612 -204 -36548
rect -140 -36612 -120 -36548
rect -224 -36628 -120 -36612
rect -224 -36692 -204 -36628
rect -140 -36692 -120 -36628
rect -224 -36708 -120 -36692
rect -224 -36772 -204 -36708
rect -140 -36772 -120 -36708
rect -224 -36788 -120 -36772
rect -224 -36852 -204 -36788
rect -140 -36852 -120 -36788
rect -224 -36868 -120 -36852
rect -224 -36932 -204 -36868
rect -140 -36932 -120 -36868
rect -224 -36948 -120 -36932
rect -224 -37012 -204 -36948
rect -140 -37012 -120 -36948
rect -224 -37028 -120 -37012
rect -5836 -37240 -5732 -37092
rect -3004 -37240 -2900 -37041
rect -224 -37092 -204 -37028
rect -140 -37092 -120 -37028
rect 199 -32148 5121 -32119
rect 199 -37012 228 -32148
rect 5092 -37012 5121 -32148
rect 199 -37041 5121 -37012
rect 5388 -32132 5408 -32068
rect 5472 -32132 5492 -32068
rect 8220 -32119 8324 -31721
rect 11000 -31772 11020 -31708
rect 11084 -31772 11104 -31708
rect 11423 -26828 16345 -26799
rect 11423 -31692 11452 -26828
rect 16316 -31692 16345 -26828
rect 11423 -31721 16345 -31692
rect 16612 -26812 16632 -26748
rect 16696 -26812 16716 -26748
rect 19444 -26799 19548 -26401
rect 22224 -26452 22244 -26388
rect 22308 -26452 22328 -26388
rect 22647 -21508 27569 -21479
rect 22647 -26372 22676 -21508
rect 27540 -26372 27569 -21508
rect 22647 -26401 27569 -26372
rect 27836 -21492 27856 -21428
rect 27920 -21492 27940 -21428
rect 30668 -21479 30772 -21081
rect 33448 -21132 33468 -21068
rect 33532 -21132 33552 -21068
rect 33871 -16188 38793 -16159
rect 33871 -21052 33900 -16188
rect 38764 -21052 38793 -16188
rect 33871 -21081 38793 -21052
rect 39060 -16172 39080 -16108
rect 39144 -16172 39164 -16108
rect 39060 -16188 39164 -16172
rect 39060 -16252 39080 -16188
rect 39144 -16252 39164 -16188
rect 39060 -16268 39164 -16252
rect 39060 -16332 39080 -16268
rect 39144 -16332 39164 -16268
rect 39060 -16348 39164 -16332
rect 39060 -16412 39080 -16348
rect 39144 -16412 39164 -16348
rect 39060 -16428 39164 -16412
rect 39060 -16492 39080 -16428
rect 39144 -16492 39164 -16428
rect 39060 -16508 39164 -16492
rect 39060 -16572 39080 -16508
rect 39144 -16572 39164 -16508
rect 39060 -16588 39164 -16572
rect 39060 -16652 39080 -16588
rect 39144 -16652 39164 -16588
rect 39060 -16668 39164 -16652
rect 39060 -16732 39080 -16668
rect 39144 -16732 39164 -16668
rect 39060 -16748 39164 -16732
rect 39060 -16812 39080 -16748
rect 39144 -16812 39164 -16748
rect 39060 -16828 39164 -16812
rect 39060 -16892 39080 -16828
rect 39144 -16892 39164 -16828
rect 39060 -16908 39164 -16892
rect 39060 -16972 39080 -16908
rect 39144 -16972 39164 -16908
rect 39060 -16988 39164 -16972
rect 39060 -17052 39080 -16988
rect 39144 -17052 39164 -16988
rect 39060 -17068 39164 -17052
rect 39060 -17132 39080 -17068
rect 39144 -17132 39164 -17068
rect 39060 -17148 39164 -17132
rect 39060 -17212 39080 -17148
rect 39144 -17212 39164 -17148
rect 39060 -17228 39164 -17212
rect 39060 -17292 39080 -17228
rect 39144 -17292 39164 -17228
rect 39060 -17308 39164 -17292
rect 39060 -17372 39080 -17308
rect 39144 -17372 39164 -17308
rect 39060 -17388 39164 -17372
rect 39060 -17452 39080 -17388
rect 39144 -17452 39164 -17388
rect 39060 -17468 39164 -17452
rect 39060 -17532 39080 -17468
rect 39144 -17532 39164 -17468
rect 39060 -17548 39164 -17532
rect 39060 -17612 39080 -17548
rect 39144 -17612 39164 -17548
rect 39060 -17628 39164 -17612
rect 39060 -17692 39080 -17628
rect 39144 -17692 39164 -17628
rect 39060 -17708 39164 -17692
rect 39060 -17772 39080 -17708
rect 39144 -17772 39164 -17708
rect 39060 -17788 39164 -17772
rect 39060 -17852 39080 -17788
rect 39144 -17852 39164 -17788
rect 39060 -17868 39164 -17852
rect 39060 -17932 39080 -17868
rect 39144 -17932 39164 -17868
rect 39060 -17948 39164 -17932
rect 39060 -18012 39080 -17948
rect 39144 -18012 39164 -17948
rect 39060 -18028 39164 -18012
rect 39060 -18092 39080 -18028
rect 39144 -18092 39164 -18028
rect 39060 -18108 39164 -18092
rect 39060 -18172 39080 -18108
rect 39144 -18172 39164 -18108
rect 39060 -18188 39164 -18172
rect 39060 -18252 39080 -18188
rect 39144 -18252 39164 -18188
rect 39060 -18268 39164 -18252
rect 39060 -18332 39080 -18268
rect 39144 -18332 39164 -18268
rect 39060 -18348 39164 -18332
rect 39060 -18412 39080 -18348
rect 39144 -18412 39164 -18348
rect 39060 -18428 39164 -18412
rect 39060 -18492 39080 -18428
rect 39144 -18492 39164 -18428
rect 39060 -18508 39164 -18492
rect 39060 -18572 39080 -18508
rect 39144 -18572 39164 -18508
rect 39060 -18588 39164 -18572
rect 39060 -18652 39080 -18588
rect 39144 -18652 39164 -18588
rect 39060 -18668 39164 -18652
rect 39060 -18732 39080 -18668
rect 39144 -18732 39164 -18668
rect 39060 -18748 39164 -18732
rect 39060 -18812 39080 -18748
rect 39144 -18812 39164 -18748
rect 39060 -18828 39164 -18812
rect 39060 -18892 39080 -18828
rect 39144 -18892 39164 -18828
rect 39060 -18908 39164 -18892
rect 39060 -18972 39080 -18908
rect 39144 -18972 39164 -18908
rect 39060 -18988 39164 -18972
rect 39060 -19052 39080 -18988
rect 39144 -19052 39164 -18988
rect 39060 -19068 39164 -19052
rect 39060 -19132 39080 -19068
rect 39144 -19132 39164 -19068
rect 39060 -19148 39164 -19132
rect 39060 -19212 39080 -19148
rect 39144 -19212 39164 -19148
rect 39060 -19228 39164 -19212
rect 39060 -19292 39080 -19228
rect 39144 -19292 39164 -19228
rect 39060 -19308 39164 -19292
rect 39060 -19372 39080 -19308
rect 39144 -19372 39164 -19308
rect 39060 -19388 39164 -19372
rect 39060 -19452 39080 -19388
rect 39144 -19452 39164 -19388
rect 39060 -19468 39164 -19452
rect 39060 -19532 39080 -19468
rect 39144 -19532 39164 -19468
rect 39060 -19548 39164 -19532
rect 39060 -19612 39080 -19548
rect 39144 -19612 39164 -19548
rect 39060 -19628 39164 -19612
rect 39060 -19692 39080 -19628
rect 39144 -19692 39164 -19628
rect 39060 -19708 39164 -19692
rect 39060 -19772 39080 -19708
rect 39144 -19772 39164 -19708
rect 39060 -19788 39164 -19772
rect 39060 -19852 39080 -19788
rect 39144 -19852 39164 -19788
rect 39060 -19868 39164 -19852
rect 39060 -19932 39080 -19868
rect 39144 -19932 39164 -19868
rect 39060 -19948 39164 -19932
rect 39060 -20012 39080 -19948
rect 39144 -20012 39164 -19948
rect 39060 -20028 39164 -20012
rect 39060 -20092 39080 -20028
rect 39144 -20092 39164 -20028
rect 39060 -20108 39164 -20092
rect 39060 -20172 39080 -20108
rect 39144 -20172 39164 -20108
rect 39060 -20188 39164 -20172
rect 39060 -20252 39080 -20188
rect 39144 -20252 39164 -20188
rect 39060 -20268 39164 -20252
rect 39060 -20332 39080 -20268
rect 39144 -20332 39164 -20268
rect 39060 -20348 39164 -20332
rect 39060 -20412 39080 -20348
rect 39144 -20412 39164 -20348
rect 39060 -20428 39164 -20412
rect 39060 -20492 39080 -20428
rect 39144 -20492 39164 -20428
rect 39060 -20508 39164 -20492
rect 39060 -20572 39080 -20508
rect 39144 -20572 39164 -20508
rect 39060 -20588 39164 -20572
rect 39060 -20652 39080 -20588
rect 39144 -20652 39164 -20588
rect 39060 -20668 39164 -20652
rect 39060 -20732 39080 -20668
rect 39144 -20732 39164 -20668
rect 39060 -20748 39164 -20732
rect 39060 -20812 39080 -20748
rect 39144 -20812 39164 -20748
rect 39060 -20828 39164 -20812
rect 39060 -20892 39080 -20828
rect 39144 -20892 39164 -20828
rect 39060 -20908 39164 -20892
rect 39060 -20972 39080 -20908
rect 39144 -20972 39164 -20908
rect 39060 -20988 39164 -20972
rect 39060 -21052 39080 -20988
rect 39144 -21052 39164 -20988
rect 39060 -21068 39164 -21052
rect 33448 -21428 33552 -21132
rect 27836 -21508 27940 -21492
rect 27836 -21572 27856 -21508
rect 27920 -21572 27940 -21508
rect 27836 -21588 27940 -21572
rect 27836 -21652 27856 -21588
rect 27920 -21652 27940 -21588
rect 27836 -21668 27940 -21652
rect 27836 -21732 27856 -21668
rect 27920 -21732 27940 -21668
rect 27836 -21748 27940 -21732
rect 27836 -21812 27856 -21748
rect 27920 -21812 27940 -21748
rect 27836 -21828 27940 -21812
rect 27836 -21892 27856 -21828
rect 27920 -21892 27940 -21828
rect 27836 -21908 27940 -21892
rect 27836 -21972 27856 -21908
rect 27920 -21972 27940 -21908
rect 27836 -21988 27940 -21972
rect 27836 -22052 27856 -21988
rect 27920 -22052 27940 -21988
rect 27836 -22068 27940 -22052
rect 27836 -22132 27856 -22068
rect 27920 -22132 27940 -22068
rect 27836 -22148 27940 -22132
rect 27836 -22212 27856 -22148
rect 27920 -22212 27940 -22148
rect 27836 -22228 27940 -22212
rect 27836 -22292 27856 -22228
rect 27920 -22292 27940 -22228
rect 27836 -22308 27940 -22292
rect 27836 -22372 27856 -22308
rect 27920 -22372 27940 -22308
rect 27836 -22388 27940 -22372
rect 27836 -22452 27856 -22388
rect 27920 -22452 27940 -22388
rect 27836 -22468 27940 -22452
rect 27836 -22532 27856 -22468
rect 27920 -22532 27940 -22468
rect 27836 -22548 27940 -22532
rect 27836 -22612 27856 -22548
rect 27920 -22612 27940 -22548
rect 27836 -22628 27940 -22612
rect 27836 -22692 27856 -22628
rect 27920 -22692 27940 -22628
rect 27836 -22708 27940 -22692
rect 27836 -22772 27856 -22708
rect 27920 -22772 27940 -22708
rect 27836 -22788 27940 -22772
rect 27836 -22852 27856 -22788
rect 27920 -22852 27940 -22788
rect 27836 -22868 27940 -22852
rect 27836 -22932 27856 -22868
rect 27920 -22932 27940 -22868
rect 27836 -22948 27940 -22932
rect 27836 -23012 27856 -22948
rect 27920 -23012 27940 -22948
rect 27836 -23028 27940 -23012
rect 27836 -23092 27856 -23028
rect 27920 -23092 27940 -23028
rect 27836 -23108 27940 -23092
rect 27836 -23172 27856 -23108
rect 27920 -23172 27940 -23108
rect 27836 -23188 27940 -23172
rect 27836 -23252 27856 -23188
rect 27920 -23252 27940 -23188
rect 27836 -23268 27940 -23252
rect 27836 -23332 27856 -23268
rect 27920 -23332 27940 -23268
rect 27836 -23348 27940 -23332
rect 27836 -23412 27856 -23348
rect 27920 -23412 27940 -23348
rect 27836 -23428 27940 -23412
rect 27836 -23492 27856 -23428
rect 27920 -23492 27940 -23428
rect 27836 -23508 27940 -23492
rect 27836 -23572 27856 -23508
rect 27920 -23572 27940 -23508
rect 27836 -23588 27940 -23572
rect 27836 -23652 27856 -23588
rect 27920 -23652 27940 -23588
rect 27836 -23668 27940 -23652
rect 27836 -23732 27856 -23668
rect 27920 -23732 27940 -23668
rect 27836 -23748 27940 -23732
rect 27836 -23812 27856 -23748
rect 27920 -23812 27940 -23748
rect 27836 -23828 27940 -23812
rect 27836 -23892 27856 -23828
rect 27920 -23892 27940 -23828
rect 27836 -23908 27940 -23892
rect 27836 -23972 27856 -23908
rect 27920 -23972 27940 -23908
rect 27836 -23988 27940 -23972
rect 27836 -24052 27856 -23988
rect 27920 -24052 27940 -23988
rect 27836 -24068 27940 -24052
rect 27836 -24132 27856 -24068
rect 27920 -24132 27940 -24068
rect 27836 -24148 27940 -24132
rect 27836 -24212 27856 -24148
rect 27920 -24212 27940 -24148
rect 27836 -24228 27940 -24212
rect 27836 -24292 27856 -24228
rect 27920 -24292 27940 -24228
rect 27836 -24308 27940 -24292
rect 27836 -24372 27856 -24308
rect 27920 -24372 27940 -24308
rect 27836 -24388 27940 -24372
rect 27836 -24452 27856 -24388
rect 27920 -24452 27940 -24388
rect 27836 -24468 27940 -24452
rect 27836 -24532 27856 -24468
rect 27920 -24532 27940 -24468
rect 27836 -24548 27940 -24532
rect 27836 -24612 27856 -24548
rect 27920 -24612 27940 -24548
rect 27836 -24628 27940 -24612
rect 27836 -24692 27856 -24628
rect 27920 -24692 27940 -24628
rect 27836 -24708 27940 -24692
rect 27836 -24772 27856 -24708
rect 27920 -24772 27940 -24708
rect 27836 -24788 27940 -24772
rect 27836 -24852 27856 -24788
rect 27920 -24852 27940 -24788
rect 27836 -24868 27940 -24852
rect 27836 -24932 27856 -24868
rect 27920 -24932 27940 -24868
rect 27836 -24948 27940 -24932
rect 27836 -25012 27856 -24948
rect 27920 -25012 27940 -24948
rect 27836 -25028 27940 -25012
rect 27836 -25092 27856 -25028
rect 27920 -25092 27940 -25028
rect 27836 -25108 27940 -25092
rect 27836 -25172 27856 -25108
rect 27920 -25172 27940 -25108
rect 27836 -25188 27940 -25172
rect 27836 -25252 27856 -25188
rect 27920 -25252 27940 -25188
rect 27836 -25268 27940 -25252
rect 27836 -25332 27856 -25268
rect 27920 -25332 27940 -25268
rect 27836 -25348 27940 -25332
rect 27836 -25412 27856 -25348
rect 27920 -25412 27940 -25348
rect 27836 -25428 27940 -25412
rect 27836 -25492 27856 -25428
rect 27920 -25492 27940 -25428
rect 27836 -25508 27940 -25492
rect 27836 -25572 27856 -25508
rect 27920 -25572 27940 -25508
rect 27836 -25588 27940 -25572
rect 27836 -25652 27856 -25588
rect 27920 -25652 27940 -25588
rect 27836 -25668 27940 -25652
rect 27836 -25732 27856 -25668
rect 27920 -25732 27940 -25668
rect 27836 -25748 27940 -25732
rect 27836 -25812 27856 -25748
rect 27920 -25812 27940 -25748
rect 27836 -25828 27940 -25812
rect 27836 -25892 27856 -25828
rect 27920 -25892 27940 -25828
rect 27836 -25908 27940 -25892
rect 27836 -25972 27856 -25908
rect 27920 -25972 27940 -25908
rect 27836 -25988 27940 -25972
rect 27836 -26052 27856 -25988
rect 27920 -26052 27940 -25988
rect 27836 -26068 27940 -26052
rect 27836 -26132 27856 -26068
rect 27920 -26132 27940 -26068
rect 27836 -26148 27940 -26132
rect 27836 -26212 27856 -26148
rect 27920 -26212 27940 -26148
rect 27836 -26228 27940 -26212
rect 27836 -26292 27856 -26228
rect 27920 -26292 27940 -26228
rect 27836 -26308 27940 -26292
rect 27836 -26372 27856 -26308
rect 27920 -26372 27940 -26308
rect 27836 -26388 27940 -26372
rect 22224 -26748 22328 -26452
rect 16612 -26828 16716 -26812
rect 16612 -26892 16632 -26828
rect 16696 -26892 16716 -26828
rect 16612 -26908 16716 -26892
rect 16612 -26972 16632 -26908
rect 16696 -26972 16716 -26908
rect 16612 -26988 16716 -26972
rect 16612 -27052 16632 -26988
rect 16696 -27052 16716 -26988
rect 16612 -27068 16716 -27052
rect 16612 -27132 16632 -27068
rect 16696 -27132 16716 -27068
rect 16612 -27148 16716 -27132
rect 16612 -27212 16632 -27148
rect 16696 -27212 16716 -27148
rect 16612 -27228 16716 -27212
rect 16612 -27292 16632 -27228
rect 16696 -27292 16716 -27228
rect 16612 -27308 16716 -27292
rect 16612 -27372 16632 -27308
rect 16696 -27372 16716 -27308
rect 16612 -27388 16716 -27372
rect 16612 -27452 16632 -27388
rect 16696 -27452 16716 -27388
rect 16612 -27468 16716 -27452
rect 16612 -27532 16632 -27468
rect 16696 -27532 16716 -27468
rect 16612 -27548 16716 -27532
rect 16612 -27612 16632 -27548
rect 16696 -27612 16716 -27548
rect 16612 -27628 16716 -27612
rect 16612 -27692 16632 -27628
rect 16696 -27692 16716 -27628
rect 16612 -27708 16716 -27692
rect 16612 -27772 16632 -27708
rect 16696 -27772 16716 -27708
rect 16612 -27788 16716 -27772
rect 16612 -27852 16632 -27788
rect 16696 -27852 16716 -27788
rect 16612 -27868 16716 -27852
rect 16612 -27932 16632 -27868
rect 16696 -27932 16716 -27868
rect 16612 -27948 16716 -27932
rect 16612 -28012 16632 -27948
rect 16696 -28012 16716 -27948
rect 16612 -28028 16716 -28012
rect 16612 -28092 16632 -28028
rect 16696 -28092 16716 -28028
rect 16612 -28108 16716 -28092
rect 16612 -28172 16632 -28108
rect 16696 -28172 16716 -28108
rect 16612 -28188 16716 -28172
rect 16612 -28252 16632 -28188
rect 16696 -28252 16716 -28188
rect 16612 -28268 16716 -28252
rect 16612 -28332 16632 -28268
rect 16696 -28332 16716 -28268
rect 16612 -28348 16716 -28332
rect 16612 -28412 16632 -28348
rect 16696 -28412 16716 -28348
rect 16612 -28428 16716 -28412
rect 16612 -28492 16632 -28428
rect 16696 -28492 16716 -28428
rect 16612 -28508 16716 -28492
rect 16612 -28572 16632 -28508
rect 16696 -28572 16716 -28508
rect 16612 -28588 16716 -28572
rect 16612 -28652 16632 -28588
rect 16696 -28652 16716 -28588
rect 16612 -28668 16716 -28652
rect 16612 -28732 16632 -28668
rect 16696 -28732 16716 -28668
rect 16612 -28748 16716 -28732
rect 16612 -28812 16632 -28748
rect 16696 -28812 16716 -28748
rect 16612 -28828 16716 -28812
rect 16612 -28892 16632 -28828
rect 16696 -28892 16716 -28828
rect 16612 -28908 16716 -28892
rect 16612 -28972 16632 -28908
rect 16696 -28972 16716 -28908
rect 16612 -28988 16716 -28972
rect 16612 -29052 16632 -28988
rect 16696 -29052 16716 -28988
rect 16612 -29068 16716 -29052
rect 16612 -29132 16632 -29068
rect 16696 -29132 16716 -29068
rect 16612 -29148 16716 -29132
rect 16612 -29212 16632 -29148
rect 16696 -29212 16716 -29148
rect 16612 -29228 16716 -29212
rect 16612 -29292 16632 -29228
rect 16696 -29292 16716 -29228
rect 16612 -29308 16716 -29292
rect 16612 -29372 16632 -29308
rect 16696 -29372 16716 -29308
rect 16612 -29388 16716 -29372
rect 16612 -29452 16632 -29388
rect 16696 -29452 16716 -29388
rect 16612 -29468 16716 -29452
rect 16612 -29532 16632 -29468
rect 16696 -29532 16716 -29468
rect 16612 -29548 16716 -29532
rect 16612 -29612 16632 -29548
rect 16696 -29612 16716 -29548
rect 16612 -29628 16716 -29612
rect 16612 -29692 16632 -29628
rect 16696 -29692 16716 -29628
rect 16612 -29708 16716 -29692
rect 16612 -29772 16632 -29708
rect 16696 -29772 16716 -29708
rect 16612 -29788 16716 -29772
rect 16612 -29852 16632 -29788
rect 16696 -29852 16716 -29788
rect 16612 -29868 16716 -29852
rect 16612 -29932 16632 -29868
rect 16696 -29932 16716 -29868
rect 16612 -29948 16716 -29932
rect 16612 -30012 16632 -29948
rect 16696 -30012 16716 -29948
rect 16612 -30028 16716 -30012
rect 16612 -30092 16632 -30028
rect 16696 -30092 16716 -30028
rect 16612 -30108 16716 -30092
rect 16612 -30172 16632 -30108
rect 16696 -30172 16716 -30108
rect 16612 -30188 16716 -30172
rect 16612 -30252 16632 -30188
rect 16696 -30252 16716 -30188
rect 16612 -30268 16716 -30252
rect 16612 -30332 16632 -30268
rect 16696 -30332 16716 -30268
rect 16612 -30348 16716 -30332
rect 16612 -30412 16632 -30348
rect 16696 -30412 16716 -30348
rect 16612 -30428 16716 -30412
rect 16612 -30492 16632 -30428
rect 16696 -30492 16716 -30428
rect 16612 -30508 16716 -30492
rect 16612 -30572 16632 -30508
rect 16696 -30572 16716 -30508
rect 16612 -30588 16716 -30572
rect 16612 -30652 16632 -30588
rect 16696 -30652 16716 -30588
rect 16612 -30668 16716 -30652
rect 16612 -30732 16632 -30668
rect 16696 -30732 16716 -30668
rect 16612 -30748 16716 -30732
rect 16612 -30812 16632 -30748
rect 16696 -30812 16716 -30748
rect 16612 -30828 16716 -30812
rect 16612 -30892 16632 -30828
rect 16696 -30892 16716 -30828
rect 16612 -30908 16716 -30892
rect 16612 -30972 16632 -30908
rect 16696 -30972 16716 -30908
rect 16612 -30988 16716 -30972
rect 16612 -31052 16632 -30988
rect 16696 -31052 16716 -30988
rect 16612 -31068 16716 -31052
rect 16612 -31132 16632 -31068
rect 16696 -31132 16716 -31068
rect 16612 -31148 16716 -31132
rect 16612 -31212 16632 -31148
rect 16696 -31212 16716 -31148
rect 16612 -31228 16716 -31212
rect 16612 -31292 16632 -31228
rect 16696 -31292 16716 -31228
rect 16612 -31308 16716 -31292
rect 16612 -31372 16632 -31308
rect 16696 -31372 16716 -31308
rect 16612 -31388 16716 -31372
rect 16612 -31452 16632 -31388
rect 16696 -31452 16716 -31388
rect 16612 -31468 16716 -31452
rect 16612 -31532 16632 -31468
rect 16696 -31532 16716 -31468
rect 16612 -31548 16716 -31532
rect 16612 -31612 16632 -31548
rect 16696 -31612 16716 -31548
rect 16612 -31628 16716 -31612
rect 16612 -31692 16632 -31628
rect 16696 -31692 16716 -31628
rect 16612 -31708 16716 -31692
rect 11000 -32068 11104 -31772
rect 5388 -32148 5492 -32132
rect 5388 -32212 5408 -32148
rect 5472 -32212 5492 -32148
rect 5388 -32228 5492 -32212
rect 5388 -32292 5408 -32228
rect 5472 -32292 5492 -32228
rect 5388 -32308 5492 -32292
rect 5388 -32372 5408 -32308
rect 5472 -32372 5492 -32308
rect 5388 -32388 5492 -32372
rect 5388 -32452 5408 -32388
rect 5472 -32452 5492 -32388
rect 5388 -32468 5492 -32452
rect 5388 -32532 5408 -32468
rect 5472 -32532 5492 -32468
rect 5388 -32548 5492 -32532
rect 5388 -32612 5408 -32548
rect 5472 -32612 5492 -32548
rect 5388 -32628 5492 -32612
rect 5388 -32692 5408 -32628
rect 5472 -32692 5492 -32628
rect 5388 -32708 5492 -32692
rect 5388 -32772 5408 -32708
rect 5472 -32772 5492 -32708
rect 5388 -32788 5492 -32772
rect 5388 -32852 5408 -32788
rect 5472 -32852 5492 -32788
rect 5388 -32868 5492 -32852
rect 5388 -32932 5408 -32868
rect 5472 -32932 5492 -32868
rect 5388 -32948 5492 -32932
rect 5388 -33012 5408 -32948
rect 5472 -33012 5492 -32948
rect 5388 -33028 5492 -33012
rect 5388 -33092 5408 -33028
rect 5472 -33092 5492 -33028
rect 5388 -33108 5492 -33092
rect 5388 -33172 5408 -33108
rect 5472 -33172 5492 -33108
rect 5388 -33188 5492 -33172
rect 5388 -33252 5408 -33188
rect 5472 -33252 5492 -33188
rect 5388 -33268 5492 -33252
rect 5388 -33332 5408 -33268
rect 5472 -33332 5492 -33268
rect 5388 -33348 5492 -33332
rect 5388 -33412 5408 -33348
rect 5472 -33412 5492 -33348
rect 5388 -33428 5492 -33412
rect 5388 -33492 5408 -33428
rect 5472 -33492 5492 -33428
rect 5388 -33508 5492 -33492
rect 5388 -33572 5408 -33508
rect 5472 -33572 5492 -33508
rect 5388 -33588 5492 -33572
rect 5388 -33652 5408 -33588
rect 5472 -33652 5492 -33588
rect 5388 -33668 5492 -33652
rect 5388 -33732 5408 -33668
rect 5472 -33732 5492 -33668
rect 5388 -33748 5492 -33732
rect 5388 -33812 5408 -33748
rect 5472 -33812 5492 -33748
rect 5388 -33828 5492 -33812
rect 5388 -33892 5408 -33828
rect 5472 -33892 5492 -33828
rect 5388 -33908 5492 -33892
rect 5388 -33972 5408 -33908
rect 5472 -33972 5492 -33908
rect 5388 -33988 5492 -33972
rect 5388 -34052 5408 -33988
rect 5472 -34052 5492 -33988
rect 5388 -34068 5492 -34052
rect 5388 -34132 5408 -34068
rect 5472 -34132 5492 -34068
rect 5388 -34148 5492 -34132
rect 5388 -34212 5408 -34148
rect 5472 -34212 5492 -34148
rect 5388 -34228 5492 -34212
rect 5388 -34292 5408 -34228
rect 5472 -34292 5492 -34228
rect 5388 -34308 5492 -34292
rect 5388 -34372 5408 -34308
rect 5472 -34372 5492 -34308
rect 5388 -34388 5492 -34372
rect 5388 -34452 5408 -34388
rect 5472 -34452 5492 -34388
rect 5388 -34468 5492 -34452
rect 5388 -34532 5408 -34468
rect 5472 -34532 5492 -34468
rect 5388 -34548 5492 -34532
rect 5388 -34612 5408 -34548
rect 5472 -34612 5492 -34548
rect 5388 -34628 5492 -34612
rect 5388 -34692 5408 -34628
rect 5472 -34692 5492 -34628
rect 5388 -34708 5492 -34692
rect 5388 -34772 5408 -34708
rect 5472 -34772 5492 -34708
rect 5388 -34788 5492 -34772
rect 5388 -34852 5408 -34788
rect 5472 -34852 5492 -34788
rect 5388 -34868 5492 -34852
rect 5388 -34932 5408 -34868
rect 5472 -34932 5492 -34868
rect 5388 -34948 5492 -34932
rect 5388 -35012 5408 -34948
rect 5472 -35012 5492 -34948
rect 5388 -35028 5492 -35012
rect 5388 -35092 5408 -35028
rect 5472 -35092 5492 -35028
rect 5388 -35108 5492 -35092
rect 5388 -35172 5408 -35108
rect 5472 -35172 5492 -35108
rect 5388 -35188 5492 -35172
rect 5388 -35252 5408 -35188
rect 5472 -35252 5492 -35188
rect 5388 -35268 5492 -35252
rect 5388 -35332 5408 -35268
rect 5472 -35332 5492 -35268
rect 5388 -35348 5492 -35332
rect 5388 -35412 5408 -35348
rect 5472 -35412 5492 -35348
rect 5388 -35428 5492 -35412
rect 5388 -35492 5408 -35428
rect 5472 -35492 5492 -35428
rect 5388 -35508 5492 -35492
rect 5388 -35572 5408 -35508
rect 5472 -35572 5492 -35508
rect 5388 -35588 5492 -35572
rect 5388 -35652 5408 -35588
rect 5472 -35652 5492 -35588
rect 5388 -35668 5492 -35652
rect 5388 -35732 5408 -35668
rect 5472 -35732 5492 -35668
rect 5388 -35748 5492 -35732
rect 5388 -35812 5408 -35748
rect 5472 -35812 5492 -35748
rect 5388 -35828 5492 -35812
rect 5388 -35892 5408 -35828
rect 5472 -35892 5492 -35828
rect 5388 -35908 5492 -35892
rect 5388 -35972 5408 -35908
rect 5472 -35972 5492 -35908
rect 5388 -35988 5492 -35972
rect 5388 -36052 5408 -35988
rect 5472 -36052 5492 -35988
rect 5388 -36068 5492 -36052
rect 5388 -36132 5408 -36068
rect 5472 -36132 5492 -36068
rect 5388 -36148 5492 -36132
rect 5388 -36212 5408 -36148
rect 5472 -36212 5492 -36148
rect 5388 -36228 5492 -36212
rect 5388 -36292 5408 -36228
rect 5472 -36292 5492 -36228
rect 5388 -36308 5492 -36292
rect 5388 -36372 5408 -36308
rect 5472 -36372 5492 -36308
rect 5388 -36388 5492 -36372
rect 5388 -36452 5408 -36388
rect 5472 -36452 5492 -36388
rect 5388 -36468 5492 -36452
rect 5388 -36532 5408 -36468
rect 5472 -36532 5492 -36468
rect 5388 -36548 5492 -36532
rect 5388 -36612 5408 -36548
rect 5472 -36612 5492 -36548
rect 5388 -36628 5492 -36612
rect 5388 -36692 5408 -36628
rect 5472 -36692 5492 -36628
rect 5388 -36708 5492 -36692
rect 5388 -36772 5408 -36708
rect 5472 -36772 5492 -36708
rect 5388 -36788 5492 -36772
rect 5388 -36852 5408 -36788
rect 5472 -36852 5492 -36788
rect 5388 -36868 5492 -36852
rect 5388 -36932 5408 -36868
rect 5472 -36932 5492 -36868
rect 5388 -36948 5492 -36932
rect 5388 -37012 5408 -36948
rect 5472 -37012 5492 -36948
rect 5388 -37028 5492 -37012
rect -224 -37240 -120 -37092
rect 2608 -37240 2712 -37041
rect 5388 -37092 5408 -37028
rect 5472 -37092 5492 -37028
rect 5811 -32148 10733 -32119
rect 5811 -37012 5840 -32148
rect 10704 -37012 10733 -32148
rect 5811 -37041 10733 -37012
rect 11000 -32132 11020 -32068
rect 11084 -32132 11104 -32068
rect 13832 -32119 13936 -31721
rect 16612 -31772 16632 -31708
rect 16696 -31772 16716 -31708
rect 17035 -26828 21957 -26799
rect 17035 -31692 17064 -26828
rect 21928 -31692 21957 -26828
rect 17035 -31721 21957 -31692
rect 22224 -26812 22244 -26748
rect 22308 -26812 22328 -26748
rect 25056 -26799 25160 -26401
rect 27836 -26452 27856 -26388
rect 27920 -26452 27940 -26388
rect 28259 -21508 33181 -21479
rect 28259 -26372 28288 -21508
rect 33152 -26372 33181 -21508
rect 28259 -26401 33181 -26372
rect 33448 -21492 33468 -21428
rect 33532 -21492 33552 -21428
rect 36280 -21479 36384 -21081
rect 39060 -21132 39080 -21068
rect 39144 -21132 39164 -21068
rect 39060 -21428 39164 -21132
rect 33448 -21508 33552 -21492
rect 33448 -21572 33468 -21508
rect 33532 -21572 33552 -21508
rect 33448 -21588 33552 -21572
rect 33448 -21652 33468 -21588
rect 33532 -21652 33552 -21588
rect 33448 -21668 33552 -21652
rect 33448 -21732 33468 -21668
rect 33532 -21732 33552 -21668
rect 33448 -21748 33552 -21732
rect 33448 -21812 33468 -21748
rect 33532 -21812 33552 -21748
rect 33448 -21828 33552 -21812
rect 33448 -21892 33468 -21828
rect 33532 -21892 33552 -21828
rect 33448 -21908 33552 -21892
rect 33448 -21972 33468 -21908
rect 33532 -21972 33552 -21908
rect 33448 -21988 33552 -21972
rect 33448 -22052 33468 -21988
rect 33532 -22052 33552 -21988
rect 33448 -22068 33552 -22052
rect 33448 -22132 33468 -22068
rect 33532 -22132 33552 -22068
rect 33448 -22148 33552 -22132
rect 33448 -22212 33468 -22148
rect 33532 -22212 33552 -22148
rect 33448 -22228 33552 -22212
rect 33448 -22292 33468 -22228
rect 33532 -22292 33552 -22228
rect 33448 -22308 33552 -22292
rect 33448 -22372 33468 -22308
rect 33532 -22372 33552 -22308
rect 33448 -22388 33552 -22372
rect 33448 -22452 33468 -22388
rect 33532 -22452 33552 -22388
rect 33448 -22468 33552 -22452
rect 33448 -22532 33468 -22468
rect 33532 -22532 33552 -22468
rect 33448 -22548 33552 -22532
rect 33448 -22612 33468 -22548
rect 33532 -22612 33552 -22548
rect 33448 -22628 33552 -22612
rect 33448 -22692 33468 -22628
rect 33532 -22692 33552 -22628
rect 33448 -22708 33552 -22692
rect 33448 -22772 33468 -22708
rect 33532 -22772 33552 -22708
rect 33448 -22788 33552 -22772
rect 33448 -22852 33468 -22788
rect 33532 -22852 33552 -22788
rect 33448 -22868 33552 -22852
rect 33448 -22932 33468 -22868
rect 33532 -22932 33552 -22868
rect 33448 -22948 33552 -22932
rect 33448 -23012 33468 -22948
rect 33532 -23012 33552 -22948
rect 33448 -23028 33552 -23012
rect 33448 -23092 33468 -23028
rect 33532 -23092 33552 -23028
rect 33448 -23108 33552 -23092
rect 33448 -23172 33468 -23108
rect 33532 -23172 33552 -23108
rect 33448 -23188 33552 -23172
rect 33448 -23252 33468 -23188
rect 33532 -23252 33552 -23188
rect 33448 -23268 33552 -23252
rect 33448 -23332 33468 -23268
rect 33532 -23332 33552 -23268
rect 33448 -23348 33552 -23332
rect 33448 -23412 33468 -23348
rect 33532 -23412 33552 -23348
rect 33448 -23428 33552 -23412
rect 33448 -23492 33468 -23428
rect 33532 -23492 33552 -23428
rect 33448 -23508 33552 -23492
rect 33448 -23572 33468 -23508
rect 33532 -23572 33552 -23508
rect 33448 -23588 33552 -23572
rect 33448 -23652 33468 -23588
rect 33532 -23652 33552 -23588
rect 33448 -23668 33552 -23652
rect 33448 -23732 33468 -23668
rect 33532 -23732 33552 -23668
rect 33448 -23748 33552 -23732
rect 33448 -23812 33468 -23748
rect 33532 -23812 33552 -23748
rect 33448 -23828 33552 -23812
rect 33448 -23892 33468 -23828
rect 33532 -23892 33552 -23828
rect 33448 -23908 33552 -23892
rect 33448 -23972 33468 -23908
rect 33532 -23972 33552 -23908
rect 33448 -23988 33552 -23972
rect 33448 -24052 33468 -23988
rect 33532 -24052 33552 -23988
rect 33448 -24068 33552 -24052
rect 33448 -24132 33468 -24068
rect 33532 -24132 33552 -24068
rect 33448 -24148 33552 -24132
rect 33448 -24212 33468 -24148
rect 33532 -24212 33552 -24148
rect 33448 -24228 33552 -24212
rect 33448 -24292 33468 -24228
rect 33532 -24292 33552 -24228
rect 33448 -24308 33552 -24292
rect 33448 -24372 33468 -24308
rect 33532 -24372 33552 -24308
rect 33448 -24388 33552 -24372
rect 33448 -24452 33468 -24388
rect 33532 -24452 33552 -24388
rect 33448 -24468 33552 -24452
rect 33448 -24532 33468 -24468
rect 33532 -24532 33552 -24468
rect 33448 -24548 33552 -24532
rect 33448 -24612 33468 -24548
rect 33532 -24612 33552 -24548
rect 33448 -24628 33552 -24612
rect 33448 -24692 33468 -24628
rect 33532 -24692 33552 -24628
rect 33448 -24708 33552 -24692
rect 33448 -24772 33468 -24708
rect 33532 -24772 33552 -24708
rect 33448 -24788 33552 -24772
rect 33448 -24852 33468 -24788
rect 33532 -24852 33552 -24788
rect 33448 -24868 33552 -24852
rect 33448 -24932 33468 -24868
rect 33532 -24932 33552 -24868
rect 33448 -24948 33552 -24932
rect 33448 -25012 33468 -24948
rect 33532 -25012 33552 -24948
rect 33448 -25028 33552 -25012
rect 33448 -25092 33468 -25028
rect 33532 -25092 33552 -25028
rect 33448 -25108 33552 -25092
rect 33448 -25172 33468 -25108
rect 33532 -25172 33552 -25108
rect 33448 -25188 33552 -25172
rect 33448 -25252 33468 -25188
rect 33532 -25252 33552 -25188
rect 33448 -25268 33552 -25252
rect 33448 -25332 33468 -25268
rect 33532 -25332 33552 -25268
rect 33448 -25348 33552 -25332
rect 33448 -25412 33468 -25348
rect 33532 -25412 33552 -25348
rect 33448 -25428 33552 -25412
rect 33448 -25492 33468 -25428
rect 33532 -25492 33552 -25428
rect 33448 -25508 33552 -25492
rect 33448 -25572 33468 -25508
rect 33532 -25572 33552 -25508
rect 33448 -25588 33552 -25572
rect 33448 -25652 33468 -25588
rect 33532 -25652 33552 -25588
rect 33448 -25668 33552 -25652
rect 33448 -25732 33468 -25668
rect 33532 -25732 33552 -25668
rect 33448 -25748 33552 -25732
rect 33448 -25812 33468 -25748
rect 33532 -25812 33552 -25748
rect 33448 -25828 33552 -25812
rect 33448 -25892 33468 -25828
rect 33532 -25892 33552 -25828
rect 33448 -25908 33552 -25892
rect 33448 -25972 33468 -25908
rect 33532 -25972 33552 -25908
rect 33448 -25988 33552 -25972
rect 33448 -26052 33468 -25988
rect 33532 -26052 33552 -25988
rect 33448 -26068 33552 -26052
rect 33448 -26132 33468 -26068
rect 33532 -26132 33552 -26068
rect 33448 -26148 33552 -26132
rect 33448 -26212 33468 -26148
rect 33532 -26212 33552 -26148
rect 33448 -26228 33552 -26212
rect 33448 -26292 33468 -26228
rect 33532 -26292 33552 -26228
rect 33448 -26308 33552 -26292
rect 33448 -26372 33468 -26308
rect 33532 -26372 33552 -26308
rect 33448 -26388 33552 -26372
rect 27836 -26748 27940 -26452
rect 22224 -26828 22328 -26812
rect 22224 -26892 22244 -26828
rect 22308 -26892 22328 -26828
rect 22224 -26908 22328 -26892
rect 22224 -26972 22244 -26908
rect 22308 -26972 22328 -26908
rect 22224 -26988 22328 -26972
rect 22224 -27052 22244 -26988
rect 22308 -27052 22328 -26988
rect 22224 -27068 22328 -27052
rect 22224 -27132 22244 -27068
rect 22308 -27132 22328 -27068
rect 22224 -27148 22328 -27132
rect 22224 -27212 22244 -27148
rect 22308 -27212 22328 -27148
rect 22224 -27228 22328 -27212
rect 22224 -27292 22244 -27228
rect 22308 -27292 22328 -27228
rect 22224 -27308 22328 -27292
rect 22224 -27372 22244 -27308
rect 22308 -27372 22328 -27308
rect 22224 -27388 22328 -27372
rect 22224 -27452 22244 -27388
rect 22308 -27452 22328 -27388
rect 22224 -27468 22328 -27452
rect 22224 -27532 22244 -27468
rect 22308 -27532 22328 -27468
rect 22224 -27548 22328 -27532
rect 22224 -27612 22244 -27548
rect 22308 -27612 22328 -27548
rect 22224 -27628 22328 -27612
rect 22224 -27692 22244 -27628
rect 22308 -27692 22328 -27628
rect 22224 -27708 22328 -27692
rect 22224 -27772 22244 -27708
rect 22308 -27772 22328 -27708
rect 22224 -27788 22328 -27772
rect 22224 -27852 22244 -27788
rect 22308 -27852 22328 -27788
rect 22224 -27868 22328 -27852
rect 22224 -27932 22244 -27868
rect 22308 -27932 22328 -27868
rect 22224 -27948 22328 -27932
rect 22224 -28012 22244 -27948
rect 22308 -28012 22328 -27948
rect 22224 -28028 22328 -28012
rect 22224 -28092 22244 -28028
rect 22308 -28092 22328 -28028
rect 22224 -28108 22328 -28092
rect 22224 -28172 22244 -28108
rect 22308 -28172 22328 -28108
rect 22224 -28188 22328 -28172
rect 22224 -28252 22244 -28188
rect 22308 -28252 22328 -28188
rect 22224 -28268 22328 -28252
rect 22224 -28332 22244 -28268
rect 22308 -28332 22328 -28268
rect 22224 -28348 22328 -28332
rect 22224 -28412 22244 -28348
rect 22308 -28412 22328 -28348
rect 22224 -28428 22328 -28412
rect 22224 -28492 22244 -28428
rect 22308 -28492 22328 -28428
rect 22224 -28508 22328 -28492
rect 22224 -28572 22244 -28508
rect 22308 -28572 22328 -28508
rect 22224 -28588 22328 -28572
rect 22224 -28652 22244 -28588
rect 22308 -28652 22328 -28588
rect 22224 -28668 22328 -28652
rect 22224 -28732 22244 -28668
rect 22308 -28732 22328 -28668
rect 22224 -28748 22328 -28732
rect 22224 -28812 22244 -28748
rect 22308 -28812 22328 -28748
rect 22224 -28828 22328 -28812
rect 22224 -28892 22244 -28828
rect 22308 -28892 22328 -28828
rect 22224 -28908 22328 -28892
rect 22224 -28972 22244 -28908
rect 22308 -28972 22328 -28908
rect 22224 -28988 22328 -28972
rect 22224 -29052 22244 -28988
rect 22308 -29052 22328 -28988
rect 22224 -29068 22328 -29052
rect 22224 -29132 22244 -29068
rect 22308 -29132 22328 -29068
rect 22224 -29148 22328 -29132
rect 22224 -29212 22244 -29148
rect 22308 -29212 22328 -29148
rect 22224 -29228 22328 -29212
rect 22224 -29292 22244 -29228
rect 22308 -29292 22328 -29228
rect 22224 -29308 22328 -29292
rect 22224 -29372 22244 -29308
rect 22308 -29372 22328 -29308
rect 22224 -29388 22328 -29372
rect 22224 -29452 22244 -29388
rect 22308 -29452 22328 -29388
rect 22224 -29468 22328 -29452
rect 22224 -29532 22244 -29468
rect 22308 -29532 22328 -29468
rect 22224 -29548 22328 -29532
rect 22224 -29612 22244 -29548
rect 22308 -29612 22328 -29548
rect 22224 -29628 22328 -29612
rect 22224 -29692 22244 -29628
rect 22308 -29692 22328 -29628
rect 22224 -29708 22328 -29692
rect 22224 -29772 22244 -29708
rect 22308 -29772 22328 -29708
rect 22224 -29788 22328 -29772
rect 22224 -29852 22244 -29788
rect 22308 -29852 22328 -29788
rect 22224 -29868 22328 -29852
rect 22224 -29932 22244 -29868
rect 22308 -29932 22328 -29868
rect 22224 -29948 22328 -29932
rect 22224 -30012 22244 -29948
rect 22308 -30012 22328 -29948
rect 22224 -30028 22328 -30012
rect 22224 -30092 22244 -30028
rect 22308 -30092 22328 -30028
rect 22224 -30108 22328 -30092
rect 22224 -30172 22244 -30108
rect 22308 -30172 22328 -30108
rect 22224 -30188 22328 -30172
rect 22224 -30252 22244 -30188
rect 22308 -30252 22328 -30188
rect 22224 -30268 22328 -30252
rect 22224 -30332 22244 -30268
rect 22308 -30332 22328 -30268
rect 22224 -30348 22328 -30332
rect 22224 -30412 22244 -30348
rect 22308 -30412 22328 -30348
rect 22224 -30428 22328 -30412
rect 22224 -30492 22244 -30428
rect 22308 -30492 22328 -30428
rect 22224 -30508 22328 -30492
rect 22224 -30572 22244 -30508
rect 22308 -30572 22328 -30508
rect 22224 -30588 22328 -30572
rect 22224 -30652 22244 -30588
rect 22308 -30652 22328 -30588
rect 22224 -30668 22328 -30652
rect 22224 -30732 22244 -30668
rect 22308 -30732 22328 -30668
rect 22224 -30748 22328 -30732
rect 22224 -30812 22244 -30748
rect 22308 -30812 22328 -30748
rect 22224 -30828 22328 -30812
rect 22224 -30892 22244 -30828
rect 22308 -30892 22328 -30828
rect 22224 -30908 22328 -30892
rect 22224 -30972 22244 -30908
rect 22308 -30972 22328 -30908
rect 22224 -30988 22328 -30972
rect 22224 -31052 22244 -30988
rect 22308 -31052 22328 -30988
rect 22224 -31068 22328 -31052
rect 22224 -31132 22244 -31068
rect 22308 -31132 22328 -31068
rect 22224 -31148 22328 -31132
rect 22224 -31212 22244 -31148
rect 22308 -31212 22328 -31148
rect 22224 -31228 22328 -31212
rect 22224 -31292 22244 -31228
rect 22308 -31292 22328 -31228
rect 22224 -31308 22328 -31292
rect 22224 -31372 22244 -31308
rect 22308 -31372 22328 -31308
rect 22224 -31388 22328 -31372
rect 22224 -31452 22244 -31388
rect 22308 -31452 22328 -31388
rect 22224 -31468 22328 -31452
rect 22224 -31532 22244 -31468
rect 22308 -31532 22328 -31468
rect 22224 -31548 22328 -31532
rect 22224 -31612 22244 -31548
rect 22308 -31612 22328 -31548
rect 22224 -31628 22328 -31612
rect 22224 -31692 22244 -31628
rect 22308 -31692 22328 -31628
rect 22224 -31708 22328 -31692
rect 16612 -32068 16716 -31772
rect 11000 -32148 11104 -32132
rect 11000 -32212 11020 -32148
rect 11084 -32212 11104 -32148
rect 11000 -32228 11104 -32212
rect 11000 -32292 11020 -32228
rect 11084 -32292 11104 -32228
rect 11000 -32308 11104 -32292
rect 11000 -32372 11020 -32308
rect 11084 -32372 11104 -32308
rect 11000 -32388 11104 -32372
rect 11000 -32452 11020 -32388
rect 11084 -32452 11104 -32388
rect 11000 -32468 11104 -32452
rect 11000 -32532 11020 -32468
rect 11084 -32532 11104 -32468
rect 11000 -32548 11104 -32532
rect 11000 -32612 11020 -32548
rect 11084 -32612 11104 -32548
rect 11000 -32628 11104 -32612
rect 11000 -32692 11020 -32628
rect 11084 -32692 11104 -32628
rect 11000 -32708 11104 -32692
rect 11000 -32772 11020 -32708
rect 11084 -32772 11104 -32708
rect 11000 -32788 11104 -32772
rect 11000 -32852 11020 -32788
rect 11084 -32852 11104 -32788
rect 11000 -32868 11104 -32852
rect 11000 -32932 11020 -32868
rect 11084 -32932 11104 -32868
rect 11000 -32948 11104 -32932
rect 11000 -33012 11020 -32948
rect 11084 -33012 11104 -32948
rect 11000 -33028 11104 -33012
rect 11000 -33092 11020 -33028
rect 11084 -33092 11104 -33028
rect 11000 -33108 11104 -33092
rect 11000 -33172 11020 -33108
rect 11084 -33172 11104 -33108
rect 11000 -33188 11104 -33172
rect 11000 -33252 11020 -33188
rect 11084 -33252 11104 -33188
rect 11000 -33268 11104 -33252
rect 11000 -33332 11020 -33268
rect 11084 -33332 11104 -33268
rect 11000 -33348 11104 -33332
rect 11000 -33412 11020 -33348
rect 11084 -33412 11104 -33348
rect 11000 -33428 11104 -33412
rect 11000 -33492 11020 -33428
rect 11084 -33492 11104 -33428
rect 11000 -33508 11104 -33492
rect 11000 -33572 11020 -33508
rect 11084 -33572 11104 -33508
rect 11000 -33588 11104 -33572
rect 11000 -33652 11020 -33588
rect 11084 -33652 11104 -33588
rect 11000 -33668 11104 -33652
rect 11000 -33732 11020 -33668
rect 11084 -33732 11104 -33668
rect 11000 -33748 11104 -33732
rect 11000 -33812 11020 -33748
rect 11084 -33812 11104 -33748
rect 11000 -33828 11104 -33812
rect 11000 -33892 11020 -33828
rect 11084 -33892 11104 -33828
rect 11000 -33908 11104 -33892
rect 11000 -33972 11020 -33908
rect 11084 -33972 11104 -33908
rect 11000 -33988 11104 -33972
rect 11000 -34052 11020 -33988
rect 11084 -34052 11104 -33988
rect 11000 -34068 11104 -34052
rect 11000 -34132 11020 -34068
rect 11084 -34132 11104 -34068
rect 11000 -34148 11104 -34132
rect 11000 -34212 11020 -34148
rect 11084 -34212 11104 -34148
rect 11000 -34228 11104 -34212
rect 11000 -34292 11020 -34228
rect 11084 -34292 11104 -34228
rect 11000 -34308 11104 -34292
rect 11000 -34372 11020 -34308
rect 11084 -34372 11104 -34308
rect 11000 -34388 11104 -34372
rect 11000 -34452 11020 -34388
rect 11084 -34452 11104 -34388
rect 11000 -34468 11104 -34452
rect 11000 -34532 11020 -34468
rect 11084 -34532 11104 -34468
rect 11000 -34548 11104 -34532
rect 11000 -34612 11020 -34548
rect 11084 -34612 11104 -34548
rect 11000 -34628 11104 -34612
rect 11000 -34692 11020 -34628
rect 11084 -34692 11104 -34628
rect 11000 -34708 11104 -34692
rect 11000 -34772 11020 -34708
rect 11084 -34772 11104 -34708
rect 11000 -34788 11104 -34772
rect 11000 -34852 11020 -34788
rect 11084 -34852 11104 -34788
rect 11000 -34868 11104 -34852
rect 11000 -34932 11020 -34868
rect 11084 -34932 11104 -34868
rect 11000 -34948 11104 -34932
rect 11000 -35012 11020 -34948
rect 11084 -35012 11104 -34948
rect 11000 -35028 11104 -35012
rect 11000 -35092 11020 -35028
rect 11084 -35092 11104 -35028
rect 11000 -35108 11104 -35092
rect 11000 -35172 11020 -35108
rect 11084 -35172 11104 -35108
rect 11000 -35188 11104 -35172
rect 11000 -35252 11020 -35188
rect 11084 -35252 11104 -35188
rect 11000 -35268 11104 -35252
rect 11000 -35332 11020 -35268
rect 11084 -35332 11104 -35268
rect 11000 -35348 11104 -35332
rect 11000 -35412 11020 -35348
rect 11084 -35412 11104 -35348
rect 11000 -35428 11104 -35412
rect 11000 -35492 11020 -35428
rect 11084 -35492 11104 -35428
rect 11000 -35508 11104 -35492
rect 11000 -35572 11020 -35508
rect 11084 -35572 11104 -35508
rect 11000 -35588 11104 -35572
rect 11000 -35652 11020 -35588
rect 11084 -35652 11104 -35588
rect 11000 -35668 11104 -35652
rect 11000 -35732 11020 -35668
rect 11084 -35732 11104 -35668
rect 11000 -35748 11104 -35732
rect 11000 -35812 11020 -35748
rect 11084 -35812 11104 -35748
rect 11000 -35828 11104 -35812
rect 11000 -35892 11020 -35828
rect 11084 -35892 11104 -35828
rect 11000 -35908 11104 -35892
rect 11000 -35972 11020 -35908
rect 11084 -35972 11104 -35908
rect 11000 -35988 11104 -35972
rect 11000 -36052 11020 -35988
rect 11084 -36052 11104 -35988
rect 11000 -36068 11104 -36052
rect 11000 -36132 11020 -36068
rect 11084 -36132 11104 -36068
rect 11000 -36148 11104 -36132
rect 11000 -36212 11020 -36148
rect 11084 -36212 11104 -36148
rect 11000 -36228 11104 -36212
rect 11000 -36292 11020 -36228
rect 11084 -36292 11104 -36228
rect 11000 -36308 11104 -36292
rect 11000 -36372 11020 -36308
rect 11084 -36372 11104 -36308
rect 11000 -36388 11104 -36372
rect 11000 -36452 11020 -36388
rect 11084 -36452 11104 -36388
rect 11000 -36468 11104 -36452
rect 11000 -36532 11020 -36468
rect 11084 -36532 11104 -36468
rect 11000 -36548 11104 -36532
rect 11000 -36612 11020 -36548
rect 11084 -36612 11104 -36548
rect 11000 -36628 11104 -36612
rect 11000 -36692 11020 -36628
rect 11084 -36692 11104 -36628
rect 11000 -36708 11104 -36692
rect 11000 -36772 11020 -36708
rect 11084 -36772 11104 -36708
rect 11000 -36788 11104 -36772
rect 11000 -36852 11020 -36788
rect 11084 -36852 11104 -36788
rect 11000 -36868 11104 -36852
rect 11000 -36932 11020 -36868
rect 11084 -36932 11104 -36868
rect 11000 -36948 11104 -36932
rect 11000 -37012 11020 -36948
rect 11084 -37012 11104 -36948
rect 11000 -37028 11104 -37012
rect 5388 -37240 5492 -37092
rect 8220 -37240 8324 -37041
rect 11000 -37092 11020 -37028
rect 11084 -37092 11104 -37028
rect 11423 -32148 16345 -32119
rect 11423 -37012 11452 -32148
rect 16316 -37012 16345 -32148
rect 11423 -37041 16345 -37012
rect 16612 -32132 16632 -32068
rect 16696 -32132 16716 -32068
rect 19444 -32119 19548 -31721
rect 22224 -31772 22244 -31708
rect 22308 -31772 22328 -31708
rect 22647 -26828 27569 -26799
rect 22647 -31692 22676 -26828
rect 27540 -31692 27569 -26828
rect 22647 -31721 27569 -31692
rect 27836 -26812 27856 -26748
rect 27920 -26812 27940 -26748
rect 30668 -26799 30772 -26401
rect 33448 -26452 33468 -26388
rect 33532 -26452 33552 -26388
rect 33871 -21508 38793 -21479
rect 33871 -26372 33900 -21508
rect 38764 -26372 38793 -21508
rect 33871 -26401 38793 -26372
rect 39060 -21492 39080 -21428
rect 39144 -21492 39164 -21428
rect 39060 -21508 39164 -21492
rect 39060 -21572 39080 -21508
rect 39144 -21572 39164 -21508
rect 39060 -21588 39164 -21572
rect 39060 -21652 39080 -21588
rect 39144 -21652 39164 -21588
rect 39060 -21668 39164 -21652
rect 39060 -21732 39080 -21668
rect 39144 -21732 39164 -21668
rect 39060 -21748 39164 -21732
rect 39060 -21812 39080 -21748
rect 39144 -21812 39164 -21748
rect 39060 -21828 39164 -21812
rect 39060 -21892 39080 -21828
rect 39144 -21892 39164 -21828
rect 39060 -21908 39164 -21892
rect 39060 -21972 39080 -21908
rect 39144 -21972 39164 -21908
rect 39060 -21988 39164 -21972
rect 39060 -22052 39080 -21988
rect 39144 -22052 39164 -21988
rect 39060 -22068 39164 -22052
rect 39060 -22132 39080 -22068
rect 39144 -22132 39164 -22068
rect 39060 -22148 39164 -22132
rect 39060 -22212 39080 -22148
rect 39144 -22212 39164 -22148
rect 39060 -22228 39164 -22212
rect 39060 -22292 39080 -22228
rect 39144 -22292 39164 -22228
rect 39060 -22308 39164 -22292
rect 39060 -22372 39080 -22308
rect 39144 -22372 39164 -22308
rect 39060 -22388 39164 -22372
rect 39060 -22452 39080 -22388
rect 39144 -22452 39164 -22388
rect 39060 -22468 39164 -22452
rect 39060 -22532 39080 -22468
rect 39144 -22532 39164 -22468
rect 39060 -22548 39164 -22532
rect 39060 -22612 39080 -22548
rect 39144 -22612 39164 -22548
rect 39060 -22628 39164 -22612
rect 39060 -22692 39080 -22628
rect 39144 -22692 39164 -22628
rect 39060 -22708 39164 -22692
rect 39060 -22772 39080 -22708
rect 39144 -22772 39164 -22708
rect 39060 -22788 39164 -22772
rect 39060 -22852 39080 -22788
rect 39144 -22852 39164 -22788
rect 39060 -22868 39164 -22852
rect 39060 -22932 39080 -22868
rect 39144 -22932 39164 -22868
rect 39060 -22948 39164 -22932
rect 39060 -23012 39080 -22948
rect 39144 -23012 39164 -22948
rect 39060 -23028 39164 -23012
rect 39060 -23092 39080 -23028
rect 39144 -23092 39164 -23028
rect 39060 -23108 39164 -23092
rect 39060 -23172 39080 -23108
rect 39144 -23172 39164 -23108
rect 39060 -23188 39164 -23172
rect 39060 -23252 39080 -23188
rect 39144 -23252 39164 -23188
rect 39060 -23268 39164 -23252
rect 39060 -23332 39080 -23268
rect 39144 -23332 39164 -23268
rect 39060 -23348 39164 -23332
rect 39060 -23412 39080 -23348
rect 39144 -23412 39164 -23348
rect 39060 -23428 39164 -23412
rect 39060 -23492 39080 -23428
rect 39144 -23492 39164 -23428
rect 39060 -23508 39164 -23492
rect 39060 -23572 39080 -23508
rect 39144 -23572 39164 -23508
rect 39060 -23588 39164 -23572
rect 39060 -23652 39080 -23588
rect 39144 -23652 39164 -23588
rect 39060 -23668 39164 -23652
rect 39060 -23732 39080 -23668
rect 39144 -23732 39164 -23668
rect 39060 -23748 39164 -23732
rect 39060 -23812 39080 -23748
rect 39144 -23812 39164 -23748
rect 39060 -23828 39164 -23812
rect 39060 -23892 39080 -23828
rect 39144 -23892 39164 -23828
rect 39060 -23908 39164 -23892
rect 39060 -23972 39080 -23908
rect 39144 -23972 39164 -23908
rect 39060 -23988 39164 -23972
rect 39060 -24052 39080 -23988
rect 39144 -24052 39164 -23988
rect 39060 -24068 39164 -24052
rect 39060 -24132 39080 -24068
rect 39144 -24132 39164 -24068
rect 39060 -24148 39164 -24132
rect 39060 -24212 39080 -24148
rect 39144 -24212 39164 -24148
rect 39060 -24228 39164 -24212
rect 39060 -24292 39080 -24228
rect 39144 -24292 39164 -24228
rect 39060 -24308 39164 -24292
rect 39060 -24372 39080 -24308
rect 39144 -24372 39164 -24308
rect 39060 -24388 39164 -24372
rect 39060 -24452 39080 -24388
rect 39144 -24452 39164 -24388
rect 39060 -24468 39164 -24452
rect 39060 -24532 39080 -24468
rect 39144 -24532 39164 -24468
rect 39060 -24548 39164 -24532
rect 39060 -24612 39080 -24548
rect 39144 -24612 39164 -24548
rect 39060 -24628 39164 -24612
rect 39060 -24692 39080 -24628
rect 39144 -24692 39164 -24628
rect 39060 -24708 39164 -24692
rect 39060 -24772 39080 -24708
rect 39144 -24772 39164 -24708
rect 39060 -24788 39164 -24772
rect 39060 -24852 39080 -24788
rect 39144 -24852 39164 -24788
rect 39060 -24868 39164 -24852
rect 39060 -24932 39080 -24868
rect 39144 -24932 39164 -24868
rect 39060 -24948 39164 -24932
rect 39060 -25012 39080 -24948
rect 39144 -25012 39164 -24948
rect 39060 -25028 39164 -25012
rect 39060 -25092 39080 -25028
rect 39144 -25092 39164 -25028
rect 39060 -25108 39164 -25092
rect 39060 -25172 39080 -25108
rect 39144 -25172 39164 -25108
rect 39060 -25188 39164 -25172
rect 39060 -25252 39080 -25188
rect 39144 -25252 39164 -25188
rect 39060 -25268 39164 -25252
rect 39060 -25332 39080 -25268
rect 39144 -25332 39164 -25268
rect 39060 -25348 39164 -25332
rect 39060 -25412 39080 -25348
rect 39144 -25412 39164 -25348
rect 39060 -25428 39164 -25412
rect 39060 -25492 39080 -25428
rect 39144 -25492 39164 -25428
rect 39060 -25508 39164 -25492
rect 39060 -25572 39080 -25508
rect 39144 -25572 39164 -25508
rect 39060 -25588 39164 -25572
rect 39060 -25652 39080 -25588
rect 39144 -25652 39164 -25588
rect 39060 -25668 39164 -25652
rect 39060 -25732 39080 -25668
rect 39144 -25732 39164 -25668
rect 39060 -25748 39164 -25732
rect 39060 -25812 39080 -25748
rect 39144 -25812 39164 -25748
rect 39060 -25828 39164 -25812
rect 39060 -25892 39080 -25828
rect 39144 -25892 39164 -25828
rect 39060 -25908 39164 -25892
rect 39060 -25972 39080 -25908
rect 39144 -25972 39164 -25908
rect 39060 -25988 39164 -25972
rect 39060 -26052 39080 -25988
rect 39144 -26052 39164 -25988
rect 39060 -26068 39164 -26052
rect 39060 -26132 39080 -26068
rect 39144 -26132 39164 -26068
rect 39060 -26148 39164 -26132
rect 39060 -26212 39080 -26148
rect 39144 -26212 39164 -26148
rect 39060 -26228 39164 -26212
rect 39060 -26292 39080 -26228
rect 39144 -26292 39164 -26228
rect 39060 -26308 39164 -26292
rect 39060 -26372 39080 -26308
rect 39144 -26372 39164 -26308
rect 39060 -26388 39164 -26372
rect 33448 -26748 33552 -26452
rect 27836 -26828 27940 -26812
rect 27836 -26892 27856 -26828
rect 27920 -26892 27940 -26828
rect 27836 -26908 27940 -26892
rect 27836 -26972 27856 -26908
rect 27920 -26972 27940 -26908
rect 27836 -26988 27940 -26972
rect 27836 -27052 27856 -26988
rect 27920 -27052 27940 -26988
rect 27836 -27068 27940 -27052
rect 27836 -27132 27856 -27068
rect 27920 -27132 27940 -27068
rect 27836 -27148 27940 -27132
rect 27836 -27212 27856 -27148
rect 27920 -27212 27940 -27148
rect 27836 -27228 27940 -27212
rect 27836 -27292 27856 -27228
rect 27920 -27292 27940 -27228
rect 27836 -27308 27940 -27292
rect 27836 -27372 27856 -27308
rect 27920 -27372 27940 -27308
rect 27836 -27388 27940 -27372
rect 27836 -27452 27856 -27388
rect 27920 -27452 27940 -27388
rect 27836 -27468 27940 -27452
rect 27836 -27532 27856 -27468
rect 27920 -27532 27940 -27468
rect 27836 -27548 27940 -27532
rect 27836 -27612 27856 -27548
rect 27920 -27612 27940 -27548
rect 27836 -27628 27940 -27612
rect 27836 -27692 27856 -27628
rect 27920 -27692 27940 -27628
rect 27836 -27708 27940 -27692
rect 27836 -27772 27856 -27708
rect 27920 -27772 27940 -27708
rect 27836 -27788 27940 -27772
rect 27836 -27852 27856 -27788
rect 27920 -27852 27940 -27788
rect 27836 -27868 27940 -27852
rect 27836 -27932 27856 -27868
rect 27920 -27932 27940 -27868
rect 27836 -27948 27940 -27932
rect 27836 -28012 27856 -27948
rect 27920 -28012 27940 -27948
rect 27836 -28028 27940 -28012
rect 27836 -28092 27856 -28028
rect 27920 -28092 27940 -28028
rect 27836 -28108 27940 -28092
rect 27836 -28172 27856 -28108
rect 27920 -28172 27940 -28108
rect 27836 -28188 27940 -28172
rect 27836 -28252 27856 -28188
rect 27920 -28252 27940 -28188
rect 27836 -28268 27940 -28252
rect 27836 -28332 27856 -28268
rect 27920 -28332 27940 -28268
rect 27836 -28348 27940 -28332
rect 27836 -28412 27856 -28348
rect 27920 -28412 27940 -28348
rect 27836 -28428 27940 -28412
rect 27836 -28492 27856 -28428
rect 27920 -28492 27940 -28428
rect 27836 -28508 27940 -28492
rect 27836 -28572 27856 -28508
rect 27920 -28572 27940 -28508
rect 27836 -28588 27940 -28572
rect 27836 -28652 27856 -28588
rect 27920 -28652 27940 -28588
rect 27836 -28668 27940 -28652
rect 27836 -28732 27856 -28668
rect 27920 -28732 27940 -28668
rect 27836 -28748 27940 -28732
rect 27836 -28812 27856 -28748
rect 27920 -28812 27940 -28748
rect 27836 -28828 27940 -28812
rect 27836 -28892 27856 -28828
rect 27920 -28892 27940 -28828
rect 27836 -28908 27940 -28892
rect 27836 -28972 27856 -28908
rect 27920 -28972 27940 -28908
rect 27836 -28988 27940 -28972
rect 27836 -29052 27856 -28988
rect 27920 -29052 27940 -28988
rect 27836 -29068 27940 -29052
rect 27836 -29132 27856 -29068
rect 27920 -29132 27940 -29068
rect 27836 -29148 27940 -29132
rect 27836 -29212 27856 -29148
rect 27920 -29212 27940 -29148
rect 27836 -29228 27940 -29212
rect 27836 -29292 27856 -29228
rect 27920 -29292 27940 -29228
rect 27836 -29308 27940 -29292
rect 27836 -29372 27856 -29308
rect 27920 -29372 27940 -29308
rect 27836 -29388 27940 -29372
rect 27836 -29452 27856 -29388
rect 27920 -29452 27940 -29388
rect 27836 -29468 27940 -29452
rect 27836 -29532 27856 -29468
rect 27920 -29532 27940 -29468
rect 27836 -29548 27940 -29532
rect 27836 -29612 27856 -29548
rect 27920 -29612 27940 -29548
rect 27836 -29628 27940 -29612
rect 27836 -29692 27856 -29628
rect 27920 -29692 27940 -29628
rect 27836 -29708 27940 -29692
rect 27836 -29772 27856 -29708
rect 27920 -29772 27940 -29708
rect 27836 -29788 27940 -29772
rect 27836 -29852 27856 -29788
rect 27920 -29852 27940 -29788
rect 27836 -29868 27940 -29852
rect 27836 -29932 27856 -29868
rect 27920 -29932 27940 -29868
rect 27836 -29948 27940 -29932
rect 27836 -30012 27856 -29948
rect 27920 -30012 27940 -29948
rect 27836 -30028 27940 -30012
rect 27836 -30092 27856 -30028
rect 27920 -30092 27940 -30028
rect 27836 -30108 27940 -30092
rect 27836 -30172 27856 -30108
rect 27920 -30172 27940 -30108
rect 27836 -30188 27940 -30172
rect 27836 -30252 27856 -30188
rect 27920 -30252 27940 -30188
rect 27836 -30268 27940 -30252
rect 27836 -30332 27856 -30268
rect 27920 -30332 27940 -30268
rect 27836 -30348 27940 -30332
rect 27836 -30412 27856 -30348
rect 27920 -30412 27940 -30348
rect 27836 -30428 27940 -30412
rect 27836 -30492 27856 -30428
rect 27920 -30492 27940 -30428
rect 27836 -30508 27940 -30492
rect 27836 -30572 27856 -30508
rect 27920 -30572 27940 -30508
rect 27836 -30588 27940 -30572
rect 27836 -30652 27856 -30588
rect 27920 -30652 27940 -30588
rect 27836 -30668 27940 -30652
rect 27836 -30732 27856 -30668
rect 27920 -30732 27940 -30668
rect 27836 -30748 27940 -30732
rect 27836 -30812 27856 -30748
rect 27920 -30812 27940 -30748
rect 27836 -30828 27940 -30812
rect 27836 -30892 27856 -30828
rect 27920 -30892 27940 -30828
rect 27836 -30908 27940 -30892
rect 27836 -30972 27856 -30908
rect 27920 -30972 27940 -30908
rect 27836 -30988 27940 -30972
rect 27836 -31052 27856 -30988
rect 27920 -31052 27940 -30988
rect 27836 -31068 27940 -31052
rect 27836 -31132 27856 -31068
rect 27920 -31132 27940 -31068
rect 27836 -31148 27940 -31132
rect 27836 -31212 27856 -31148
rect 27920 -31212 27940 -31148
rect 27836 -31228 27940 -31212
rect 27836 -31292 27856 -31228
rect 27920 -31292 27940 -31228
rect 27836 -31308 27940 -31292
rect 27836 -31372 27856 -31308
rect 27920 -31372 27940 -31308
rect 27836 -31388 27940 -31372
rect 27836 -31452 27856 -31388
rect 27920 -31452 27940 -31388
rect 27836 -31468 27940 -31452
rect 27836 -31532 27856 -31468
rect 27920 -31532 27940 -31468
rect 27836 -31548 27940 -31532
rect 27836 -31612 27856 -31548
rect 27920 -31612 27940 -31548
rect 27836 -31628 27940 -31612
rect 27836 -31692 27856 -31628
rect 27920 -31692 27940 -31628
rect 27836 -31708 27940 -31692
rect 22224 -32068 22328 -31772
rect 16612 -32148 16716 -32132
rect 16612 -32212 16632 -32148
rect 16696 -32212 16716 -32148
rect 16612 -32228 16716 -32212
rect 16612 -32292 16632 -32228
rect 16696 -32292 16716 -32228
rect 16612 -32308 16716 -32292
rect 16612 -32372 16632 -32308
rect 16696 -32372 16716 -32308
rect 16612 -32388 16716 -32372
rect 16612 -32452 16632 -32388
rect 16696 -32452 16716 -32388
rect 16612 -32468 16716 -32452
rect 16612 -32532 16632 -32468
rect 16696 -32532 16716 -32468
rect 16612 -32548 16716 -32532
rect 16612 -32612 16632 -32548
rect 16696 -32612 16716 -32548
rect 16612 -32628 16716 -32612
rect 16612 -32692 16632 -32628
rect 16696 -32692 16716 -32628
rect 16612 -32708 16716 -32692
rect 16612 -32772 16632 -32708
rect 16696 -32772 16716 -32708
rect 16612 -32788 16716 -32772
rect 16612 -32852 16632 -32788
rect 16696 -32852 16716 -32788
rect 16612 -32868 16716 -32852
rect 16612 -32932 16632 -32868
rect 16696 -32932 16716 -32868
rect 16612 -32948 16716 -32932
rect 16612 -33012 16632 -32948
rect 16696 -33012 16716 -32948
rect 16612 -33028 16716 -33012
rect 16612 -33092 16632 -33028
rect 16696 -33092 16716 -33028
rect 16612 -33108 16716 -33092
rect 16612 -33172 16632 -33108
rect 16696 -33172 16716 -33108
rect 16612 -33188 16716 -33172
rect 16612 -33252 16632 -33188
rect 16696 -33252 16716 -33188
rect 16612 -33268 16716 -33252
rect 16612 -33332 16632 -33268
rect 16696 -33332 16716 -33268
rect 16612 -33348 16716 -33332
rect 16612 -33412 16632 -33348
rect 16696 -33412 16716 -33348
rect 16612 -33428 16716 -33412
rect 16612 -33492 16632 -33428
rect 16696 -33492 16716 -33428
rect 16612 -33508 16716 -33492
rect 16612 -33572 16632 -33508
rect 16696 -33572 16716 -33508
rect 16612 -33588 16716 -33572
rect 16612 -33652 16632 -33588
rect 16696 -33652 16716 -33588
rect 16612 -33668 16716 -33652
rect 16612 -33732 16632 -33668
rect 16696 -33732 16716 -33668
rect 16612 -33748 16716 -33732
rect 16612 -33812 16632 -33748
rect 16696 -33812 16716 -33748
rect 16612 -33828 16716 -33812
rect 16612 -33892 16632 -33828
rect 16696 -33892 16716 -33828
rect 16612 -33908 16716 -33892
rect 16612 -33972 16632 -33908
rect 16696 -33972 16716 -33908
rect 16612 -33988 16716 -33972
rect 16612 -34052 16632 -33988
rect 16696 -34052 16716 -33988
rect 16612 -34068 16716 -34052
rect 16612 -34132 16632 -34068
rect 16696 -34132 16716 -34068
rect 16612 -34148 16716 -34132
rect 16612 -34212 16632 -34148
rect 16696 -34212 16716 -34148
rect 16612 -34228 16716 -34212
rect 16612 -34292 16632 -34228
rect 16696 -34292 16716 -34228
rect 16612 -34308 16716 -34292
rect 16612 -34372 16632 -34308
rect 16696 -34372 16716 -34308
rect 16612 -34388 16716 -34372
rect 16612 -34452 16632 -34388
rect 16696 -34452 16716 -34388
rect 16612 -34468 16716 -34452
rect 16612 -34532 16632 -34468
rect 16696 -34532 16716 -34468
rect 16612 -34548 16716 -34532
rect 16612 -34612 16632 -34548
rect 16696 -34612 16716 -34548
rect 16612 -34628 16716 -34612
rect 16612 -34692 16632 -34628
rect 16696 -34692 16716 -34628
rect 16612 -34708 16716 -34692
rect 16612 -34772 16632 -34708
rect 16696 -34772 16716 -34708
rect 16612 -34788 16716 -34772
rect 16612 -34852 16632 -34788
rect 16696 -34852 16716 -34788
rect 16612 -34868 16716 -34852
rect 16612 -34932 16632 -34868
rect 16696 -34932 16716 -34868
rect 16612 -34948 16716 -34932
rect 16612 -35012 16632 -34948
rect 16696 -35012 16716 -34948
rect 16612 -35028 16716 -35012
rect 16612 -35092 16632 -35028
rect 16696 -35092 16716 -35028
rect 16612 -35108 16716 -35092
rect 16612 -35172 16632 -35108
rect 16696 -35172 16716 -35108
rect 16612 -35188 16716 -35172
rect 16612 -35252 16632 -35188
rect 16696 -35252 16716 -35188
rect 16612 -35268 16716 -35252
rect 16612 -35332 16632 -35268
rect 16696 -35332 16716 -35268
rect 16612 -35348 16716 -35332
rect 16612 -35412 16632 -35348
rect 16696 -35412 16716 -35348
rect 16612 -35428 16716 -35412
rect 16612 -35492 16632 -35428
rect 16696 -35492 16716 -35428
rect 16612 -35508 16716 -35492
rect 16612 -35572 16632 -35508
rect 16696 -35572 16716 -35508
rect 16612 -35588 16716 -35572
rect 16612 -35652 16632 -35588
rect 16696 -35652 16716 -35588
rect 16612 -35668 16716 -35652
rect 16612 -35732 16632 -35668
rect 16696 -35732 16716 -35668
rect 16612 -35748 16716 -35732
rect 16612 -35812 16632 -35748
rect 16696 -35812 16716 -35748
rect 16612 -35828 16716 -35812
rect 16612 -35892 16632 -35828
rect 16696 -35892 16716 -35828
rect 16612 -35908 16716 -35892
rect 16612 -35972 16632 -35908
rect 16696 -35972 16716 -35908
rect 16612 -35988 16716 -35972
rect 16612 -36052 16632 -35988
rect 16696 -36052 16716 -35988
rect 16612 -36068 16716 -36052
rect 16612 -36132 16632 -36068
rect 16696 -36132 16716 -36068
rect 16612 -36148 16716 -36132
rect 16612 -36212 16632 -36148
rect 16696 -36212 16716 -36148
rect 16612 -36228 16716 -36212
rect 16612 -36292 16632 -36228
rect 16696 -36292 16716 -36228
rect 16612 -36308 16716 -36292
rect 16612 -36372 16632 -36308
rect 16696 -36372 16716 -36308
rect 16612 -36388 16716 -36372
rect 16612 -36452 16632 -36388
rect 16696 -36452 16716 -36388
rect 16612 -36468 16716 -36452
rect 16612 -36532 16632 -36468
rect 16696 -36532 16716 -36468
rect 16612 -36548 16716 -36532
rect 16612 -36612 16632 -36548
rect 16696 -36612 16716 -36548
rect 16612 -36628 16716 -36612
rect 16612 -36692 16632 -36628
rect 16696 -36692 16716 -36628
rect 16612 -36708 16716 -36692
rect 16612 -36772 16632 -36708
rect 16696 -36772 16716 -36708
rect 16612 -36788 16716 -36772
rect 16612 -36852 16632 -36788
rect 16696 -36852 16716 -36788
rect 16612 -36868 16716 -36852
rect 16612 -36932 16632 -36868
rect 16696 -36932 16716 -36868
rect 16612 -36948 16716 -36932
rect 16612 -37012 16632 -36948
rect 16696 -37012 16716 -36948
rect 16612 -37028 16716 -37012
rect 11000 -37240 11104 -37092
rect 13832 -37240 13936 -37041
rect 16612 -37092 16632 -37028
rect 16696 -37092 16716 -37028
rect 17035 -32148 21957 -32119
rect 17035 -37012 17064 -32148
rect 21928 -37012 21957 -32148
rect 17035 -37041 21957 -37012
rect 22224 -32132 22244 -32068
rect 22308 -32132 22328 -32068
rect 25056 -32119 25160 -31721
rect 27836 -31772 27856 -31708
rect 27920 -31772 27940 -31708
rect 28259 -26828 33181 -26799
rect 28259 -31692 28288 -26828
rect 33152 -31692 33181 -26828
rect 28259 -31721 33181 -31692
rect 33448 -26812 33468 -26748
rect 33532 -26812 33552 -26748
rect 36280 -26799 36384 -26401
rect 39060 -26452 39080 -26388
rect 39144 -26452 39164 -26388
rect 39060 -26748 39164 -26452
rect 33448 -26828 33552 -26812
rect 33448 -26892 33468 -26828
rect 33532 -26892 33552 -26828
rect 33448 -26908 33552 -26892
rect 33448 -26972 33468 -26908
rect 33532 -26972 33552 -26908
rect 33448 -26988 33552 -26972
rect 33448 -27052 33468 -26988
rect 33532 -27052 33552 -26988
rect 33448 -27068 33552 -27052
rect 33448 -27132 33468 -27068
rect 33532 -27132 33552 -27068
rect 33448 -27148 33552 -27132
rect 33448 -27212 33468 -27148
rect 33532 -27212 33552 -27148
rect 33448 -27228 33552 -27212
rect 33448 -27292 33468 -27228
rect 33532 -27292 33552 -27228
rect 33448 -27308 33552 -27292
rect 33448 -27372 33468 -27308
rect 33532 -27372 33552 -27308
rect 33448 -27388 33552 -27372
rect 33448 -27452 33468 -27388
rect 33532 -27452 33552 -27388
rect 33448 -27468 33552 -27452
rect 33448 -27532 33468 -27468
rect 33532 -27532 33552 -27468
rect 33448 -27548 33552 -27532
rect 33448 -27612 33468 -27548
rect 33532 -27612 33552 -27548
rect 33448 -27628 33552 -27612
rect 33448 -27692 33468 -27628
rect 33532 -27692 33552 -27628
rect 33448 -27708 33552 -27692
rect 33448 -27772 33468 -27708
rect 33532 -27772 33552 -27708
rect 33448 -27788 33552 -27772
rect 33448 -27852 33468 -27788
rect 33532 -27852 33552 -27788
rect 33448 -27868 33552 -27852
rect 33448 -27932 33468 -27868
rect 33532 -27932 33552 -27868
rect 33448 -27948 33552 -27932
rect 33448 -28012 33468 -27948
rect 33532 -28012 33552 -27948
rect 33448 -28028 33552 -28012
rect 33448 -28092 33468 -28028
rect 33532 -28092 33552 -28028
rect 33448 -28108 33552 -28092
rect 33448 -28172 33468 -28108
rect 33532 -28172 33552 -28108
rect 33448 -28188 33552 -28172
rect 33448 -28252 33468 -28188
rect 33532 -28252 33552 -28188
rect 33448 -28268 33552 -28252
rect 33448 -28332 33468 -28268
rect 33532 -28332 33552 -28268
rect 33448 -28348 33552 -28332
rect 33448 -28412 33468 -28348
rect 33532 -28412 33552 -28348
rect 33448 -28428 33552 -28412
rect 33448 -28492 33468 -28428
rect 33532 -28492 33552 -28428
rect 33448 -28508 33552 -28492
rect 33448 -28572 33468 -28508
rect 33532 -28572 33552 -28508
rect 33448 -28588 33552 -28572
rect 33448 -28652 33468 -28588
rect 33532 -28652 33552 -28588
rect 33448 -28668 33552 -28652
rect 33448 -28732 33468 -28668
rect 33532 -28732 33552 -28668
rect 33448 -28748 33552 -28732
rect 33448 -28812 33468 -28748
rect 33532 -28812 33552 -28748
rect 33448 -28828 33552 -28812
rect 33448 -28892 33468 -28828
rect 33532 -28892 33552 -28828
rect 33448 -28908 33552 -28892
rect 33448 -28972 33468 -28908
rect 33532 -28972 33552 -28908
rect 33448 -28988 33552 -28972
rect 33448 -29052 33468 -28988
rect 33532 -29052 33552 -28988
rect 33448 -29068 33552 -29052
rect 33448 -29132 33468 -29068
rect 33532 -29132 33552 -29068
rect 33448 -29148 33552 -29132
rect 33448 -29212 33468 -29148
rect 33532 -29212 33552 -29148
rect 33448 -29228 33552 -29212
rect 33448 -29292 33468 -29228
rect 33532 -29292 33552 -29228
rect 33448 -29308 33552 -29292
rect 33448 -29372 33468 -29308
rect 33532 -29372 33552 -29308
rect 33448 -29388 33552 -29372
rect 33448 -29452 33468 -29388
rect 33532 -29452 33552 -29388
rect 33448 -29468 33552 -29452
rect 33448 -29532 33468 -29468
rect 33532 -29532 33552 -29468
rect 33448 -29548 33552 -29532
rect 33448 -29612 33468 -29548
rect 33532 -29612 33552 -29548
rect 33448 -29628 33552 -29612
rect 33448 -29692 33468 -29628
rect 33532 -29692 33552 -29628
rect 33448 -29708 33552 -29692
rect 33448 -29772 33468 -29708
rect 33532 -29772 33552 -29708
rect 33448 -29788 33552 -29772
rect 33448 -29852 33468 -29788
rect 33532 -29852 33552 -29788
rect 33448 -29868 33552 -29852
rect 33448 -29932 33468 -29868
rect 33532 -29932 33552 -29868
rect 33448 -29948 33552 -29932
rect 33448 -30012 33468 -29948
rect 33532 -30012 33552 -29948
rect 33448 -30028 33552 -30012
rect 33448 -30092 33468 -30028
rect 33532 -30092 33552 -30028
rect 33448 -30108 33552 -30092
rect 33448 -30172 33468 -30108
rect 33532 -30172 33552 -30108
rect 33448 -30188 33552 -30172
rect 33448 -30252 33468 -30188
rect 33532 -30252 33552 -30188
rect 33448 -30268 33552 -30252
rect 33448 -30332 33468 -30268
rect 33532 -30332 33552 -30268
rect 33448 -30348 33552 -30332
rect 33448 -30412 33468 -30348
rect 33532 -30412 33552 -30348
rect 33448 -30428 33552 -30412
rect 33448 -30492 33468 -30428
rect 33532 -30492 33552 -30428
rect 33448 -30508 33552 -30492
rect 33448 -30572 33468 -30508
rect 33532 -30572 33552 -30508
rect 33448 -30588 33552 -30572
rect 33448 -30652 33468 -30588
rect 33532 -30652 33552 -30588
rect 33448 -30668 33552 -30652
rect 33448 -30732 33468 -30668
rect 33532 -30732 33552 -30668
rect 33448 -30748 33552 -30732
rect 33448 -30812 33468 -30748
rect 33532 -30812 33552 -30748
rect 33448 -30828 33552 -30812
rect 33448 -30892 33468 -30828
rect 33532 -30892 33552 -30828
rect 33448 -30908 33552 -30892
rect 33448 -30972 33468 -30908
rect 33532 -30972 33552 -30908
rect 33448 -30988 33552 -30972
rect 33448 -31052 33468 -30988
rect 33532 -31052 33552 -30988
rect 33448 -31068 33552 -31052
rect 33448 -31132 33468 -31068
rect 33532 -31132 33552 -31068
rect 33448 -31148 33552 -31132
rect 33448 -31212 33468 -31148
rect 33532 -31212 33552 -31148
rect 33448 -31228 33552 -31212
rect 33448 -31292 33468 -31228
rect 33532 -31292 33552 -31228
rect 33448 -31308 33552 -31292
rect 33448 -31372 33468 -31308
rect 33532 -31372 33552 -31308
rect 33448 -31388 33552 -31372
rect 33448 -31452 33468 -31388
rect 33532 -31452 33552 -31388
rect 33448 -31468 33552 -31452
rect 33448 -31532 33468 -31468
rect 33532 -31532 33552 -31468
rect 33448 -31548 33552 -31532
rect 33448 -31612 33468 -31548
rect 33532 -31612 33552 -31548
rect 33448 -31628 33552 -31612
rect 33448 -31692 33468 -31628
rect 33532 -31692 33552 -31628
rect 33448 -31708 33552 -31692
rect 27836 -32068 27940 -31772
rect 22224 -32148 22328 -32132
rect 22224 -32212 22244 -32148
rect 22308 -32212 22328 -32148
rect 22224 -32228 22328 -32212
rect 22224 -32292 22244 -32228
rect 22308 -32292 22328 -32228
rect 22224 -32308 22328 -32292
rect 22224 -32372 22244 -32308
rect 22308 -32372 22328 -32308
rect 22224 -32388 22328 -32372
rect 22224 -32452 22244 -32388
rect 22308 -32452 22328 -32388
rect 22224 -32468 22328 -32452
rect 22224 -32532 22244 -32468
rect 22308 -32532 22328 -32468
rect 22224 -32548 22328 -32532
rect 22224 -32612 22244 -32548
rect 22308 -32612 22328 -32548
rect 22224 -32628 22328 -32612
rect 22224 -32692 22244 -32628
rect 22308 -32692 22328 -32628
rect 22224 -32708 22328 -32692
rect 22224 -32772 22244 -32708
rect 22308 -32772 22328 -32708
rect 22224 -32788 22328 -32772
rect 22224 -32852 22244 -32788
rect 22308 -32852 22328 -32788
rect 22224 -32868 22328 -32852
rect 22224 -32932 22244 -32868
rect 22308 -32932 22328 -32868
rect 22224 -32948 22328 -32932
rect 22224 -33012 22244 -32948
rect 22308 -33012 22328 -32948
rect 22224 -33028 22328 -33012
rect 22224 -33092 22244 -33028
rect 22308 -33092 22328 -33028
rect 22224 -33108 22328 -33092
rect 22224 -33172 22244 -33108
rect 22308 -33172 22328 -33108
rect 22224 -33188 22328 -33172
rect 22224 -33252 22244 -33188
rect 22308 -33252 22328 -33188
rect 22224 -33268 22328 -33252
rect 22224 -33332 22244 -33268
rect 22308 -33332 22328 -33268
rect 22224 -33348 22328 -33332
rect 22224 -33412 22244 -33348
rect 22308 -33412 22328 -33348
rect 22224 -33428 22328 -33412
rect 22224 -33492 22244 -33428
rect 22308 -33492 22328 -33428
rect 22224 -33508 22328 -33492
rect 22224 -33572 22244 -33508
rect 22308 -33572 22328 -33508
rect 22224 -33588 22328 -33572
rect 22224 -33652 22244 -33588
rect 22308 -33652 22328 -33588
rect 22224 -33668 22328 -33652
rect 22224 -33732 22244 -33668
rect 22308 -33732 22328 -33668
rect 22224 -33748 22328 -33732
rect 22224 -33812 22244 -33748
rect 22308 -33812 22328 -33748
rect 22224 -33828 22328 -33812
rect 22224 -33892 22244 -33828
rect 22308 -33892 22328 -33828
rect 22224 -33908 22328 -33892
rect 22224 -33972 22244 -33908
rect 22308 -33972 22328 -33908
rect 22224 -33988 22328 -33972
rect 22224 -34052 22244 -33988
rect 22308 -34052 22328 -33988
rect 22224 -34068 22328 -34052
rect 22224 -34132 22244 -34068
rect 22308 -34132 22328 -34068
rect 22224 -34148 22328 -34132
rect 22224 -34212 22244 -34148
rect 22308 -34212 22328 -34148
rect 22224 -34228 22328 -34212
rect 22224 -34292 22244 -34228
rect 22308 -34292 22328 -34228
rect 22224 -34308 22328 -34292
rect 22224 -34372 22244 -34308
rect 22308 -34372 22328 -34308
rect 22224 -34388 22328 -34372
rect 22224 -34452 22244 -34388
rect 22308 -34452 22328 -34388
rect 22224 -34468 22328 -34452
rect 22224 -34532 22244 -34468
rect 22308 -34532 22328 -34468
rect 22224 -34548 22328 -34532
rect 22224 -34612 22244 -34548
rect 22308 -34612 22328 -34548
rect 22224 -34628 22328 -34612
rect 22224 -34692 22244 -34628
rect 22308 -34692 22328 -34628
rect 22224 -34708 22328 -34692
rect 22224 -34772 22244 -34708
rect 22308 -34772 22328 -34708
rect 22224 -34788 22328 -34772
rect 22224 -34852 22244 -34788
rect 22308 -34852 22328 -34788
rect 22224 -34868 22328 -34852
rect 22224 -34932 22244 -34868
rect 22308 -34932 22328 -34868
rect 22224 -34948 22328 -34932
rect 22224 -35012 22244 -34948
rect 22308 -35012 22328 -34948
rect 22224 -35028 22328 -35012
rect 22224 -35092 22244 -35028
rect 22308 -35092 22328 -35028
rect 22224 -35108 22328 -35092
rect 22224 -35172 22244 -35108
rect 22308 -35172 22328 -35108
rect 22224 -35188 22328 -35172
rect 22224 -35252 22244 -35188
rect 22308 -35252 22328 -35188
rect 22224 -35268 22328 -35252
rect 22224 -35332 22244 -35268
rect 22308 -35332 22328 -35268
rect 22224 -35348 22328 -35332
rect 22224 -35412 22244 -35348
rect 22308 -35412 22328 -35348
rect 22224 -35428 22328 -35412
rect 22224 -35492 22244 -35428
rect 22308 -35492 22328 -35428
rect 22224 -35508 22328 -35492
rect 22224 -35572 22244 -35508
rect 22308 -35572 22328 -35508
rect 22224 -35588 22328 -35572
rect 22224 -35652 22244 -35588
rect 22308 -35652 22328 -35588
rect 22224 -35668 22328 -35652
rect 22224 -35732 22244 -35668
rect 22308 -35732 22328 -35668
rect 22224 -35748 22328 -35732
rect 22224 -35812 22244 -35748
rect 22308 -35812 22328 -35748
rect 22224 -35828 22328 -35812
rect 22224 -35892 22244 -35828
rect 22308 -35892 22328 -35828
rect 22224 -35908 22328 -35892
rect 22224 -35972 22244 -35908
rect 22308 -35972 22328 -35908
rect 22224 -35988 22328 -35972
rect 22224 -36052 22244 -35988
rect 22308 -36052 22328 -35988
rect 22224 -36068 22328 -36052
rect 22224 -36132 22244 -36068
rect 22308 -36132 22328 -36068
rect 22224 -36148 22328 -36132
rect 22224 -36212 22244 -36148
rect 22308 -36212 22328 -36148
rect 22224 -36228 22328 -36212
rect 22224 -36292 22244 -36228
rect 22308 -36292 22328 -36228
rect 22224 -36308 22328 -36292
rect 22224 -36372 22244 -36308
rect 22308 -36372 22328 -36308
rect 22224 -36388 22328 -36372
rect 22224 -36452 22244 -36388
rect 22308 -36452 22328 -36388
rect 22224 -36468 22328 -36452
rect 22224 -36532 22244 -36468
rect 22308 -36532 22328 -36468
rect 22224 -36548 22328 -36532
rect 22224 -36612 22244 -36548
rect 22308 -36612 22328 -36548
rect 22224 -36628 22328 -36612
rect 22224 -36692 22244 -36628
rect 22308 -36692 22328 -36628
rect 22224 -36708 22328 -36692
rect 22224 -36772 22244 -36708
rect 22308 -36772 22328 -36708
rect 22224 -36788 22328 -36772
rect 22224 -36852 22244 -36788
rect 22308 -36852 22328 -36788
rect 22224 -36868 22328 -36852
rect 22224 -36932 22244 -36868
rect 22308 -36932 22328 -36868
rect 22224 -36948 22328 -36932
rect 22224 -37012 22244 -36948
rect 22308 -37012 22328 -36948
rect 22224 -37028 22328 -37012
rect 16612 -37240 16716 -37092
rect 19444 -37240 19548 -37041
rect 22224 -37092 22244 -37028
rect 22308 -37092 22328 -37028
rect 22647 -32148 27569 -32119
rect 22647 -37012 22676 -32148
rect 27540 -37012 27569 -32148
rect 22647 -37041 27569 -37012
rect 27836 -32132 27856 -32068
rect 27920 -32132 27940 -32068
rect 30668 -32119 30772 -31721
rect 33448 -31772 33468 -31708
rect 33532 -31772 33552 -31708
rect 33871 -26828 38793 -26799
rect 33871 -31692 33900 -26828
rect 38764 -31692 38793 -26828
rect 33871 -31721 38793 -31692
rect 39060 -26812 39080 -26748
rect 39144 -26812 39164 -26748
rect 39060 -26828 39164 -26812
rect 39060 -26892 39080 -26828
rect 39144 -26892 39164 -26828
rect 39060 -26908 39164 -26892
rect 39060 -26972 39080 -26908
rect 39144 -26972 39164 -26908
rect 39060 -26988 39164 -26972
rect 39060 -27052 39080 -26988
rect 39144 -27052 39164 -26988
rect 39060 -27068 39164 -27052
rect 39060 -27132 39080 -27068
rect 39144 -27132 39164 -27068
rect 39060 -27148 39164 -27132
rect 39060 -27212 39080 -27148
rect 39144 -27212 39164 -27148
rect 39060 -27228 39164 -27212
rect 39060 -27292 39080 -27228
rect 39144 -27292 39164 -27228
rect 39060 -27308 39164 -27292
rect 39060 -27372 39080 -27308
rect 39144 -27372 39164 -27308
rect 39060 -27388 39164 -27372
rect 39060 -27452 39080 -27388
rect 39144 -27452 39164 -27388
rect 39060 -27468 39164 -27452
rect 39060 -27532 39080 -27468
rect 39144 -27532 39164 -27468
rect 39060 -27548 39164 -27532
rect 39060 -27612 39080 -27548
rect 39144 -27612 39164 -27548
rect 39060 -27628 39164 -27612
rect 39060 -27692 39080 -27628
rect 39144 -27692 39164 -27628
rect 39060 -27708 39164 -27692
rect 39060 -27772 39080 -27708
rect 39144 -27772 39164 -27708
rect 39060 -27788 39164 -27772
rect 39060 -27852 39080 -27788
rect 39144 -27852 39164 -27788
rect 39060 -27868 39164 -27852
rect 39060 -27932 39080 -27868
rect 39144 -27932 39164 -27868
rect 39060 -27948 39164 -27932
rect 39060 -28012 39080 -27948
rect 39144 -28012 39164 -27948
rect 39060 -28028 39164 -28012
rect 39060 -28092 39080 -28028
rect 39144 -28092 39164 -28028
rect 39060 -28108 39164 -28092
rect 39060 -28172 39080 -28108
rect 39144 -28172 39164 -28108
rect 39060 -28188 39164 -28172
rect 39060 -28252 39080 -28188
rect 39144 -28252 39164 -28188
rect 39060 -28268 39164 -28252
rect 39060 -28332 39080 -28268
rect 39144 -28332 39164 -28268
rect 39060 -28348 39164 -28332
rect 39060 -28412 39080 -28348
rect 39144 -28412 39164 -28348
rect 39060 -28428 39164 -28412
rect 39060 -28492 39080 -28428
rect 39144 -28492 39164 -28428
rect 39060 -28508 39164 -28492
rect 39060 -28572 39080 -28508
rect 39144 -28572 39164 -28508
rect 39060 -28588 39164 -28572
rect 39060 -28652 39080 -28588
rect 39144 -28652 39164 -28588
rect 39060 -28668 39164 -28652
rect 39060 -28732 39080 -28668
rect 39144 -28732 39164 -28668
rect 39060 -28748 39164 -28732
rect 39060 -28812 39080 -28748
rect 39144 -28812 39164 -28748
rect 39060 -28828 39164 -28812
rect 39060 -28892 39080 -28828
rect 39144 -28892 39164 -28828
rect 39060 -28908 39164 -28892
rect 39060 -28972 39080 -28908
rect 39144 -28972 39164 -28908
rect 39060 -28988 39164 -28972
rect 39060 -29052 39080 -28988
rect 39144 -29052 39164 -28988
rect 39060 -29068 39164 -29052
rect 39060 -29132 39080 -29068
rect 39144 -29132 39164 -29068
rect 39060 -29148 39164 -29132
rect 39060 -29212 39080 -29148
rect 39144 -29212 39164 -29148
rect 39060 -29228 39164 -29212
rect 39060 -29292 39080 -29228
rect 39144 -29292 39164 -29228
rect 39060 -29308 39164 -29292
rect 39060 -29372 39080 -29308
rect 39144 -29372 39164 -29308
rect 39060 -29388 39164 -29372
rect 39060 -29452 39080 -29388
rect 39144 -29452 39164 -29388
rect 39060 -29468 39164 -29452
rect 39060 -29532 39080 -29468
rect 39144 -29532 39164 -29468
rect 39060 -29548 39164 -29532
rect 39060 -29612 39080 -29548
rect 39144 -29612 39164 -29548
rect 39060 -29628 39164 -29612
rect 39060 -29692 39080 -29628
rect 39144 -29692 39164 -29628
rect 39060 -29708 39164 -29692
rect 39060 -29772 39080 -29708
rect 39144 -29772 39164 -29708
rect 39060 -29788 39164 -29772
rect 39060 -29852 39080 -29788
rect 39144 -29852 39164 -29788
rect 39060 -29868 39164 -29852
rect 39060 -29932 39080 -29868
rect 39144 -29932 39164 -29868
rect 39060 -29948 39164 -29932
rect 39060 -30012 39080 -29948
rect 39144 -30012 39164 -29948
rect 39060 -30028 39164 -30012
rect 39060 -30092 39080 -30028
rect 39144 -30092 39164 -30028
rect 39060 -30108 39164 -30092
rect 39060 -30172 39080 -30108
rect 39144 -30172 39164 -30108
rect 39060 -30188 39164 -30172
rect 39060 -30252 39080 -30188
rect 39144 -30252 39164 -30188
rect 39060 -30268 39164 -30252
rect 39060 -30332 39080 -30268
rect 39144 -30332 39164 -30268
rect 39060 -30348 39164 -30332
rect 39060 -30412 39080 -30348
rect 39144 -30412 39164 -30348
rect 39060 -30428 39164 -30412
rect 39060 -30492 39080 -30428
rect 39144 -30492 39164 -30428
rect 39060 -30508 39164 -30492
rect 39060 -30572 39080 -30508
rect 39144 -30572 39164 -30508
rect 39060 -30588 39164 -30572
rect 39060 -30652 39080 -30588
rect 39144 -30652 39164 -30588
rect 39060 -30668 39164 -30652
rect 39060 -30732 39080 -30668
rect 39144 -30732 39164 -30668
rect 39060 -30748 39164 -30732
rect 39060 -30812 39080 -30748
rect 39144 -30812 39164 -30748
rect 39060 -30828 39164 -30812
rect 39060 -30892 39080 -30828
rect 39144 -30892 39164 -30828
rect 39060 -30908 39164 -30892
rect 39060 -30972 39080 -30908
rect 39144 -30972 39164 -30908
rect 39060 -30988 39164 -30972
rect 39060 -31052 39080 -30988
rect 39144 -31052 39164 -30988
rect 39060 -31068 39164 -31052
rect 39060 -31132 39080 -31068
rect 39144 -31132 39164 -31068
rect 39060 -31148 39164 -31132
rect 39060 -31212 39080 -31148
rect 39144 -31212 39164 -31148
rect 39060 -31228 39164 -31212
rect 39060 -31292 39080 -31228
rect 39144 -31292 39164 -31228
rect 39060 -31308 39164 -31292
rect 39060 -31372 39080 -31308
rect 39144 -31372 39164 -31308
rect 39060 -31388 39164 -31372
rect 39060 -31452 39080 -31388
rect 39144 -31452 39164 -31388
rect 39060 -31468 39164 -31452
rect 39060 -31532 39080 -31468
rect 39144 -31532 39164 -31468
rect 39060 -31548 39164 -31532
rect 39060 -31612 39080 -31548
rect 39144 -31612 39164 -31548
rect 39060 -31628 39164 -31612
rect 39060 -31692 39080 -31628
rect 39144 -31692 39164 -31628
rect 39060 -31708 39164 -31692
rect 33448 -32068 33552 -31772
rect 27836 -32148 27940 -32132
rect 27836 -32212 27856 -32148
rect 27920 -32212 27940 -32148
rect 27836 -32228 27940 -32212
rect 27836 -32292 27856 -32228
rect 27920 -32292 27940 -32228
rect 27836 -32308 27940 -32292
rect 27836 -32372 27856 -32308
rect 27920 -32372 27940 -32308
rect 27836 -32388 27940 -32372
rect 27836 -32452 27856 -32388
rect 27920 -32452 27940 -32388
rect 27836 -32468 27940 -32452
rect 27836 -32532 27856 -32468
rect 27920 -32532 27940 -32468
rect 27836 -32548 27940 -32532
rect 27836 -32612 27856 -32548
rect 27920 -32612 27940 -32548
rect 27836 -32628 27940 -32612
rect 27836 -32692 27856 -32628
rect 27920 -32692 27940 -32628
rect 27836 -32708 27940 -32692
rect 27836 -32772 27856 -32708
rect 27920 -32772 27940 -32708
rect 27836 -32788 27940 -32772
rect 27836 -32852 27856 -32788
rect 27920 -32852 27940 -32788
rect 27836 -32868 27940 -32852
rect 27836 -32932 27856 -32868
rect 27920 -32932 27940 -32868
rect 27836 -32948 27940 -32932
rect 27836 -33012 27856 -32948
rect 27920 -33012 27940 -32948
rect 27836 -33028 27940 -33012
rect 27836 -33092 27856 -33028
rect 27920 -33092 27940 -33028
rect 27836 -33108 27940 -33092
rect 27836 -33172 27856 -33108
rect 27920 -33172 27940 -33108
rect 27836 -33188 27940 -33172
rect 27836 -33252 27856 -33188
rect 27920 -33252 27940 -33188
rect 27836 -33268 27940 -33252
rect 27836 -33332 27856 -33268
rect 27920 -33332 27940 -33268
rect 27836 -33348 27940 -33332
rect 27836 -33412 27856 -33348
rect 27920 -33412 27940 -33348
rect 27836 -33428 27940 -33412
rect 27836 -33492 27856 -33428
rect 27920 -33492 27940 -33428
rect 27836 -33508 27940 -33492
rect 27836 -33572 27856 -33508
rect 27920 -33572 27940 -33508
rect 27836 -33588 27940 -33572
rect 27836 -33652 27856 -33588
rect 27920 -33652 27940 -33588
rect 27836 -33668 27940 -33652
rect 27836 -33732 27856 -33668
rect 27920 -33732 27940 -33668
rect 27836 -33748 27940 -33732
rect 27836 -33812 27856 -33748
rect 27920 -33812 27940 -33748
rect 27836 -33828 27940 -33812
rect 27836 -33892 27856 -33828
rect 27920 -33892 27940 -33828
rect 27836 -33908 27940 -33892
rect 27836 -33972 27856 -33908
rect 27920 -33972 27940 -33908
rect 27836 -33988 27940 -33972
rect 27836 -34052 27856 -33988
rect 27920 -34052 27940 -33988
rect 27836 -34068 27940 -34052
rect 27836 -34132 27856 -34068
rect 27920 -34132 27940 -34068
rect 27836 -34148 27940 -34132
rect 27836 -34212 27856 -34148
rect 27920 -34212 27940 -34148
rect 27836 -34228 27940 -34212
rect 27836 -34292 27856 -34228
rect 27920 -34292 27940 -34228
rect 27836 -34308 27940 -34292
rect 27836 -34372 27856 -34308
rect 27920 -34372 27940 -34308
rect 27836 -34388 27940 -34372
rect 27836 -34452 27856 -34388
rect 27920 -34452 27940 -34388
rect 27836 -34468 27940 -34452
rect 27836 -34532 27856 -34468
rect 27920 -34532 27940 -34468
rect 27836 -34548 27940 -34532
rect 27836 -34612 27856 -34548
rect 27920 -34612 27940 -34548
rect 27836 -34628 27940 -34612
rect 27836 -34692 27856 -34628
rect 27920 -34692 27940 -34628
rect 27836 -34708 27940 -34692
rect 27836 -34772 27856 -34708
rect 27920 -34772 27940 -34708
rect 27836 -34788 27940 -34772
rect 27836 -34852 27856 -34788
rect 27920 -34852 27940 -34788
rect 27836 -34868 27940 -34852
rect 27836 -34932 27856 -34868
rect 27920 -34932 27940 -34868
rect 27836 -34948 27940 -34932
rect 27836 -35012 27856 -34948
rect 27920 -35012 27940 -34948
rect 27836 -35028 27940 -35012
rect 27836 -35092 27856 -35028
rect 27920 -35092 27940 -35028
rect 27836 -35108 27940 -35092
rect 27836 -35172 27856 -35108
rect 27920 -35172 27940 -35108
rect 27836 -35188 27940 -35172
rect 27836 -35252 27856 -35188
rect 27920 -35252 27940 -35188
rect 27836 -35268 27940 -35252
rect 27836 -35332 27856 -35268
rect 27920 -35332 27940 -35268
rect 27836 -35348 27940 -35332
rect 27836 -35412 27856 -35348
rect 27920 -35412 27940 -35348
rect 27836 -35428 27940 -35412
rect 27836 -35492 27856 -35428
rect 27920 -35492 27940 -35428
rect 27836 -35508 27940 -35492
rect 27836 -35572 27856 -35508
rect 27920 -35572 27940 -35508
rect 27836 -35588 27940 -35572
rect 27836 -35652 27856 -35588
rect 27920 -35652 27940 -35588
rect 27836 -35668 27940 -35652
rect 27836 -35732 27856 -35668
rect 27920 -35732 27940 -35668
rect 27836 -35748 27940 -35732
rect 27836 -35812 27856 -35748
rect 27920 -35812 27940 -35748
rect 27836 -35828 27940 -35812
rect 27836 -35892 27856 -35828
rect 27920 -35892 27940 -35828
rect 27836 -35908 27940 -35892
rect 27836 -35972 27856 -35908
rect 27920 -35972 27940 -35908
rect 27836 -35988 27940 -35972
rect 27836 -36052 27856 -35988
rect 27920 -36052 27940 -35988
rect 27836 -36068 27940 -36052
rect 27836 -36132 27856 -36068
rect 27920 -36132 27940 -36068
rect 27836 -36148 27940 -36132
rect 27836 -36212 27856 -36148
rect 27920 -36212 27940 -36148
rect 27836 -36228 27940 -36212
rect 27836 -36292 27856 -36228
rect 27920 -36292 27940 -36228
rect 27836 -36308 27940 -36292
rect 27836 -36372 27856 -36308
rect 27920 -36372 27940 -36308
rect 27836 -36388 27940 -36372
rect 27836 -36452 27856 -36388
rect 27920 -36452 27940 -36388
rect 27836 -36468 27940 -36452
rect 27836 -36532 27856 -36468
rect 27920 -36532 27940 -36468
rect 27836 -36548 27940 -36532
rect 27836 -36612 27856 -36548
rect 27920 -36612 27940 -36548
rect 27836 -36628 27940 -36612
rect 27836 -36692 27856 -36628
rect 27920 -36692 27940 -36628
rect 27836 -36708 27940 -36692
rect 27836 -36772 27856 -36708
rect 27920 -36772 27940 -36708
rect 27836 -36788 27940 -36772
rect 27836 -36852 27856 -36788
rect 27920 -36852 27940 -36788
rect 27836 -36868 27940 -36852
rect 27836 -36932 27856 -36868
rect 27920 -36932 27940 -36868
rect 27836 -36948 27940 -36932
rect 27836 -37012 27856 -36948
rect 27920 -37012 27940 -36948
rect 27836 -37028 27940 -37012
rect 22224 -37240 22328 -37092
rect 25056 -37240 25160 -37041
rect 27836 -37092 27856 -37028
rect 27920 -37092 27940 -37028
rect 28259 -32148 33181 -32119
rect 28259 -37012 28288 -32148
rect 33152 -37012 33181 -32148
rect 28259 -37041 33181 -37012
rect 33448 -32132 33468 -32068
rect 33532 -32132 33552 -32068
rect 36280 -32119 36384 -31721
rect 39060 -31772 39080 -31708
rect 39144 -31772 39164 -31708
rect 39060 -32068 39164 -31772
rect 33448 -32148 33552 -32132
rect 33448 -32212 33468 -32148
rect 33532 -32212 33552 -32148
rect 33448 -32228 33552 -32212
rect 33448 -32292 33468 -32228
rect 33532 -32292 33552 -32228
rect 33448 -32308 33552 -32292
rect 33448 -32372 33468 -32308
rect 33532 -32372 33552 -32308
rect 33448 -32388 33552 -32372
rect 33448 -32452 33468 -32388
rect 33532 -32452 33552 -32388
rect 33448 -32468 33552 -32452
rect 33448 -32532 33468 -32468
rect 33532 -32532 33552 -32468
rect 33448 -32548 33552 -32532
rect 33448 -32612 33468 -32548
rect 33532 -32612 33552 -32548
rect 33448 -32628 33552 -32612
rect 33448 -32692 33468 -32628
rect 33532 -32692 33552 -32628
rect 33448 -32708 33552 -32692
rect 33448 -32772 33468 -32708
rect 33532 -32772 33552 -32708
rect 33448 -32788 33552 -32772
rect 33448 -32852 33468 -32788
rect 33532 -32852 33552 -32788
rect 33448 -32868 33552 -32852
rect 33448 -32932 33468 -32868
rect 33532 -32932 33552 -32868
rect 33448 -32948 33552 -32932
rect 33448 -33012 33468 -32948
rect 33532 -33012 33552 -32948
rect 33448 -33028 33552 -33012
rect 33448 -33092 33468 -33028
rect 33532 -33092 33552 -33028
rect 33448 -33108 33552 -33092
rect 33448 -33172 33468 -33108
rect 33532 -33172 33552 -33108
rect 33448 -33188 33552 -33172
rect 33448 -33252 33468 -33188
rect 33532 -33252 33552 -33188
rect 33448 -33268 33552 -33252
rect 33448 -33332 33468 -33268
rect 33532 -33332 33552 -33268
rect 33448 -33348 33552 -33332
rect 33448 -33412 33468 -33348
rect 33532 -33412 33552 -33348
rect 33448 -33428 33552 -33412
rect 33448 -33492 33468 -33428
rect 33532 -33492 33552 -33428
rect 33448 -33508 33552 -33492
rect 33448 -33572 33468 -33508
rect 33532 -33572 33552 -33508
rect 33448 -33588 33552 -33572
rect 33448 -33652 33468 -33588
rect 33532 -33652 33552 -33588
rect 33448 -33668 33552 -33652
rect 33448 -33732 33468 -33668
rect 33532 -33732 33552 -33668
rect 33448 -33748 33552 -33732
rect 33448 -33812 33468 -33748
rect 33532 -33812 33552 -33748
rect 33448 -33828 33552 -33812
rect 33448 -33892 33468 -33828
rect 33532 -33892 33552 -33828
rect 33448 -33908 33552 -33892
rect 33448 -33972 33468 -33908
rect 33532 -33972 33552 -33908
rect 33448 -33988 33552 -33972
rect 33448 -34052 33468 -33988
rect 33532 -34052 33552 -33988
rect 33448 -34068 33552 -34052
rect 33448 -34132 33468 -34068
rect 33532 -34132 33552 -34068
rect 33448 -34148 33552 -34132
rect 33448 -34212 33468 -34148
rect 33532 -34212 33552 -34148
rect 33448 -34228 33552 -34212
rect 33448 -34292 33468 -34228
rect 33532 -34292 33552 -34228
rect 33448 -34308 33552 -34292
rect 33448 -34372 33468 -34308
rect 33532 -34372 33552 -34308
rect 33448 -34388 33552 -34372
rect 33448 -34452 33468 -34388
rect 33532 -34452 33552 -34388
rect 33448 -34468 33552 -34452
rect 33448 -34532 33468 -34468
rect 33532 -34532 33552 -34468
rect 33448 -34548 33552 -34532
rect 33448 -34612 33468 -34548
rect 33532 -34612 33552 -34548
rect 33448 -34628 33552 -34612
rect 33448 -34692 33468 -34628
rect 33532 -34692 33552 -34628
rect 33448 -34708 33552 -34692
rect 33448 -34772 33468 -34708
rect 33532 -34772 33552 -34708
rect 33448 -34788 33552 -34772
rect 33448 -34852 33468 -34788
rect 33532 -34852 33552 -34788
rect 33448 -34868 33552 -34852
rect 33448 -34932 33468 -34868
rect 33532 -34932 33552 -34868
rect 33448 -34948 33552 -34932
rect 33448 -35012 33468 -34948
rect 33532 -35012 33552 -34948
rect 33448 -35028 33552 -35012
rect 33448 -35092 33468 -35028
rect 33532 -35092 33552 -35028
rect 33448 -35108 33552 -35092
rect 33448 -35172 33468 -35108
rect 33532 -35172 33552 -35108
rect 33448 -35188 33552 -35172
rect 33448 -35252 33468 -35188
rect 33532 -35252 33552 -35188
rect 33448 -35268 33552 -35252
rect 33448 -35332 33468 -35268
rect 33532 -35332 33552 -35268
rect 33448 -35348 33552 -35332
rect 33448 -35412 33468 -35348
rect 33532 -35412 33552 -35348
rect 33448 -35428 33552 -35412
rect 33448 -35492 33468 -35428
rect 33532 -35492 33552 -35428
rect 33448 -35508 33552 -35492
rect 33448 -35572 33468 -35508
rect 33532 -35572 33552 -35508
rect 33448 -35588 33552 -35572
rect 33448 -35652 33468 -35588
rect 33532 -35652 33552 -35588
rect 33448 -35668 33552 -35652
rect 33448 -35732 33468 -35668
rect 33532 -35732 33552 -35668
rect 33448 -35748 33552 -35732
rect 33448 -35812 33468 -35748
rect 33532 -35812 33552 -35748
rect 33448 -35828 33552 -35812
rect 33448 -35892 33468 -35828
rect 33532 -35892 33552 -35828
rect 33448 -35908 33552 -35892
rect 33448 -35972 33468 -35908
rect 33532 -35972 33552 -35908
rect 33448 -35988 33552 -35972
rect 33448 -36052 33468 -35988
rect 33532 -36052 33552 -35988
rect 33448 -36068 33552 -36052
rect 33448 -36132 33468 -36068
rect 33532 -36132 33552 -36068
rect 33448 -36148 33552 -36132
rect 33448 -36212 33468 -36148
rect 33532 -36212 33552 -36148
rect 33448 -36228 33552 -36212
rect 33448 -36292 33468 -36228
rect 33532 -36292 33552 -36228
rect 33448 -36308 33552 -36292
rect 33448 -36372 33468 -36308
rect 33532 -36372 33552 -36308
rect 33448 -36388 33552 -36372
rect 33448 -36452 33468 -36388
rect 33532 -36452 33552 -36388
rect 33448 -36468 33552 -36452
rect 33448 -36532 33468 -36468
rect 33532 -36532 33552 -36468
rect 33448 -36548 33552 -36532
rect 33448 -36612 33468 -36548
rect 33532 -36612 33552 -36548
rect 33448 -36628 33552 -36612
rect 33448 -36692 33468 -36628
rect 33532 -36692 33552 -36628
rect 33448 -36708 33552 -36692
rect 33448 -36772 33468 -36708
rect 33532 -36772 33552 -36708
rect 33448 -36788 33552 -36772
rect 33448 -36852 33468 -36788
rect 33532 -36852 33552 -36788
rect 33448 -36868 33552 -36852
rect 33448 -36932 33468 -36868
rect 33532 -36932 33552 -36868
rect 33448 -36948 33552 -36932
rect 33448 -37012 33468 -36948
rect 33532 -37012 33552 -36948
rect 33448 -37028 33552 -37012
rect 27836 -37240 27940 -37092
rect 30668 -37240 30772 -37041
rect 33448 -37092 33468 -37028
rect 33532 -37092 33552 -37028
rect 33871 -32148 38793 -32119
rect 33871 -37012 33900 -32148
rect 38764 -37012 38793 -32148
rect 33871 -37041 38793 -37012
rect 39060 -32132 39080 -32068
rect 39144 -32132 39164 -32068
rect 39060 -32148 39164 -32132
rect 39060 -32212 39080 -32148
rect 39144 -32212 39164 -32148
rect 39060 -32228 39164 -32212
rect 39060 -32292 39080 -32228
rect 39144 -32292 39164 -32228
rect 39060 -32308 39164 -32292
rect 39060 -32372 39080 -32308
rect 39144 -32372 39164 -32308
rect 39060 -32388 39164 -32372
rect 39060 -32452 39080 -32388
rect 39144 -32452 39164 -32388
rect 39060 -32468 39164 -32452
rect 39060 -32532 39080 -32468
rect 39144 -32532 39164 -32468
rect 39060 -32548 39164 -32532
rect 39060 -32612 39080 -32548
rect 39144 -32612 39164 -32548
rect 39060 -32628 39164 -32612
rect 39060 -32692 39080 -32628
rect 39144 -32692 39164 -32628
rect 39060 -32708 39164 -32692
rect 39060 -32772 39080 -32708
rect 39144 -32772 39164 -32708
rect 39060 -32788 39164 -32772
rect 39060 -32852 39080 -32788
rect 39144 -32852 39164 -32788
rect 39060 -32868 39164 -32852
rect 39060 -32932 39080 -32868
rect 39144 -32932 39164 -32868
rect 39060 -32948 39164 -32932
rect 39060 -33012 39080 -32948
rect 39144 -33012 39164 -32948
rect 39060 -33028 39164 -33012
rect 39060 -33092 39080 -33028
rect 39144 -33092 39164 -33028
rect 39060 -33108 39164 -33092
rect 39060 -33172 39080 -33108
rect 39144 -33172 39164 -33108
rect 39060 -33188 39164 -33172
rect 39060 -33252 39080 -33188
rect 39144 -33252 39164 -33188
rect 39060 -33268 39164 -33252
rect 39060 -33332 39080 -33268
rect 39144 -33332 39164 -33268
rect 39060 -33348 39164 -33332
rect 39060 -33412 39080 -33348
rect 39144 -33412 39164 -33348
rect 39060 -33428 39164 -33412
rect 39060 -33492 39080 -33428
rect 39144 -33492 39164 -33428
rect 39060 -33508 39164 -33492
rect 39060 -33572 39080 -33508
rect 39144 -33572 39164 -33508
rect 39060 -33588 39164 -33572
rect 39060 -33652 39080 -33588
rect 39144 -33652 39164 -33588
rect 39060 -33668 39164 -33652
rect 39060 -33732 39080 -33668
rect 39144 -33732 39164 -33668
rect 39060 -33748 39164 -33732
rect 39060 -33812 39080 -33748
rect 39144 -33812 39164 -33748
rect 39060 -33828 39164 -33812
rect 39060 -33892 39080 -33828
rect 39144 -33892 39164 -33828
rect 39060 -33908 39164 -33892
rect 39060 -33972 39080 -33908
rect 39144 -33972 39164 -33908
rect 39060 -33988 39164 -33972
rect 39060 -34052 39080 -33988
rect 39144 -34052 39164 -33988
rect 39060 -34068 39164 -34052
rect 39060 -34132 39080 -34068
rect 39144 -34132 39164 -34068
rect 39060 -34148 39164 -34132
rect 39060 -34212 39080 -34148
rect 39144 -34212 39164 -34148
rect 39060 -34228 39164 -34212
rect 39060 -34292 39080 -34228
rect 39144 -34292 39164 -34228
rect 39060 -34308 39164 -34292
rect 39060 -34372 39080 -34308
rect 39144 -34372 39164 -34308
rect 39060 -34388 39164 -34372
rect 39060 -34452 39080 -34388
rect 39144 -34452 39164 -34388
rect 39060 -34468 39164 -34452
rect 39060 -34532 39080 -34468
rect 39144 -34532 39164 -34468
rect 39060 -34548 39164 -34532
rect 39060 -34612 39080 -34548
rect 39144 -34612 39164 -34548
rect 39060 -34628 39164 -34612
rect 39060 -34692 39080 -34628
rect 39144 -34692 39164 -34628
rect 39060 -34708 39164 -34692
rect 39060 -34772 39080 -34708
rect 39144 -34772 39164 -34708
rect 39060 -34788 39164 -34772
rect 39060 -34852 39080 -34788
rect 39144 -34852 39164 -34788
rect 39060 -34868 39164 -34852
rect 39060 -34932 39080 -34868
rect 39144 -34932 39164 -34868
rect 39060 -34948 39164 -34932
rect 39060 -35012 39080 -34948
rect 39144 -35012 39164 -34948
rect 39060 -35028 39164 -35012
rect 39060 -35092 39080 -35028
rect 39144 -35092 39164 -35028
rect 39060 -35108 39164 -35092
rect 39060 -35172 39080 -35108
rect 39144 -35172 39164 -35108
rect 39060 -35188 39164 -35172
rect 39060 -35252 39080 -35188
rect 39144 -35252 39164 -35188
rect 39060 -35268 39164 -35252
rect 39060 -35332 39080 -35268
rect 39144 -35332 39164 -35268
rect 39060 -35348 39164 -35332
rect 39060 -35412 39080 -35348
rect 39144 -35412 39164 -35348
rect 39060 -35428 39164 -35412
rect 39060 -35492 39080 -35428
rect 39144 -35492 39164 -35428
rect 39060 -35508 39164 -35492
rect 39060 -35572 39080 -35508
rect 39144 -35572 39164 -35508
rect 39060 -35588 39164 -35572
rect 39060 -35652 39080 -35588
rect 39144 -35652 39164 -35588
rect 39060 -35668 39164 -35652
rect 39060 -35732 39080 -35668
rect 39144 -35732 39164 -35668
rect 39060 -35748 39164 -35732
rect 39060 -35812 39080 -35748
rect 39144 -35812 39164 -35748
rect 39060 -35828 39164 -35812
rect 39060 -35892 39080 -35828
rect 39144 -35892 39164 -35828
rect 39060 -35908 39164 -35892
rect 39060 -35972 39080 -35908
rect 39144 -35972 39164 -35908
rect 39060 -35988 39164 -35972
rect 39060 -36052 39080 -35988
rect 39144 -36052 39164 -35988
rect 39060 -36068 39164 -36052
rect 39060 -36132 39080 -36068
rect 39144 -36132 39164 -36068
rect 39060 -36148 39164 -36132
rect 39060 -36212 39080 -36148
rect 39144 -36212 39164 -36148
rect 39060 -36228 39164 -36212
rect 39060 -36292 39080 -36228
rect 39144 -36292 39164 -36228
rect 39060 -36308 39164 -36292
rect 39060 -36372 39080 -36308
rect 39144 -36372 39164 -36308
rect 39060 -36388 39164 -36372
rect 39060 -36452 39080 -36388
rect 39144 -36452 39164 -36388
rect 39060 -36468 39164 -36452
rect 39060 -36532 39080 -36468
rect 39144 -36532 39164 -36468
rect 39060 -36548 39164 -36532
rect 39060 -36612 39080 -36548
rect 39144 -36612 39164 -36548
rect 39060 -36628 39164 -36612
rect 39060 -36692 39080 -36628
rect 39144 -36692 39164 -36628
rect 39060 -36708 39164 -36692
rect 39060 -36772 39080 -36708
rect 39144 -36772 39164 -36708
rect 39060 -36788 39164 -36772
rect 39060 -36852 39080 -36788
rect 39144 -36852 39164 -36788
rect 39060 -36868 39164 -36852
rect 39060 -36932 39080 -36868
rect 39144 -36932 39164 -36868
rect 39060 -36948 39164 -36932
rect 39060 -37012 39080 -36948
rect 39144 -37012 39164 -36948
rect 39060 -37028 39164 -37012
rect 33448 -37240 33552 -37092
rect 36280 -37240 36384 -37041
rect 39060 -37092 39080 -37028
rect 39144 -37092 39164 -37028
rect 39060 -37240 39164 -37092
<< properties >>
string FIXED_BBOX 33792 32040 38872 37120
<< end >>
