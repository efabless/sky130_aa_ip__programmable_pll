magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect 0 322 1209 587
rect 1040 314 1208 322
rect -101 5 1 258
rect 1491 211 1496 329
rect 94 5 194 38
rect 252 5 352 37
rect 410 5 510 40
rect 568 5 668 40
rect 856 9 955 44
rect 1014 9 1113 49
rect 1208 9 1496 211
rect 761 5 1496 9
rect -341 -125 -340 -6
rect -101 -66 1496 5
rect -101 -389 1 -66
rect 94 -104 194 -66
rect 252 -105 352 -66
rect 410 -102 510 -66
rect 568 -102 668 -66
rect 856 -108 955 -66
rect 1014 -103 1113 -66
rect 1208 -390 1491 -66
<< pwell >>
rect -323 -2079 1428 -1936
<< psubdiff >>
rect -297 -1991 1402 -1962
rect -297 -2025 -257 -1991
rect -223 -2025 -189 -1991
rect -155 -2025 -121 -1991
rect -87 -2025 -53 -1991
rect -19 -2025 15 -1991
rect 49 -2025 83 -1991
rect 117 -2025 151 -1991
rect 185 -2025 219 -1991
rect 253 -2025 287 -1991
rect 321 -2025 355 -1991
rect 389 -2025 423 -1991
rect 457 -2025 491 -1991
rect 525 -2025 559 -1991
rect 593 -2025 627 -1991
rect 661 -2025 695 -1991
rect 729 -2025 763 -1991
rect 797 -2025 831 -1991
rect 865 -2025 899 -1991
rect 933 -2025 967 -1991
rect 1001 -2025 1035 -1991
rect 1069 -2025 1103 -1991
rect 1137 -2025 1171 -1991
rect 1205 -2025 1239 -1991
rect 1273 -2025 1307 -1991
rect 1341 -2025 1402 -1991
rect -297 -2053 1402 -2025
<< nsubdiff >>
rect 50 517 1118 551
rect 50 483 106 517
rect 140 483 174 517
rect 208 483 242 517
rect 276 483 310 517
rect 344 483 378 517
rect 412 483 446 517
rect 480 483 514 517
rect 548 483 582 517
rect 616 483 650 517
rect 684 483 718 517
rect 752 483 786 517
rect 820 483 854 517
rect 888 483 922 517
rect 956 483 990 517
rect 1024 483 1118 517
rect 50 452 1118 483
<< psubdiffcont >>
rect -257 -2025 -223 -1991
rect -189 -2025 -155 -1991
rect -121 -2025 -87 -1991
rect -53 -2025 -19 -1991
rect 15 -2025 49 -1991
rect 83 -2025 117 -1991
rect 151 -2025 185 -1991
rect 219 -2025 253 -1991
rect 287 -2025 321 -1991
rect 355 -2025 389 -1991
rect 423 -2025 457 -1991
rect 491 -2025 525 -1991
rect 559 -2025 593 -1991
rect 627 -2025 661 -1991
rect 695 -2025 729 -1991
rect 763 -2025 797 -1991
rect 831 -2025 865 -1991
rect 899 -2025 933 -1991
rect 967 -2025 1001 -1991
rect 1035 -2025 1069 -1991
rect 1103 -2025 1137 -1991
rect 1171 -2025 1205 -1991
rect 1239 -2025 1273 -1991
rect 1307 -2025 1341 -1991
<< nsubdiffcont >>
rect 106 483 140 517
rect 174 483 208 517
rect 242 483 276 517
rect 310 483 344 517
rect 378 483 412 517
rect 446 483 480 517
rect 514 483 548 517
rect 582 483 616 517
rect 650 483 684 517
rect 718 483 752 517
rect 786 483 820 517
rect 854 483 888 517
rect 922 483 956 517
rect 990 483 1024 517
<< poly >>
rect 10 386 194 407
rect 10 352 24 386
rect 58 385 194 386
rect 58 352 102 385
rect 10 351 102 352
rect 136 351 194 385
rect 10 315 194 351
rect -340 292 -147 311
rect -340 290 -212 292
rect -340 256 -288 290
rect -254 258 -212 290
rect -178 258 -147 292
rect 94 274 194 315
rect 1014 372 1208 400
rect 1014 338 1066 372
rect 1100 338 1146 372
rect 1180 338 1208 372
rect 1014 314 1208 338
rect 1298 380 1444 401
rect 1298 346 1311 380
rect 1345 346 1386 380
rect 1420 346 1444 380
rect 1298 328 1444 346
rect 1014 292 1114 314
rect 1298 293 1398 328
rect -254 256 -147 258
rect -340 242 -147 256
rect -294 221 -194 242
rect 856 43 955 44
rect 94 -18 194 38
rect 252 -18 352 37
rect 410 -18 510 40
rect 568 -18 668 40
rect 856 -18 956 43
rect 1288 16 1412 50
rect -294 -105 -194 -29
rect 94 -70 956 -18
rect 94 -104 194 -70
rect 252 -105 352 -70
rect 410 -102 510 -70
rect 568 -102 668 -70
rect 856 -101 956 -70
rect 1014 -21 1232 -4
rect 1014 -27 1132 -21
rect 1014 -61 1042 -27
rect 1076 -55 1132 -27
rect 1166 -55 1232 -21
rect 1076 -61 1232 -55
rect 1014 -73 1232 -61
rect 1303 -68 1400 16
rect 856 -108 955 -101
rect 1014 -104 1114 -73
rect 1290 -102 1414 -68
rect 239 -579 931 -524
rect 239 -633 497 -579
rect 831 -631 931 -579
rect 890 -865 931 -863
rect -199 -1086 -99 -878
rect 81 -904 181 -870
rect 81 -938 116 -904
rect 150 -938 181 -904
rect 81 -950 181 -938
rect 554 -907 655 -874
rect 554 -941 577 -907
rect 611 -941 655 -907
rect 831 -909 931 -865
rect 554 -954 655 -941
rect 728 -950 931 -909
rect 1107 -937 1207 -879
rect 728 -997 769 -950
rect 1060 -957 1237 -937
rect 1060 -958 1174 -957
rect 1060 -992 1087 -958
rect 1121 -991 1174 -958
rect 1208 -991 1237 -957
rect 1121 -992 1237 -991
rect 81 -1038 769 -997
rect 831 -1019 931 -992
rect 1060 -1017 1237 -992
rect 81 -1109 181 -1038
rect 555 -1109 655 -1038
rect 831 -1053 871 -1019
rect 905 -1053 931 -1019
rect 831 -1081 931 -1053
rect 1106 -1082 1206 -1017
rect -199 -1330 -99 -1328
rect -211 -1348 -53 -1330
rect -211 -1382 -190 -1348
rect -156 -1382 -109 -1348
rect -75 -1382 -53 -1348
rect -211 -1401 -53 -1382
rect 81 -1416 181 -1323
rect -12 -1430 181 -1416
rect -12 -1464 8 -1430
rect 42 -1464 89 -1430
rect 123 -1464 181 -1430
rect -12 -1471 181 -1464
rect 239 -1443 497 -1328
rect 831 -1443 931 -1331
rect -12 -1486 152 -1471
rect 239 -1476 931 -1443
rect -524 -1535 -332 -1521
rect -524 -1536 -406 -1535
rect -524 -1570 -491 -1536
rect -457 -1569 -406 -1536
rect -372 -1569 -332 -1535
rect -457 -1570 -332 -1569
rect -524 -1593 -332 -1570
rect -206 -1592 1316 -1551
rect -280 -1854 -106 -1836
rect -294 -1875 -106 -1854
rect -294 -1909 -272 -1875
rect -238 -1876 -106 -1875
rect -238 -1909 -195 -1876
rect -294 -1910 -195 -1909
rect -161 -1899 -106 -1876
rect 1454 -1861 1634 -1836
rect 1454 -1864 1565 -1861
rect 1454 -1898 1474 -1864
rect 1508 -1895 1565 -1864
rect 1599 -1895 1634 -1861
rect 1508 -1898 1634 -1895
rect -161 -1910 -141 -1899
rect -294 -1928 -141 -1910
rect 1454 -1914 1634 -1898
<< polycont >>
rect 24 352 58 386
rect 102 351 136 385
rect -288 256 -254 290
rect -212 258 -178 292
rect 1066 338 1100 372
rect 1146 338 1180 372
rect 1311 346 1345 380
rect 1386 346 1420 380
rect 1042 -61 1076 -27
rect 1132 -55 1166 -21
rect 116 -938 150 -904
rect 577 -941 611 -907
rect 1087 -992 1121 -958
rect 1174 -991 1208 -957
rect 871 -1053 905 -1019
rect -190 -1382 -156 -1348
rect -109 -1382 -75 -1348
rect 8 -1464 42 -1430
rect 89 -1464 123 -1430
rect -491 -1570 -457 -1536
rect -406 -1569 -372 -1535
rect -272 -1909 -238 -1875
rect -195 -1910 -161 -1876
rect 1474 -1898 1508 -1864
rect 1565 -1895 1599 -1861
<< locali >>
rect 71 519 1072 532
rect -340 517 1072 519
rect -340 485 106 517
rect -340 311 -306 485
rect 71 483 106 485
rect 140 483 174 517
rect 208 483 242 517
rect 276 483 310 517
rect 344 483 378 517
rect 412 483 446 517
rect 480 483 514 517
rect 548 483 582 517
rect 616 483 650 517
rect 684 483 718 517
rect 752 483 786 517
rect 820 483 854 517
rect 888 483 922 517
rect 956 483 990 517
rect 1024 514 1072 517
rect 1024 483 1444 514
rect 71 480 1444 483
rect 71 467 1072 480
rect 2 386 158 407
rect 275 388 316 467
rect 671 388 712 467
rect 1410 401 1444 480
rect 2 384 24 386
rect -53 352 24 384
rect 58 385 158 386
rect 58 352 102 385
rect -53 351 102 352
rect 136 351 158 385
rect -53 345 158 351
rect 2 330 158 345
rect 206 354 1002 388
rect -340 292 -147 311
rect -340 290 -212 292
rect -340 256 -288 290
rect -254 258 -212 290
rect -178 258 -147 292
rect 206 264 240 354
rect 522 264 556 354
rect 968 262 1002 354
rect 1040 372 1208 400
rect 1040 338 1066 372
rect 1100 338 1146 372
rect 1180 338 1208 372
rect 1040 314 1208 338
rect 1298 380 1444 401
rect 1298 346 1311 380
rect 1345 346 1386 380
rect 1420 346 1444 380
rect 1298 328 1444 346
rect 1410 269 1444 328
rect -254 256 -147 258
rect -340 242 -147 256
rect -340 196 -306 242
rect -182 200 -148 242
rect 48 24 82 60
rect 680 24 714 61
rect 1126 24 1160 65
rect -340 -125 -306 -6
rect -182 -124 -148 -7
rect -61 -17 1742 24
rect -61 -505 -20 -17
rect 364 -126 398 -17
rect 810 -125 844 -17
rect 1014 -21 1742 -17
rect 1014 -27 1132 -21
rect 1014 -61 1042 -27
rect 1076 -55 1132 -27
rect 1166 -55 1742 -21
rect 1076 -61 1742 -55
rect 1014 -73 1742 -61
rect 1745 -373 1786 -350
rect 1199 -387 1786 -373
rect 1199 -391 1297 -387
rect 1199 -425 1212 -391
rect 1246 -421 1297 -391
rect 1331 -421 1786 -387
rect 1246 -425 1786 -421
rect 1199 -439 1786 -425
rect -61 -511 1009 -505
rect -554 -549 1009 -511
rect -929 -807 -611 -789
rect -994 -824 -611 -807
rect -994 -858 -908 -824
rect -874 -825 -611 -824
rect -874 -858 -730 -825
rect -994 -859 -730 -858
rect -696 -859 -611 -825
rect -994 -872 -611 -859
rect -929 -889 -611 -872
rect -554 -1023 -516 -549
rect -61 -580 1009 -549
rect -61 -596 69 -580
rect 35 -652 69 -596
rect 667 -654 701 -580
rect -406 -789 -334 -760
rect -406 -823 -393 -789
rect -359 -823 -334 -789
rect -406 -872 -334 -823
rect -406 -906 -392 -872
rect -358 -906 -334 -872
rect -406 -910 -334 -906
rect 98 -904 169 -900
rect 98 -910 116 -904
rect -406 -938 116 -910
rect 150 -910 169 -904
rect 558 -907 636 -899
rect 558 -910 577 -907
rect 150 -938 577 -910
rect -406 -941 577 -938
rect 611 -910 636 -907
rect 611 -941 972 -910
rect 1061 -937 1095 -862
rect 1219 -937 1253 -860
rect -406 -977 972 -941
rect 1040 -957 1275 -937
rect 1040 -958 1174 -957
rect 855 -1019 924 -977
rect 1040 -992 1087 -958
rect 1121 -991 1174 -958
rect 1208 -991 1275 -957
rect 1121 -992 1275 -991
rect 1040 -1018 1275 -992
rect 1310 -938 1385 -926
rect 1310 -972 1329 -938
rect 1363 -972 1385 -938
rect -554 -1060 819 -1023
rect 351 -1104 385 -1060
rect 785 -1118 819 -1060
rect 855 -1053 871 -1019
rect 905 -1053 924 -1019
rect 855 -1071 924 -1053
rect 1060 -1103 1094 -1018
rect 1218 -1104 1252 -1018
rect 1310 -1023 1385 -972
rect 1310 -1057 1329 -1023
rect 1363 -1057 1385 -1023
rect 1310 -1074 1385 -1057
rect -87 -1309 -53 -1306
rect -245 -1348 -53 -1309
rect 35 -1345 69 -1307
rect 667 -1345 701 -1309
rect 1329 -1345 1366 -1074
rect -245 -1382 -190 -1348
rect -156 -1382 -109 -1348
rect -75 -1382 -53 -1348
rect 8 -1382 1366 -1345
rect -245 -1392 -53 -1382
rect -12 -1428 152 -1416
rect -985 -1430 152 -1428
rect -985 -1464 8 -1430
rect 42 -1464 89 -1430
rect 123 -1464 152 -1430
rect -985 -1469 152 -1464
rect -12 -1486 152 -1469
rect -524 -1535 -332 -1521
rect -524 -1536 -406 -1535
rect -524 -1570 -491 -1536
rect -457 -1569 -406 -1536
rect -372 -1569 -332 -1535
rect -457 -1570 -332 -1569
rect -524 -1593 -332 -1570
rect -524 -1615 -490 -1593
rect -366 -1618 -332 -1593
rect -524 -1986 -490 -1822
rect -294 -1873 -141 -1854
rect -332 -1875 -141 -1873
rect -332 -1909 -272 -1875
rect -238 -1876 -141 -1875
rect -238 -1909 -195 -1876
rect -332 -1910 -195 -1909
rect -161 -1910 -141 -1876
rect -332 -1916 -141 -1910
rect -294 -1928 -141 -1916
rect -94 -1977 -60 -1817
rect 222 -1977 256 -1819
rect 538 -1977 572 -1817
rect 854 -1977 888 -1817
rect 1170 -1977 1204 -1817
rect 1445 -1836 1479 -1818
rect 1603 -1836 1637 -1818
rect 1445 -1861 1637 -1836
rect 1445 -1864 1565 -1861
rect 1445 -1898 1474 -1864
rect 1508 -1895 1565 -1864
rect 1599 -1895 1637 -1861
rect 1508 -1898 1637 -1895
rect 1445 -1927 1637 -1898
rect 1528 -1977 1586 -1927
rect -280 -1986 1586 -1977
rect -524 -1991 1586 -1986
rect -524 -2020 -257 -1991
rect -280 -2025 -257 -2020
rect -223 -2025 -189 -1991
rect -155 -2025 -121 -1991
rect -87 -2025 -53 -1991
rect -19 -2025 15 -1991
rect 49 -2025 83 -1991
rect 117 -2025 151 -1991
rect 185 -2025 219 -1991
rect 253 -2025 287 -1991
rect 321 -2025 355 -1991
rect 389 -2025 423 -1991
rect 457 -2025 491 -1991
rect 525 -2025 559 -1991
rect 593 -2025 627 -1991
rect 661 -2025 695 -1991
rect 729 -2025 763 -1991
rect 797 -2025 831 -1991
rect 865 -2025 899 -1991
rect 933 -2025 967 -1991
rect 1001 -2025 1035 -1991
rect 1069 -2025 1103 -1991
rect 1137 -2025 1171 -1991
rect 1205 -2025 1239 -1991
rect 1273 -2025 1307 -1991
rect 1341 -2025 1586 -1991
rect -280 -2035 1586 -2025
<< viali >>
rect 1066 338 1100 372
rect 1146 338 1180 372
rect 1212 -425 1246 -391
rect 1297 -421 1331 -387
rect -908 -858 -874 -824
rect -730 -859 -696 -825
rect -393 -823 -359 -789
rect -392 -906 -358 -872
rect 1329 -972 1363 -938
rect 1329 -1057 1363 -1023
<< metal1 >>
rect 1130 384 1208 400
rect 1014 372 1208 384
rect 1014 358 1066 372
rect -45 338 1066 358
rect 1100 338 1146 372
rect 1180 338 1208 372
rect -45 329 1208 338
rect -45 -390 -7 329
rect 358 261 404 329
rect 804 266 850 329
rect 200 -128 246 65
rect 516 -128 562 65
rect 962 -128 1008 93
rect 1246 5 1292 68
rect 1404 5 1450 68
rect 1225 -41 1485 5
rect 1250 -128 1296 -41
rect 1408 -129 1454 -41
rect 42 -390 88 -305
rect 674 -390 720 -323
rect 1120 -388 1166 -325
rect 1199 -387 1354 -373
rect 1199 -388 1297 -387
rect 1120 -390 1297 -388
rect -45 -391 1297 -390
rect -45 -425 1212 -391
rect 1246 -421 1297 -391
rect 1331 -421 1354 -387
rect 1246 -425 1354 -421
rect -45 -427 1354 -425
rect -45 -499 1155 -427
rect 1199 -439 1354 -427
rect 345 -658 391 -499
rect 779 -656 825 -499
rect 1063 -569 1385 -499
rect -406 -789 -334 -760
rect -929 -809 -611 -789
rect -406 -809 -393 -789
rect -929 -823 -393 -809
rect -359 -823 -334 -789
rect -929 -824 -334 -823
rect -929 -858 -908 -824
rect -874 -825 -334 -824
rect -874 -858 -730 -825
rect -929 -859 -730 -858
rect -696 -859 -334 -825
rect -929 -872 -334 -859
rect -929 -874 -392 -872
rect -929 -889 -611 -874
rect -406 -906 -392 -874
rect -358 -906 -334 -872
rect -406 -929 -334 -906
rect -251 -1109 -205 -850
rect -93 -1107 -47 -831
rect 187 -1106 233 -856
rect 503 -1106 549 -856
rect 937 -1106 983 -856
rect 1310 -938 1385 -569
rect 1310 -972 1329 -938
rect 1363 -972 1385 -938
rect 1310 -1023 1385 -972
rect 1310 -1057 1329 -1023
rect 1363 -1057 1385 -1023
rect 1310 -1074 1385 -1057
rect -251 -1397 -205 -1299
rect -372 -1443 -205 -1397
rect 187 -1425 233 -1302
rect 503 -1425 549 -1299
rect 937 -1425 983 -1298
rect -372 -1619 -326 -1443
rect 1 -1471 995 -1425
rect 1212 -1426 1258 -1300
rect 186 -1551 232 -1471
rect 503 -1551 549 -1471
rect 934 -1551 980 -1471
rect 1212 -1472 1485 -1426
rect -261 -1580 1374 -1551
rect -258 -1617 -212 -1580
rect 58 -1617 104 -1580
rect 186 -1584 232 -1580
rect 374 -1616 420 -1580
rect 690 -1617 736 -1580
rect 1006 -1617 1052 -1580
rect 1322 -1617 1368 -1580
rect 1439 -1619 1485 -1472
use sky130_fd_pr__nfet_01v8_N7QDUL  sky130_fd_pr__nfet_01v8_N7QDUL_0 paramcells
timestamp 1726359333
transform 1 0 555 0 1 -1716
box -845 -126 845 126
use sky130_fd_pr__nfet_01v8_QAG9NA  sky130_fd_pr__nfet_01v8_QAG9NA_0 paramcells
timestamp 1726359333
transform 1 0 881 0 1 -1206
box -134 -126 134 126
use sky130_fd_pr__nfet_01v8_QAG9NA  sky130_fd_pr__nfet_01v8_QAG9NA_1
timestamp 1726359333
transform 1 0 881 0 1 -756
box -134 -126 134 126
use sky130_fd_pr__nfet_01v8_QAG9NA  sky130_fd_pr__nfet_01v8_QAG9NA_2
timestamp 1726359333
transform 1 0 1156 0 1 -1206
box -134 -126 134 126
use sky130_fd_pr__nfet_01v8_QAG9NA  sky130_fd_pr__nfet_01v8_QAG9NA_3
timestamp 1726359333
transform 1 0 1157 0 1 -758
box -134 -126 134 126
use sky130_fd_pr__nfet_01v8_QAG9NA  sky130_fd_pr__nfet_01v8_QAG9NA_4
timestamp 1726359333
transform 1 0 -149 0 1 -754
box -134 -126 134 126
use sky130_fd_pr__nfet_01v8_QAG9NA  sky130_fd_pr__nfet_01v8_QAG9NA_5
timestamp 1726359333
transform 1 0 -149 0 1 -1206
box -134 -126 134 126
use sky130_fd_pr__nfet_01v8_QAG9NA  sky130_fd_pr__nfet_01v8_QAG9NA_6
timestamp 1726359333
transform 1 0 1541 0 1 -1716
box -134 -126 134 126
use sky130_fd_pr__nfet_01v8_QAG9NA  sky130_fd_pr__nfet_01v8_QAG9NA_7
timestamp 1726359333
transform 1 0 -428 0 1 -1718
box -134 -126 134 126
use sky130_fd_pr__nfet_01v8_SMD9NL  sky130_fd_pr__nfet_01v8_SMD9NL_0 paramcells
timestamp 1726359333
transform 1 0 368 0 1 -1206
box -371 -126 371 126
use sky130_fd_pr__nfet_01v8_SMD9NL  sky130_fd_pr__nfet_01v8_SMD9NL_1
timestamp 1726359333
transform 1 0 368 0 1 -756
box -371 -126 371 126
use sky130_fd_pr__pfet_01v8_ES6JVF  sky130_fd_pr__pfet_01v8_ES6JVF_0 paramcells
timestamp 1726359333
transform 1 0 -244 0 1 -227
box -144 -162 144 162
use sky130_fd_pr__pfet_01v8_ES6JVF  sky130_fd_pr__pfet_01v8_ES6JVF_1
timestamp 1726359333
transform 1 0 1348 0 1 167
box -144 -162 144 162
use sky130_fd_pr__pfet_01v8_ES6JVF  sky130_fd_pr__pfet_01v8_ES6JVF_2
timestamp 1726359333
transform 1 0 -244 0 1 96
box -144 -162 144 162
use sky130_fd_pr__pfet_01v8_ES6JVF  sky130_fd_pr__pfet_01v8_ES6JVF_3
timestamp 1726359333
transform 1 0 1352 0 1 -228
box -144 -162 144 162
use sky130_fd_pr__pfet_01v8_ES28UG  sky130_fd_pr__pfet_01v8_ES28UG_0 paramcells
timestamp 1726359333
transform 1 0 381 0 1 -227
box -381 -162 381 162
use sky130_fd_pr__pfet_01v8_ES28UG  sky130_fd_pr__pfet_01v8_ES28UG_1
timestamp 1726359333
transform 1 0 381 0 1 162
box -381 -162 381 162
use sky130_fd_pr__pfet_01v8_ESSCXF  sky130_fd_pr__pfet_01v8_ESSCXF_0 paramcells
timestamp 1726359333
transform 1 0 985 0 1 167
box -223 -162 223 162
use sky130_fd_pr__pfet_01v8_ESSCXF  sky130_fd_pr__pfet_01v8_ESSCXF_1
timestamp 1726359333
transform 1 0 985 0 1 -227
box -223 -162 223 162
<< labels >>
flabel locali s 1735 3 1735 3 0 FreeSans 1250 0 0 0 OUT
flabel locali s 1762 -360 1762 -360 0 FreeSans 1250 0 0 0 OUTB
flabel locali s -972 -1452 -972 -1452 0 FreeSans 1250 0 0 0 INB
flabel locali s 351 -2017 351 -2017 0 FreeSans 1250 0 0 0 VSS
flabel locali s -322 -1894 -322 -1894 0 FreeSans 1250 0 0 0 VCTRL2
flabel locali s 523 509 523 509 0 FreeSans 1250 0 0 0 VDD
flabel locali s -41 370 -41 370 0 FreeSans 1250 0 0 0 VCTRL
flabel locali s -966 -845 -966 -845 0 FreeSans 1250 0 0 0 IN
<< end >>
