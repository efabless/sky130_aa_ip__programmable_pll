magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< pwell >>
rect -4196 1479 -4108 1522
rect -3565 1454 -3532 1497
<< psubdiff >>
rect -4196 1479 -4108 1522
rect -3565 1454 -3532 1497
<< locali >>
rect -4820 43957 -3786 44102
rect -4820 42551 -4707 43957
rect -3915 42551 -3786 43957
rect -4820 42470 -3786 42551
rect -2105 43973 -746 44258
rect -2105 42567 -1815 43973
rect -1023 42567 -746 43973
rect -3742 40415 -2527 40571
rect -3742 39539 -3598 40415
rect -2667 39539 -2527 40415
rect -3742 39356 -2527 39539
rect -16160 8555 -16024 8692
rect -15790 8555 -15654 8720
rect -15496 8555 -15355 8722
rect -16182 8440 -15355 8555
rect -16182 8117 -16077 8440
rect -15564 8210 -15355 8440
rect -15564 8117 -15367 8210
rect -16182 8044 -15367 8117
rect -15205 7856 -15069 8692
rect -19000 7720 -15069 7856
rect -14950 7153 -14814 8692
rect -19851 7017 -14814 7153
rect -14717 5489 -14581 8724
rect -19980 5353 -14581 5489
rect -14717 5310 -14581 5353
rect -14518 4472 -14382 8692
rect -9654 7738 -9468 9038
rect -2105 8544 -746 42567
rect 3428 9172 14566 9807
rect -20516 4336 -14382 4472
rect -13709 7552 -9468 7738
rect -6647 8398 -745 8544
rect -13709 2685 -13523 7552
rect -6647 7393 -6475 8398
rect -5556 7393 -745 8398
rect 3428 8200 4063 9172
rect 14586 8869 14773 8899
rect 14586 8763 14599 8869
rect 14739 8817 14773 8869
rect 14739 8764 15071 8817
rect 14739 8763 14773 8764
rect 6966 8732 7312 8756
rect 14586 8746 14773 8763
rect 6966 8509 7009 8732
rect 7275 8691 7312 8732
rect 15942 8691 15978 8805
rect 16226 8722 16396 8743
rect 7275 8530 16005 8691
rect 16226 8621 16254 8722
rect 16384 8621 16396 8722
rect 16226 8605 16396 8621
rect 7275 8509 7312 8530
rect 6966 8466 7312 8509
rect 7289 8267 7635 8307
rect 3375 8071 4103 8200
rect 3375 7636 3492 8071
rect 3927 7918 4103 8071
rect 7289 8056 7332 8267
rect 7560 8261 7635 8267
rect 16722 8261 16775 8824
rect 26753 8650 38073 8844
rect 7560 8079 16799 8261
rect 7560 8056 7635 8079
rect 7289 8017 7635 8056
rect 3927 7659 8854 7918
rect 14552 7821 14795 7846
rect 14552 7815 16664 7821
rect 14552 7666 14591 7815
rect 14740 7685 16664 7815
rect 14740 7666 14795 7685
rect 3927 7636 4103 7659
rect 14552 7642 14795 7666
rect 3375 7565 4103 7636
rect 26753 7762 27003 8650
rect 37629 7762 38073 8650
rect 26753 7623 38073 7762
rect -6647 7185 -745 7393
rect -12975 6803 -11404 6943
rect -12975 6743 -2388 6803
rect -12975 5686 -12802 6743
rect -11669 6690 -2388 6743
rect -11669 5746 -3482 6690
rect -2539 5746 -2388 6690
rect -11669 5686 -2388 5746
rect -12975 5558 -2388 5686
rect -12975 5372 -11404 5558
rect -2105 4551 -746 7185
rect 19201 6996 19643 7085
rect 14997 6931 15211 6970
rect 19201 6931 19300 6996
rect 14997 6913 19300 6931
rect 14997 6801 15031 6913
rect 15166 6807 19300 6913
rect 15166 6801 15211 6807
rect 14997 6756 15211 6801
rect 19201 6709 19300 6807
rect 19588 6931 19643 6996
rect 22939 6995 23303 7116
rect 22939 6931 23009 6995
rect 19588 6807 23009 6931
rect 19588 6709 19643 6807
rect 16227 6583 16406 6623
rect 19201 6620 19643 6709
rect 22939 6735 23009 6807
rect 23217 6735 23303 6995
rect 22939 6666 23303 6735
rect 16227 6562 16261 6583
rect 12164 6481 16261 6562
rect 16370 6481 16406 6583
rect 12164 6480 16406 6481
rect 16227 6444 16406 6480
rect 14443 6192 14691 6213
rect 14443 6151 14484 6192
rect 12023 6047 14484 6151
rect 14639 6047 14691 6192
rect 12023 6038 14691 6047
rect 12023 5692 12136 6038
rect 14443 6016 14691 6038
rect 13866 5937 14130 5964
rect 13866 5898 13908 5937
rect 12465 5734 13908 5898
rect 14090 5734 14130 5937
rect 12465 5641 14130 5734
rect 12470 5556 12504 5641
rect 18791 5539 19168 5573
rect 18791 5255 18835 5539
rect 19139 5255 19168 5539
rect 18791 5216 19168 5255
rect 23929 4733 61121 4741
rect 2866 4551 3250 4560
rect -2197 4480 12654 4551
rect -2197 4186 2911 4480
rect 3195 4186 12654 4480
rect -2197 4085 12654 4186
rect 23929 4322 41705 4733
rect 44546 4367 61121 4733
rect 44546 4322 98798 4367
rect 23929 4290 98798 4322
rect 15817 4168 16331 4171
rect 23929 4168 24380 4290
rect 14819 4127 24380 4168
rect 14819 3748 15869 4127
rect 16252 3748 24380 4127
rect 14819 3717 24380 3748
rect 26583 3817 38866 3886
rect 14819 3692 15270 3717
rect -13207 3577 15270 3692
rect -13207 3529 3558 3577
rect -13207 3359 -13070 3529
rect -9285 3359 3558 3529
rect -13207 3328 3558 3359
rect 3807 3328 15270 3577
rect 21388 3567 21612 3717
rect 26583 3540 26668 3817
rect 38672 3540 38866 3817
rect 26583 3483 38866 3540
rect -13207 3241 15270 3328
rect -5845 2730 -5539 2764
rect -5845 2685 -5811 2730
rect -13709 2548 -5811 2685
rect -5845 2515 -5811 2548
rect -5591 2515 -5539 2730
rect -5845 2483 -5539 2515
rect -2198 2241 -1747 3241
rect 6011 2400 6354 3241
rect 11748 2486 12550 3241
rect 41815 3211 44205 3238
rect 51135 3226 51730 4290
rect 53312 3230 53907 4290
rect 55261 3230 55856 4290
rect 18156 3163 18330 3181
rect 18156 3007 18170 3163
rect 18307 3110 18330 3163
rect 41815 3154 41845 3211
rect 44154 3154 44205 3211
rect 57618 3209 58213 4290
rect 18307 3036 19662 3110
rect 41815 3072 44205 3154
rect 18307 3007 18330 3036
rect 18156 2985 18330 3007
rect 22316 2881 22554 2900
rect 19567 2877 19632 2878
rect 19341 2565 19481 2579
rect 18629 2540 18739 2549
rect 19341 2540 19368 2565
rect 18629 2449 18635 2540
rect 18734 2458 19368 2540
rect 19468 2458 19481 2565
rect 18734 2449 19481 2458
rect 18629 2447 19481 2449
rect 18629 2441 18739 2447
rect 19341 2444 19481 2447
rect 7054 2052 7303 2079
rect 3222 1884 4073 1923
rect 3500 1609 3875 1654
rect 4034 1638 4073 1884
rect 7054 1856 7079 2052
rect 7277 1856 7303 2052
rect 7054 1845 7303 1856
rect 3500 1574 3539 1609
rect -4212 1522 -4099 1535
rect -5642 1514 -5574 1521
rect -22664 1391 -13491 1425
rect -5779 1365 -5761 1514
rect -5593 1365 -5574 1514
rect -4212 1479 -4196 1522
rect -4108 1479 -4099 1522
rect -4212 1461 -4099 1479
rect -5779 1352 -5574 1365
rect -5779 1299 -5642 1352
rect -4187 680 -4102 1461
rect -3565 1454 -3532 1497
rect 2935 1331 3539 1574
rect 3817 1331 3875 1609
rect 3990 1625 4106 1638
rect 3990 1517 4005 1625
rect 4087 1517 4106 1625
rect 4626 1517 4768 1644
rect 7096 1568 7234 1845
rect 15522 1804 15742 1833
rect 15522 1707 15548 1804
rect 7337 1661 7470 1680
rect 15184 1673 15548 1707
rect 7337 1586 7355 1661
rect 7442 1586 7470 1661
rect 15522 1631 15548 1673
rect 15711 1631 15742 1804
rect 15522 1597 15742 1631
rect 7029 1526 7278 1568
rect 7337 1562 7470 1586
rect 3990 1499 4106 1517
rect 2935 1319 3875 1331
rect 3500 1279 3875 1319
rect 4196 1496 4326 1504
rect 4196 1401 4211 1496
rect 4314 1401 4326 1496
rect -6175 595 -4102 680
rect -18039 544 -17604 565
rect -18039 457 -18015 544
rect -22512 346 -18015 457
rect -17624 457 -17604 544
rect -6543 457 -5591 465
rect -17624 444 -5591 457
rect -17624 346 -6513 444
rect -22512 320 -6513 346
rect -6543 312 -6513 320
rect -5616 312 -5591 444
rect -6543 299 -5591 312
rect -3695 212 -3643 1090
rect 3563 1027 3725 1039
rect 3563 978 3581 1027
rect 3231 939 3581 978
rect 3563 901 3581 939
rect 3707 901 3725 1027
rect 3563 885 3725 901
rect -2404 576 -2375 608
rect 4196 595 4326 1401
rect 4600 1494 4817 1517
rect 4600 1409 4620 1494
rect 4785 1409 4817 1494
rect 4600 1392 4817 1409
rect 7029 1380 7096 1526
rect 7253 1380 7278 1526
rect 7029 1334 7278 1380
rect 4415 1243 4467 1266
rect 4388 1218 4549 1243
rect 19567 1242 19632 2800
rect 22316 2725 22360 2881
rect 22516 2725 22554 2881
rect 22316 2711 22554 2725
rect 26688 2858 26963 2876
rect 26688 2849 28014 2858
rect 22376 2297 22532 2711
rect 26688 2685 26714 2849
rect 26932 2685 28014 2849
rect 26688 2669 28014 2685
rect 26688 2653 26963 2669
rect 58711 2553 58930 2597
rect 58711 2484 58755 2553
rect 50510 2422 50749 2467
rect 58493 2450 58755 2484
rect 25061 2326 25333 2372
rect 25061 2297 25084 2326
rect 22376 2141 25084 2297
rect 25061 2124 25084 2141
rect 25279 2124 25333 2326
rect 25061 2085 25333 2124
rect 26111 2145 27166 2273
rect 50510 2243 50542 2422
rect 50721 2243 50749 2422
rect 58711 2386 58755 2450
rect 58904 2386 58930 2553
rect 58711 2334 58930 2386
rect 50510 2215 50749 2243
rect 46637 1940 46961 1997
rect 4388 1086 4409 1218
rect 4532 1086 4549 1218
rect 4388 1066 4549 1086
rect 19404 1241 19736 1242
rect 19404 1182 19770 1241
rect 5730 762 6208 775
rect 5730 698 5743 762
rect 6186 698 6208 762
rect 8203 744 8571 936
rect 9394 744 9762 971
rect 19404 969 19503 1182
rect 19720 969 19770 1182
rect 10640 744 11008 885
rect 12204 744 12572 911
rect 13329 744 13697 920
rect 14498 744 14866 947
rect 19404 943 19770 969
rect 19404 744 19742 943
rect 5730 686 6208 698
rect 8089 595 19742 744
rect -2404 364 -2075 576
rect 3030 382 19742 595
rect -22962 160 -3643 212
rect -3192 35 -2075 364
rect 15818 275 16268 345
rect 5857 272 16268 275
rect 3985 241 4186 265
rect 3985 213 4009 241
rect -1806 100 4009 213
rect -13197 -194 -7163 -135
rect -3192 -153 -2863 35
rect -13197 -393 -13067 -194
rect -7302 -274 -7163 -194
rect -7302 -285 -5720 -274
rect -7302 -357 -6033 -285
rect -5757 -357 -5720 -285
rect -7302 -378 -5720 -357
rect -7302 -393 -7163 -378
rect -13197 -453 -7163 -393
rect -25553 -685 -25165 -654
rect -22114 -677 -5221 -603
rect -25553 -973 -25491 -685
rect -25219 -806 -25165 -685
rect -5976 -806 -5800 -784
rect -25219 -943 -5950 -806
rect -25219 -973 -25165 -943
rect -25553 -1050 -25165 -973
rect -5976 -986 -5950 -943
rect -5822 -986 -5800 -806
rect -5976 -1005 -5800 -986
rect -1806 -1962 -1693 100
rect 3985 92 4009 100
rect 4158 92 4186 241
rect 3985 76 4186 92
rect 5857 182 15862 272
rect 4383 -36 4585 -15
rect -1577 -40 4585 -36
rect -1577 -85 4399 -40
rect -1581 -109 4399 -85
rect -1581 -303 -1561 -109
rect -1357 -175 4399 -109
rect -1357 -303 -1323 -175
rect 4383 -189 4399 -175
rect 4556 -189 4585 -40
rect 5857 -107 5908 182
rect 6180 -107 15862 182
rect 5857 -126 15862 -107
rect 16220 -126 16268 272
rect 21288 224 21541 1919
rect 21915 199 22067 1925
rect 46637 1720 46667 1940
rect 46883 1720 46961 1940
rect 46637 1686 46961 1720
rect 47896 1963 48216 1992
rect 47896 1693 47931 1963
rect 48166 1900 48216 1963
rect 50541 1900 50720 2215
rect 48166 1721 50720 1900
rect 48166 1693 48216 1721
rect 47896 1636 48216 1693
rect 22419 1250 25673 1356
rect 22419 924 22484 1250
rect 22810 924 25673 1250
rect 22419 876 25673 924
rect 51870 824 52157 1672
rect 60670 1398 98798 4290
rect 60670 1310 61121 1398
rect 47592 537 52157 824
rect 53362 859 64533 1310
rect 53362 326 54000 859
rect 54759 326 55397 859
rect 56173 343 56811 859
rect 57259 326 57897 859
rect 5857 -176 16268 -126
rect 4383 -213 4585 -189
rect 5877 -291 6211 -176
rect 8303 -302 8754 -176
rect 9891 -302 10342 -176
rect -1581 -342 -1323 -303
rect 11432 -321 11883 -176
rect 12650 -283 13101 -176
rect 13848 -283 14299 -176
rect 15818 -209 16268 -176
rect 60613 -363 61078 -338
rect 60613 -427 60637 -363
rect 58332 -445 60637 -427
rect 50434 -572 50725 -478
rect 47758 -586 50725 -572
rect 3281 -685 3574 -645
rect 3281 -890 3332 -685
rect 3556 -745 3574 -685
rect 47758 -719 47770 -586
rect 47930 -632 50725 -586
rect 58324 -618 60637 -445
rect 47930 -719 50588 -632
rect 60613 -650 60637 -618
rect 61047 -650 61078 -363
rect 60613 -669 61078 -650
rect 47758 -726 50588 -719
rect 3556 -819 4361 -745
rect 47758 -752 47953 -726
rect 3556 -890 3574 -819
rect 3281 -911 3574 -890
rect 16101 -922 16445 -871
rect 16101 -1021 16127 -922
rect 7334 -1105 7443 -1093
rect 7334 -1190 7348 -1105
rect 7431 -1190 7443 -1105
rect 15047 -1127 16127 -1021
rect 7334 -1207 7443 -1190
rect 16101 -1183 16127 -1127
rect 16382 -1183 16445 -922
rect 16101 -1228 16445 -1183
rect 19836 -1038 20098 -916
rect 19836 -1236 19863 -1038
rect 20055 -1129 20098 -1038
rect 20055 -1236 20093 -1129
rect 19836 -1279 20093 -1236
rect -26391 -2075 -1693 -1962
rect 8336 -1966 8557 -1837
rect 9274 -1966 9547 -1837
rect 10255 -1966 10528 -1871
rect 11457 -1966 11730 -1845
rect 12412 -1966 12685 -1879
rect 13206 -1966 13479 -1845
rect 13931 -1966 14204 -1845
rect 26281 -1966 26638 -1361
rect 4310 -2185 4465 -2171
rect 4310 -2204 4329 -2185
rect -26307 -2295 4329 -2204
rect 4444 -2295 4465 -2185
rect -26307 -2300 4465 -2295
rect 4310 -2309 4465 -2300
rect 8168 -2323 26638 -1966
rect 46864 -1737 47369 -1268
rect 52463 -1737 52968 -1175
rect 55332 -1517 55783 -1516
rect 56669 -1517 57120 -1516
rect 57856 -1517 58307 -1516
rect 64082 -1517 64533 859
rect 46864 -2104 52968 -1737
rect -1585 -2389 -1283 -2369
rect -1585 -2393 -1565 -2389
rect -26253 -2533 -1565 -2393
rect -1585 -2555 -1565 -2533
rect -1322 -2555 -1283 -2389
rect 46864 -2436 46922 -2104
rect 47268 -2242 52968 -2104
rect 53892 -1968 64533 -1517
rect 47268 -2436 47369 -2242
rect 46864 -2515 47369 -2436
rect -1585 -2584 -1283 -2555
rect 3196 -2577 3624 -2539
rect 3196 -2628 3272 -2577
rect -26211 -2865 3272 -2628
rect 3578 -2865 3624 -2577
rect 53892 -2712 54343 -1968
rect 55332 -2712 55783 -1968
rect 56669 -2731 57120 -1968
rect 57856 -2731 58307 -1968
rect 64082 -2655 64533 -1968
rect -26211 -2873 3624 -2865
rect 3196 -2900 3624 -2873
rect 15440 -2934 15853 -2842
rect -26114 -2937 15853 -2934
rect -26114 -3174 15509 -2937
rect 15772 -3174 15853 -2937
rect -26114 -3188 15853 -3174
rect 15440 -3211 15853 -3188
rect 87785 -3270 88210 -3189
rect 87785 -3288 87922 -3270
rect 16088 -3296 16483 -3292
rect -26140 -3330 16483 -3296
rect -26140 -3560 16127 -3330
rect 16439 -3560 16483 -3330
rect 65127 -3352 87922 -3288
rect -26140 -3586 16483 -3560
rect 16088 -3623 16483 -3586
rect 48966 -3400 49277 -3371
rect 48966 -3654 49001 -3400
rect 49228 -3547 49277 -3400
rect 62387 -3378 62911 -3375
rect 62387 -3380 62884 -3378
rect 61873 -3419 62067 -3407
rect 61873 -3432 61891 -3419
rect 58166 -3456 61891 -3432
rect 58163 -3490 61891 -3456
rect 58332 -3498 61891 -3490
rect 62043 -3474 62067 -3419
rect 62387 -3424 62407 -3380
rect 62387 -3428 62884 -3424
rect 62908 -3428 62911 -3378
rect 62387 -3436 62911 -3428
rect 65127 -3454 65203 -3352
rect 65314 -3454 87922 -3352
rect 62043 -3498 62096 -3474
rect 58332 -3508 62096 -3498
rect 65127 -3477 87922 -3454
rect 88155 -3477 88210 -3270
rect 65127 -3507 88210 -3477
rect 61873 -3516 62067 -3508
rect 49228 -3608 50651 -3547
rect 87785 -3581 88210 -3507
rect 49228 -3654 49277 -3608
rect 48966 -3697 49277 -3654
rect 62432 -3819 62779 -3786
rect 62432 -4119 62459 -3819
rect 62739 -4119 62779 -3819
rect 62432 -4139 62779 -4119
rect 17293 -4336 17906 -4235
rect 16975 -4354 17387 -4336
rect -26205 -4748 17387 -4354
rect 17851 -4748 17906 -4336
rect -26205 -4766 17906 -4748
rect 17293 -4848 17906 -4766
rect 46778 -4698 47398 -4670
rect 52571 -4698 53148 -4252
rect 95829 -4698 98798 1398
rect 46778 -4756 92959 -4698
rect 17978 -4983 18468 -4849
rect 17978 -5013 18041 -4983
rect -26311 -5366 18041 -5013
rect 18388 -5366 18468 -4983
rect 46778 -5188 46893 -4756
rect 47282 -4819 92959 -4756
rect 47282 -4968 61311 -4819
rect 61459 -4968 92959 -4819
rect 47282 -5041 92959 -4968
rect 47282 -5188 90356 -5041
rect 46778 -5275 90356 -5188
rect 46778 -5304 47412 -5275
rect -26311 -5399 18468 -5366
rect 17978 -5437 18468 -5399
rect -26321 -6062 18534 -5664
rect -26321 -6098 18704 -6062
rect 18949 -6346 19611 -6293
rect -26653 -6399 19611 -6346
rect -26653 -6756 19096 -6399
rect 19485 -6756 19611 -6399
rect -26653 -6787 19611 -6756
rect 18949 -6850 19611 -6787
rect 19665 -7100 20295 -7025
rect -26746 -7105 20295 -7100
rect -26746 -7533 19761 -7105
rect 20205 -7533 20295 -7105
rect -26746 -7593 20295 -7533
rect 19665 -7634 20295 -7593
rect 70077 -7278 90356 -5275
rect 92687 -7278 92959 -5041
rect 70077 -7667 92959 -7278
rect 95743 -7667 98798 -4698
rect 70077 -7803 73046 -7667
rect 81551 -7803 84520 -7667
rect -31467 -8957 -30570 -8797
rect -31467 -9060 -31403 -8957
rect -34283 -9713 -31403 -9060
rect -31467 -9854 -31403 -9713
rect -30698 -9060 -30570 -8957
rect 58913 -8995 59860 -8831
rect 58913 -9060 59141 -8995
rect -30698 -9713 59141 -9060
rect -30698 -9854 -30570 -9713
rect -31467 -10014 -30570 -9854
rect 58913 -9746 59141 -9713
rect 59762 -9746 59860 -8995
rect 58913 -9909 59860 -9746
rect 60423 -9800 61454 -9617
rect -29173 -9983 -28472 -9982
rect 60423 -9983 60606 -9800
rect -29347 -10522 60606 -9983
rect -29564 -10565 60606 -10522
rect 61337 -10565 61454 -9800
rect -29564 -10681 61454 -10565
rect -29564 -10684 -28286 -10681
rect -29564 -11622 -29386 -10684
rect -28448 -11622 -28286 -10684
rect 60423 -10731 61454 -10681
rect -29564 -11751 -28286 -11622
rect -26907 -11088 -25983 -10980
rect -24373 -11046 -23278 -10959
rect -24373 -11088 -24163 -11046
rect -29173 -12595 -28472 -11751
rect -26907 -11775 -26778 -11088
rect -26091 -11688 -24163 -11088
rect -23436 -11688 -23278 -11046
rect -26091 -11732 -23278 -11688
rect -26091 -11775 -25983 -11732
rect -26907 -11904 -25983 -11775
rect -24373 -11840 -23278 -11732
rect -6611 -11233 -5937 -11153
rect -6611 -11841 -6545 -11233
rect -6016 -11274 -5937 -11233
rect 61366 -11260 62272 -11116
rect 61366 -11274 61603 -11260
rect -6016 -11734 61603 -11274
rect 62208 -11734 62272 -11260
rect -6016 -11839 62272 -11734
rect -6016 -11841 -5937 -11839
rect -6611 -11894 -5937 -11841
rect 61366 -11971 62272 -11839
rect 62246 -12546 63072 -12441
rect -34369 -13296 -28472 -12595
rect -26996 -12580 63072 -12546
rect -26996 -13054 62379 -12580
rect 62984 -13054 63072 -12580
rect 95829 -12668 98798 -7667
rect -26996 -13121 63072 -13054
rect -26996 -13991 -26421 -13121
rect 62246 -13180 63072 -13121
rect -34505 -14566 -26421 -13991
rect -25931 -14188 -24870 -14108
rect -25931 -14334 -7185 -14188
rect -25931 -14763 -25660 -14334
rect -25005 -14763 -7185 -14334
rect -25931 -14808 -7185 -14763
rect -25931 -14876 -24870 -14808
rect -12874 -15031 -7870 -14969
rect -12874 -15176 -12812 -15031
rect -7984 -15176 -7870 -15031
rect -12874 -15238 -7870 -15176
rect -34293 -15952 -15114 -15892
rect -7536 -15913 -7185 -14808
rect 81378 -15816 98798 -12668
rect -34293 -15986 -15075 -15952
rect -34293 -16022 -15114 -15986
rect -14106 -18273 -13756 -16708
rect -11883 -18273 -11533 -16708
rect -9810 -18248 -9410 -16724
rect 81378 -16770 84526 -15816
rect 90329 -17718 91702 -17504
rect 90329 -18041 90543 -17718
rect 88428 -18579 90543 -18041
rect 90329 -18603 90543 -18579
rect 91459 -18603 91702 -17718
rect 90329 -18877 91702 -18603
rect -25664 -22879 -25039 -22779
rect -25664 -23304 -25539 -22879
rect -25139 -22999 -25039 -22879
rect -25139 -23185 -24246 -22999
rect -25139 -23304 -25039 -23185
rect -25664 -23404 -25039 -23304
rect -32565 -28049 -24427 -27913
rect -32538 -28248 -24481 -28112
rect 95829 -28339 98798 -15816
rect -32538 -28481 -24400 -28345
rect -32592 -28736 -24400 -28600
rect -33001 -29027 -24533 -28886
rect -32755 -29321 -24481 -29185
rect -32917 -29691 -24454 -29555
rect 83333 -31308 98798 -28339
rect -32225 -33190 -26140 -32972
rect -26347 -33893 -26140 -33190
rect 83333 -33215 86302 -31308
rect 90604 -34254 92221 -33888
rect 90604 -34632 90878 -34254
rect 88763 -35139 90878 -34632
rect 91794 -35139 92221 -34254
rect 88763 -35170 92221 -35139
rect 90604 -35414 92221 -35170
rect -25408 -35732 -23381 -35460
rect -25408 -36532 -23381 -36260
rect -27604 -37041 -27464 -37004
rect -27604 -41124 -27597 -37041
rect -27494 -37174 -27464 -37041
rect -27494 -37351 -26938 -37174
rect -27494 -37685 -27464 -37351
rect -25408 -37593 -23381 -37321
rect -27494 -37862 -26953 -37685
rect -27494 -38300 -27464 -37862
rect -27494 -38477 -26975 -38300
rect -27494 -39092 -27464 -38477
rect -20537 -38893 -20422 -38680
rect -24450 -39008 -20422 -38893
rect -27494 -39269 -26953 -39092
rect -27494 -39973 -27464 -39269
rect -27494 -40150 -26953 -39973
rect -27494 -40795 -27464 -40150
rect -27494 -40972 -26953 -40795
rect -27494 -41124 -27464 -40972
rect -27604 -41184 -27464 -41124
rect -26388 -41420 -26202 -41401
rect -26388 -44174 -26195 -41420
rect -25977 -42828 -25639 -42789
rect -25977 -43047 -25900 -42828
rect -25681 -42872 -25639 -42828
rect -24450 -42872 -24335 -39008
rect -25681 -42987 -24335 -42872
rect -25681 -43047 -25639 -42987
rect -25977 -43127 -25639 -43047
rect -23728 -44174 -23542 -39590
rect -26388 -44360 -23542 -44174
rect -32434 -44640 -16322 -44504
rect -32450 -44839 -16322 -44703
rect -32458 -45072 -15025 -44936
rect -32482 -45327 -16322 -45191
rect -29580 -46364 -29447 -45411
rect -28280 -46364 -28157 -45411
rect -24214 -45613 -14730 -45477
rect -24214 -45618 -24059 -45613
rect -24214 -45776 -24078 -45618
rect -24214 -45912 -16322 -45776
rect -24214 -46146 -24078 -45912
rect 95829 -46113 98798 -31308
rect -24214 -46282 -16322 -46146
rect -29580 -46390 -28157 -46364
rect -29580 -46526 -16322 -46390
rect 83333 -49082 98798 -46113
rect -32776 -50847 -27886 -50668
rect -28065 -52016 -27886 -50847
rect 83333 -51532 86302 -49082
rect 91309 -52469 92592 -52202
rect 91309 -52743 91488 -52469
rect 89400 -53281 91488 -52743
rect 91309 -53354 91488 -53281
rect 92404 -53354 92592 -52469
rect 91309 -53546 92592 -53354
rect -27203 -54080 -22678 -53808
rect -29448 -54826 -29178 -54761
rect -29448 -58999 -29398 -54826
rect -29235 -54911 -29178 -54826
rect -27217 -54866 -22678 -54594
rect -29235 -55189 -28800 -54911
rect -29235 -56093 -29178 -55189
rect -27203 -55600 -22678 -55328
rect -29235 -56371 -28814 -56093
rect -29235 -57168 -29178 -56371
rect -19804 -57056 -19689 -56823
rect -29235 -57446 -28793 -57168
rect -26527 -57171 -19689 -57056
rect -29235 -58329 -29178 -57446
rect -29235 -58607 -28821 -58329
rect -29235 -58999 -29178 -58607
rect -29448 -59163 -29178 -58999
rect -28147 -62311 -28010 -59815
rect -26527 -60736 -26412 -57171
rect -26896 -60851 -26412 -60736
rect -23096 -62272 -22910 -57701
rect -23449 -62311 -22910 -62272
rect -28147 -62448 -22910 -62311
rect -23449 -62458 -22910 -62448
rect -33062 -62751 -16322 -62615
rect -33463 -62950 -16322 -62814
rect -32991 -63183 -16322 -63047
rect -32976 -63438 -16322 -63302
rect -31679 -63836 -30520 -63625
rect -23846 -63729 -23123 -63588
rect -31679 -64772 -31540 -63836
rect -30673 -64501 -30522 -63836
rect -23846 -63887 -23710 -63729
rect -23846 -64023 -22771 -63887
rect -23846 -64257 -23710 -64023
rect -23846 -64393 -23184 -64257
rect -30673 -64637 -22352 -64501
rect -30673 -64772 -30522 -64637
rect -31679 -64865 -30522 -64772
<< viali >>
rect -4707 42551 -3915 43957
rect -1815 42567 -1023 43973
rect -3598 39539 -2667 40415
rect -16077 8117 -15564 8440
rect -6475 7393 -5556 8398
rect 14599 8763 14739 8869
rect 7009 8509 7275 8732
rect 16254 8621 16384 8722
rect 3492 7636 3927 8071
rect 7332 8056 7560 8267
rect 14591 7666 14740 7815
rect 16664 7621 16961 7884
rect 27003 7762 37629 8650
rect -12802 5686 -11669 6743
rect -3482 5746 -2539 6690
rect 15031 6801 15166 6913
rect 19300 6709 19588 6996
rect 23009 6735 23217 6995
rect 16261 6481 16370 6583
rect 14484 6047 14639 6192
rect 13908 5734 14090 5937
rect 18835 5255 19139 5539
rect 2911 4186 3195 4480
rect 41705 4322 44546 4733
rect 15869 3748 16252 4127
rect -13070 3359 -9285 3529
rect 3558 3328 3807 3577
rect 26668 3540 38672 3817
rect -5811 2515 -5591 2730
rect -13326 2173 -9322 2305
rect 18170 3007 18307 3163
rect 41845 3154 44154 3211
rect 19563 2800 19636 2877
rect 18635 2449 18734 2540
rect 19368 2458 19468 2565
rect 7079 1856 7277 2052
rect -5761 1365 -5593 1514
rect -4196 1479 -4108 1522
rect -13321 581 -6175 692
rect -3532 1458 -3098 1493
rect 3539 1331 3817 1609
rect 4005 1517 4087 1625
rect 7355 1586 7442 1661
rect 15548 1631 15711 1804
rect 4211 1401 4314 1496
rect -18015 346 -17624 544
rect -6513 312 -5616 444
rect 3581 901 3707 1027
rect 4620 1409 4785 1494
rect 7096 1380 7253 1526
rect 19826 2796 20301 2844
rect 22360 2725 22516 2881
rect 26714 2685 26932 2849
rect 25084 2124 25279 2326
rect 25955 2116 26111 2333
rect 50542 2243 50721 2422
rect 58755 2386 58904 2553
rect 4409 1086 4532 1218
rect 5743 698 6186 762
rect 19503 969 19720 1182
rect -13067 -393 -7302 -194
rect -6033 -357 -5757 -285
rect -25491 -973 -25219 -685
rect -5950 -986 -5822 -806
rect -5038 -916 -4568 -869
rect -4169 -1070 -4077 -1007
rect 4009 92 4158 241
rect -1561 -303 -1357 -109
rect 4399 -189 4556 -40
rect 5908 -107 6180 182
rect 15862 -126 16220 272
rect 46667 1720 46883 1940
rect 47931 1693 48166 1963
rect 22484 924 22810 1250
rect 19992 -557 20496 -512
rect 3332 -890 3556 -685
rect 47770 -719 47930 -586
rect 60637 -650 61047 -363
rect 4545 -1058 4984 -1020
rect 7348 -1190 7431 -1105
rect 16127 -1183 16382 -922
rect 19863 -1236 20055 -1038
rect 4329 -2295 4444 -2185
rect -1565 -2555 -1322 -2389
rect 46922 -2436 47268 -2104
rect 3272 -2865 3578 -2577
rect 15509 -3174 15772 -2937
rect 16127 -3560 16439 -3330
rect 49001 -3654 49228 -3400
rect 61891 -3498 62043 -3419
rect 62407 -3424 62884 -3380
rect 65203 -3454 65314 -3352
rect 87922 -3477 88155 -3270
rect 62459 -4119 62739 -3819
rect 17387 -4748 17851 -4336
rect 18041 -5366 18388 -4983
rect 46893 -5188 47282 -4756
rect 61311 -4968 61459 -4819
rect 18534 -6062 18990 -5587
rect 19096 -6756 19485 -6399
rect 19761 -7533 20205 -7105
rect 90356 -7278 92687 -5041
rect -31403 -9854 -30698 -8957
rect 59141 -9746 59762 -8995
rect 60606 -10565 61337 -9800
rect -29386 -11622 -28448 -10684
rect -26778 -11775 -26091 -11088
rect -24163 -11688 -23436 -11046
rect -6545 -11841 -6016 -11233
rect 61603 -11734 62208 -11260
rect 62379 -13054 62984 -12580
rect -25660 -14763 -25005 -14334
rect -12812 -15176 -7984 -15031
rect 90543 -18603 91459 -17718
rect -25539 -23304 -25139 -22879
rect 90878 -35139 91794 -34254
rect -27597 -41124 -27494 -37041
rect -25900 -43047 -25681 -42828
rect -29447 -46364 -28280 -45411
rect 91488 -53354 92404 -52469
rect -29398 -58999 -29235 -54826
rect -27236 -60993 -26896 -60567
rect -31540 -64772 -30673 -63836
<< metal1 >>
rect -4820 44054 -3786 44102
rect -1993 44054 -862 44070
rect -4820 43973 -797 44054
rect -4820 43957 -1815 43973
rect -4820 42551 -4707 43957
rect -3915 42567 -1815 43957
rect -1023 42567 -797 43973
rect -3915 42551 -797 42567
rect -4820 42503 -797 42551
rect -4820 42470 -3786 42503
rect -1993 42470 -862 42503
rect -3742 40415 -2527 40571
rect -3742 39539 -3598 40415
rect -2667 40236 -2527 40415
rect -2667 39539 -2367 40236
rect -3742 39356 -2367 39539
rect -17836 9129 -15919 9265
rect -17836 565 -17700 9129
rect -16277 8494 -5438 8555
rect -16277 8440 -5433 8494
rect -16277 8117 -16077 8440
rect -15564 8398 -5433 8440
rect -15564 8117 -6475 8398
rect -16277 8032 -6475 8117
rect -6540 7393 -6475 8032
rect -5556 7393 -5433 8398
rect -6540 7273 -5433 7393
rect -12975 6743 -11404 6943
rect -12975 5686 -12802 6743
rect -11669 5686 -11404 6743
rect -12975 3566 -11404 5686
rect -3582 6690 -2367 39356
rect 13898 8915 14773 8919
rect 13898 8869 14775 8915
rect 13898 8763 14599 8869
rect 14739 8763 14775 8869
rect 6966 8732 7312 8756
rect 6966 8509 7009 8732
rect 7275 8509 7312 8732
rect 6966 8466 7312 8509
rect 13898 8737 14775 8763
rect 3375 8071 4103 8200
rect 3375 7636 3492 8071
rect 3927 7636 4103 8071
rect 3375 7565 4103 7636
rect -3582 5746 -3482 6690
rect -2539 5746 -2367 6690
rect -3582 5554 -2367 5746
rect 2866 4480 3250 4560
rect 2866 4186 2911 4480
rect 3195 4186 3250 4480
rect 2866 4116 3250 4186
rect -13122 3529 -8953 3566
rect -13122 3359 -13070 3529
rect -9285 3359 -8953 3529
rect -13122 3329 -8953 3359
rect -13011 2361 -12663 3329
rect -11909 2361 -11561 3329
rect -11015 2361 -10667 3329
rect -10239 2361 -9891 3329
rect -9633 2361 -9285 3329
rect -5845 2730 -5539 2764
rect -5845 2515 -5811 2730
rect -5591 2515 -5539 2730
rect -5845 2483 -5539 2515
rect -613 2710 538 2816
rect -13395 2305 -9226 2361
rect -13395 2173 -13326 2305
rect -9322 2173 -9226 2305
rect -13395 2124 -9226 2173
rect -5742 1521 -5581 2483
rect -613 1575 -456 2710
rect 3061 2090 3235 4116
rect 3500 3577 3875 7565
rect 3500 3328 3558 3577
rect 3807 3328 3875 3577
rect -4212 1522 -4099 1535
rect -5774 1514 -5574 1521
rect -5774 1365 -5761 1514
rect -5593 1415 -5574 1514
rect -4212 1479 -4196 1522
rect -4108 1498 -4099 1522
rect -3572 1498 -3060 1502
rect -4108 1493 -3060 1498
rect -4108 1479 -3532 1493
rect -4212 1461 -3532 1479
rect -3572 1458 -3532 1461
rect -3098 1458 -3060 1493
rect -3572 1449 -3060 1458
rect -1188 1423 -456 1575
rect 3500 1609 3875 3328
rect 7080 2079 7229 8466
rect 7289 8267 7635 8307
rect 7289 8056 7332 8267
rect 7560 8056 7635 8267
rect 7289 8017 7635 8056
rect 7054 2052 7303 2079
rect 7054 1856 7079 2052
rect 7277 1856 7303 2052
rect 7054 1845 7303 1856
rect 7341 1680 7460 8017
rect 13898 5964 14080 8737
rect 14547 8736 14775 8737
rect 14484 7856 14591 7858
rect 14484 7815 14796 7856
rect 14484 7666 14591 7815
rect 14740 7749 14796 7815
rect 14740 7666 14795 7749
rect 14484 7642 14795 7666
rect 14484 6213 14653 7642
rect 15079 6970 15125 8735
rect 16226 8722 16396 8743
rect 16226 8621 16254 8722
rect 16384 8621 16396 8722
rect 16226 8605 16396 8621
rect 26753 8650 38073 8844
rect 14997 6913 15211 6970
rect 14997 6801 15031 6913
rect 15166 6801 15211 6913
rect 14997 6756 15211 6801
rect 16250 6623 16388 8605
rect 16519 7884 17132 8006
rect 16519 7621 16664 7884
rect 16961 7621 17132 7884
rect 26753 7762 27003 8650
rect 37629 7762 38073 8650
rect 26753 7623 38073 7762
rect 16227 6583 16406 6623
rect 16227 6481 16261 6583
rect 16370 6481 16406 6583
rect 16227 6444 16406 6481
rect 14443 6192 14691 6213
rect 14443 6047 14484 6192
rect 14639 6047 14691 6192
rect 14443 6016 14691 6047
rect 13866 5937 14130 5964
rect 13866 5734 13908 5937
rect 14090 5734 14130 5937
rect 13866 5703 14130 5734
rect 15814 4127 16331 4171
rect 15814 3748 15869 4127
rect 16252 3748 16331 4127
rect 15814 3722 16331 3748
rect 15522 1804 15742 1833
rect 7337 1670 7470 1680
rect 6982 1661 7470 1670
rect -5593 1371 -3699 1415
rect -5593 1365 -5574 1371
rect -5774 1352 -5574 1365
rect 3500 1331 3539 1609
rect 3817 1331 3875 1609
rect 3990 1625 4106 1638
rect 3990 1517 4005 1625
rect 4087 1591 4106 1625
rect 6982 1624 7355 1661
rect 4087 1547 4392 1591
rect 7337 1586 7355 1624
rect 7442 1586 7470 1661
rect 15522 1631 15548 1804
rect 15711 1631 15742 1804
rect 15522 1597 15742 1631
rect 7337 1562 7470 1586
rect 4087 1517 4106 1547
rect 7061 1526 7270 1554
rect 3990 1499 4106 1517
rect 4186 1496 4963 1519
rect 4186 1401 4211 1496
rect 4314 1494 4963 1496
rect 4314 1409 4620 1494
rect 4785 1409 4963 1494
rect 4314 1401 4963 1409
rect 4186 1385 4963 1401
rect 4580 1384 4827 1385
rect 7061 1380 7096 1526
rect 7253 1380 7270 1526
rect 7061 1355 7270 1380
rect 3500 1279 3875 1331
rect 4064 1310 4362 1354
rect -5243 1073 -3681 1219
rect 3161 1101 3899 1159
rect -13350 692 -6080 721
rect -13350 581 -13321 692
rect -6175 581 -6080 692
rect -18039 544 -17604 565
rect -13350 548 -6080 581
rect -18039 346 -18015 544
rect -17624 346 -17604 544
rect -18039 321 -17604 346
rect -12759 -135 -12272 548
rect -11199 -135 -10712 548
rect -10006 -135 -9519 548
rect -8823 -135 -8336 548
rect -7809 -135 -7322 548
rect -5243 473 -5078 1073
rect 3563 1027 3725 1039
rect 3563 901 3581 1027
rect 3707 973 3725 1027
rect 3707 929 3812 973
rect 3707 901 3725 929
rect 3563 885 3725 901
rect -6599 444 -5077 473
rect -6599 389 -6513 444
rect -6600 312 -6513 389
rect -5616 312 -5077 444
rect -6600 308 -5077 312
rect -6600 257 -5078 308
rect -6601 224 -5078 257
rect -13197 -194 -7163 -135
rect -13197 -393 -13067 -194
rect -7302 -393 -7163 -194
rect -13197 -453 -7163 -393
rect -25553 -685 -25165 -654
rect -25553 -973 -25491 -685
rect -25219 -973 -25165 -685
rect -25553 -1050 -25165 -973
rect -31679 -8957 -30522 -8679
rect -31679 -9854 -31403 -8957
rect -30698 -9854 -30522 -8957
rect -31679 -62597 -30522 -9854
rect -29580 -10684 -28157 -10506
rect -29580 -11622 -29386 -10684
rect -28448 -11622 -28157 -10684
rect -26907 -11088 -25983 -10980
rect -26907 -11153 -26778 -11088
rect -29580 -45411 -28157 -11622
rect -27809 -11705 -26778 -11153
rect -27809 -37041 -27257 -11705
rect -26907 -11775 -26778 -11705
rect -26091 -11775 -25983 -11088
rect -26907 -11904 -25983 -11775
rect -25501 -14108 -25219 -1050
rect -12865 -10939 -11924 -453
rect -24248 -11046 -11923 -10939
rect -24248 -11688 -24163 -11046
rect -23436 -11688 -11923 -11046
rect -24248 -11880 -11923 -11688
rect -25931 -14334 -24870 -14108
rect -25931 -14763 -25660 -14334
rect -25005 -14763 -24870 -14334
rect -25931 -14876 -24870 -14763
rect -25501 -22779 -25219 -14876
rect -12865 -14969 -11924 -11880
rect -10614 -14969 -9673 -453
rect -8935 -14969 -7994 -453
rect -6601 -11153 -6294 224
rect -2521 0 182 106
rect -6059 -285 -5507 -276
rect -6059 -357 -6033 -285
rect -5757 -357 -5507 -285
rect -6059 -378 -5507 -357
rect -5976 -806 -5800 -784
rect -5976 -986 -5950 -806
rect -5822 -957 -5800 -806
rect -5544 -873 -5507 -378
rect -2521 -665 -2415 0
rect -1581 -109 -1323 -85
rect -1581 -303 -1561 -109
rect -1357 -303 -1323 -109
rect -1581 -342 -1323 -303
rect -2521 -779 -2422 -665
rect -5056 -869 -4533 -861
rect -5056 -873 -5038 -869
rect -5544 -910 -5038 -873
rect -5056 -916 -5038 -910
rect -4568 -916 -4533 -869
rect -2650 -887 -2422 -779
rect -5056 -922 -4533 -916
rect -2598 -924 -2422 -887
rect -5822 -986 -5194 -957
rect -5976 -1001 -5194 -986
rect -5976 -1005 -5800 -1001
rect -4185 -1007 -4062 -989
rect -4185 -1070 -4169 -1007
rect -4077 -1070 -4062 -1007
rect -4185 -1079 -4062 -1070
rect -4182 -1094 -4138 -1079
rect -1517 -2369 -1361 -342
rect 3281 -685 3574 -645
rect 3281 -890 3332 -685
rect 3556 -890 3574 -685
rect 3281 -911 3574 -890
rect -1585 -2389 -1283 -2369
rect -1585 -2555 -1565 -2389
rect -1322 -2555 -1283 -2389
rect 3313 -2539 3558 -911
rect 3768 -1099 3812 929
rect 3841 -1011 3899 1101
rect 4064 265 4108 1310
rect 4388 1218 4549 1243
rect 4388 1086 4409 1218
rect 4532 1086 4549 1218
rect 4388 1066 4549 1086
rect 3985 241 4186 265
rect 3985 92 4009 241
rect 4158 92 4186 241
rect 3985 76 4186 92
rect 4408 -15 4507 1066
rect 5730 762 6208 775
rect 5730 698 5743 762
rect 6186 698 6208 762
rect 5730 686 6208 698
rect 5943 223 6135 686
rect 5891 182 6236 223
rect 4383 -40 4585 -15
rect 4383 -189 4399 -40
rect 4556 -189 4585 -40
rect 5891 -107 5908 182
rect 6180 -107 6236 182
rect 5891 -122 6236 -107
rect 4383 -213 4585 -189
rect 3841 -1020 4999 -1011
rect 7131 -1020 7230 1355
rect 3841 -1058 4545 -1020
rect 4984 -1058 4999 -1020
rect 3841 -1066 4999 -1058
rect 6997 -1066 7412 -1020
rect 3841 -1069 4601 -1066
rect 7334 -1093 7412 -1066
rect 3768 -1143 4387 -1099
rect 7334 -1105 7443 -1093
rect 7334 -1190 7348 -1105
rect 7431 -1190 7443 -1105
rect 7334 -1207 7443 -1190
rect 4353 -2171 4397 -1336
rect 4310 -2185 4465 -2171
rect 4310 -2295 4329 -2185
rect 4444 -2295 4465 -2185
rect 4310 -2309 4465 -2295
rect -1585 -2584 -1283 -2555
rect 3196 -2577 3624 -2539
rect 3196 -2865 3272 -2577
rect 3578 -2865 3624 -2577
rect 15547 -2842 15703 1597
rect 15814 272 16329 3722
rect 16519 909 17132 7621
rect 19201 6996 19643 7085
rect 19201 6709 19300 6996
rect 19588 6709 19643 6996
rect 19201 6620 19643 6709
rect 22939 6995 23303 7116
rect 22939 6735 23009 6995
rect 23217 6735 23303 6995
rect 22939 6666 23303 6735
rect 18791 5539 19168 5573
rect 18791 5255 18835 5539
rect 19139 5255 19168 5539
rect 18791 5216 19168 5255
rect 18137 3181 18324 3184
rect 18137 3163 18330 3181
rect 18137 3007 18170 3163
rect 18307 3007 18330 3163
rect 18137 2985 18330 3007
rect 16519 296 17906 909
rect 15814 -126 15862 272
rect 16220 -126 16329 272
rect 15814 -255 16329 -126
rect 16101 -922 16445 -871
rect 16101 -1183 16127 -922
rect 16382 -1183 16445 -922
rect 16101 -1228 16445 -1183
rect 3196 -2900 3624 -2865
rect 15440 -2937 15853 -2842
rect 15440 -3174 15509 -2937
rect 15772 -3174 15853 -2937
rect 15440 -3211 15853 -3174
rect 16133 -3292 16375 -1228
rect 16088 -3330 16483 -3292
rect 16088 -3560 16127 -3330
rect 16439 -3560 16483 -3330
rect 16088 -3623 16483 -3560
rect 17293 -4336 17906 296
rect 17293 -4748 17387 -4336
rect 17851 -4748 17906 -4336
rect 17293 -4848 17906 -4748
rect 18137 -4849 18324 2985
rect 18621 2540 18758 2557
rect 18621 2449 18635 2540
rect 18734 2449 18758 2540
rect 17978 -4983 18468 -4849
rect 17978 -5366 18041 -4983
rect 18388 -5366 18468 -4983
rect 17978 -5437 18468 -5366
rect 18621 -5532 18758 2449
rect 18861 -594 19153 5216
rect 19341 2756 19470 6620
rect 19552 2877 19650 2892
rect 19552 2800 19563 2877
rect 19636 2862 19650 2877
rect 22316 2881 22554 2900
rect 22316 2875 22360 2881
rect 19636 2858 19659 2862
rect 19636 2844 20314 2858
rect 19636 2800 19826 2844
rect 19552 2796 19826 2800
rect 20301 2796 20314 2844
rect 19552 2787 20314 2796
rect 19341 2712 19648 2756
rect 22188 2745 22360 2875
rect 22316 2725 22360 2745
rect 22516 2725 22554 2881
rect 19341 2700 19470 2712
rect 22316 2711 22554 2725
rect 19341 2565 19481 2579
rect 19341 2458 19368 2565
rect 19468 2519 19481 2565
rect 19468 2475 19671 2519
rect 19468 2458 19481 2475
rect 19341 2444 19481 2458
rect 22436 1250 22925 1317
rect 22436 1241 22484 1250
rect 19472 1182 22484 1241
rect 19472 969 19503 1182
rect 19720 969 22484 1182
rect 19472 943 22484 969
rect 19472 -496 19542 943
rect 22436 924 22484 943
rect 22810 924 22925 1250
rect 22436 895 22925 924
rect 22358 -353 22513 -345
rect 23046 -353 23217 6666
rect 26836 3886 28029 7623
rect 29111 3886 30304 7623
rect 31275 3886 32468 7623
rect 33884 3886 35077 7623
rect 36381 3886 37574 7623
rect 41672 4733 44640 4844
rect 41672 4322 41705 4733
rect 44546 4322 44640 4733
rect 41672 4185 44640 4322
rect 26583 3817 38866 3886
rect 26583 3540 26668 3817
rect 38672 3540 38866 3817
rect 26583 3483 38866 3540
rect 41865 3233 42195 4185
rect 42554 3233 42884 4185
rect 43243 3233 43573 4185
rect 43752 3233 44082 4185
rect 41827 3211 44196 3233
rect 41827 3154 41845 3211
rect 44154 3154 44196 3211
rect 41827 3129 44196 3154
rect 26688 2849 26963 2876
rect 26688 2685 26714 2849
rect 26932 2685 26963 2849
rect 26688 2653 26963 2685
rect 25061 2326 25333 2372
rect 25061 2124 25084 2326
rect 25279 2295 25333 2326
rect 25947 2333 26150 2357
rect 25947 2295 25955 2333
rect 25279 2124 25955 2295
rect 25061 2085 25333 2124
rect 25947 2116 25955 2124
rect 26111 2116 26150 2333
rect 25947 2092 26150 2116
rect 26762 646 26890 2653
rect 58706 2553 59616 2704
rect 50510 2422 50749 2467
rect 50510 2243 50542 2422
rect 50721 2243 50749 2422
rect 58706 2386 58755 2553
rect 58904 2386 59616 2553
rect 58706 2260 59616 2386
rect 50510 2215 50749 2243
rect 46637 1940 46961 1997
rect 46637 1720 46667 1940
rect 46883 1917 46961 1940
rect 47896 1963 48216 1992
rect 47896 1917 47931 1963
rect 46883 1738 47931 1917
rect 46883 1720 46961 1738
rect 46637 1686 46961 1720
rect 47896 1693 47931 1738
rect 48166 1884 48216 1963
rect 50542 1917 50721 2215
rect 48166 1705 49256 1884
rect 48166 1693 48216 1705
rect 47896 1636 48216 1693
rect 26762 518 27180 646
rect 27052 -166 27180 518
rect 19472 -512 20517 -496
rect 19472 -557 19992 -512
rect 20496 -557 20517 -512
rect 22342 -524 23217 -353
rect 22358 -525 22513 -524
rect 19472 -566 20517 -557
rect 22433 -561 22513 -525
rect 18861 -638 19820 -594
rect 46227 -632 46301 1314
rect 47758 -586 47953 -572
rect 47758 -632 47770 -586
rect 46227 -706 47770 -632
rect 47758 -719 47770 -706
rect 47930 -719 47953 -586
rect 47758 -752 47953 -719
rect 19212 -831 19359 -829
rect 19212 -875 20074 -831
rect 18424 -5587 19081 -5532
rect 18424 -6062 18534 -5587
rect 18990 -6062 19081 -5587
rect 18424 -6171 19081 -6062
rect 19212 -6293 19542 -875
rect 19836 -1038 20093 -990
rect 19836 -1236 19863 -1038
rect 20055 -1236 20093 -1038
rect 19836 -1279 20093 -1236
rect 18949 -6399 19611 -6293
rect 18949 -6756 19096 -6399
rect 19485 -6756 19611 -6399
rect 18949 -6850 19611 -6756
rect 19868 -7025 20066 -1279
rect 46850 -2104 47412 -1960
rect 46850 -2436 46922 -2104
rect 47268 -2436 47412 -2104
rect 46850 -4670 47412 -2436
rect 49077 -3371 49256 1705
rect 48966 -3400 49277 -3371
rect 48966 -3654 49001 -3400
rect 49228 -3654 49277 -3400
rect 48966 -3697 49277 -3654
rect 46778 -4756 47412 -4670
rect 46778 -5188 46893 -4756
rect 47282 -5188 47412 -4756
rect 46778 -5304 47412 -5188
rect 19665 -7105 20295 -7025
rect 19665 -7533 19761 -7105
rect 20205 -7533 20295 -7105
rect 19665 -7634 20295 -7533
rect 59172 -8831 59616 2260
rect 60549 -363 61159 -228
rect 60549 -650 60637 -363
rect 61047 -650 61159 -363
rect 58913 -8995 59860 -8831
rect 58913 -9746 59141 -8995
rect 59762 -9746 59860 -8995
rect 60549 -9617 61159 -650
rect 61353 -3293 62176 -3228
rect 61353 -4779 61418 -3293
rect 62111 -3360 62176 -3293
rect 87785 -3270 88210 -3189
rect 65187 -3352 65330 -3337
rect 62111 -3380 62910 -3360
rect 61873 -3419 62067 -3407
rect 61873 -3498 61891 -3419
rect 62043 -3460 62067 -3419
rect 62111 -3424 62407 -3380
rect 62884 -3424 62910 -3380
rect 65187 -3381 65203 -3352
rect 62111 -3425 62910 -3424
rect 62387 -3431 62910 -3425
rect 64860 -3427 65203 -3381
rect 65187 -3454 65203 -3427
rect 65314 -3454 65330 -3352
rect 62043 -3498 62250 -3460
rect 65187 -3468 65330 -3454
rect 61873 -3504 62250 -3498
rect 87785 -3477 87922 -3270
rect 88155 -3477 88210 -3270
rect 61873 -3516 62067 -3504
rect 87785 -3581 88210 -3477
rect 61655 -3741 62267 -3697
rect 61261 -4819 61482 -4779
rect 61261 -4968 61311 -4819
rect 61459 -4968 61482 -4819
rect 61261 -5041 61482 -4968
rect 58913 -9909 59860 -9746
rect 60423 -9800 61454 -9617
rect 60423 -10565 60606 -9800
rect 61337 -10565 61454 -9800
rect 60423 -10731 61454 -10565
rect 61655 -11116 62108 -3741
rect 62432 -3819 62779 -3786
rect 62432 -4119 62459 -3819
rect 62739 -4119 62779 -3819
rect 62432 -4139 62779 -4119
rect -6611 -11233 -5937 -11153
rect -6611 -11841 -6545 -11233
rect -6016 -11841 -5937 -11233
rect -6611 -11894 -5937 -11841
rect 61366 -11260 62272 -11116
rect 61366 -11734 61603 -11260
rect 62208 -11734 62272 -11260
rect 61366 -11971 62272 -11734
rect 62465 -12441 62732 -4139
rect 62246 -12580 63072 -12441
rect 62246 -13054 62379 -12580
rect 62984 -13054 63072 -12580
rect 62246 -13180 63072 -13054
rect -12874 -15031 -7870 -14969
rect -12874 -15176 -12812 -15031
rect -7984 -15176 -7870 -15031
rect -12874 -15238 -7870 -15176
rect -12865 -15240 -11924 -15238
rect -25664 -22879 -25039 -22779
rect -25664 -23304 -25539 -22879
rect -25139 -23304 -25039 -22879
rect -25664 -23404 -25039 -23304
rect 87916 -26943 88161 -3581
rect 89990 -5041 92959 -4698
rect 89990 -7278 90356 -5041
rect 92687 -7278 92959 -5041
rect 89990 -7667 92959 -7278
rect 84040 -27188 88161 -26943
rect 90119 -17718 92731 -7667
rect 90119 -18603 90543 -17718
rect 91459 -18603 92731 -17718
rect 84612 -27482 84857 -27188
rect 80867 -27727 84857 -27482
rect -27809 -41124 -27597 -37041
rect -27494 -41124 -27257 -37041
rect -27809 -42856 -27257 -41124
rect 90119 -34254 92731 -18603
rect 90119 -35139 90878 -34254
rect 91794 -35139 92731 -34254
rect -25977 -42828 -25639 -42789
rect -25977 -42856 -25900 -42828
rect -27809 -43047 -25900 -42856
rect -25681 -43047 -25639 -42828
rect -22415 -42924 -22111 -42864
rect -27809 -43351 -27257 -43047
rect -25977 -43127 -25639 -43047
rect -29580 -46364 -29447 -45411
rect -28280 -46364 -28157 -45411
rect -29580 -46472 -28157 -46364
rect 90119 -52469 92731 -35139
rect -29536 -54826 -29081 -52616
rect 90119 -53354 91488 -52469
rect 92404 -53354 92731 -52469
rect 90119 -54278 92731 -53354
rect -29536 -58999 -29398 -54826
rect -29235 -58999 -29081 -54826
rect -29536 -60594 -29081 -58999
rect -27322 -60567 -26810 -60453
rect -27322 -60594 -27236 -60567
rect -29536 -60993 -27236 -60594
rect -26896 -60993 -26810 -60567
rect -29536 -61049 -26810 -60993
rect -21712 -61035 -21354 -60975
rect -27322 -61078 -26810 -61049
rect -31679 -63836 -30520 -62597
rect -31679 -64772 -31540 -63836
rect -30673 -64772 -30522 -63836
rect -31679 -64865 -30522 -64772
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_0
timestamp 1717691374
transform 1 0 5174 0 1 -1085
box -887 -901 1869 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_1
timestamp 1717691374
transform 1 0 -2940 0 1 1429
box -887 -901 1869 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_2
timestamp 1717691374
transform 1 0 -4408 0 1 -943
box -887 -901 1869 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_3
timestamp 1717691374
transform 1 0 20610 0 1 -580
box -887 -901 1869 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_4
timestamp 1717691374
transform 1 0 5159 0 1 1605
box -887 -901 1869 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_5
timestamp 1717691374
transform 1 0 20438 0 1 2770
box -887 -901 1869 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_6
timestamp 1717691374
transform 1 0 63037 0 1 -3446
box -887 -901 1869 842
use CP  CP_0
timestamp 1717691374
transform 0 -1 14952 1 0 9056
box -3766 -80648 80252 15106
use divider_top  divider_top_0
timestamp 1717691374
transform 1 0 9841 0 1 -30857
box -34598 -95 78026 15696
use divider_top  divider_top_1
timestamp 1717691374
transform 1 0 10539 0 1 -47448
box -34598 -95 78026 15696
use divider_top  divider_top_2
timestamp 1717691374
transform 0 1 -17326 1 0 43154
box -34598 -95 78026 15696
use divider_top  divider_top_3
timestamp 1717691374
transform 1 0 11242 0 1 -65559
box -34598 -95 78026 15696
use mirror_mag  mirror_mag_0
timestamp 1717691374
transform -1 0 14294 0 1 4889
box 1529 -557 6212 3030
use PFD  PFD_0
timestamp 1717691374
transform 1 0 540 0 1 474
box -539 -474 2730 2342
use Tapered_Buffer_mag  Tapered_Buffer_mag_0
timestamp 1717691374
transform -1 0 -5857 0 1 1513
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_1
timestamp 1717691374
transform 1 0 7529 0 1 -961
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_2
timestamp 1717691374
transform -1 0 -7497 0 -1 -16074
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_3
timestamp 1717691374
transform 1 0 50645 0 1 -3386
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_4
timestamp 1717691374
transform 1 0 50848 0 1 2572
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_5
timestamp 1717691374
transform 1 0 50645 0 1 -339
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_6
timestamp 1717691374
transform 1 0 7570 0 1 1795
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_7
timestamp 1717691374
transform 0 1 -27894 1 0 -59716
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_8
timestamp 1717691374
transform 0 1 -26074 1 0 -41571
box -156 -982 7721 769
use VCO  VCO_0
timestamp 1717691374
transform 1 0 33690 0 1 -975
box -8117 -475 13984 4754
<< labels >>
flabel locali -32843 -63367 -32843 -63367 0 FreeSans 1600 0 0 0 D19
port 44 nsew
flabel locali -32912 -63121 -32912 -63121 0 FreeSans 1600 0 0 0 D18
port 43 nsew
flabel locali -33364 -62901 -33364 -62901 0 FreeSans 1600 0 0 0 D17
port 42 nsew
flabel locali -32966 -62696 -32966 -62696 0 FreeSans 1600 0 0 0 D16
port 41 nsew
flabel locali -18882 7776 -18882 7776 0 FreeSans 1600 0 0 0 D10
port 40 nsew
flabel locali -19736 7109 -19736 7109 0 FreeSans 1600 0 0 0 D9
port 39 nsew
flabel locali -19883 5428 -19883 5428 0 FreeSans 1600 0 0 0 D8
port 38 nsew
flabel locali -20443 4401 -20443 4401 0 FreeSans 1600 0 0 0 D7
port 37 nsew
flabel locali -32808 -29624 -32808 -29624 0 FreeSans 1600 0 0 0 D6
port 36 nsew
flabel locali -32684 -29264 -32684 -29264 0 FreeSans 1600 0 0 0 D5
port 35 nsew
flabel locali -32907 -28960 -32907 -28960 0 FreeSans 1600 0 0 0 D4
port 34 nsew
flabel locali -32504 -28656 -32504 -28656 0 FreeSans 1600 0 0 0 D3
port 33 nsew
flabel locali -32417 -28414 -32417 -28414 0 FreeSans 1600 0 0 0 D2
port 32 nsew
flabel locali -32448 -28196 -32448 -28196 0 FreeSans 1600 0 0 0 D1
port 31 nsew
flabel locali -32479 -27992 -32479 -27992 0 FreeSans 1600 0 0 0 D0
port 30 nsew
flabel locali -22154 405 -22154 405 0 FreeSans 1600 0 0 0 F_IN
port 29 nsew
flabel locali -26050 -4594 -26050 -4594 0 FreeSans 1600 0 0 0 ITAIL
port 11 nsew
flabel locali -32390 -45265 -32390 -45265 0 FreeSans 1600 0 0 0 D15
port 28 nsew
flabel locali -32390 -45015 -32390 -45015 0 FreeSans 1600 0 0 0 D14
port 27 nsew
flabel locali -32366 -44780 -32366 -44780 0 FreeSans 1600 0 0 0 D13
port 26 nsew
flabel locali -32358 -44578 -32358 -44578 0 FreeSans 1600 0 0 0 D12
port 25 nsew
flabel locali -32436 -50788 -32436 -50788 0 FreeSans 1600 0 0 0 OUT_USB
port 24 nsew
flabel locali -32043 -33050 -32043 -33050 0 FreeSans 1600 0 0 0 OUT_CORE
port 23 nsew
flabel locali -26457 -7358 -26457 -7358 0 FreeSans 1600 0 0 0 S5
port 15 nsew
flabel locali -26433 -6567 -26433 -6567 0 FreeSans 1600 0 0 0 LF_OFFCHIP
port 14 nsew
flabel locali -26146 -6015 -26146 -6015 0 FreeSans 1600 0 0 0 VCTRL_IN
port 13 nsew
flabel locali -26022 -5307 -26022 -5307 0 FreeSans 1600 0 0 0 S4
port 12 nsew
flabel locali -26013 -3482 -26013 -3482 0 FreeSans 1600 0 0 0 DN_OUT
port 9 nsew
flabel locali -25937 -3111 -25937 -3111 0 FreeSans 1600 0 0 0 UP_OUT
port 8 nsew
flabel locali -26089 -2778 -26089 -2778 0 FreeSans 1600 0 0 0 S3
port 7 nsew
flabel locali -26048 -2492 -26048 -2492 0 FreeSans 1600 0 0 0 S2
port 6 nsew
flabel locali -26267 -2271 -26267 -2271 0 FreeSans 1600 0 0 0 DN_INPUT
port 5 nsew
flabel locali -26239 -2019 -26239 -2019 0 FreeSans 1600 0 0 0 UP_INPUT
port 4 nsew
flabel locali -21980 -628 -21980 -628 0 FreeSans 1600 0 0 0 S6
port 3 nsew
flabel locali -33957 -9382 -33957 -9382 0 FreeSans 1600 0 0 0 OUTB
port 47 nsew
flabel locali -34119 -12958 -34119 -12958 0 FreeSans 1600 0 0 0 OUT
port 48 nsew
flabel locali -22650 1410 -22650 1410 0 FreeSans 1600 0 0 0 PRE_SCALAR
port 49 nsew
flabel locali -22938 181 -22938 181 0 FreeSans 1600 0 0 0 S1
port 50 nsew
flabel locali -34376 -14319 -34376 -14319 0 FreeSans 1600 0 0 0 S7
port 51 nsew
flabel locali -34232 -15974 -34232 -15974 0 FreeSans 1600 0 0 0 DIV_OUT
port 52 nsew
flabel locali 97170 -15073 97170 -15073 0 FreeSans 16000 0 0 0 VDD
port 53 nsew
flabel locali 79409 -6079 79409 -6079 0 FreeSans 16000 0 0 0 VSS
port 55 nsew
<< end >>
