magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< locali >>
rect 2073 2833 2367 2894
rect 3565 1673 3968 1790
rect 5244 1738 6364 1860
rect 3002 1663 3100 1666
rect 3565 1663 3682 1673
rect 3002 1656 3682 1663
rect 2774 1618 2836 1646
rect 2650 1616 2836 1618
rect 2650 1582 2788 1616
rect 2822 1582 2836 1616
rect 2650 1566 2836 1582
rect 2774 1552 2836 1566
rect 3002 1622 3034 1656
rect 3068 1622 3682 1656
rect 3002 1584 3682 1622
rect 3002 1550 3034 1584
rect 3068 1550 3682 1584
rect 3002 1546 3682 1550
rect 3002 1540 3100 1546
rect -191 967 37 1003
rect 249 -259 325 900
rect 3406 889 3808 923
rect 3406 570 3449 889
rect 5165 836 5219 849
rect 5165 832 5175 836
rect 5079 802 5175 832
rect 5209 802 5219 836
rect 5079 798 5219 802
rect 5165 790 5219 798
rect 3642 754 3846 788
rect 3642 627 3714 754
rect 5280 642 5572 680
rect 3642 618 3726 627
rect 3647 604 3726 618
rect 3647 570 3669 604
rect 3703 570 3726 604
rect 3647 548 3726 570
rect 3396 127 4007 195
rect 1740 82 4007 127
rect 1740 14 3509 82
rect 5534 -253 5572 642
rect 249 -335 3559 -259
rect 249 -517 325 -335
rect 3009 -452 3411 -386
rect 249 -593 391 -517
rect 315 -1091 391 -593
rect 580 -1870 1427 -1717
rect 1695 -1741 1854 -1735
rect 1695 -1847 1721 -1741
rect 1827 -1847 1854 -1741
rect 3009 -1753 3075 -452
rect 3133 -557 3225 -531
rect 3133 -591 3162 -557
rect 3196 -591 3225 -557
rect 3133 -616 3225 -591
rect 1695 -1853 1854 -1847
rect 2992 -1757 3076 -1753
rect 2992 -1791 3017 -1757
rect 3051 -1791 3076 -1757
rect 2992 -1829 3076 -1791
rect 2992 -1863 3017 -1829
rect 3051 -1863 3076 -1829
rect 2992 -1866 3076 -1863
rect -145 -2486 205 -2450
rect 38 -3513 174 -2486
rect 3156 -2591 3199 -616
rect 3345 -1782 3411 -452
rect 3483 -1039 3559 -335
rect 3785 -291 5572 -253
rect 3785 -669 3823 -291
rect 6242 -659 6364 1738
rect 3762 -679 3835 -669
rect 3762 -713 3781 -679
rect 3815 -713 3835 -679
rect 3762 -723 3835 -713
rect 6242 -781 6874 -659
rect 3483 -1115 4091 -1039
rect 4015 -1213 4091 -1115
rect 6752 -1777 6874 -781
rect 3345 -1848 4275 -1782
rect 6412 -1809 6491 -1792
rect 6412 -1823 6434 -1809
rect 6312 -1843 6434 -1823
rect 6468 -1843 6491 -1809
rect 6312 -1881 6491 -1843
rect 6312 -1906 6434 -1881
rect 6412 -1915 6434 -1906
rect 6468 -1915 6491 -1881
rect 6412 -1931 6491 -1915
rect 6662 -1808 6874 -1777
rect 6662 -1914 6678 -1808
rect 6784 -1914 6874 -1808
rect 6662 -1916 6874 -1914
rect 6662 -1944 6801 -1916
rect 3156 -2634 3441 -2591
rect 3398 -2883 3441 -2634
rect 3637 -3513 3773 -2481
rect 7060 -2914 7387 -2871
rect 38 -3649 3773 -3513
<< viali >>
rect 2788 1582 2822 1616
rect 3034 1622 3068 1656
rect 3034 1550 3068 1584
rect 5175 802 5209 836
rect 3669 570 3703 604
rect 1721 -1847 1827 -1741
rect 3162 -591 3196 -557
rect 3017 -1791 3051 -1757
rect 3017 -1863 3051 -1829
rect 3781 -713 3815 -679
rect 6434 -1843 6468 -1809
rect 6434 -1915 6468 -1881
rect 6678 -1914 6784 -1808
<< metal1 >>
rect -149 2761 156 2815
rect 2768 1642 2842 1658
rect 2996 1656 3106 1678
rect 2996 1642 3034 1656
rect 2768 1622 3034 1642
rect 3068 1622 3106 1656
rect 2768 1616 3106 1622
rect 2768 1582 2788 1616
rect 2822 1584 3106 1616
rect 2822 1582 3034 1584
rect 2768 1550 3034 1582
rect 3068 1550 3106 1584
rect 2768 1546 3106 1550
rect 2768 1540 2842 1546
rect 2996 1528 3106 1546
rect 5159 849 5225 861
rect 5159 836 6781 849
rect 5159 802 5175 836
rect 5209 802 6781 836
rect 5159 787 6781 802
rect 5159 778 5225 787
rect 3635 604 3738 633
rect 3635 570 3669 604
rect 3703 570 3738 604
rect 3635 542 3738 570
rect -305 -692 148 -638
rect 2804 -1129 2917 128
rect 3647 -91 3726 542
rect 3147 -170 3726 -91
rect 3147 -525 3226 -170
rect 3121 -557 3237 -525
rect 3121 -591 3162 -557
rect 3196 -591 3237 -557
rect 3121 -622 3237 -591
rect 3750 -679 3847 -663
rect 3750 -713 3781 -679
rect 3815 -713 3847 -679
rect 3750 -729 3847 -713
rect 1683 -1741 1866 -1729
rect 1683 -1847 1721 -1741
rect 1827 -1770 1866 -1741
rect 2986 -1757 3082 -1741
rect 2986 -1770 3017 -1757
rect 1827 -1791 3017 -1770
rect 3051 -1791 3082 -1757
rect 1827 -1829 3082 -1791
rect 1827 -1847 3017 -1829
rect 1683 -1852 3017 -1847
rect 1683 -1859 1866 -1852
rect 2986 -1863 3017 -1852
rect 3051 -1863 3082 -1829
rect 2986 -1878 3082 -1863
rect 6406 -1792 6497 -1780
rect 6656 -1792 6807 -1765
rect 6406 -1808 6807 -1792
rect 6406 -1809 6678 -1808
rect 6406 -1843 6434 -1809
rect 6468 -1843 6678 -1809
rect 6406 -1881 6678 -1843
rect 6406 -1915 6434 -1881
rect 6468 -1914 6678 -1881
rect 6784 -1914 6807 -1808
rect 6468 -1915 6807 -1914
rect 6406 -1931 6807 -1915
rect 6406 -1943 6497 -1931
rect 6656 -1956 6807 -1931
rect 2610 -3470 6564 -3357
use MUX_1  MUX_1_0
timestamp 1726359333
transform 1 0 88 0 1 399
box -88 -432 3425 2692
use MUX_1  MUX_1_1
timestamp 1726359333
transform 1 0 80 0 1 -3054
box -88 -432 3425 2692
use MUX_1  MUX_1_2
timestamp 1726359333
transform 1 0 3748 0 1 -3085
box -88 -432 3425 2692
use TSPC_MAGIC_1  TSPC_MAGIC_1_0
timestamp 1726359333
transform 1 0 3893 0 1 1023
box -119 -1019 1471 877
<< labels >>
flabel metal1 s -98 2790 -98 2790 0 FreeSans 3125 0 0 0 CLK
flabel locali s -162 982 -162 982 0 FreeSans 3125 0 0 0 G-CLK
flabel metal1 s -278 -672 -278 -672 0 FreeSans 3125 0 0 0 D1
flabel locali s -120 -2470 -120 -2470 0 FreeSans 3125 0 0 0 DATA
flabel locali s 258 -29 258 -29 0 FreeSans 3125 0 0 0 LD
flabel locali s 7327 -2896 7327 -2896 0 FreeSans 3125 0 0 0 Q
flabel locali s 2263 2857 2263 2857 0 FreeSans 3125 0 0 0 VSS
flabel locali s 963 -1807 963 -1807 0 FreeSans 3125 0 0 0 VDD
flabel metal1 s 6703 812 6703 812 0 FreeSans 3125 0 0 0 QB
<< end >>
