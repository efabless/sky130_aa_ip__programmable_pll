magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect -114 -362 114 362
<< pmos >>
rect -20 -300 20 300
<< pdiff >>
rect -78 255 -20 300
rect -78 221 -66 255
rect -32 221 -20 255
rect -78 187 -20 221
rect -78 153 -66 187
rect -32 153 -20 187
rect -78 119 -20 153
rect -78 85 -66 119
rect -32 85 -20 119
rect -78 51 -20 85
rect -78 17 -66 51
rect -32 17 -20 51
rect -78 -17 -20 17
rect -78 -51 -66 -17
rect -32 -51 -20 -17
rect -78 -85 -20 -51
rect -78 -119 -66 -85
rect -32 -119 -20 -85
rect -78 -153 -20 -119
rect -78 -187 -66 -153
rect -32 -187 -20 -153
rect -78 -221 -20 -187
rect -78 -255 -66 -221
rect -32 -255 -20 -221
rect -78 -300 -20 -255
rect 20 255 78 300
rect 20 221 32 255
rect 66 221 78 255
rect 20 187 78 221
rect 20 153 32 187
rect 66 153 78 187
rect 20 119 78 153
rect 20 85 32 119
rect 66 85 78 119
rect 20 51 78 85
rect 20 17 32 51
rect 66 17 78 51
rect 20 -17 78 17
rect 20 -51 32 -17
rect 66 -51 78 -17
rect 20 -85 78 -51
rect 20 -119 32 -85
rect 66 -119 78 -85
rect 20 -153 78 -119
rect 20 -187 32 -153
rect 66 -187 78 -153
rect 20 -221 78 -187
rect 20 -255 32 -221
rect 66 -255 78 -221
rect 20 -300 78 -255
<< pdiffc >>
rect -66 221 -32 255
rect -66 153 -32 187
rect -66 85 -32 119
rect -66 17 -32 51
rect -66 -51 -32 -17
rect -66 -119 -32 -85
rect -66 -187 -32 -153
rect -66 -255 -32 -221
rect 32 221 66 255
rect 32 153 66 187
rect 32 85 66 119
rect 32 17 66 51
rect 32 -51 66 -17
rect 32 -119 66 -85
rect 32 -187 66 -153
rect 32 -255 66 -221
<< poly >>
rect -20 300 20 326
rect -20 -326 20 -300
<< locali >>
rect -66 269 -32 304
rect -66 197 -32 221
rect -66 125 -32 153
rect -66 53 -32 85
rect -66 -17 -32 17
rect -66 -85 -32 -53
rect -66 -153 -32 -125
rect -66 -221 -32 -197
rect -66 -304 -32 -269
rect 32 269 66 304
rect 32 197 66 221
rect 32 125 66 153
rect 32 53 66 85
rect 32 -17 66 17
rect 32 -85 66 -53
rect 32 -153 66 -125
rect 32 -221 66 -197
rect 32 -304 66 -269
<< viali >>
rect -66 255 -32 269
rect -66 235 -32 255
rect -66 187 -32 197
rect -66 163 -32 187
rect -66 119 -32 125
rect -66 91 -32 119
rect -66 51 -32 53
rect -66 19 -32 51
rect -66 -51 -32 -19
rect -66 -53 -32 -51
rect -66 -119 -32 -91
rect -66 -125 -32 -119
rect -66 -187 -32 -163
rect -66 -197 -32 -187
rect -66 -255 -32 -235
rect -66 -269 -32 -255
rect 32 255 66 269
rect 32 235 66 255
rect 32 187 66 197
rect 32 163 66 187
rect 32 119 66 125
rect 32 91 66 119
rect 32 51 66 53
rect 32 19 66 51
rect 32 -51 66 -19
rect 32 -53 66 -51
rect 32 -119 66 -91
rect 32 -125 66 -119
rect 32 -187 66 -163
rect 32 -197 66 -187
rect 32 -255 66 -235
rect 32 -269 66 -255
<< metal1 >>
rect -72 269 -26 300
rect -72 235 -66 269
rect -32 235 -26 269
rect -72 197 -26 235
rect -72 163 -66 197
rect -32 163 -26 197
rect -72 125 -26 163
rect -72 91 -66 125
rect -32 91 -26 125
rect -72 53 -26 91
rect -72 19 -66 53
rect -32 19 -26 53
rect -72 -19 -26 19
rect -72 -53 -66 -19
rect -32 -53 -26 -19
rect -72 -91 -26 -53
rect -72 -125 -66 -91
rect -32 -125 -26 -91
rect -72 -163 -26 -125
rect -72 -197 -66 -163
rect -32 -197 -26 -163
rect -72 -235 -26 -197
rect -72 -269 -66 -235
rect -32 -269 -26 -235
rect -72 -300 -26 -269
rect 26 269 72 300
rect 26 235 32 269
rect 66 235 72 269
rect 26 197 72 235
rect 26 163 32 197
rect 66 163 72 197
rect 26 125 72 163
rect 26 91 32 125
rect 66 91 72 125
rect 26 53 72 91
rect 26 19 32 53
rect 66 19 72 53
rect 26 -19 72 19
rect 26 -53 32 -19
rect 66 -53 72 -19
rect 26 -91 72 -53
rect 26 -125 32 -91
rect 66 -125 72 -91
rect 26 -163 72 -125
rect 26 -197 32 -163
rect 66 -197 72 -163
rect 26 -235 72 -197
rect 26 -269 32 -235
rect 66 -269 72 -235
rect 26 -300 72 -269
<< end >>
