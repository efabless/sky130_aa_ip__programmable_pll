magic
tech sky130A
magscale 1 2
timestamp 1717685973
<< pwell >>
rect -134 -126 134 126
<< nmos >>
rect -50 -100 50 100
<< ndiff >>
rect -108 85 -50 100
rect -108 51 -96 85
rect -62 51 -50 85
rect -108 17 -50 51
rect -108 -17 -96 17
rect -62 -17 -50 17
rect -108 -51 -50 -17
rect -108 -85 -96 -51
rect -62 -85 -50 -51
rect -108 -100 -50 -85
rect 50 85 108 100
rect 50 51 62 85
rect 96 51 108 85
rect 50 17 108 51
rect 50 -17 62 17
rect 96 -17 108 17
rect 50 -51 108 -17
rect 50 -85 62 -51
rect 96 -85 108 -51
rect 50 -100 108 -85
<< ndiffc >>
rect -96 51 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -51
rect 62 51 96 85
rect 62 -17 96 17
rect 62 -85 96 -51
<< poly >>
rect -50 100 50 126
rect -50 -126 50 -100
<< locali >>
rect -96 85 -62 104
rect -96 17 -62 19
rect -96 -19 -62 -17
rect -96 -104 -62 -85
rect 62 85 96 104
rect 62 17 96 19
rect 62 -19 96 -17
rect 62 -104 96 -85
<< viali >>
rect -96 51 -62 53
rect -96 19 -62 51
rect -96 -51 -62 -19
rect -96 -53 -62 -51
rect 62 51 96 53
rect 62 19 96 51
rect 62 -51 96 -19
rect 62 -53 96 -51
<< metal1 >>
rect -102 53 -56 100
rect -102 19 -96 53
rect -62 19 -56 53
rect -102 -19 -56 19
rect -102 -53 -96 -19
rect -62 -53 -56 -19
rect -102 -100 -56 -53
rect 56 53 102 100
rect 56 19 62 53
rect 96 19 102 53
rect 56 -19 102 19
rect 56 -53 62 -19
rect 96 -53 102 -19
rect 56 -100 102 -53
<< properties >>
string GDS_END 29578
string GDS_FILE /home/shahid/Sky130Projects/top_layout/VCO.gds
string GDS_START 28486
<< end >>
