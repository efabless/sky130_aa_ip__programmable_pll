magic
tech sky130A
magscale 1 2
timestamp 1726363496
<< nwell >>
rect -11141 119923 -10767 119955
rect -12101 119237 -10767 119923
rect -12101 119150 -10760 119237
rect -12101 119076 -10566 119150
rect -11696 118858 -10566 119076
rect -11689 118628 -10566 118858
rect -11689 118373 -10581 118628
rect -11689 118238 -10537 118373
rect -11696 118151 -10537 118238
rect -11890 117655 -10537 118151
rect -11890 117629 -10947 117655
rect -8375 117408 -7502 118885
rect -11110 116255 -10736 116287
rect -7657 116263 -7283 116295
rect -12070 115569 -10736 116255
rect -12070 115482 -10729 115569
rect -12070 115408 -10535 115482
rect -11665 115190 -10535 115408
rect -11658 114960 -10535 115190
rect -8617 115577 -7283 116263
rect -8617 115490 -7276 115577
rect -8617 115416 -7082 115490
rect -8212 115198 -7082 115416
rect -11658 114705 -10550 114960
rect -11658 114570 -10506 114705
rect -8205 114968 -7082 115198
rect -8205 114713 -7097 114968
rect -11665 114483 -10506 114570
rect -11859 113987 -10506 114483
rect -8205 114578 -7053 114713
rect -8212 114491 -7053 114578
rect -11859 113961 -10916 113987
rect -8406 113995 -7053 114491
rect -8406 113969 -7463 113995
rect -11179 110559 -10805 110591
rect -12139 109873 -10805 110559
rect -12139 109786 -10798 109873
rect -12139 109712 -10604 109786
rect -11734 109494 -10604 109712
rect -11727 109264 -10604 109494
rect -11727 109009 -10619 109264
rect -11727 108874 -10575 109009
rect -11734 108787 -10575 108874
rect -11928 108291 -10575 108787
rect -11928 108265 -10985 108291
rect -8413 108044 -7540 109521
rect -11148 106891 -10774 106923
rect -7695 106899 -7321 106931
rect -12108 106205 -10774 106891
rect -12108 106118 -10767 106205
rect -12108 106044 -10573 106118
rect -11703 105826 -10573 106044
rect -11696 105596 -10573 105826
rect -8655 106213 -7321 106899
rect -8655 106126 -7314 106213
rect -8655 106052 -7120 106126
rect -8250 105834 -7120 106052
rect -11696 105341 -10588 105596
rect -11696 105206 -10544 105341
rect -8243 105604 -7120 105834
rect -8243 105349 -7135 105604
rect -11703 105119 -10544 105206
rect -11897 104623 -10544 105119
rect -8243 105214 -7091 105349
rect -8250 105127 -7091 105214
rect -11897 104597 -10954 104623
rect -8444 104631 -7091 105127
rect -8444 104605 -7501 104631
rect -11196 101406 -10822 101438
rect -12156 100720 -10822 101406
rect -12156 100633 -10815 100720
rect -12156 100559 -10621 100633
rect -11751 100341 -10621 100559
rect -11744 100111 -10621 100341
rect -11744 99856 -10636 100111
rect -11744 99721 -10592 99856
rect -11751 99634 -10592 99721
rect -11945 99138 -10592 99634
rect -11945 99112 -11002 99138
rect -8430 98891 -7557 100368
rect -11165 97738 -10791 97770
rect -7712 97746 -7338 97778
rect -12125 97052 -10791 97738
rect -12125 96965 -10784 97052
rect -12125 96891 -10590 96965
rect -11720 96673 -10590 96891
rect -11713 96443 -10590 96673
rect -8672 97060 -7338 97746
rect -8672 96973 -7331 97060
rect -8672 96899 -7137 96973
rect -8267 96681 -7137 96899
rect -11713 96188 -10605 96443
rect -11713 96053 -10561 96188
rect -8260 96451 -7137 96681
rect -8260 96196 -7152 96451
rect -11720 95966 -10561 96053
rect -11914 95470 -10561 95966
rect -8260 96061 -7108 96196
rect -8267 95974 -7108 96061
rect -11914 95444 -10971 95470
rect -8461 95478 -7108 95974
rect -8461 95452 -7518 95478
rect -11262 92652 -10888 92684
rect -12222 91966 -10888 92652
rect -12222 91879 -10881 91966
rect -12222 91805 -10687 91879
rect -11817 91587 -10687 91805
rect -11810 91357 -10687 91587
rect -11810 91102 -10702 91357
rect -11810 90967 -10658 91102
rect -11817 90880 -10658 90967
rect -12011 90384 -10658 90880
rect -12011 90358 -11068 90384
rect -8496 90137 -7623 91614
rect -11231 88984 -10857 89016
rect -7778 88992 -7404 89024
rect -12191 88298 -10857 88984
rect -12191 88211 -10850 88298
rect -12191 88137 -10656 88211
rect -11786 87919 -10656 88137
rect -11779 87689 -10656 87919
rect -8738 88306 -7404 88992
rect -8738 88219 -7397 88306
rect -8738 88145 -7203 88219
rect -8333 87927 -7203 88145
rect -11779 87434 -10671 87689
rect -11779 87299 -10627 87434
rect -8326 87697 -7203 87927
rect -8326 87442 -7218 87697
rect -11786 87212 -10627 87299
rect -11980 86716 -10627 87212
rect -8326 87307 -7174 87442
rect -8333 87220 -7174 87307
rect -11980 86690 -11037 86716
rect -8527 86724 -7174 87220
rect -8527 86698 -7584 86724
rect -11296 83454 -10922 83486
rect -12256 82768 -10922 83454
rect -12256 82681 -10915 82768
rect -12256 82607 -10721 82681
rect -11851 82389 -10721 82607
rect -11844 82159 -10721 82389
rect -11844 81904 -10736 82159
rect -11844 81769 -10692 81904
rect -11851 81682 -10692 81769
rect -12045 81186 -10692 81682
rect -12045 81160 -11102 81186
rect -8530 80939 -7657 82416
rect -11265 79786 -10891 79818
rect -7812 79794 -7438 79826
rect -12225 79100 -10891 79786
rect -12225 79013 -10884 79100
rect -12225 78939 -10690 79013
rect -11820 78721 -10690 78939
rect -11813 78491 -10690 78721
rect -8772 79108 -7438 79794
rect -8772 79021 -7431 79108
rect -8772 78947 -7237 79021
rect -8367 78729 -7237 78947
rect -11813 78236 -10705 78491
rect -11813 78101 -10661 78236
rect -8360 78499 -7237 78729
rect -8360 78244 -7252 78499
rect -11820 78014 -10661 78101
rect -12014 77518 -10661 78014
rect -8360 78109 -7208 78244
rect -8367 78022 -7208 78109
rect -12014 77492 -11071 77518
rect -8561 77526 -7208 78022
rect -8561 77500 -7618 77526
rect -11257 74591 -10883 74623
rect -12217 73905 -10883 74591
rect -12217 73818 -10876 73905
rect -12217 73744 -10682 73818
rect -11812 73526 -10682 73744
rect -11805 73296 -10682 73526
rect -11805 73041 -10697 73296
rect -11805 72906 -10653 73041
rect -11812 72819 -10653 72906
rect -12006 72323 -10653 72819
rect -12006 72297 -11063 72323
rect -8491 72076 -7618 73553
rect -11226 70923 -10852 70955
rect -7773 70931 -7399 70963
rect -12186 70237 -10852 70923
rect -12186 70150 -10845 70237
rect -12186 70076 -10651 70150
rect -11781 69858 -10651 70076
rect -11774 69628 -10651 69858
rect -8733 70245 -7399 70931
rect -8733 70158 -7392 70245
rect -8733 70084 -7198 70158
rect -8328 69866 -7198 70084
rect -11774 69373 -10666 69628
rect -11774 69238 -10622 69373
rect -8321 69636 -7198 69866
rect -8321 69381 -7213 69636
rect -11781 69151 -10622 69238
rect -11975 68655 -10622 69151
rect -8321 69246 -7169 69381
rect -8328 69159 -7169 69246
rect -11975 68629 -11032 68655
rect -8522 68663 -7169 69159
rect -8522 68637 -7579 68663
rect -11246 66151 -10872 66183
rect -12206 65465 -10872 66151
rect -12206 65378 -10865 65465
rect -12206 65304 -10671 65378
rect -11801 65086 -10671 65304
rect -11794 64856 -10671 65086
rect -11794 64601 -10686 64856
rect -11794 64466 -10642 64601
rect -11801 64379 -10642 64466
rect -11995 63883 -10642 64379
rect -11995 63857 -11052 63883
rect -8480 63636 -7607 65113
rect -11215 62483 -10841 62515
rect -7762 62491 -7388 62523
rect -12175 61797 -10841 62483
rect -12175 61710 -10834 61797
rect -12175 61636 -10640 61710
rect -11770 61418 -10640 61636
rect -11763 61188 -10640 61418
rect -8722 61805 -7388 62491
rect -8722 61718 -7381 61805
rect -8722 61644 -7187 61718
rect -8317 61426 -7187 61644
rect -11763 60933 -10655 61188
rect -11763 60798 -10611 60933
rect -8310 61196 -7187 61426
rect -8310 60941 -7202 61196
rect -11770 60711 -10611 60798
rect -11964 60215 -10611 60711
rect -8310 60806 -7158 60941
rect -8317 60719 -7158 60806
rect -11964 60189 -11021 60215
rect -8511 60223 -7158 60719
rect -8511 60197 -7568 60223
rect -11543 55240 -10511 57966
rect -9283 55187 -8829 57923
rect -7835 55209 -7381 57910
rect -11535 54360 -11082 54980
rect -9282 54932 -8829 55187
rect -10105 54410 -8829 54932
rect -7841 55174 -7381 55209
rect -9551 54399 -8829 54410
rect -11547 53926 -11089 53957
rect -11548 52501 -11089 53926
rect -9282 52910 -8829 54399
rect -7841 54368 -7382 55174
rect -9282 52569 -8818 52910
rect -7835 52848 -7382 54368
rect -11536 51585 -10855 52220
rect -9282 51589 -8829 52569
rect -11536 50639 -10855 51274
rect -9282 50644 -8309 51589
rect -9282 50643 -8829 50644
rect -13839 47081 -13385 49782
rect -13839 47046 -13379 47081
rect -13838 46240 -13379 47046
rect -12391 47059 -11937 49795
rect -13838 44720 -13385 46240
rect -12391 44782 -11938 47059
rect -12402 44441 -11938 44782
rect -12391 43837 -11938 44441
rect -14023 38820 -13548 40737
rect -14023 38819 -13621 38820
rect -14023 35820 -13548 37737
rect -11772 36822 -11297 40747
rect -7585 36822 -7110 40747
rect -5334 38820 -4859 40737
rect -5261 38819 -4859 38820
rect -11772 36300 -11183 36822
rect -7699 36300 -7110 36822
rect -11772 36213 -11377 36300
rect -7505 36213 -7110 36300
rect -14023 35819 -13621 35820
rect -14023 33320 -13548 35237
rect -11772 35217 -11384 36213
rect -7498 35217 -7110 36213
rect -5334 35820 -4859 37737
rect -5261 35819 -4859 35820
rect -11772 34695 -11185 35217
rect -7697 34695 -7110 35217
rect -11772 34608 -11379 34695
rect -7503 34608 -7110 34695
rect -11772 33613 -11386 34608
rect -7496 33613 -7110 34608
rect -14023 33319 -13621 33320
rect -14023 30820 -13548 32737
rect -11772 31627 -11299 33613
rect -11772 31341 -11316 31627
rect -11772 31000 -11305 31341
rect -7583 31627 -7110 33613
rect -5334 33320 -4859 35237
rect -5261 33319 -4859 33320
rect -7566 31341 -7110 31627
rect -14023 30819 -13621 30820
rect -14023 28320 -13548 30237
rect -14023 28319 -13621 28320
rect -14023 25820 -13548 27737
rect -11772 25987 -11316 31000
rect -10322 29542 -9869 31062
rect -10328 28736 -9869 29542
rect -9013 29542 -8560 31062
rect -7577 31000 -7110 31341
rect -9013 28736 -8554 29542
rect -10328 28701 -9868 28736
rect -10322 26000 -9868 28701
rect -9014 28701 -8554 28736
rect -9014 26000 -8560 28701
rect -7566 25987 -7110 31000
rect -5334 30820 -4859 32737
rect -5261 30819 -4859 30820
rect -5334 28320 -4859 30237
rect -5261 28319 -4859 28320
rect -6792 26257 -6339 26877
rect -5334 25820 -4859 27737
rect -14023 25819 -13621 25820
rect -5261 25819 -4859 25820
rect -10472 24417 -9595 25264
rect -5538 24390 -4661 25237
rect -11502 23467 -11049 24071
rect -11502 23126 -11038 23467
rect -6575 23467 -6122 24071
rect -11502 20849 -11049 23126
rect -10055 21668 -9602 23188
rect -11503 18113 -11049 20849
rect -10061 20862 -9602 21668
rect -6575 23126 -6111 23467
rect -8774 21445 -8400 21477
rect -10061 20827 -9601 20862
rect -10055 18126 -9601 20827
rect -8774 20759 -7440 21445
rect -8781 20672 -7440 20759
rect -8975 20598 -7440 20672
rect -6575 20849 -6122 23126
rect -5128 21668 -4675 23188
rect -8975 20380 -7845 20598
rect -8975 20150 -7852 20380
rect -8960 19895 -7852 20150
rect -9004 19760 -7852 19895
rect -9004 19673 -7845 19760
rect -9004 19177 -7651 19673
rect -8594 19151 -7651 19177
rect -6576 18113 -6122 20849
rect -5134 20862 -4675 21668
rect -5134 20827 -4674 20862
rect -5128 18126 -4674 20827
rect -12798 16456 -12424 16488
rect -7798 16456 -7424 16488
rect -12798 15770 -11464 16456
rect -12805 15683 -11464 15770
rect -12999 15609 -11464 15683
rect -7798 15770 -6464 16456
rect -7805 15683 -6464 15770
rect -12999 15391 -11869 15609
rect -12999 15161 -11876 15391
rect -12984 14906 -11876 15161
rect -13028 14771 -11876 14906
rect -7999 15609 -6464 15683
rect -7999 15391 -6869 15609
rect -7999 15161 -6876 15391
rect -7984 14906 -6876 15161
rect -13028 14684 -11869 14771
rect -13028 14188 -11675 14684
rect -12618 14162 -11675 14188
rect -8028 14771 -6876 14906
rect -8028 14684 -6869 14771
rect -8028 14188 -6675 14684
rect -7618 14162 -6675 14188
rect -7851 13782 -7393 13813
rect -11270 12760 -10589 13395
rect -11269 11855 -10588 12490
rect -7851 12357 -7392 13782
rect -5936 13135 -5562 13853
rect -5943 13048 -5562 13135
rect -6137 12526 -5562 13048
rect -5915 11952 -5457 11983
rect -14093 10343 -13634 11768
rect -11540 10649 -10595 11594
rect -7845 11193 -7471 11911
rect -7852 11106 -7471 11193
rect -8046 10584 -7471 11106
rect -5915 10527 -5456 11952
rect -14092 10312 -13634 10343
rect 14469 9053 15950 10215
rect 15664 8806 15948 9053
rect 8096 6634 12765 7919
rect 8190 6589 12714 6634
rect 19746 3116 22156 3612
rect -13457 1513 -5857 2282
rect -3632 1775 -1222 2271
rect 4467 1951 6877 2447
rect 1717 1883 1921 1927
rect 577 1881 913 1883
rect 1717 1881 2979 1883
rect -2782 528 -1222 1024
rect 577 981 2979 1881
rect 7570 1795 15170 2564
rect 20596 1869 22156 2365
rect 577 979 913 981
rect 1717 979 2979 981
rect 1717 935 1921 979
rect 5317 704 6877 1200
rect -5100 -597 -2690 -101
rect 4482 -739 6892 -243
rect 7529 -961 15129 -192
rect 19918 -234 22328 262
rect -4250 -1844 -2690 -1348
rect 5332 -1986 6892 -1490
rect 20768 -1481 22328 -985
rect 42360 3126 45096 3127
rect 39138 2673 45096 3126
rect 39742 2662 40083 2673
rect 28061 2124 29270 2382
rect 28061 2053 29557 2124
rect 32916 2117 34125 2375
rect 27673 1406 29557 2053
rect 32916 2046 34412 2117
rect 29269 1405 29557 1406
rect 30282 378 31676 1902
rect 32528 1399 34412 2046
rect 34124 1398 34412 1399
rect 35017 401 36411 1924
rect 36738 444 38132 1881
rect 41541 1679 42382 1685
rect 40021 1226 45083 1679
rect 45531 1316 46151 1769
rect 42347 1225 45083 1226
rect 50848 2572 58448 3341
rect 50645 -339 58245 430
rect 50645 -3386 58245 -2617
rect 62345 -3100 64755 -2604
rect 63195 -4347 64755 -3851
rect -15097 -16843 -7497 -16074
rect -15187 -18206 -12451 -18205
rect -15187 -18659 -10125 -18206
rect -12486 -18665 -11645 -18659
rect -22786 -18988 -21361 -18987
rect -22786 -19446 -21330 -18988
rect -8923 -19069 -8076 -18192
rect -7494 -18792 -5576 -18390
rect -4994 -18792 -3076 -18390
rect -2494 -18792 -576 -18390
rect 6 -18792 1924 -18390
rect 2506 -18792 4424 -18390
rect 5506 -18792 7424 -18390
rect -7493 -18865 -5576 -18792
rect -4993 -18865 -3076 -18792
rect -2493 -18865 -576 -18792
rect 7 -18865 1924 -18792
rect 2507 -18865 4424 -18792
rect 5507 -18865 7424 -18792
rect -20787 -19467 -19460 -19093
rect -20787 -19474 -20178 -19467
rect -20787 -19668 -20265 -19474
rect -10187 -19653 -9846 -19642
rect -19151 -20400 -18629 -20206
rect -17704 -20400 -16857 -19995
rect -15200 -20106 -9242 -19653
rect -15200 -20107 -12464 -20106
rect -7056 -20323 -6436 -19870
rect -19151 -20407 -18542 -20400
rect -17922 -20407 -16857 -20400
rect -20956 -20924 -19531 -20923
rect -22729 -21376 -21402 -21002
rect -22729 -21383 -22120 -21376
rect -20956 -21382 -19500 -20924
rect -19151 -20955 -16857 -20407
rect -19151 -21149 -16825 -20955
rect -19125 -21329 -16825 -21149
rect -19125 -21336 -17543 -21329
rect -22729 -21577 -22207 -21383
rect -19125 -21515 -17630 -21336
rect -19125 -21559 -18407 -21515
rect -18152 -21530 -17630 -21515
rect -14162 -21376 -13640 -21182
rect -12715 -21376 -11868 -20971
rect -7326 -21027 7434 -20641
rect 26910 -20733 27628 -20689
rect 27883 -20733 28405 -20718
rect 26910 -20912 28405 -20733
rect 35350 -20744 36068 -20700
rect 36323 -20744 36845 -20729
rect 21861 -20913 24597 -20912
rect -7326 -21097 300 -21027
rect 1295 -21029 7434 -21027
rect 1295 -21034 1904 -21029
rect -2313 -21108 -1972 -21097
rect -1686 -21114 300 -21097
rect -14162 -21383 -13553 -21376
rect -12933 -21383 -11868 -21376
rect -14162 -21931 -11868 -21383
rect 1382 -21228 1904 -21034
rect 2900 -21036 7434 -21029
rect 2987 -21116 7434 -21036
rect 2987 -21230 3509 -21116
rect -14162 -22125 -11836 -21931
rect 19535 -21366 24597 -20913
rect 26910 -20919 28492 -20912
rect 26910 -21099 29210 -20919
rect 26884 -21293 29210 -21099
rect 35350 -20923 36845 -20744
rect 44213 -20783 44931 -20739
rect 45186 -20783 45708 -20768
rect 53411 -20749 54129 -20705
rect 54384 -20749 54906 -20734
rect 62165 -20683 62883 -20639
rect 63138 -20683 63660 -20668
rect 71318 -20666 72036 -20622
rect 72291 -20666 72813 -20651
rect 80682 -20628 81400 -20584
rect 81655 -20628 82177 -20613
rect 35350 -20930 36932 -20923
rect 35350 -21110 37650 -20930
rect 21055 -21372 21896 -21366
rect -4612 -22091 -3771 -22085
rect -14136 -22305 -11836 -22125
rect -14136 -22312 -12554 -22305
rect -14136 -22491 -12641 -22312
rect -14136 -22535 -13418 -22491
rect -13163 -22506 -12641 -22491
rect -7313 -22544 -2251 -22091
rect 17331 -22360 18276 -21840
rect 26884 -21841 29178 -21293
rect 26884 -21848 27493 -21841
rect 28113 -21848 29178 -21841
rect 26884 -22042 27406 -21848
rect 19256 -22360 19597 -22349
rect -7313 -22545 -4577 -22544
rect 17330 -22813 24610 -22360
rect 28331 -22253 29178 -21848
rect 30323 -22011 31800 -21138
rect 35324 -21304 37650 -21110
rect 44213 -20962 45708 -20783
rect 53411 -20928 54906 -20749
rect 62165 -20862 63660 -20683
rect 71318 -20845 72813 -20666
rect 80682 -20807 82177 -20628
rect 80682 -20814 82264 -20807
rect 71318 -20852 72900 -20845
rect 62165 -20869 63747 -20862
rect 53411 -20935 54993 -20928
rect 44213 -20969 45795 -20962
rect 44213 -21149 46513 -20969
rect 53411 -21115 55711 -20935
rect 62165 -21049 64465 -20869
rect 71318 -21032 73618 -20852
rect 80682 -20994 82982 -20814
rect 35324 -21852 37618 -21304
rect 35324 -21859 35933 -21852
rect 36553 -21859 37618 -21852
rect 35324 -22053 35846 -21859
rect 21086 -23082 21619 -22813
rect 21874 -22814 24610 -22813
rect 36771 -22264 37618 -21859
rect 38763 -22022 40240 -21149
rect 44187 -21343 46513 -21149
rect 44187 -21891 46481 -21343
rect 44187 -21898 44796 -21891
rect 45416 -21898 46481 -21891
rect 44187 -22092 44709 -21898
rect -15187 -23133 -12451 -23132
rect -15187 -23586 -10125 -23133
rect -12486 -23592 -11645 -23586
rect -8896 -24003 -8049 -23126
rect -7313 -23400 -4577 -23399
rect -7313 -23853 -2251 -23400
rect 21097 -23636 21619 -23082
rect 45634 -22303 46481 -21898
rect 47626 -22061 49103 -21188
rect 53385 -21309 55711 -21115
rect 53385 -21857 55679 -21309
rect 53385 -21864 53994 -21857
rect 54614 -21864 55679 -21857
rect 53385 -22058 53907 -21864
rect 54832 -22269 55679 -21864
rect 56824 -22027 58301 -21154
rect 62139 -21243 64465 -21049
rect 62139 -21791 64433 -21243
rect 62139 -21798 62748 -21791
rect 63368 -21798 64433 -21791
rect 62139 -21992 62661 -21798
rect 63586 -22203 64433 -21798
rect 65578 -21961 67055 -21088
rect 71292 -21226 73618 -21032
rect 71292 -21774 73586 -21226
rect 71292 -21781 71901 -21774
rect 72521 -21781 73586 -21774
rect 71292 -21975 71814 -21781
rect 72739 -22186 73586 -21781
rect 74731 -21944 76208 -21071
rect 80656 -21188 82982 -20994
rect 80656 -21736 82950 -21188
rect 80656 -21743 81265 -21736
rect 81885 -21743 82950 -21736
rect 80656 -21937 81178 -21743
rect 82103 -22148 82950 -21743
rect 84095 -21906 85572 -21033
rect -4612 -23859 -3771 -23853
rect -22664 -25071 -21719 -24126
rect -21458 -24800 -20823 -24119
rect -20553 -24801 -19918 -24120
rect -10187 -24580 -9846 -24569
rect -19151 -25400 -18629 -25206
rect -17704 -25400 -16857 -24995
rect -15200 -25033 -9242 -24580
rect -2313 -24847 -1972 -24836
rect -1686 -24847 300 -24830
rect -7326 -24917 300 -24847
rect 1382 -24910 1904 -24716
rect 2987 -24828 3509 -24714
rect 2987 -24908 7434 -24828
rect 1295 -24915 1904 -24910
rect 2900 -24915 7434 -24908
rect 1295 -24917 7434 -24915
rect -15200 -25034 -12464 -25033
rect -7326 -25303 7434 -24917
rect 17326 -25067 17961 -24386
rect 18272 -25067 18907 -24386
rect 19188 -25078 20644 -24620
rect 21047 -25066 21667 -24613
rect 21927 -25074 24653 -24042
rect 26902 -24186 27620 -24142
rect 27875 -24186 28397 -24171
rect 26902 -24365 28397 -24186
rect 30570 -24217 31288 -24173
rect 31543 -24217 32065 -24202
rect 35342 -24197 36060 -24153
rect 36315 -24197 36837 -24182
rect 26902 -24372 28484 -24365
rect 26902 -24552 29202 -24372
rect 26876 -24746 29202 -24552
rect 30570 -24396 32065 -24217
rect 35342 -24376 36837 -24197
rect 39010 -24228 39728 -24184
rect 39983 -24228 40505 -24213
rect 35342 -24383 36924 -24376
rect 30570 -24403 32152 -24396
rect 30570 -24583 32870 -24403
rect 35342 -24563 37642 -24383
rect 19188 -25079 20613 -25078
rect 26876 -25294 29170 -24746
rect 26876 -25301 27485 -25294
rect 28105 -25301 29170 -25294
rect -19151 -25407 -18542 -25400
rect -17922 -25407 -16857 -25400
rect -19151 -25955 -16857 -25407
rect 13746 -25469 16482 -25468
rect 10524 -25922 16482 -25469
rect 26876 -25495 27398 -25301
rect 11128 -25933 11469 -25922
rect -19151 -26149 -16825 -25955
rect 28323 -25706 29170 -25301
rect 30544 -24777 32870 -24583
rect 35316 -24757 37642 -24563
rect 39010 -24407 40505 -24228
rect 44205 -24236 44923 -24192
rect 45178 -24236 45700 -24221
rect 39010 -24414 40592 -24407
rect 39010 -24594 41310 -24414
rect 30544 -25325 32838 -24777
rect 30544 -25332 31153 -25325
rect 31773 -25332 32838 -25325
rect 30544 -25526 31066 -25332
rect -19125 -26329 -16825 -26149
rect 31991 -25737 32838 -25332
rect 35316 -25305 37610 -24757
rect 35316 -25312 35925 -25305
rect 36545 -25312 37610 -25305
rect 35316 -25506 35838 -25312
rect 36763 -25717 37610 -25312
rect 38984 -24788 41310 -24594
rect 44205 -24415 45700 -24236
rect 47873 -24267 48591 -24223
rect 48846 -24267 49368 -24252
rect 53403 -24202 54121 -24158
rect 54376 -24202 54898 -24187
rect 44205 -24422 45787 -24415
rect 44205 -24602 46505 -24422
rect 38984 -25336 41278 -24788
rect 38984 -25343 39593 -25336
rect 40213 -25343 41278 -25336
rect 38984 -25537 39506 -25343
rect 40431 -25748 41278 -25343
rect 44179 -24796 46505 -24602
rect 47873 -24446 49368 -24267
rect 53403 -24381 54898 -24202
rect 57071 -24233 57789 -24189
rect 58044 -24233 58566 -24218
rect 62157 -24136 62875 -24092
rect 63130 -24136 63652 -24121
rect 53403 -24388 54985 -24381
rect 47873 -24453 49455 -24446
rect 47873 -24633 50173 -24453
rect 53403 -24568 55703 -24388
rect 44179 -25344 46473 -24796
rect 44179 -25351 44788 -25344
rect 45408 -25351 46473 -25344
rect 44179 -25545 44701 -25351
rect 45626 -25756 46473 -25351
rect 47847 -24827 50173 -24633
rect 53377 -24762 55703 -24568
rect 57071 -24412 58566 -24233
rect 62157 -24315 63652 -24136
rect 65825 -24167 66543 -24123
rect 66798 -24167 67320 -24152
rect 71310 -24119 72028 -24075
rect 72283 -24119 72805 -24104
rect 62157 -24322 63739 -24315
rect 57071 -24419 58653 -24412
rect 57071 -24599 59371 -24419
rect 62157 -24502 64457 -24322
rect 47847 -25375 50141 -24827
rect 47847 -25382 48456 -25375
rect 49076 -25382 50141 -25375
rect 47847 -25576 48369 -25382
rect -19125 -26336 -17543 -26329
rect 49294 -25787 50141 -25382
rect 53377 -25310 55671 -24762
rect 53377 -25317 53986 -25310
rect 54606 -25317 55671 -25310
rect 53377 -25511 53899 -25317
rect -19125 -26515 -17630 -26336
rect -19125 -26559 -18407 -26515
rect -18152 -26530 -17630 -26515
rect 54824 -25722 55671 -25317
rect 57045 -24793 59371 -24599
rect 62131 -24696 64457 -24502
rect 65825 -24346 67320 -24167
rect 71310 -24298 72805 -24119
rect 74978 -24150 75696 -24106
rect 75951 -24150 76473 -24135
rect 80674 -24081 81392 -24037
rect 81647 -24081 82169 -24066
rect 71310 -24305 72892 -24298
rect 65825 -24353 67407 -24346
rect 65825 -24533 68125 -24353
rect 71310 -24485 73610 -24305
rect 57045 -25341 59339 -24793
rect 57045 -25348 57654 -25341
rect 58274 -25348 59339 -25341
rect 57045 -25542 57567 -25348
rect 58492 -25753 59339 -25348
rect 62131 -25244 64425 -24696
rect 62131 -25251 62740 -25244
rect 63360 -25251 64425 -25244
rect 62131 -25445 62653 -25251
rect 63578 -25656 64425 -25251
rect 65799 -24727 68125 -24533
rect 71284 -24679 73610 -24485
rect 74978 -24329 76473 -24150
rect 80674 -24260 82169 -24081
rect 84342 -24112 85060 -24068
rect 85315 -24112 85837 -24097
rect 80674 -24267 82256 -24260
rect 74978 -24336 76560 -24329
rect 74978 -24516 77278 -24336
rect 80674 -24447 82974 -24267
rect 65799 -25275 68093 -24727
rect 65799 -25282 66408 -25275
rect 67028 -25282 68093 -25275
rect 65799 -25476 66321 -25282
rect 67246 -25687 68093 -25282
rect 71284 -25227 73578 -24679
rect 71284 -25234 71893 -25227
rect 72513 -25234 73578 -25227
rect 71284 -25428 71806 -25234
rect 72731 -25639 73578 -25234
rect 74952 -24710 77278 -24516
rect 80648 -24641 82974 -24447
rect 84342 -24291 85837 -24112
rect 84342 -24298 85924 -24291
rect 84342 -24478 86642 -24298
rect 74952 -25258 77246 -24710
rect 74952 -25265 75561 -25258
rect 76181 -25265 77246 -25258
rect 74952 -25459 75474 -25265
rect 76399 -25670 77246 -25265
rect 80648 -25189 82942 -24641
rect 80648 -25196 81257 -25189
rect 81877 -25196 82942 -25189
rect 80648 -25390 81170 -25196
rect 82095 -25601 82942 -25196
rect 84316 -24672 86642 -24478
rect 84316 -25220 86610 -24672
rect 84316 -25227 84925 -25220
rect 85545 -25227 86610 -25220
rect 84316 -25421 84838 -25227
rect 85763 -25632 86610 -25227
rect 12927 -26916 13768 -26910
rect -7493 -27152 -5576 -27079
rect -4993 -27152 -3076 -27079
rect -2493 -27152 -576 -27079
rect 7 -27152 1924 -27079
rect 2507 -27152 4424 -27079
rect 5507 -27152 7424 -27079
rect -23001 -27623 -21545 -27165
rect -7494 -27554 -5576 -27152
rect -4994 -27554 -3076 -27152
rect -2494 -27554 -576 -27152
rect 6 -27554 1924 -27152
rect 2506 -27554 4424 -27152
rect 5506 -27554 7424 -27152
rect 11407 -27369 16469 -26916
rect 13733 -27370 16469 -27369
rect -22970 -27624 -21545 -27623
rect -26074 -41571 -25305 -33971
rect -14489 -34797 -11753 -34796
rect -14489 -35250 -9427 -34797
rect -11788 -35256 -10947 -35250
rect -22088 -35579 -20663 -35578
rect -22088 -36037 -20632 -35579
rect -8225 -35660 -7378 -34783
rect -6796 -35383 -4878 -34981
rect -4296 -35383 -2378 -34981
rect -1796 -35383 122 -34981
rect 704 -35383 2622 -34981
rect 3204 -35383 5122 -34981
rect 6204 -35383 8122 -34981
rect -6795 -35456 -4878 -35383
rect -4295 -35456 -2378 -35383
rect -1795 -35456 122 -35383
rect 705 -35456 2622 -35383
rect 3205 -35456 5122 -35383
rect 6205 -35456 8122 -35383
rect -20089 -36058 -18762 -35684
rect -20089 -36065 -19480 -36058
rect -20089 -36259 -19567 -36065
rect -9489 -36244 -9148 -36233
rect -18453 -36991 -17931 -36797
rect -17006 -36991 -16159 -36586
rect -14502 -36697 -8544 -36244
rect -14502 -36698 -11766 -36697
rect -6358 -36914 -5738 -36461
rect -18453 -36998 -17844 -36991
rect -17224 -36998 -16159 -36991
rect -20258 -37515 -18833 -37514
rect -22031 -37967 -20704 -37593
rect -22031 -37974 -21422 -37967
rect -20258 -37973 -18802 -37515
rect -18453 -37546 -16159 -36998
rect -18453 -37740 -16127 -37546
rect -18427 -37920 -16127 -37740
rect -18427 -37927 -16845 -37920
rect -22031 -38168 -21509 -37974
rect -18427 -38106 -16932 -37927
rect -18427 -38150 -17709 -38106
rect -17454 -38121 -16932 -38106
rect -13464 -37967 -12942 -37773
rect -12017 -37967 -11170 -37562
rect -6628 -37618 8132 -37232
rect 27608 -37324 28326 -37280
rect 28581 -37324 29103 -37309
rect 27608 -37503 29103 -37324
rect 36048 -37335 36766 -37291
rect 37021 -37335 37543 -37320
rect 22559 -37504 25295 -37503
rect -6628 -37688 998 -37618
rect 1993 -37620 8132 -37618
rect 1993 -37625 2602 -37620
rect -1615 -37699 -1274 -37688
rect -988 -37705 998 -37688
rect -13464 -37974 -12855 -37967
rect -12235 -37974 -11170 -37967
rect -13464 -38522 -11170 -37974
rect 2080 -37819 2602 -37625
rect 3598 -37627 8132 -37620
rect 3685 -37707 8132 -37627
rect 3685 -37821 4207 -37707
rect -13464 -38716 -11138 -38522
rect 20233 -37957 25295 -37504
rect 27608 -37510 29190 -37503
rect 27608 -37690 29908 -37510
rect 27582 -37884 29908 -37690
rect 36048 -37514 37543 -37335
rect 44911 -37374 45629 -37330
rect 45884 -37374 46406 -37359
rect 54109 -37340 54827 -37296
rect 55082 -37340 55604 -37325
rect 62863 -37274 63581 -37230
rect 63836 -37274 64358 -37259
rect 72016 -37257 72734 -37213
rect 72989 -37257 73511 -37242
rect 81380 -37219 82098 -37175
rect 82353 -37219 82875 -37204
rect 36048 -37521 37630 -37514
rect 36048 -37701 38348 -37521
rect 21753 -37963 22594 -37957
rect -3914 -38682 -3073 -38676
rect -13438 -38896 -11138 -38716
rect -13438 -38903 -11856 -38896
rect -13438 -39082 -11943 -38903
rect -13438 -39126 -12720 -39082
rect -12465 -39097 -11943 -39082
rect -6615 -39135 -1553 -38682
rect 18029 -38951 18974 -38431
rect 27582 -38432 29876 -37884
rect 27582 -38439 28191 -38432
rect 28811 -38439 29876 -38432
rect 27582 -38633 28104 -38439
rect 19954 -38951 20295 -38940
rect -6615 -39136 -3879 -39135
rect 18028 -39404 25308 -38951
rect 29029 -38844 29876 -38439
rect 31021 -38602 32498 -37729
rect 36022 -37895 38348 -37701
rect 44911 -37553 46406 -37374
rect 54109 -37519 55604 -37340
rect 62863 -37453 64358 -37274
rect 72016 -37436 73511 -37257
rect 81380 -37398 82875 -37219
rect 81380 -37405 82962 -37398
rect 72016 -37443 73598 -37436
rect 62863 -37460 64445 -37453
rect 54109 -37526 55691 -37519
rect 44911 -37560 46493 -37553
rect 44911 -37740 47211 -37560
rect 54109 -37706 56409 -37526
rect 62863 -37640 65163 -37460
rect 72016 -37623 74316 -37443
rect 81380 -37585 83680 -37405
rect 36022 -38443 38316 -37895
rect 36022 -38450 36631 -38443
rect 37251 -38450 38316 -38443
rect 36022 -38644 36544 -38450
rect 21784 -39673 22317 -39404
rect 22572 -39405 25308 -39404
rect 37469 -38855 38316 -38450
rect 39461 -38613 40938 -37740
rect 44885 -37934 47211 -37740
rect 44885 -38482 47179 -37934
rect 44885 -38489 45494 -38482
rect 46114 -38489 47179 -38482
rect 44885 -38683 45407 -38489
rect -14489 -39724 -11753 -39723
rect -14489 -40177 -9427 -39724
rect -11788 -40183 -10947 -40177
rect -8198 -40594 -7351 -39717
rect -6615 -39991 -3879 -39990
rect -6615 -40444 -1553 -39991
rect 21795 -40227 22317 -39673
rect 46332 -38894 47179 -38489
rect 48324 -38652 49801 -37779
rect 54083 -37900 56409 -37706
rect 54083 -38448 56377 -37900
rect 54083 -38455 54692 -38448
rect 55312 -38455 56377 -38448
rect 54083 -38649 54605 -38455
rect 55530 -38860 56377 -38455
rect 57522 -38618 58999 -37745
rect 62837 -37834 65163 -37640
rect 62837 -38382 65131 -37834
rect 62837 -38389 63446 -38382
rect 64066 -38389 65131 -38382
rect 62837 -38583 63359 -38389
rect 64284 -38794 65131 -38389
rect 66276 -38552 67753 -37679
rect 71990 -37817 74316 -37623
rect 71990 -38365 74284 -37817
rect 71990 -38372 72599 -38365
rect 73219 -38372 74284 -38365
rect 71990 -38566 72512 -38372
rect 73437 -38777 74284 -38372
rect 75429 -38535 76906 -37662
rect 81354 -37779 83680 -37585
rect 81354 -38327 83648 -37779
rect 81354 -38334 81963 -38327
rect 82583 -38334 83648 -38327
rect 81354 -38528 81876 -38334
rect 82801 -38739 83648 -38334
rect 84793 -38497 86270 -37624
rect -3914 -40450 -3073 -40444
rect -21966 -41662 -21021 -40717
rect -20760 -41391 -20125 -40710
rect -19855 -41392 -19220 -40711
rect -9489 -41171 -9148 -41160
rect -18453 -41991 -17931 -41797
rect -17006 -41991 -16159 -41586
rect -14502 -41624 -8544 -41171
rect -1615 -41438 -1274 -41427
rect -988 -41438 998 -41421
rect -6628 -41508 998 -41438
rect 2080 -41501 2602 -41307
rect 3685 -41419 4207 -41305
rect 3685 -41499 8132 -41419
rect 1993 -41506 2602 -41501
rect 3598 -41506 8132 -41499
rect 1993 -41508 8132 -41506
rect -14502 -41625 -11766 -41624
rect -6628 -41894 8132 -41508
rect 18024 -41658 18659 -40977
rect 18970 -41658 19605 -40977
rect 19886 -41669 21342 -41211
rect 21745 -41657 22365 -41204
rect 22625 -41665 25351 -40633
rect 27600 -40777 28318 -40733
rect 28573 -40777 29095 -40762
rect 27600 -40956 29095 -40777
rect 31268 -40808 31986 -40764
rect 32241 -40808 32763 -40793
rect 36040 -40788 36758 -40744
rect 37013 -40788 37535 -40773
rect 27600 -40963 29182 -40956
rect 27600 -41143 29900 -40963
rect 27574 -41337 29900 -41143
rect 31268 -40987 32763 -40808
rect 36040 -40967 37535 -40788
rect 39708 -40819 40426 -40775
rect 40681 -40819 41203 -40804
rect 36040 -40974 37622 -40967
rect 31268 -40994 32850 -40987
rect 31268 -41174 33568 -40994
rect 36040 -41154 38340 -40974
rect 19886 -41670 21311 -41669
rect 27574 -41885 29868 -41337
rect 27574 -41892 28183 -41885
rect 28803 -41892 29868 -41885
rect -18453 -41998 -17844 -41991
rect -17224 -41998 -16159 -41991
rect -18453 -42546 -16159 -41998
rect 14444 -42060 17180 -42059
rect 11222 -42513 17180 -42060
rect 27574 -42086 28096 -41892
rect 11826 -42524 12167 -42513
rect -18453 -42740 -16127 -42546
rect 29021 -42297 29868 -41892
rect 31242 -41368 33568 -41174
rect 36014 -41348 38340 -41154
rect 39708 -40998 41203 -40819
rect 44903 -40827 45621 -40783
rect 45876 -40827 46398 -40812
rect 39708 -41005 41290 -40998
rect 39708 -41185 42008 -41005
rect 31242 -41916 33536 -41368
rect 31242 -41923 31851 -41916
rect 32471 -41923 33536 -41916
rect 31242 -42117 31764 -41923
rect -18427 -42920 -16127 -42740
rect 32689 -42328 33536 -41923
rect 36014 -41896 38308 -41348
rect 36014 -41903 36623 -41896
rect 37243 -41903 38308 -41896
rect 36014 -42097 36536 -41903
rect 37461 -42308 38308 -41903
rect 39682 -41379 42008 -41185
rect 44903 -41006 46398 -40827
rect 48571 -40858 49289 -40814
rect 49544 -40858 50066 -40843
rect 54101 -40793 54819 -40749
rect 55074 -40793 55596 -40778
rect 44903 -41013 46485 -41006
rect 44903 -41193 47203 -41013
rect 39682 -41927 41976 -41379
rect 39682 -41934 40291 -41927
rect 40911 -41934 41976 -41927
rect 39682 -42128 40204 -41934
rect 41129 -42339 41976 -41934
rect 44877 -41387 47203 -41193
rect 48571 -41037 50066 -40858
rect 54101 -40972 55596 -40793
rect 57769 -40824 58487 -40780
rect 58742 -40824 59264 -40809
rect 62855 -40727 63573 -40683
rect 63828 -40727 64350 -40712
rect 54101 -40979 55683 -40972
rect 48571 -41044 50153 -41037
rect 48571 -41224 50871 -41044
rect 54101 -41159 56401 -40979
rect 44877 -41935 47171 -41387
rect 44877 -41942 45486 -41935
rect 46106 -41942 47171 -41935
rect 44877 -42136 45399 -41942
rect 46324 -42347 47171 -41942
rect 48545 -41418 50871 -41224
rect 54075 -41353 56401 -41159
rect 57769 -41003 59264 -40824
rect 62855 -40906 64350 -40727
rect 66523 -40758 67241 -40714
rect 67496 -40758 68018 -40743
rect 72008 -40710 72726 -40666
rect 72981 -40710 73503 -40695
rect 62855 -40913 64437 -40906
rect 57769 -41010 59351 -41003
rect 57769 -41190 60069 -41010
rect 62855 -41093 65155 -40913
rect 48545 -41966 50839 -41418
rect 48545 -41973 49154 -41966
rect 49774 -41973 50839 -41966
rect 48545 -42167 49067 -41973
rect -18427 -42927 -16845 -42920
rect 49992 -42378 50839 -41973
rect 54075 -41901 56369 -41353
rect 54075 -41908 54684 -41901
rect 55304 -41908 56369 -41901
rect 54075 -42102 54597 -41908
rect -18427 -43106 -16932 -42927
rect -18427 -43150 -17709 -43106
rect -17454 -43121 -16932 -43106
rect 55522 -42313 56369 -41908
rect 57743 -41384 60069 -41190
rect 62829 -41287 65155 -41093
rect 66523 -40937 68018 -40758
rect 72008 -40889 73503 -40710
rect 75676 -40741 76394 -40697
rect 76649 -40741 77171 -40726
rect 81372 -40672 82090 -40628
rect 82345 -40672 82867 -40657
rect 72008 -40896 73590 -40889
rect 66523 -40944 68105 -40937
rect 66523 -41124 68823 -40944
rect 72008 -41076 74308 -40896
rect 57743 -41932 60037 -41384
rect 57743 -41939 58352 -41932
rect 58972 -41939 60037 -41932
rect 57743 -42133 58265 -41939
rect 59190 -42344 60037 -41939
rect 62829 -41835 65123 -41287
rect 62829 -41842 63438 -41835
rect 64058 -41842 65123 -41835
rect 62829 -42036 63351 -41842
rect 64276 -42247 65123 -41842
rect 66497 -41318 68823 -41124
rect 71982 -41270 74308 -41076
rect 75676 -40920 77171 -40741
rect 81372 -40851 82867 -40672
rect 85040 -40703 85758 -40659
rect 86013 -40703 86535 -40688
rect 81372 -40858 82954 -40851
rect 75676 -40927 77258 -40920
rect 75676 -41107 77976 -40927
rect 81372 -41038 83672 -40858
rect 66497 -41866 68791 -41318
rect 66497 -41873 67106 -41866
rect 67726 -41873 68791 -41866
rect 66497 -42067 67019 -41873
rect 67944 -42278 68791 -41873
rect 71982 -41818 74276 -41270
rect 71982 -41825 72591 -41818
rect 73211 -41825 74276 -41818
rect 71982 -42019 72504 -41825
rect 73429 -42230 74276 -41825
rect 75650 -41301 77976 -41107
rect 81346 -41232 83672 -41038
rect 85040 -40882 86535 -40703
rect 85040 -40889 86622 -40882
rect 85040 -41069 87340 -40889
rect 75650 -41849 77944 -41301
rect 75650 -41856 76259 -41849
rect 76879 -41856 77944 -41849
rect 75650 -42050 76172 -41856
rect 77097 -42261 77944 -41856
rect 81346 -41780 83640 -41232
rect 81346 -41787 81955 -41780
rect 82575 -41787 83640 -41780
rect 81346 -41981 81868 -41787
rect 82793 -42192 83640 -41787
rect 85014 -41263 87340 -41069
rect 85014 -41811 87308 -41263
rect 85014 -41818 85623 -41811
rect 86243 -41818 87308 -41811
rect 85014 -42012 85536 -41818
rect 86461 -42223 87308 -41818
rect 13625 -43507 14466 -43501
rect -6795 -43743 -4878 -43670
rect -4295 -43743 -2378 -43670
rect -1795 -43743 122 -43670
rect 705 -43743 2622 -43670
rect 3205 -43743 5122 -43670
rect 6205 -43743 8122 -43670
rect -22303 -44214 -20847 -43756
rect -6796 -44145 -4878 -43743
rect -4296 -44145 -2378 -43743
rect -1796 -44145 122 -43743
rect 704 -44145 2622 -43743
rect 3204 -44145 5122 -43743
rect 6204 -44145 8122 -43743
rect 12105 -43960 17167 -43507
rect 14431 -43961 17167 -43960
rect -22272 -44215 -20847 -44214
rect -27894 -59716 -27125 -52116
rect -13786 -52908 -11050 -52907
rect -13786 -53361 -8724 -52908
rect -11085 -53367 -10244 -53361
rect -21385 -53690 -19960 -53689
rect -21385 -54148 -19929 -53690
rect -7522 -53771 -6675 -52894
rect -6093 -53494 -4175 -53092
rect -3593 -53494 -1675 -53092
rect -1093 -53494 825 -53092
rect 1407 -53494 3325 -53092
rect 3907 -53494 5825 -53092
rect 6907 -53494 8825 -53092
rect -6092 -53567 -4175 -53494
rect -3592 -53567 -1675 -53494
rect -1092 -53567 825 -53494
rect 1408 -53567 3325 -53494
rect 3908 -53567 5825 -53494
rect 6908 -53567 8825 -53494
rect -19386 -54169 -18059 -53795
rect -19386 -54176 -18777 -54169
rect -19386 -54370 -18864 -54176
rect -8786 -54355 -8445 -54344
rect -17750 -55102 -17228 -54908
rect -16303 -55102 -15456 -54697
rect -13799 -54808 -7841 -54355
rect -13799 -54809 -11063 -54808
rect -5655 -55025 -5035 -54572
rect -17750 -55109 -17141 -55102
rect -16521 -55109 -15456 -55102
rect -19555 -55626 -18130 -55625
rect -21328 -56078 -20001 -55704
rect -21328 -56085 -20719 -56078
rect -19555 -56084 -18099 -55626
rect -17750 -55657 -15456 -55109
rect -17750 -55851 -15424 -55657
rect -17724 -56031 -15424 -55851
rect -17724 -56038 -16142 -56031
rect -21328 -56279 -20806 -56085
rect -17724 -56217 -16229 -56038
rect -17724 -56261 -17006 -56217
rect -16751 -56232 -16229 -56217
rect -12761 -56078 -12239 -55884
rect -11314 -56078 -10467 -55673
rect -5925 -55729 8835 -55343
rect 28311 -55435 29029 -55391
rect 29284 -55435 29806 -55420
rect 28311 -55614 29806 -55435
rect 36751 -55446 37469 -55402
rect 37724 -55446 38246 -55431
rect 23262 -55615 25998 -55614
rect -5925 -55799 1701 -55729
rect 2696 -55731 8835 -55729
rect 2696 -55736 3305 -55731
rect -912 -55810 -571 -55799
rect -285 -55816 1701 -55799
rect -12761 -56085 -12152 -56078
rect -11532 -56085 -10467 -56078
rect -12761 -56633 -10467 -56085
rect 2783 -55930 3305 -55736
rect 4301 -55738 8835 -55731
rect 4388 -55818 8835 -55738
rect 4388 -55932 4910 -55818
rect -12761 -56827 -10435 -56633
rect 20936 -56068 25998 -55615
rect 28311 -55621 29893 -55614
rect 28311 -55801 30611 -55621
rect 28285 -55995 30611 -55801
rect 36751 -55625 38246 -55446
rect 45614 -55485 46332 -55441
rect 46587 -55485 47109 -55470
rect 54812 -55451 55530 -55407
rect 55785 -55451 56307 -55436
rect 63566 -55385 64284 -55341
rect 64539 -55385 65061 -55370
rect 72719 -55368 73437 -55324
rect 73692 -55368 74214 -55353
rect 82083 -55330 82801 -55286
rect 83056 -55330 83578 -55315
rect 36751 -55632 38333 -55625
rect 36751 -55812 39051 -55632
rect 22456 -56074 23297 -56068
rect -3211 -56793 -2370 -56787
rect -12735 -57007 -10435 -56827
rect -12735 -57014 -11153 -57007
rect -12735 -57193 -11240 -57014
rect -12735 -57237 -12017 -57193
rect -11762 -57208 -11240 -57193
rect -5912 -57246 -850 -56793
rect 18732 -57062 19677 -56542
rect 28285 -56543 30579 -55995
rect 28285 -56550 28894 -56543
rect 29514 -56550 30579 -56543
rect 28285 -56744 28807 -56550
rect 20657 -57062 20998 -57051
rect -5912 -57247 -3176 -57246
rect 18731 -57515 26011 -57062
rect 29732 -56955 30579 -56550
rect 31724 -56713 33201 -55840
rect 36725 -56006 39051 -55812
rect 45614 -55664 47109 -55485
rect 54812 -55630 56307 -55451
rect 63566 -55564 65061 -55385
rect 72719 -55547 74214 -55368
rect 82083 -55509 83578 -55330
rect 82083 -55516 83665 -55509
rect 72719 -55554 74301 -55547
rect 63566 -55571 65148 -55564
rect 54812 -55637 56394 -55630
rect 45614 -55671 47196 -55664
rect 45614 -55851 47914 -55671
rect 54812 -55817 57112 -55637
rect 63566 -55751 65866 -55571
rect 72719 -55734 75019 -55554
rect 82083 -55696 84383 -55516
rect 36725 -56554 39019 -56006
rect 36725 -56561 37334 -56554
rect 37954 -56561 39019 -56554
rect 36725 -56755 37247 -56561
rect 22487 -57784 23020 -57515
rect 23275 -57516 26011 -57515
rect 38172 -56966 39019 -56561
rect 40164 -56724 41641 -55851
rect 45588 -56045 47914 -55851
rect 45588 -56593 47882 -56045
rect 45588 -56600 46197 -56593
rect 46817 -56600 47882 -56593
rect 45588 -56794 46110 -56600
rect -13786 -57835 -11050 -57834
rect -13786 -58288 -8724 -57835
rect -11085 -58294 -10244 -58288
rect -7495 -58705 -6648 -57828
rect -5912 -58102 -3176 -58101
rect -5912 -58555 -850 -58102
rect 22498 -58338 23020 -57784
rect 47035 -57005 47882 -56600
rect 49027 -56763 50504 -55890
rect 54786 -56011 57112 -55817
rect 54786 -56559 57080 -56011
rect 54786 -56566 55395 -56559
rect 56015 -56566 57080 -56559
rect 54786 -56760 55308 -56566
rect 56233 -56971 57080 -56566
rect 58225 -56729 59702 -55856
rect 63540 -55945 65866 -55751
rect 63540 -56493 65834 -55945
rect 63540 -56500 64149 -56493
rect 64769 -56500 65834 -56493
rect 63540 -56694 64062 -56500
rect 64987 -56905 65834 -56500
rect 66979 -56663 68456 -55790
rect 72693 -55928 75019 -55734
rect 72693 -56476 74987 -55928
rect 72693 -56483 73302 -56476
rect 73922 -56483 74987 -56476
rect 72693 -56677 73215 -56483
rect 74140 -56888 74987 -56483
rect 76132 -56646 77609 -55773
rect 82057 -55890 84383 -55696
rect 82057 -56438 84351 -55890
rect 82057 -56445 82666 -56438
rect 83286 -56445 84351 -56438
rect 82057 -56639 82579 -56445
rect 83504 -56850 84351 -56445
rect 85496 -56608 86973 -55735
rect -3211 -58561 -2370 -58555
rect -21263 -59773 -20318 -58828
rect -20057 -59502 -19422 -58821
rect -19152 -59503 -18517 -58822
rect -8786 -59282 -8445 -59271
rect -17750 -60102 -17228 -59908
rect -16303 -60102 -15456 -59697
rect -13799 -59735 -7841 -59282
rect -912 -59549 -571 -59538
rect -285 -59549 1701 -59532
rect -5925 -59619 1701 -59549
rect 2783 -59612 3305 -59418
rect 4388 -59530 4910 -59416
rect 4388 -59610 8835 -59530
rect 2696 -59617 3305 -59612
rect 4301 -59617 8835 -59610
rect 2696 -59619 8835 -59617
rect -13799 -59736 -11063 -59735
rect -5925 -60005 8835 -59619
rect 18727 -59769 19362 -59088
rect 19673 -59769 20308 -59088
rect 20589 -59780 22045 -59322
rect 22448 -59768 23068 -59315
rect 23328 -59776 26054 -58744
rect 28303 -58888 29021 -58844
rect 29276 -58888 29798 -58873
rect 28303 -59067 29798 -58888
rect 31971 -58919 32689 -58875
rect 32944 -58919 33466 -58904
rect 36743 -58899 37461 -58855
rect 37716 -58899 38238 -58884
rect 28303 -59074 29885 -59067
rect 28303 -59254 30603 -59074
rect 28277 -59448 30603 -59254
rect 31971 -59098 33466 -58919
rect 36743 -59078 38238 -58899
rect 40411 -58930 41129 -58886
rect 41384 -58930 41906 -58915
rect 36743 -59085 38325 -59078
rect 31971 -59105 33553 -59098
rect 31971 -59285 34271 -59105
rect 36743 -59265 39043 -59085
rect 20589 -59781 22014 -59780
rect 28277 -59996 30571 -59448
rect 28277 -60003 28886 -59996
rect 29506 -60003 30571 -59996
rect -17750 -60109 -17141 -60102
rect -16521 -60109 -15456 -60102
rect -17750 -60657 -15456 -60109
rect 15147 -60171 17883 -60170
rect 11925 -60624 17883 -60171
rect 28277 -60197 28799 -60003
rect 12529 -60635 12870 -60624
rect -17750 -60851 -15424 -60657
rect 29724 -60408 30571 -60003
rect 31945 -59479 34271 -59285
rect 36717 -59459 39043 -59265
rect 40411 -59109 41906 -58930
rect 45606 -58938 46324 -58894
rect 46579 -58938 47101 -58923
rect 40411 -59116 41993 -59109
rect 40411 -59296 42711 -59116
rect 31945 -60027 34239 -59479
rect 31945 -60034 32554 -60027
rect 33174 -60034 34239 -60027
rect 31945 -60228 32467 -60034
rect -17724 -61031 -15424 -60851
rect 33392 -60439 34239 -60034
rect 36717 -60007 39011 -59459
rect 36717 -60014 37326 -60007
rect 37946 -60014 39011 -60007
rect 36717 -60208 37239 -60014
rect 38164 -60419 39011 -60014
rect 40385 -59490 42711 -59296
rect 45606 -59117 47101 -58938
rect 49274 -58969 49992 -58925
rect 50247 -58969 50769 -58954
rect 54804 -58904 55522 -58860
rect 55777 -58904 56299 -58889
rect 45606 -59124 47188 -59117
rect 45606 -59304 47906 -59124
rect 40385 -60038 42679 -59490
rect 40385 -60045 40994 -60038
rect 41614 -60045 42679 -60038
rect 40385 -60239 40907 -60045
rect 41832 -60450 42679 -60045
rect 45580 -59498 47906 -59304
rect 49274 -59148 50769 -58969
rect 54804 -59083 56299 -58904
rect 58472 -58935 59190 -58891
rect 59445 -58935 59967 -58920
rect 63558 -58838 64276 -58794
rect 64531 -58838 65053 -58823
rect 54804 -59090 56386 -59083
rect 49274 -59155 50856 -59148
rect 49274 -59335 51574 -59155
rect 54804 -59270 57104 -59090
rect 45580 -60046 47874 -59498
rect 45580 -60053 46189 -60046
rect 46809 -60053 47874 -60046
rect 45580 -60247 46102 -60053
rect 47027 -60458 47874 -60053
rect 49248 -59529 51574 -59335
rect 54778 -59464 57104 -59270
rect 58472 -59114 59967 -58935
rect 63558 -59017 65053 -58838
rect 67226 -58869 67944 -58825
rect 68199 -58869 68721 -58854
rect 72711 -58821 73429 -58777
rect 73684 -58821 74206 -58806
rect 63558 -59024 65140 -59017
rect 58472 -59121 60054 -59114
rect 58472 -59301 60772 -59121
rect 63558 -59204 65858 -59024
rect 49248 -60077 51542 -59529
rect 49248 -60084 49857 -60077
rect 50477 -60084 51542 -60077
rect 49248 -60278 49770 -60084
rect -17724 -61038 -16142 -61031
rect 50695 -60489 51542 -60084
rect 54778 -60012 57072 -59464
rect 54778 -60019 55387 -60012
rect 56007 -60019 57072 -60012
rect 54778 -60213 55300 -60019
rect -17724 -61217 -16229 -61038
rect -17724 -61261 -17006 -61217
rect -16751 -61232 -16229 -61217
rect 56225 -60424 57072 -60019
rect 58446 -59495 60772 -59301
rect 63532 -59398 65858 -59204
rect 67226 -59048 68721 -58869
rect 72711 -59000 74206 -58821
rect 76379 -58852 77097 -58808
rect 77352 -58852 77874 -58837
rect 82075 -58783 82793 -58739
rect 83048 -58783 83570 -58768
rect 72711 -59007 74293 -59000
rect 67226 -59055 68808 -59048
rect 67226 -59235 69526 -59055
rect 72711 -59187 75011 -59007
rect 58446 -60043 60740 -59495
rect 58446 -60050 59055 -60043
rect 59675 -60050 60740 -60043
rect 58446 -60244 58968 -60050
rect 59893 -60455 60740 -60050
rect 63532 -59946 65826 -59398
rect 63532 -59953 64141 -59946
rect 64761 -59953 65826 -59946
rect 63532 -60147 64054 -59953
rect 64979 -60358 65826 -59953
rect 67200 -59429 69526 -59235
rect 72685 -59381 75011 -59187
rect 76379 -59031 77874 -58852
rect 82075 -58962 83570 -58783
rect 85743 -58814 86461 -58770
rect 86716 -58814 87238 -58799
rect 82075 -58969 83657 -58962
rect 76379 -59038 77961 -59031
rect 76379 -59218 78679 -59038
rect 82075 -59149 84375 -58969
rect 67200 -59977 69494 -59429
rect 67200 -59984 67809 -59977
rect 68429 -59984 69494 -59977
rect 67200 -60178 67722 -59984
rect 68647 -60389 69494 -59984
rect 72685 -59929 74979 -59381
rect 72685 -59936 73294 -59929
rect 73914 -59936 74979 -59929
rect 72685 -60130 73207 -59936
rect 74132 -60341 74979 -59936
rect 76353 -59412 78679 -59218
rect 82049 -59343 84375 -59149
rect 85743 -58993 87238 -58814
rect 85743 -59000 87325 -58993
rect 85743 -59180 88043 -59000
rect 76353 -59960 78647 -59412
rect 76353 -59967 76962 -59960
rect 77582 -59967 78647 -59960
rect 76353 -60161 76875 -59967
rect 77800 -60372 78647 -59967
rect 82049 -59891 84343 -59343
rect 82049 -59898 82658 -59891
rect 83278 -59898 84343 -59891
rect 82049 -60092 82571 -59898
rect 83496 -60303 84343 -59898
rect 85717 -59374 88043 -59180
rect 85717 -59922 88011 -59374
rect 85717 -59929 86326 -59922
rect 86946 -59929 88011 -59922
rect 85717 -60123 86239 -59929
rect 87164 -60334 88011 -59929
rect 14328 -61618 15169 -61612
rect -6092 -61854 -4175 -61781
rect -3592 -61854 -1675 -61781
rect -1092 -61854 825 -61781
rect 1408 -61854 3325 -61781
rect 3908 -61854 5825 -61781
rect 6908 -61854 8825 -61781
rect -21600 -62325 -20144 -61867
rect -6093 -62256 -4175 -61854
rect -3593 -62256 -1675 -61854
rect -1093 -62256 825 -61854
rect 1407 -62256 3325 -61854
rect 3907 -62256 5825 -61854
rect 6907 -62256 8825 -61854
rect 12808 -62071 17870 -61618
rect 15134 -62072 17870 -62071
rect -21569 -62326 -20144 -62325
<< pwell >>
rect -12868 119107 -12734 119906
rect -12677 119622 -12325 119830
rect -12677 119184 -12325 119490
rect -10724 119345 -10572 119749
rect -10570 119273 -10439 119854
rect -12017 118274 -11886 118855
rect -11884 118346 -11732 118750
rect -10417 118638 -10065 119140
rect -10061 118630 -9948 119131
rect -12508 117631 -12395 118132
rect -12391 117639 -12039 118141
rect -10495 117763 -10243 118167
rect -10241 117691 -10110 118272
rect -9398 117352 -9185 118877
rect -9135 118665 -8783 118873
rect -9135 118339 -8583 118645
rect -9135 118111 -8583 118319
rect -9135 117888 -8583 118096
rect -9135 117418 -8783 117626
rect -12837 115439 -12703 116238
rect -12646 115954 -12294 116162
rect -12646 115516 -12294 115822
rect -10693 115677 -10541 116081
rect -10539 115605 -10408 116186
rect -11986 114606 -11855 115187
rect -11853 114678 -11701 115082
rect -10386 114970 -10034 115472
rect -10030 114962 -9917 115463
rect -9384 115447 -9250 116246
rect -9193 115962 -8841 116170
rect -9193 115524 -8841 115830
rect -7240 115685 -7088 116089
rect -7086 115613 -6955 116194
rect -8533 114614 -8402 115195
rect -8400 114686 -8248 115090
rect -6933 114978 -6581 115480
rect -6577 114970 -6464 115471
rect -12477 113963 -12364 114464
rect -12360 113971 -12008 114473
rect -10464 114095 -10212 114499
rect -10210 114023 -10079 114604
rect -9024 113971 -8911 114472
rect -8907 113979 -8555 114481
rect -7011 114103 -6759 114507
rect -6757 114031 -6626 114612
rect -12906 109743 -12772 110542
rect -12715 110258 -12363 110466
rect -12715 109820 -12363 110126
rect -10762 109981 -10610 110385
rect -10608 109909 -10477 110490
rect -12055 108910 -11924 109491
rect -11922 108982 -11770 109386
rect -10455 109274 -10103 109776
rect -10099 109266 -9986 109767
rect -12546 108267 -12433 108768
rect -12429 108275 -12077 108777
rect -10533 108399 -10281 108803
rect -10279 108327 -10148 108908
rect -9436 107988 -9223 109513
rect -9173 109301 -8821 109509
rect -9173 108975 -8621 109281
rect -9173 108747 -8621 108955
rect -9173 108524 -8621 108732
rect -9173 108054 -8821 108262
rect -12875 106075 -12741 106874
rect -12684 106590 -12332 106798
rect -12684 106152 -12332 106458
rect -10731 106313 -10579 106717
rect -10577 106241 -10446 106822
rect -12024 105242 -11893 105823
rect -11891 105314 -11739 105718
rect -10424 105606 -10072 106108
rect -10068 105598 -9955 106099
rect -9422 106083 -9288 106882
rect -9231 106598 -8879 106806
rect -9231 106160 -8879 106466
rect -7278 106321 -7126 106725
rect -7124 106249 -6993 106830
rect -8571 105250 -8440 105831
rect -8438 105322 -8286 105726
rect -6971 105614 -6619 106116
rect -6615 105606 -6502 106107
rect -12515 104599 -12402 105100
rect -12398 104607 -12046 105109
rect -10502 104731 -10250 105135
rect -10248 104659 -10117 105240
rect -9062 104607 -8949 105108
rect -8945 104615 -8593 105117
rect -7049 104739 -6797 105143
rect -6795 104667 -6664 105248
rect -12923 100590 -12789 101389
rect -12732 101105 -12380 101313
rect -12732 100667 -12380 100973
rect -10779 100828 -10627 101232
rect -10625 100756 -10494 101337
rect -12072 99757 -11941 100338
rect -11939 99829 -11787 100233
rect -10472 100121 -10120 100623
rect -10116 100113 -10003 100614
rect -12563 99114 -12450 99615
rect -12446 99122 -12094 99624
rect -10550 99246 -10298 99650
rect -10296 99174 -10165 99755
rect -9453 98835 -9240 100360
rect -9190 100148 -8838 100356
rect -9190 99822 -8638 100128
rect -9190 99594 -8638 99802
rect -9190 99371 -8638 99579
rect -9190 98901 -8838 99109
rect -12892 96922 -12758 97721
rect -12701 97437 -12349 97645
rect -12701 96999 -12349 97305
rect -10748 97160 -10596 97564
rect -10594 97088 -10463 97669
rect -12041 96089 -11910 96670
rect -11908 96161 -11756 96565
rect -10441 96453 -10089 96955
rect -10085 96445 -9972 96946
rect -9439 96930 -9305 97729
rect -9248 97445 -8896 97653
rect -9248 97007 -8896 97313
rect -7295 97168 -7143 97572
rect -7141 97096 -7010 97677
rect -8588 96097 -8457 96678
rect -8455 96169 -8303 96573
rect -6988 96461 -6636 96963
rect -6632 96453 -6519 96954
rect -12532 95446 -12419 95947
rect -12415 95454 -12063 95956
rect -10519 95578 -10267 95982
rect -10265 95506 -10134 96087
rect -9079 95454 -8966 95955
rect -8962 95462 -8610 95964
rect -7066 95586 -6814 95990
rect -6812 95514 -6681 96095
rect -12989 91836 -12855 92635
rect -12798 92351 -12446 92559
rect -12798 91913 -12446 92219
rect -10845 92074 -10693 92478
rect -10691 92002 -10560 92583
rect -12138 91003 -12007 91584
rect -12005 91075 -11853 91479
rect -10538 91367 -10186 91869
rect -10182 91359 -10069 91860
rect -12629 90360 -12516 90861
rect -12512 90368 -12160 90870
rect -10616 90492 -10364 90896
rect -10362 90420 -10231 91001
rect -9519 90081 -9306 91606
rect -9256 91394 -8904 91602
rect -9256 91068 -8704 91374
rect -9256 90840 -8704 91048
rect -9256 90617 -8704 90825
rect -9256 90147 -8904 90355
rect -12958 88168 -12824 88967
rect -12767 88683 -12415 88891
rect -12767 88245 -12415 88551
rect -10814 88406 -10662 88810
rect -10660 88334 -10529 88915
rect -12107 87335 -11976 87916
rect -11974 87407 -11822 87811
rect -10507 87699 -10155 88201
rect -10151 87691 -10038 88192
rect -9505 88176 -9371 88975
rect -9314 88691 -8962 88899
rect -9314 88253 -8962 88559
rect -7361 88414 -7209 88818
rect -7207 88342 -7076 88923
rect -8654 87343 -8523 87924
rect -8521 87415 -8369 87819
rect -7054 87707 -6702 88209
rect -6698 87699 -6585 88200
rect -12598 86692 -12485 87193
rect -12481 86700 -12129 87202
rect -10585 86824 -10333 87228
rect -10331 86752 -10200 87333
rect -9145 86700 -9032 87201
rect -9028 86708 -8676 87210
rect -7132 86832 -6880 87236
rect -6878 86760 -6747 87341
rect -13023 82638 -12889 83437
rect -12832 83153 -12480 83361
rect -12832 82715 -12480 83021
rect -10879 82876 -10727 83280
rect -10725 82804 -10594 83385
rect -12172 81805 -12041 82386
rect -12039 81877 -11887 82281
rect -10572 82169 -10220 82671
rect -10216 82161 -10103 82662
rect -12663 81162 -12550 81663
rect -12546 81170 -12194 81672
rect -10650 81294 -10398 81698
rect -10396 81222 -10265 81803
rect -9553 80883 -9340 82408
rect -9290 82196 -8938 82404
rect -9290 81870 -8738 82176
rect -9290 81642 -8738 81850
rect -9290 81419 -8738 81627
rect -9290 80949 -8938 81157
rect -12992 78970 -12858 79769
rect -12801 79485 -12449 79693
rect -12801 79047 -12449 79353
rect -10848 79208 -10696 79612
rect -10694 79136 -10563 79717
rect -12141 78137 -12010 78718
rect -12008 78209 -11856 78613
rect -10541 78501 -10189 79003
rect -10185 78493 -10072 78994
rect -9539 78978 -9405 79777
rect -9348 79493 -8996 79701
rect -9348 79055 -8996 79361
rect -7395 79216 -7243 79620
rect -7241 79144 -7110 79725
rect -8688 78145 -8557 78726
rect -8555 78217 -8403 78621
rect -7088 78509 -6736 79011
rect -6732 78501 -6619 79002
rect -12632 77494 -12519 77995
rect -12515 77502 -12163 78004
rect -10619 77626 -10367 78030
rect -10365 77554 -10234 78135
rect -9179 77502 -9066 78003
rect -9062 77510 -8710 78012
rect -7166 77634 -6914 78038
rect -6912 77562 -6781 78143
rect -12984 73775 -12850 74574
rect -12793 74290 -12441 74498
rect -12793 73852 -12441 74158
rect -10840 74013 -10688 74417
rect -10686 73941 -10555 74522
rect -12133 72942 -12002 73523
rect -12000 73014 -11848 73418
rect -10533 73306 -10181 73808
rect -10177 73298 -10064 73799
rect -12624 72299 -12511 72800
rect -12507 72307 -12155 72809
rect -10611 72431 -10359 72835
rect -10357 72359 -10226 72940
rect -9514 72020 -9301 73545
rect -9251 73333 -8899 73541
rect -9251 73007 -8699 73313
rect -9251 72779 -8699 72987
rect -9251 72556 -8699 72764
rect -9251 72086 -8899 72294
rect -12953 70107 -12819 70906
rect -12762 70622 -12410 70830
rect -12762 70184 -12410 70490
rect -10809 70345 -10657 70749
rect -10655 70273 -10524 70854
rect -12102 69274 -11971 69855
rect -11969 69346 -11817 69750
rect -10502 69638 -10150 70140
rect -10146 69630 -10033 70131
rect -9500 70115 -9366 70914
rect -9309 70630 -8957 70838
rect -9309 70192 -8957 70498
rect -7356 70353 -7204 70757
rect -7202 70281 -7071 70862
rect -8649 69282 -8518 69863
rect -8516 69354 -8364 69758
rect -7049 69646 -6697 70148
rect -6693 69638 -6580 70139
rect -12593 68631 -12480 69132
rect -12476 68639 -12124 69141
rect -10580 68763 -10328 69167
rect -10326 68691 -10195 69272
rect -9140 68639 -9027 69140
rect -9023 68647 -8671 69149
rect -7127 68771 -6875 69175
rect -6873 68699 -6742 69280
rect -12973 65335 -12839 66134
rect -12782 65850 -12430 66058
rect -12782 65412 -12430 65718
rect -10829 65573 -10677 65977
rect -10675 65501 -10544 66082
rect -12122 64502 -11991 65083
rect -11989 64574 -11837 64978
rect -10522 64866 -10170 65368
rect -10166 64858 -10053 65359
rect -12613 63859 -12500 64360
rect -12496 63867 -12144 64369
rect -10600 63991 -10348 64395
rect -10346 63919 -10215 64500
rect -9503 63580 -9290 65105
rect -9240 64893 -8888 65101
rect -9240 64567 -8688 64873
rect -9240 64339 -8688 64547
rect -9240 64116 -8688 64324
rect -9240 63646 -8888 63854
rect -12942 61667 -12808 62466
rect -12751 62182 -12399 62390
rect -12751 61744 -12399 62050
rect -10798 61905 -10646 62309
rect -10644 61833 -10513 62414
rect -12091 60834 -11960 61415
rect -11958 60906 -11806 61310
rect -10491 61198 -10139 61700
rect -10135 61190 -10022 61691
rect -9489 61675 -9355 62474
rect -9298 62190 -8946 62398
rect -9298 61752 -8946 62058
rect -7345 61913 -7193 62317
rect -7191 61841 -7060 62422
rect -8638 60842 -8507 61423
rect -8505 60914 -8353 61318
rect -7038 61206 -6686 61708
rect -6682 61198 -6569 61699
rect -12582 60191 -12469 60692
rect -12465 60199 -12113 60701
rect -10569 60323 -10317 60727
rect -10315 60251 -10184 60832
rect -9129 60199 -9016 60700
rect -9012 60207 -8660 60709
rect -7116 60331 -6864 60735
rect -6862 60259 -6731 60840
rect -10414 57650 -9662 57858
rect -10414 57250 -9662 57458
rect -10414 56650 -9662 56858
rect -10414 56250 -9662 56458
rect -10414 55650 -9662 55858
rect -10414 55250 -9662 55458
rect -9597 55165 -9448 57944
rect -8737 57300 -8585 57900
rect -8582 57303 -8462 57889
rect -8202 57311 -8082 57897
rect -8079 57300 -7927 57900
rect -8687 56266 -8535 57062
rect -8202 56474 -8082 57060
rect -8079 56463 -7927 57063
rect -8737 55557 -8585 56157
rect -8582 55560 -8462 56146
rect -8129 55558 -7977 56354
rect -10990 54370 -10838 54970
rect -10835 54373 -10715 54959
rect -10712 54399 -10579 54930
rect -10523 54630 -10271 54838
rect -10523 54420 -10271 54628
rect -8737 54600 -8585 55200
rect -8582 54603 -8462 55189
rect -8202 54611 -8082 55197
rect -8079 54600 -7927 55200
rect -10669 53641 -10417 53849
rect -10769 53130 -10417 53436
rect -10769 52821 -10417 53127
rect -10770 52511 -10418 52817
rect -10277 52523 -10160 53849
rect -8687 53566 -8535 54362
rect -8202 53774 -8082 54360
rect -8079 53763 -7927 54363
rect -8737 52857 -8585 53457
rect -8582 52860 -8462 53446
rect -8129 52858 -7977 53654
rect -10651 51693 -10399 51999
rect -10344 51572 -10203 52221
rect -8737 51975 -8585 52575
rect -8582 51978 -8462 52564
rect -10651 50747 -10399 51053
rect -10344 50626 -10203 51275
rect -8033 50752 -7781 51156
rect -7720 50655 -7562 51564
rect -13293 49172 -13141 49772
rect -13138 49183 -13018 49769
rect -12758 49175 -12638 49761
rect -12635 49172 -12483 49772
rect -13293 48335 -13141 48935
rect -13138 48346 -13018 48932
rect -13243 47430 -13091 48226
rect -12685 48138 -12533 48934
rect -12758 47432 -12638 48018
rect -12635 47429 -12483 48029
rect -13293 46472 -13141 47072
rect -13138 46483 -13018 47069
rect -12758 46475 -12638 47061
rect -12635 46472 -12483 47072
rect -13293 45635 -13141 46235
rect -13138 45646 -13018 46232
rect -13243 44730 -13091 45526
rect -12685 45438 -12533 46234
rect -12758 44732 -12638 45318
rect -12635 44729 -12483 45329
rect -12758 43850 -12638 44436
rect -12635 43847 -12483 44447
rect -13230 40519 -12978 40727
rect -13230 40210 -12978 40418
rect -13230 39900 -12978 40108
rect -12949 40039 -12801 40723
rect -13230 39606 -12978 39814
rect -13230 39244 -12978 39452
rect -13230 38830 -12978 39038
rect -13230 37519 -12978 37727
rect -13230 37210 -12978 37418
rect -13230 36900 -12978 37108
rect -12949 37039 -12801 37723
rect -10979 40529 -10727 40737
rect -10979 40220 -10727 40428
rect -10979 39910 -10727 40118
rect -10698 40049 -10550 40733
rect -8332 40049 -8184 40733
rect -8155 40529 -7903 40737
rect -8155 40220 -7903 40428
rect -8155 39910 -7903 40118
rect -10979 39616 -10727 39824
rect -8155 39616 -7903 39824
rect -10979 39254 -10727 39462
rect -8155 39254 -7903 39462
rect -10979 38840 -10727 39048
rect -8155 38840 -7903 39048
rect -10989 38259 -10637 38565
rect -10988 37949 -10636 38255
rect -10988 37640 -10636 37946
rect -10888 37227 -10636 37435
rect -10496 37227 -10379 38553
rect -8503 37227 -8386 38553
rect -8245 38259 -7893 38565
rect -8246 37949 -7894 38255
rect -8246 37640 -7894 37946
rect -8246 37227 -7994 37435
rect -6081 40039 -5933 40723
rect -5904 40519 -5652 40727
rect -5904 40210 -5652 40418
rect -5904 39900 -5652 40108
rect -5904 39606 -5652 39814
rect -5904 39244 -5652 39452
rect -5904 38830 -5652 39038
rect -6081 37039 -5933 37723
rect -5904 37519 -5652 37727
rect -5904 37210 -5652 37418
rect -5904 36900 -5652 37108
rect -13230 36606 -12978 36814
rect -13230 36244 -12978 36452
rect -11034 36310 -10682 36812
rect -10678 36319 -10565 36820
rect -8317 36319 -8204 36820
rect -8200 36310 -7848 36812
rect -5904 36606 -5652 36814
rect -5904 36244 -5652 36452
rect -13230 35830 -12978 36038
rect -13230 35019 -12978 35227
rect -13230 34710 -12978 34918
rect -13230 34400 -12978 34608
rect -12949 34539 -12801 35223
rect -11341 35701 -11189 36105
rect -11187 35596 -11056 36177
rect -7826 35596 -7695 36177
rect -7693 35701 -7541 36105
rect -5904 35830 -5652 36038
rect -11036 34705 -10684 35207
rect -10680 34714 -10567 35215
rect -8315 34714 -8202 35215
rect -8198 34705 -7846 35207
rect -13230 34106 -12978 34314
rect -13230 33744 -12978 33952
rect -11343 34096 -11191 34500
rect -11189 33991 -11058 34572
rect -7824 33991 -7693 34572
rect -7691 34096 -7539 34500
rect -6081 34539 -5933 35223
rect -5904 35019 -5652 35227
rect -5904 34710 -5652 34918
rect -5904 34400 -5652 34608
rect -5904 34106 -5652 34314
rect -5904 33744 -5652 33952
rect -13230 33330 -12978 33538
rect -13230 32519 -12978 32727
rect -13230 32210 -12978 32418
rect -13230 31900 -12978 32108
rect -12949 32039 -12801 32723
rect -13230 31606 -12978 31814
rect -10980 33297 -10628 33603
rect -10979 32987 -10627 33293
rect -10979 32678 -10627 32984
rect -10879 32265 -10627 32473
rect -10487 32265 -10370 33591
rect -8512 32265 -8395 33591
rect -8254 33297 -7902 33603
rect -8255 32987 -7903 33293
rect -8255 32678 -7903 32984
rect -8255 32265 -8003 32473
rect -13230 31244 -12978 31452
rect -13230 30830 -12978 31038
rect -11224 31335 -11072 31935
rect -11069 31346 -10949 31932
rect -7933 31346 -7813 31932
rect -7810 31335 -7658 31935
rect -5904 33330 -5652 33538
rect -6081 32039 -5933 32723
rect -5904 32519 -5652 32727
rect -5904 32210 -5652 32418
rect -5904 31900 -5652 32108
rect -5904 31606 -5652 31814
rect -13230 30019 -12978 30227
rect -13230 29710 -12978 29918
rect -13230 29400 -12978 29608
rect -12949 29539 -12801 30223
rect -13230 29106 -12978 29314
rect -13230 28744 -12978 28952
rect -13230 28330 -12978 28538
rect -13230 27519 -12978 27727
rect -13230 27210 -12978 27418
rect -13230 26900 -12978 27108
rect -12949 27039 -12801 27723
rect -13230 26606 -12978 26814
rect -13230 26244 -12978 26452
rect -13230 25830 -12978 26038
rect -11224 30453 -11072 31053
rect -11069 30464 -10949 31050
rect -11174 29548 -11022 30344
rect -10616 30256 -10464 31052
rect -10689 29550 -10569 30136
rect -10566 29547 -10414 30147
rect -11224 28710 -11072 29310
rect -11069 28721 -10949 29307
rect -10689 28713 -10569 29299
rect -10566 28710 -10414 29310
rect -8418 30256 -8266 31052
rect -7933 30464 -7813 31050
rect -7810 30453 -7658 31053
rect -5904 31244 -5652 31452
rect -8468 29547 -8316 30147
rect -8313 29550 -8193 30136
rect -7860 29548 -7708 30344
rect -11224 27753 -11072 28353
rect -11069 27764 -10949 28350
rect -11174 26848 -11022 27644
rect -10616 27556 -10464 28352
rect -10689 26850 -10569 27436
rect -10566 26847 -10414 27447
rect -11224 26010 -11072 26610
rect -11069 26021 -10949 26607
rect -10689 26013 -10569 26599
rect -10566 26010 -10414 26610
rect -8468 28710 -8316 29310
rect -8313 28713 -8193 29299
rect -7933 28721 -7813 29307
rect -7810 28710 -7658 29310
rect -8418 27556 -8266 28352
rect -7933 27764 -7813 28350
rect -7810 27753 -7658 28353
rect -8468 26847 -8316 27447
rect -8313 26850 -8193 27436
rect -7860 26848 -7708 27644
rect -8468 26010 -8316 26610
rect -8313 26013 -8193 26599
rect -7933 26021 -7813 26607
rect -7810 26010 -7658 26610
rect -5904 30830 -5652 31038
rect -6081 29539 -5933 30223
rect -5904 30019 -5652 30227
rect -5904 29710 -5652 29918
rect -5904 29400 -5652 29608
rect -5904 29106 -5652 29314
rect -5904 28744 -5652 28952
rect -5904 28330 -5652 28538
rect -6081 27039 -5933 27723
rect -5904 27519 -5652 27727
rect -5904 27210 -5652 27418
rect -5904 26900 -5652 27108
rect -6247 26267 -6095 26867
rect -6092 26270 -5972 26856
rect -5904 26606 -5652 26814
rect -5904 26244 -5652 26452
rect -5904 25830 -5652 26038
rect -11239 24434 -11105 25233
rect -11048 24850 -10696 25156
rect -11048 24510 -10696 24718
rect -6305 24407 -6171 25206
rect -6114 24823 -5762 25129
rect -6114 24483 -5762 24691
rect -10957 23461 -10805 24061
rect -10802 23472 -10682 24058
rect -10957 22579 -10805 23179
rect -10802 22590 -10682 23176
rect -10907 21674 -10755 22470
rect -10349 22382 -10197 23178
rect -10422 21676 -10302 22262
rect -10299 21673 -10147 22273
rect -10957 20836 -10805 21436
rect -10802 20847 -10682 21433
rect -10422 20839 -10302 21425
rect -10299 20836 -10147 21436
rect -6030 23461 -5878 24061
rect -5875 23472 -5755 24058
rect -10957 19879 -10805 20479
rect -10802 19890 -10682 20476
rect -10907 18974 -10755 19770
rect -10349 19682 -10197 20478
rect -10422 18976 -10302 19562
rect -10299 18973 -10147 19573
rect -10957 18136 -10805 18736
rect -10802 18147 -10682 18733
rect -10422 18139 -10302 18725
rect -10299 18136 -10147 18736
rect -9102 20795 -8971 21376
rect -8969 20867 -8817 21271
rect -7216 21144 -6864 21352
rect -7216 20706 -6864 21012
rect -9593 20152 -9480 20653
rect -9476 20160 -9124 20662
rect -6807 20629 -6673 21428
rect -6030 22579 -5878 23179
rect -5875 22590 -5755 23176
rect -5980 21674 -5828 22470
rect -5422 22382 -5270 23178
rect -5495 21676 -5375 22262
rect -5372 21673 -5220 22273
rect -9431 19213 -9300 19794
rect -7809 19868 -7657 20272
rect -7655 19796 -7524 20377
rect -9298 19285 -9046 19689
rect -7502 19161 -7150 19663
rect -7146 19153 -7033 19654
rect -6030 20836 -5878 21436
rect -5875 20847 -5755 21433
rect -5495 20839 -5375 21425
rect -5372 20836 -5220 21436
rect -6030 19879 -5878 20479
rect -5875 19890 -5755 20476
rect -5980 18974 -5828 19770
rect -5422 19682 -5270 20478
rect -5495 18976 -5375 19562
rect -5372 18973 -5220 19573
rect -6030 18136 -5878 18736
rect -5875 18147 -5755 18733
rect -5495 18139 -5375 18725
rect -5372 18136 -5220 18736
rect -13126 15806 -12995 16387
rect -12993 15878 -12841 16282
rect -11240 16155 -10888 16363
rect -11240 15717 -10888 16023
rect -13617 15163 -13504 15664
rect -13500 15171 -13148 15673
rect -10831 15640 -10697 16439
rect -8126 15806 -7995 16387
rect -7993 15878 -7841 16282
rect -6240 16155 -5888 16363
rect -6240 15717 -5888 16023
rect -13455 14224 -13324 14805
rect -11833 14879 -11681 15283
rect -11679 14807 -11548 15388
rect -8617 15163 -8504 15664
rect -8500 15171 -8148 15673
rect -5831 15640 -5697 16439
rect -13322 14296 -13070 14700
rect -11526 14172 -11174 14674
rect -11170 14164 -11057 14665
rect -8455 14224 -8324 14805
rect -6833 14879 -6681 15283
rect -6679 14807 -6548 15388
rect -8322 14296 -8070 14700
rect -6526 14172 -6174 14674
rect -6170 14164 -6057 14665
rect -11922 12747 -11781 13396
rect -11726 12868 -11474 13174
rect -11921 11842 -11780 12491
rect -11725 11963 -11473 12269
rect -8780 12379 -8663 13705
rect -8523 13497 -8271 13705
rect -8523 12986 -8171 13292
rect -8523 12677 -8171 12983
rect -8522 12367 -8170 12673
rect -6264 13171 -6133 13752
rect -6131 13243 -5979 13647
rect -6755 12528 -6642 13029
rect -6638 12536 -6286 13038
rect -13315 11452 -12963 11758
rect -13314 11142 -12962 11448
rect -13314 10833 -12962 11139
rect -13214 10420 -12962 10628
rect -12822 10420 -12705 11746
rect -12287 10660 -12129 11569
rect -12068 10757 -11816 11161
rect -8173 11229 -8042 11810
rect -8040 11301 -7888 11705
rect -8664 10586 -8551 11087
rect -8547 10594 -8195 11096
rect -6844 10549 -6727 11875
rect -6587 11667 -6335 11875
rect -6587 11156 -6235 11462
rect -6587 10847 -6235 11153
rect -6586 10537 -6234 10843
rect 15992 9068 16244 10210
rect 16392 9068 16644 10210
rect 16792 9068 17044 10210
rect 16007 8816 16143 9044
rect 17109 8966 17341 10210
rect 69208 9612 92372 10082
rect 8142 5617 11684 6469
rect 8142 4617 12542 5469
rect 8082 4332 12576 4530
rect 25581 3506 47660 3753
rect 19756 2872 20356 3024
rect 20606 2872 21206 3024
rect 19759 2749 20345 2869
rect 20609 2749 21195 2869
rect 21252 2806 22146 3058
rect 20609 2612 21195 2732
rect 2794 2393 3125 2534
rect 539 2260 3125 2393
rect 539 2246 1153 2260
rect 1535 2248 3125 2260
rect 1535 2246 2991 2248
rect 565 2146 818 2246
rect 587 1975 785 2111
rect 833 1964 1473 2136
rect 1477 1969 1763 2141
rect 1791 1976 2373 2148
rect 2429 2146 2991 2246
rect 2462 1975 2660 2111
rect 2771 1975 2969 2111
rect -4222 1453 -4082 1548
rect -3622 1531 -3022 1683
rect -2772 1531 -2172 1683
rect -3619 1408 -3033 1528
rect -2769 1408 -2183 1528
rect -2126 1465 -1232 1717
rect -2769 1271 -2183 1391
rect -13349 741 -6159 1193
rect -2772 1116 -2172 1268
rect -2126 1082 -1232 1334
rect -13376 531 -6123 709
rect 4477 1707 5077 1859
rect 5327 1707 5927 1859
rect 4480 1584 5066 1704
rect 5330 1584 5916 1704
rect 5973 1641 6867 1893
rect 20606 2457 21206 2609
rect 21252 2423 22146 2675
rect 5330 1447 5916 1567
rect 5327 1292 5927 1444
rect 5973 1258 6867 1510
rect 587 751 785 887
rect 833 726 1473 898
rect 1477 721 1763 893
rect 565 616 818 716
rect 1791 714 2373 886
rect 2462 751 2660 887
rect 2771 751 2969 887
rect 2429 616 2991 716
rect 7872 1023 15062 1475
rect 7836 813 15089 991
rect 539 602 1153 616
rect 1535 602 2991 616
rect 539 469 2991 602
rect -5090 -841 -4490 -689
rect -4240 -841 -3640 -689
rect -5087 -964 -4501 -844
rect -4237 -964 -3651 -844
rect -3594 -907 -2700 -655
rect -4237 -1101 -3651 -981
rect 4492 -983 5092 -831
rect 5342 -983 5942 -831
rect -4240 -1256 -3640 -1104
rect -3594 -1290 -2700 -1038
rect 4495 -1106 5081 -986
rect 5345 -1106 5931 -986
rect 5988 -1049 6882 -797
rect 19928 -478 20528 -326
rect 20778 -478 21378 -326
rect 19931 -601 20517 -481
rect 20781 -601 21367 -481
rect 21424 -544 22318 -292
rect 20781 -738 21367 -618
rect 20778 -893 21378 -741
rect 21424 -927 22318 -675
rect 5345 -1243 5931 -1123
rect 5342 -1398 5942 -1246
rect 5988 -1432 6882 -1180
rect 7831 -1733 15021 -1281
rect 25581 -1203 25828 3506
rect 30279 2628 31667 2805
rect 35014 2650 36402 2827
rect 36735 2607 38123 2784
rect 30292 2070 31666 2522
rect 35027 2092 36401 2544
rect 36748 2049 38122 2501
rect 39148 2429 39748 2581
rect 40030 2429 40630 2581
rect 39151 2306 39737 2426
rect 40033 2306 40619 2426
rect 40739 2379 41535 2531
rect 41773 2429 42373 2581
rect 42730 2429 43330 2581
rect 41776 2306 42362 2426
rect 42733 2306 43319 2426
rect 43439 2379 44235 2531
rect 44473 2429 45073 2581
rect 44476 2306 45062 2426
rect 27778 915 28046 1167
rect 28058 913 28800 1165
rect 28808 913 29076 1165
rect 29084 911 29352 1163
rect 27778 463 28046 715
rect 28058 463 28800 715
rect 28808 463 29076 715
rect 29083 463 29351 715
rect 32633 908 32901 1160
rect 32913 906 33655 1158
rect 33663 906 33931 1158
rect 33939 904 34207 1156
rect 32633 456 32901 708
rect 32913 456 33655 708
rect 33663 456 33931 708
rect 33938 456 34206 708
rect 40031 1821 40827 1973
rect 40947 1926 41533 2046
rect 41784 1926 42370 2046
rect 40936 1771 41536 1923
rect 41773 1771 42373 1923
rect 42731 1821 43527 1973
rect 43647 1926 44233 2046
rect 44484 1926 45070 2046
rect 45544 2016 46130 2136
rect 43636 1771 44236 1923
rect 44473 1771 45073 1923
rect 45541 1861 46141 2013
rect 27499 -49 27767 203
rect 27771 -47 29461 205
rect 29468 -47 29736 205
rect 27738 -284 29489 -141
rect 30292 -242 31666 210
rect 32354 -56 32622 196
rect 32626 -54 34316 198
rect 34323 -54 34591 198
rect 32593 -291 34344 -148
rect 35027 -219 36401 233
rect 36748 -176 38122 276
rect 30279 -525 31667 -348
rect 35014 -502 36402 -325
rect 36735 -459 38123 -282
rect 47413 -1203 47660 3506
rect 51150 1800 58340 2252
rect 51114 1590 58367 1768
rect 50947 -1111 58137 -659
rect 25581 -1450 47660 -1203
rect 50911 -1321 58164 -1143
rect 7795 -1943 15048 -1765
rect 62355 -3344 62955 -3192
rect 63205 -3344 63805 -3192
rect 62358 -3467 62944 -3347
rect 63208 -3467 63794 -3347
rect 63851 -3410 64745 -3158
rect 63208 -3604 63794 -3484
rect 50947 -4158 58137 -3706
rect 63205 -3759 63805 -3607
rect 63851 -3793 64745 -3541
rect 50911 -4368 58164 -4190
rect -15016 -15270 -7763 -15092
rect -14989 -15754 -7799 -15302
rect -15177 -18903 -14577 -18751
rect -14340 -18903 -13740 -18751
rect -15174 -19026 -14588 -18906
rect -14337 -19026 -13751 -18906
rect -13631 -18953 -12835 -18801
rect -12477 -18903 -11877 -18751
rect -11640 -18903 -11040 -18751
rect -12474 -19026 -11888 -18906
rect -11637 -19026 -11051 -18906
rect -10931 -18953 -10135 -18801
rect -17673 -19362 -16874 -19228
rect -15166 -19406 -14580 -19286
rect -20070 -19662 -19666 -19510
rect -22776 -20117 -22470 -19765
rect -22466 -20118 -22160 -19766
rect -22157 -20118 -21851 -19766
rect -20142 -19795 -19561 -19664
rect -19149 -19701 -18648 -19588
rect -21646 -20118 -21438 -19866
rect -20777 -20169 -20275 -19817
rect -19141 -20057 -18639 -19705
rect -17596 -19771 -17290 -19419
rect -17158 -19771 -16950 -19419
rect -15177 -19561 -14577 -19409
rect -14339 -19511 -13543 -19359
rect -13423 -19406 -12837 -19286
rect -12466 -19406 -11880 -19286
rect -13434 -19561 -12834 -19409
rect -12477 -19561 -11877 -19409
rect -11639 -19511 -10843 -19359
rect -10723 -19406 -10137 -19286
rect -9841 -19406 -9255 -19286
rect -10734 -19561 -10134 -19409
rect -9852 -19561 -9252 -19409
rect -8830 -19645 -8622 -19293
rect -8490 -19645 -8184 -19293
rect -7483 -19435 -7275 -19183
rect -7069 -19435 -6861 -19183
rect -6707 -19435 -6499 -19183
rect -6413 -19435 -6205 -19183
rect -6103 -19435 -5895 -19183
rect -5794 -19435 -5586 -19183
rect -4983 -19435 -4775 -19183
rect -4569 -19435 -4361 -19183
rect -4207 -19435 -3999 -19183
rect -3913 -19435 -3705 -19183
rect -3603 -19435 -3395 -19183
rect -3294 -19435 -3086 -19183
rect -2483 -19435 -2275 -19183
rect -2069 -19435 -1861 -19183
rect -1707 -19435 -1499 -19183
rect -1413 -19435 -1205 -19183
rect -1103 -19435 -895 -19183
rect -794 -19435 -586 -19183
rect 17 -19435 225 -19183
rect 431 -19435 639 -19183
rect 793 -19435 1001 -19183
rect 1087 -19435 1295 -19183
rect 1397 -19435 1605 -19183
rect 1706 -19435 1914 -19183
rect 2517 -19435 2725 -19183
rect 2931 -19435 3139 -19183
rect 3293 -19435 3501 -19183
rect 3587 -19435 3795 -19183
rect 3897 -19435 4105 -19183
rect 4206 -19435 4414 -19183
rect 5517 -19435 5725 -19183
rect 5931 -19435 6139 -19183
rect 6293 -19435 6501 -19183
rect 6587 -19435 6795 -19183
rect 6897 -19435 7105 -19183
rect 7206 -19435 7414 -19183
rect -7043 -19623 -6457 -19503
rect -6274 -19612 -5590 -19464
rect -3774 -19612 -3090 -19464
rect -1274 -19612 -590 -19464
rect 1226 -19612 1910 -19464
rect 3726 -19612 4410 -19464
rect 6726 -19612 7410 -19464
rect -22764 -20375 -21438 -20258
rect -20785 -20286 -20284 -20173
rect -18506 -20210 -17925 -20079
rect -18434 -20364 -18030 -20212
rect -8906 -19836 -8107 -19702
rect -7046 -19778 -6446 -19626
rect -12684 -20338 -11885 -20204
rect 27885 -20213 28386 -20100
rect 26946 -20393 27527 -20262
rect -14160 -20677 -13659 -20564
rect -14152 -21033 -13650 -20681
rect -12607 -20747 -12301 -20395
rect -12169 -20747 -11961 -20395
rect -22012 -21571 -21608 -21419
rect -17435 -21524 -17031 -21372
rect -13517 -21186 -12936 -21055
rect -13445 -21340 -13041 -21188
rect 27018 -20647 27422 -20395
rect 27893 -20569 28395 -20217
rect 36325 -20224 36826 -20111
rect 35386 -20404 35967 -20273
rect 28528 -20722 29109 -20591
rect 35458 -20658 35862 -20406
rect 36333 -20580 36835 -20228
rect 45188 -20263 45689 -20150
rect 54386 -20229 54887 -20116
rect 63140 -20163 63641 -20050
rect 72293 -20146 72794 -20033
rect 81657 -20108 82158 -19995
rect 44249 -20443 44830 -20312
rect 28600 -20876 29004 -20724
rect 36968 -20733 37549 -20602
rect 44321 -20697 44725 -20445
rect 45196 -20619 45698 -20267
rect 53447 -20409 54028 -20278
rect -7303 -21341 -6703 -21189
rect -22084 -21704 -21503 -21573
rect -22719 -22078 -22217 -21726
rect -20946 -22053 -20640 -21701
rect -20636 -22054 -20330 -21702
rect -20327 -22054 -20021 -21702
rect -19816 -22054 -19608 -21802
rect -19017 -21853 -18613 -21601
rect -17507 -21657 -16926 -21526
rect -19089 -21986 -18508 -21855
rect -18142 -22031 -17640 -21679
rect -7292 -21464 -6706 -21344
rect -6465 -21391 -5669 -21239
rect -5560 -21341 -4960 -21189
rect -4603 -21341 -4003 -21189
rect -5549 -21464 -4963 -21344
rect -4592 -21464 -4006 -21344
rect -3765 -21391 -2969 -21239
rect -2860 -21341 -2260 -21189
rect -1978 -21341 -1378 -21189
rect 783 -21222 1187 -21070
rect -2849 -21464 -2263 -21344
rect -1967 -21464 -1381 -21344
rect 678 -21355 1259 -21224
rect 2388 -21224 2792 -21072
rect 2283 -21357 2864 -21226
rect 17342 -21251 18251 -21093
rect -7300 -21844 -6714 -21724
rect -6463 -21844 -5877 -21724
rect -22727 -22195 -22226 -22082
rect -18150 -22148 -17649 -22035
rect -7303 -21999 -6703 -21847
rect -6466 -21999 -5866 -21847
rect -5757 -21949 -4961 -21797
rect -4600 -21844 -4014 -21724
rect -3763 -21844 -3177 -21724
rect -1048 -21786 -840 -21534
rect -635 -21786 -329 -21434
rect -326 -21786 -20 -21434
rect -16 -21785 290 -21433
rect 1392 -21729 1894 -21377
rect 2997 -21731 3499 -21379
rect -4603 -21999 -4003 -21847
rect -3766 -21999 -3166 -21847
rect -3057 -21949 -2261 -21797
rect 1401 -21846 1902 -21733
rect 3006 -21848 3507 -21735
rect 3914 -21777 4122 -21525
rect 4327 -21777 4633 -21425
rect 4636 -21777 4942 -21425
rect 4946 -21776 5252 -21424
rect 5527 -21686 5735 -21434
rect 5941 -21686 6149 -21434
rect 6303 -21686 6511 -21434
rect 6597 -21686 6805 -21434
rect 6907 -21686 7115 -21434
rect 7216 -21686 7424 -21434
rect 17439 -21564 17843 -21312
rect 37040 -20887 37444 -20735
rect 45831 -20772 46412 -20641
rect 53519 -20663 53923 -20411
rect 54394 -20585 54896 -20233
rect 62201 -20343 62782 -20212
rect 62273 -20597 62677 -20345
rect 63148 -20519 63650 -20167
rect 71354 -20326 71935 -20195
rect 55029 -20738 55610 -20607
rect 63783 -20672 64364 -20541
rect 71426 -20580 71830 -20328
rect 72301 -20502 72803 -20150
rect 80718 -20288 81299 -20157
rect 72936 -20655 73517 -20524
rect 80790 -20542 81194 -20290
rect 81665 -20464 82167 -20112
rect 82300 -20617 82881 -20486
rect 19545 -21660 20341 -21508
rect 20450 -21610 21050 -21458
rect 21287 -21610 21887 -21458
rect 6736 -21863 7420 -21715
rect 20461 -21733 21047 -21613
rect 21298 -21733 21884 -21613
rect 22245 -21660 23041 -21508
rect 23150 -21610 23750 -21458
rect 23987 -21610 24587 -21458
rect 23161 -21733 23747 -21613
rect 23998 -21733 24584 -21613
rect -1048 -22043 278 -21926
rect 3914 -22034 5240 -21917
rect -20934 -22311 -19608 -22194
rect -12446 -22500 -12042 -22348
rect -14028 -22829 -13624 -22577
rect -12518 -22633 -11937 -22502
rect 18665 -22113 19251 -21993
rect 19547 -22113 20133 -21993
rect 18662 -22268 19262 -22116
rect 19544 -22268 20144 -22116
rect 20253 -22218 21049 -22066
rect 21290 -22113 21876 -21993
rect 22247 -22113 22833 -21993
rect 21287 -22268 21887 -22116
rect 22244 -22268 22844 -22116
rect 22953 -22218 23749 -22066
rect 23990 -22113 24576 -21993
rect 27601 -22036 28005 -21884
rect 23987 -22268 24587 -22116
rect 27529 -22169 28110 -22038
rect -14100 -22962 -13519 -22831
rect -13153 -23007 -12651 -22655
rect 26894 -22543 27396 -22191
rect 45903 -20926 46307 -20774
rect 55101 -20892 55505 -20740
rect 63855 -20826 64259 -20674
rect 73008 -20809 73412 -20657
rect 82372 -20771 82776 -20619
rect 36041 -22047 36445 -21895
rect 35969 -22180 36550 -22049
rect 26886 -22660 27387 -22547
rect -13161 -23124 -12660 -23011
rect 28439 -22829 28745 -22477
rect 28877 -22829 29085 -22477
rect 30333 -22771 30541 -22419
rect 30803 -22771 31011 -22219
rect 31026 -22771 31234 -22219
rect 31254 -22771 31560 -22219
rect 31580 -22771 31788 -22419
rect 35334 -22554 35836 -22202
rect 44904 -22086 45308 -21934
rect 44832 -22219 45413 -22088
rect 35326 -22671 35827 -22558
rect -15177 -23830 -14577 -23678
rect -14340 -23830 -13740 -23678
rect -15174 -23953 -14588 -23833
rect -14337 -23953 -13751 -23833
rect -13631 -23880 -12835 -23728
rect -12477 -23830 -11877 -23678
rect -11640 -23830 -11040 -23678
rect -12474 -23953 -11888 -23833
rect -11637 -23953 -11051 -23833
rect -10931 -23880 -10135 -23728
rect 21852 -23128 24631 -22979
rect 28362 -23020 29161 -22886
rect 30267 -23034 31792 -22821
rect 36879 -22840 37185 -22488
rect 37317 -22840 37525 -22488
rect 38773 -22782 38981 -22430
rect 39243 -22782 39451 -22230
rect 39466 -22782 39674 -22230
rect 39694 -22782 40000 -22230
rect 40020 -22782 40228 -22430
rect 44197 -22593 44699 -22241
rect 54102 -22052 54506 -21900
rect 54030 -22185 54611 -22054
rect 44189 -22710 44690 -22597
rect 36802 -23031 37601 -22897
rect 38707 -23045 40232 -22832
rect 45742 -22879 46048 -22527
rect 46180 -22879 46388 -22527
rect 47636 -22821 47844 -22469
rect 48106 -22821 48314 -22269
rect 48329 -22821 48537 -22269
rect 48557 -22821 48863 -22269
rect 48883 -22821 49091 -22469
rect 53395 -22559 53897 -22207
rect 62856 -21986 63260 -21834
rect 62784 -22119 63365 -21988
rect 53387 -22676 53888 -22563
rect 54940 -22845 55246 -22493
rect 55378 -22845 55586 -22493
rect 56834 -22787 57042 -22435
rect 57304 -22787 57512 -22235
rect 57527 -22787 57735 -22235
rect 57755 -22787 58061 -22235
rect 58081 -22787 58289 -22435
rect 62149 -22493 62651 -22141
rect 72009 -21969 72413 -21817
rect 71937 -22102 72518 -21971
rect 62141 -22610 62642 -22497
rect 63694 -22779 64000 -22427
rect 64132 -22779 64340 -22427
rect 65588 -22721 65796 -22369
rect 66058 -22721 66266 -22169
rect 66281 -22721 66489 -22169
rect 66509 -22721 66815 -22169
rect 66835 -22721 67043 -22369
rect 71302 -22476 71804 -22124
rect 81373 -21931 81777 -21779
rect 81301 -22064 81882 -21933
rect 71294 -22593 71795 -22480
rect 72847 -22762 73153 -22410
rect 73285 -22762 73493 -22410
rect 74741 -22704 74949 -22352
rect 75211 -22704 75419 -22152
rect 75434 -22704 75642 -22152
rect 75662 -22704 75968 -22152
rect 75988 -22704 76196 -22352
rect 80666 -22438 81168 -22086
rect 80658 -22555 81159 -22442
rect 82211 -22724 82517 -22372
rect 82649 -22724 82857 -22372
rect 84105 -22666 84313 -22314
rect 84575 -22666 84783 -22114
rect 84798 -22666 85006 -22114
rect 85026 -22666 85332 -22114
rect 85352 -22666 85560 -22314
rect 45665 -23070 46464 -22936
rect 47570 -23084 49095 -22871
rect 54863 -23036 55662 -22902
rect 56768 -23050 58293 -22837
rect 63617 -22970 64416 -22836
rect 65522 -22984 67047 -22771
rect 72770 -22953 73569 -22819
rect 74675 -22967 76200 -22754
rect 82134 -22915 82933 -22781
rect 84039 -22929 85564 -22716
rect 17313 -23875 17962 -23734
rect 18259 -23875 18908 -23734
rect 19210 -23808 20536 -23691
rect -7303 -24097 -6703 -23945
rect -6466 -24097 -5866 -23945
rect -17673 -24362 -16874 -24228
rect -15166 -24333 -14580 -24213
rect -19149 -24701 -18648 -24588
rect -21350 -25256 -21044 -25004
rect -20445 -25257 -20139 -25005
rect -19141 -25057 -18639 -24705
rect -17596 -24771 -17290 -24419
rect -17158 -24771 -16950 -24419
rect -15177 -24488 -14577 -24336
rect -14339 -24438 -13543 -24286
rect -13423 -24333 -12837 -24213
rect -12466 -24333 -11880 -24213
rect -13434 -24488 -12834 -24336
rect -12477 -24488 -11877 -24336
rect -11639 -24438 -10843 -24286
rect -10723 -24333 -10137 -24213
rect -9841 -24333 -9255 -24213
rect -7300 -24220 -6714 -24100
rect -6463 -24220 -5877 -24100
rect -5757 -24147 -4961 -23995
rect -4603 -24097 -4003 -23945
rect -3766 -24097 -3166 -23945
rect -4600 -24220 -4014 -24100
rect -3763 -24220 -3177 -24100
rect -3057 -24147 -2261 -23995
rect -1048 -24018 278 -23901
rect 3914 -24027 5240 -23910
rect -10734 -24488 -10134 -24336
rect -9852 -24488 -9252 -24336
rect -8803 -24579 -8595 -24227
rect -8463 -24579 -8157 -24227
rect -1048 -24410 -840 -24158
rect -22556 -25599 -22152 -25347
rect -21471 -25452 -20822 -25311
rect -20566 -25453 -19917 -25312
rect -18506 -25210 -17925 -25079
rect -18434 -25364 -18030 -25212
rect -7292 -24600 -6706 -24480
rect -8879 -24770 -8080 -24636
rect -7303 -24755 -6703 -24603
rect -6465 -24705 -5669 -24553
rect -5549 -24600 -4963 -24480
rect -4592 -24600 -4006 -24480
rect -5560 -24755 -4960 -24603
rect -4603 -24755 -4003 -24603
rect -3765 -24705 -2969 -24553
rect -2849 -24600 -2263 -24480
rect -1967 -24600 -1381 -24480
rect -635 -24510 -329 -24158
rect -326 -24510 -20 -24158
rect -16 -24511 290 -24159
rect 1401 -24211 1902 -24098
rect 3006 -24209 3507 -24096
rect 1392 -24567 1894 -24215
rect 2997 -24565 3499 -24213
rect 3914 -24419 4122 -24167
rect 4327 -24519 4633 -24167
rect 4636 -24519 4942 -24167
rect 4946 -24520 5252 -24168
rect 6736 -24229 7420 -24081
rect 17434 -24182 17740 -23930
rect 18380 -24182 18686 -23930
rect 5527 -24510 5735 -24258
rect 5941 -24510 6149 -24258
rect 6303 -24510 6511 -24258
rect 6597 -24510 6805 -24258
rect 6907 -24510 7115 -24258
rect 7216 -24510 7424 -24258
rect 19198 -24301 19504 -23949
rect 19508 -24300 19814 -23948
rect 19817 -24300 20123 -23948
rect 20328 -24200 20536 -23948
rect 21107 -24054 21315 -23802
rect 21317 -24054 21525 -23802
rect 21937 -23945 22145 -23193
rect 22337 -23945 22545 -23193
rect 22937 -23945 23145 -23193
rect 23337 -23945 23545 -23193
rect 23937 -23945 24145 -23193
rect 24337 -23945 24545 -23193
rect 27877 -23666 28378 -23553
rect 26938 -23846 27519 -23715
rect 21086 -24243 21617 -24110
rect 21060 -24366 21646 -24246
rect -2860 -24755 -2260 -24603
rect -1978 -24755 -1378 -24603
rect 678 -24720 1259 -24589
rect 783 -24874 1187 -24722
rect 2283 -24718 2864 -24587
rect 2388 -24872 2792 -24720
rect 21057 -24521 21657 -24369
rect 27010 -24100 27414 -23848
rect 27885 -24022 28387 -23670
rect 31545 -23697 32046 -23584
rect 36317 -23677 36818 -23564
rect 30606 -23877 31187 -23746
rect 28520 -24175 29101 -24044
rect 30678 -24131 31082 -23879
rect 31553 -24053 32055 -23701
rect 35378 -23857 35959 -23726
rect 28592 -24329 28996 -24177
rect 32188 -24206 32769 -24075
rect 35450 -24111 35854 -23859
rect 36325 -24033 36827 -23681
rect 39985 -23708 40486 -23595
rect 39046 -23888 39627 -23757
rect 36960 -24186 37541 -24055
rect 39118 -24142 39522 -23890
rect 39993 -24064 40495 -23712
rect 45180 -23716 45681 -23603
rect 44241 -23896 44822 -23765
rect 32260 -24360 32664 -24208
rect 37032 -24340 37436 -24188
rect 40628 -24217 41209 -24086
rect 44313 -24150 44717 -23898
rect 45188 -24072 45690 -23720
rect 48848 -23747 49349 -23634
rect 54378 -23682 54879 -23569
rect 47909 -23927 48490 -23796
rect -22653 -25818 -21744 -25660
rect 27593 -25489 27997 -25337
rect 27521 -25622 28102 -25491
rect 26886 -25996 27388 -25644
rect 40700 -24371 41104 -24219
rect 45823 -24225 46404 -24094
rect 47981 -24181 48385 -23929
rect 48856 -24103 49358 -23751
rect 53439 -23862 54020 -23731
rect 53511 -24116 53915 -23864
rect 54386 -24038 54888 -23686
rect 58046 -23713 58547 -23600
rect 63132 -23616 63633 -23503
rect 57107 -23893 57688 -23762
rect 31261 -25520 31665 -25368
rect 31189 -25653 31770 -25522
rect -22893 -26353 -21567 -26236
rect 10534 -26166 11134 -26014
rect 11416 -26166 12016 -26014
rect 10537 -26289 11123 -26169
rect 11419 -26289 12005 -26169
rect 12125 -26216 12921 -26064
rect 13159 -26166 13759 -26014
rect 14116 -26166 14716 -26014
rect 13162 -26289 13748 -26169
rect 14119 -26289 14705 -26169
rect 14825 -26216 15621 -26064
rect 15859 -26166 16459 -26014
rect 26878 -26113 27379 -26000
rect 15862 -26289 16448 -26169
rect 28431 -26282 28737 -25930
rect 28869 -26282 29077 -25930
rect 30554 -26027 31056 -25675
rect 36033 -25500 36437 -25348
rect 35961 -25633 36542 -25502
rect 30546 -26144 31047 -26031
rect 32099 -26313 32405 -25961
rect 32537 -26313 32745 -25961
rect 35326 -26007 35828 -25655
rect 45895 -24379 46299 -24227
rect 49491 -24256 50072 -24125
rect 55021 -24191 55602 -24060
rect 57179 -24147 57583 -23895
rect 58054 -24069 58556 -23717
rect 62193 -23796 62774 -23665
rect 62265 -24050 62669 -23798
rect 63140 -23972 63642 -23620
rect 66800 -23647 67301 -23534
rect 72285 -23599 72786 -23486
rect 65861 -23827 66442 -23696
rect 39701 -25531 40105 -25379
rect 39629 -25664 40210 -25533
rect 35318 -26124 35819 -26011
rect 36871 -26293 37177 -25941
rect 37309 -26293 37517 -25941
rect 38994 -26038 39496 -25686
rect 49563 -24410 49967 -24258
rect 55093 -24345 55497 -24193
rect 58689 -24222 59270 -24091
rect 63775 -24125 64356 -23994
rect 65933 -24081 66337 -23829
rect 66808 -24003 67310 -23651
rect 71346 -23779 71927 -23648
rect 44896 -25539 45300 -25387
rect 44824 -25672 45405 -25541
rect 38986 -26155 39487 -26042
rect 40539 -26324 40845 -25972
rect 40977 -26324 41185 -25972
rect 44189 -26046 44691 -25694
rect 58761 -24376 59165 -24224
rect 63847 -24279 64251 -24127
rect 67443 -24156 68024 -24025
rect 71418 -24033 71822 -23781
rect 72293 -23955 72795 -23603
rect 75953 -23630 76454 -23517
rect 81649 -23561 82150 -23448
rect 75014 -23810 75595 -23679
rect 72928 -24108 73509 -23977
rect 75086 -24064 75490 -23812
rect 75961 -23986 76463 -23634
rect 80710 -23741 81291 -23610
rect 80782 -23995 81186 -23743
rect 81657 -23917 82159 -23565
rect 85317 -23592 85818 -23479
rect 84378 -23772 84959 -23641
rect 48564 -25570 48968 -25418
rect 48492 -25703 49073 -25572
rect 44181 -26163 44682 -26050
rect 45734 -26332 46040 -25980
rect 46172 -26332 46380 -25980
rect 47857 -26077 48359 -25725
rect 54094 -25505 54498 -25353
rect 54022 -25638 54603 -25507
rect 47849 -26194 48350 -26081
rect -22893 -26745 -22685 -26493
rect -22480 -26845 -22174 -26493
rect -22171 -26845 -21865 -26493
rect -21861 -26846 -21555 -26494
rect -17435 -26524 -17031 -26372
rect -6274 -26480 -5590 -26332
rect -3774 -26480 -3090 -26332
rect -1274 -26480 -590 -26332
rect 1226 -26480 1910 -26332
rect 3726 -26480 4410 -26332
rect 6726 -26480 7410 -26332
rect 28354 -26473 29153 -26339
rect 32022 -26504 32821 -26370
rect 36794 -26484 37593 -26350
rect 49402 -26363 49708 -26011
rect 49840 -26363 50048 -26011
rect 53387 -26012 53889 -25660
rect 67515 -24310 67919 -24158
rect 73000 -24262 73404 -24110
rect 76596 -24139 77177 -24008
rect 82292 -24070 82873 -23939
rect 84450 -24026 84854 -23774
rect 85325 -23948 85827 -23596
rect 57762 -25536 58166 -25384
rect 57690 -25669 58271 -25538
rect 53379 -26129 53880 -26016
rect 54932 -26298 55238 -25946
rect 55370 -26298 55578 -25946
rect 57055 -26043 57557 -25691
rect 62848 -25439 63252 -25287
rect 62776 -25572 63357 -25441
rect 62141 -25946 62643 -25594
rect 76668 -24293 77072 -24141
rect 82364 -24224 82768 -24072
rect 85960 -24101 86541 -23970
rect 66516 -25470 66920 -25318
rect 66444 -25603 67025 -25472
rect 57047 -26160 57548 -26047
rect 58600 -26329 58906 -25977
rect 59038 -26329 59246 -25977
rect 62133 -26063 62634 -25950
rect 63686 -26232 63992 -25880
rect 64124 -26232 64332 -25880
rect 65809 -25977 66311 -25625
rect 72001 -25422 72405 -25270
rect 71929 -25555 72510 -25424
rect 65801 -26094 66302 -25981
rect 67354 -26263 67660 -25911
rect 67792 -26263 68000 -25911
rect 71294 -25929 71796 -25577
rect 86032 -24255 86436 -24103
rect 75669 -25453 76073 -25301
rect 75597 -25586 76178 -25455
rect 71286 -26046 71787 -25933
rect 72839 -26215 73145 -25863
rect 73277 -26215 73485 -25863
rect 74962 -25960 75464 -25608
rect 81365 -25384 81769 -25232
rect 81293 -25517 81874 -25386
rect 80658 -25891 81160 -25539
rect 85033 -25415 85437 -25263
rect 84961 -25548 85542 -25417
rect 74954 -26077 75455 -25964
rect 76507 -26246 76813 -25894
rect 76945 -26246 77153 -25894
rect 80650 -26008 81151 -25895
rect 82203 -26177 82509 -25825
rect 82641 -26177 82849 -25825
rect 84326 -25922 84828 -25570
rect 84318 -26039 84819 -25926
rect 85871 -26208 86177 -25856
rect 86309 -26208 86517 -25856
rect -19017 -26853 -18613 -26601
rect -17507 -26657 -16926 -26526
rect -19089 -26986 -18508 -26855
rect -18142 -27031 -17640 -26679
rect -7483 -26761 -7275 -26509
rect -7069 -26761 -6861 -26509
rect -6707 -26761 -6499 -26509
rect -6413 -26761 -6205 -26509
rect -6103 -26761 -5895 -26509
rect -5794 -26761 -5586 -26509
rect -4983 -26761 -4775 -26509
rect -4569 -26761 -4361 -26509
rect -4207 -26761 -3999 -26509
rect -3913 -26761 -3705 -26509
rect -3603 -26761 -3395 -26509
rect -3294 -26761 -3086 -26509
rect -2483 -26761 -2275 -26509
rect -2069 -26761 -1861 -26509
rect -1707 -26761 -1499 -26509
rect -1413 -26761 -1205 -26509
rect -1103 -26761 -895 -26509
rect -794 -26761 -586 -26509
rect 17 -26761 225 -26509
rect 431 -26761 639 -26509
rect 793 -26761 1001 -26509
rect 1087 -26761 1295 -26509
rect 1397 -26761 1605 -26509
rect 1706 -26761 1914 -26509
rect 2517 -26761 2725 -26509
rect 2931 -26761 3139 -26509
rect 3293 -26761 3501 -26509
rect 3587 -26761 3795 -26509
rect 3897 -26761 4105 -26509
rect 4206 -26761 4414 -26509
rect 5517 -26761 5725 -26509
rect 5931 -26761 6139 -26509
rect 6293 -26761 6501 -26509
rect 6587 -26761 6795 -26509
rect 6897 -26761 7105 -26509
rect 7206 -26761 7414 -26509
rect 40462 -26515 41261 -26381
rect 45657 -26523 46456 -26389
rect 11417 -26774 12213 -26622
rect 12333 -26669 12919 -26549
rect 13170 -26669 13756 -26549
rect 12322 -26824 12922 -26672
rect 13159 -26824 13759 -26672
rect 14117 -26774 14913 -26622
rect 15033 -26669 15619 -26549
rect 15870 -26669 16456 -26549
rect 49325 -26554 50124 -26420
rect 54855 -26489 55654 -26355
rect 58523 -26520 59322 -26386
rect 63609 -26423 64408 -26289
rect 67277 -26454 68076 -26320
rect 72762 -26406 73561 -26272
rect 76430 -26437 77229 -26303
rect 82126 -26368 82925 -26234
rect 85794 -26399 86593 -26265
rect 15022 -26824 15622 -26672
rect 15859 -26824 16459 -26672
rect -18150 -27148 -17649 -27035
rect -27056 -41305 -26878 -34052
rect -26846 -41269 -26394 -34079
rect -14479 -35494 -13879 -35342
rect -13642 -35494 -13042 -35342
rect -14476 -35617 -13890 -35497
rect -13639 -35617 -13053 -35497
rect -12933 -35544 -12137 -35392
rect -11779 -35494 -11179 -35342
rect -10942 -35494 -10342 -35342
rect -11776 -35617 -11190 -35497
rect -10939 -35617 -10353 -35497
rect -10233 -35544 -9437 -35392
rect -16975 -35953 -16176 -35819
rect -14468 -35997 -13882 -35877
rect -19372 -36253 -18968 -36101
rect -22078 -36708 -21772 -36356
rect -21768 -36709 -21462 -36357
rect -21459 -36709 -21153 -36357
rect -19444 -36386 -18863 -36255
rect -18451 -36292 -17950 -36179
rect -20948 -36709 -20740 -36457
rect -20079 -36760 -19577 -36408
rect -18443 -36648 -17941 -36296
rect -16898 -36362 -16592 -36010
rect -16460 -36362 -16252 -36010
rect -14479 -36152 -13879 -36000
rect -13641 -36102 -12845 -35950
rect -12725 -35997 -12139 -35877
rect -11768 -35997 -11182 -35877
rect -12736 -36152 -12136 -36000
rect -11779 -36152 -11179 -36000
rect -10941 -36102 -10145 -35950
rect -10025 -35997 -9439 -35877
rect -9143 -35997 -8557 -35877
rect -10036 -36152 -9436 -36000
rect -9154 -36152 -8554 -36000
rect -8132 -36236 -7924 -35884
rect -7792 -36236 -7486 -35884
rect -6785 -36026 -6577 -35774
rect -6371 -36026 -6163 -35774
rect -6009 -36026 -5801 -35774
rect -5715 -36026 -5507 -35774
rect -5405 -36026 -5197 -35774
rect -5096 -36026 -4888 -35774
rect -4285 -36026 -4077 -35774
rect -3871 -36026 -3663 -35774
rect -3509 -36026 -3301 -35774
rect -3215 -36026 -3007 -35774
rect -2905 -36026 -2697 -35774
rect -2596 -36026 -2388 -35774
rect -1785 -36026 -1577 -35774
rect -1371 -36026 -1163 -35774
rect -1009 -36026 -801 -35774
rect -715 -36026 -507 -35774
rect -405 -36026 -197 -35774
rect -96 -36026 112 -35774
rect 715 -36026 923 -35774
rect 1129 -36026 1337 -35774
rect 1491 -36026 1699 -35774
rect 1785 -36026 1993 -35774
rect 2095 -36026 2303 -35774
rect 2404 -36026 2612 -35774
rect 3215 -36026 3423 -35774
rect 3629 -36026 3837 -35774
rect 3991 -36026 4199 -35774
rect 4285 -36026 4493 -35774
rect 4595 -36026 4803 -35774
rect 4904 -36026 5112 -35774
rect 6215 -36026 6423 -35774
rect 6629 -36026 6837 -35774
rect 6991 -36026 7199 -35774
rect 7285 -36026 7493 -35774
rect 7595 -36026 7803 -35774
rect 7904 -36026 8112 -35774
rect -6345 -36214 -5759 -36094
rect -5576 -36203 -4892 -36055
rect -3076 -36203 -2392 -36055
rect -576 -36203 108 -36055
rect 1924 -36203 2608 -36055
rect 4424 -36203 5108 -36055
rect 7424 -36203 8108 -36055
rect -22066 -36966 -20740 -36849
rect -20087 -36877 -19586 -36764
rect -17808 -36801 -17227 -36670
rect -17736 -36955 -17332 -36803
rect -8208 -36427 -7409 -36293
rect -6348 -36369 -5748 -36217
rect -11986 -36929 -11187 -36795
rect 28583 -36804 29084 -36691
rect 27644 -36984 28225 -36853
rect -13462 -37268 -12961 -37155
rect -13454 -37624 -12952 -37272
rect -11909 -37338 -11603 -36986
rect -11471 -37338 -11263 -36986
rect -21314 -38162 -20910 -38010
rect -16737 -38115 -16333 -37963
rect -12819 -37777 -12238 -37646
rect -12747 -37931 -12343 -37779
rect 27716 -37238 28120 -36986
rect 28591 -37160 29093 -36808
rect 37023 -36815 37524 -36702
rect 36084 -36995 36665 -36864
rect 29226 -37313 29807 -37182
rect 36156 -37249 36560 -36997
rect 37031 -37171 37533 -36819
rect 45886 -36854 46387 -36741
rect 55084 -36820 55585 -36707
rect 63838 -36754 64339 -36641
rect 72991 -36737 73492 -36624
rect 82355 -36699 82856 -36586
rect 44947 -37034 45528 -36903
rect 29298 -37467 29702 -37315
rect 37666 -37324 38247 -37193
rect 45019 -37288 45423 -37036
rect 45894 -37210 46396 -36858
rect 54145 -37000 54726 -36869
rect -6605 -37932 -6005 -37780
rect -21386 -38295 -20805 -38164
rect -22021 -38669 -21519 -38317
rect -20248 -38644 -19942 -38292
rect -19938 -38645 -19632 -38293
rect -19629 -38645 -19323 -38293
rect -19118 -38645 -18910 -38393
rect -18319 -38444 -17915 -38192
rect -16809 -38248 -16228 -38117
rect -18391 -38577 -17810 -38446
rect -17444 -38622 -16942 -38270
rect -6594 -38055 -6008 -37935
rect -5767 -37982 -4971 -37830
rect -4862 -37932 -4262 -37780
rect -3905 -37932 -3305 -37780
rect -4851 -38055 -4265 -37935
rect -3894 -38055 -3308 -37935
rect -3067 -37982 -2271 -37830
rect -2162 -37932 -1562 -37780
rect -1280 -37932 -680 -37780
rect 1481 -37813 1885 -37661
rect -2151 -38055 -1565 -37935
rect -1269 -38055 -683 -37935
rect 1376 -37946 1957 -37815
rect 3086 -37815 3490 -37663
rect 2981 -37948 3562 -37817
rect 18040 -37842 18949 -37684
rect -6602 -38435 -6016 -38315
rect -5765 -38435 -5179 -38315
rect -22029 -38786 -21528 -38673
rect -17452 -38739 -16951 -38626
rect -6605 -38590 -6005 -38438
rect -5768 -38590 -5168 -38438
rect -5059 -38540 -4263 -38388
rect -3902 -38435 -3316 -38315
rect -3065 -38435 -2479 -38315
rect -350 -38377 -142 -38125
rect 63 -38377 369 -38025
rect 372 -38377 678 -38025
rect 682 -38376 988 -38024
rect 2090 -38320 2592 -37968
rect 3695 -38322 4197 -37970
rect -3905 -38590 -3305 -38438
rect -3068 -38590 -2468 -38438
rect -2359 -38540 -1563 -38388
rect 2099 -38437 2600 -38324
rect 3704 -38439 4205 -38326
rect 4612 -38368 4820 -38116
rect 5025 -38368 5331 -38016
rect 5334 -38368 5640 -38016
rect 5644 -38367 5950 -38015
rect 6225 -38277 6433 -38025
rect 6639 -38277 6847 -38025
rect 7001 -38277 7209 -38025
rect 7295 -38277 7503 -38025
rect 7605 -38277 7813 -38025
rect 7914 -38277 8122 -38025
rect 18137 -38155 18541 -37903
rect 37738 -37478 38142 -37326
rect 46529 -37363 47110 -37232
rect 54217 -37254 54621 -37002
rect 55092 -37176 55594 -36824
rect 62899 -36934 63480 -36803
rect 62971 -37188 63375 -36936
rect 63846 -37110 64348 -36758
rect 72052 -36917 72633 -36786
rect 55727 -37329 56308 -37198
rect 64481 -37263 65062 -37132
rect 72124 -37171 72528 -36919
rect 72999 -37093 73501 -36741
rect 81416 -36879 81997 -36748
rect 73634 -37246 74215 -37115
rect 81488 -37133 81892 -36881
rect 82363 -37055 82865 -36703
rect 82998 -37208 83579 -37077
rect 20243 -38251 21039 -38099
rect 21148 -38201 21748 -38049
rect 21985 -38201 22585 -38049
rect 7434 -38454 8118 -38306
rect 21159 -38324 21745 -38204
rect 21996 -38324 22582 -38204
rect 22943 -38251 23739 -38099
rect 23848 -38201 24448 -38049
rect 24685 -38201 25285 -38049
rect 23859 -38324 24445 -38204
rect 24696 -38324 25282 -38204
rect -350 -38634 976 -38517
rect 4612 -38625 5938 -38508
rect -20236 -38902 -18910 -38785
rect -11748 -39091 -11344 -38939
rect -13330 -39420 -12926 -39168
rect -11820 -39224 -11239 -39093
rect 19363 -38704 19949 -38584
rect 20245 -38704 20831 -38584
rect 19360 -38859 19960 -38707
rect 20242 -38859 20842 -38707
rect 20951 -38809 21747 -38657
rect 21988 -38704 22574 -38584
rect 22945 -38704 23531 -38584
rect 21985 -38859 22585 -38707
rect 22942 -38859 23542 -38707
rect 23651 -38809 24447 -38657
rect 24688 -38704 25274 -38584
rect 28299 -38627 28703 -38475
rect 24685 -38859 25285 -38707
rect 28227 -38760 28808 -38629
rect -13402 -39553 -12821 -39422
rect -12455 -39598 -11953 -39246
rect 27592 -39134 28094 -38782
rect 46601 -37517 47005 -37365
rect 55799 -37483 56203 -37331
rect 64553 -37417 64957 -37265
rect 73706 -37400 74110 -37248
rect 83070 -37362 83474 -37210
rect 36739 -38638 37143 -38486
rect 36667 -38771 37248 -38640
rect 27584 -39251 28085 -39138
rect -12463 -39715 -11962 -39602
rect 29137 -39420 29443 -39068
rect 29575 -39420 29783 -39068
rect 31031 -39362 31239 -39010
rect 31501 -39362 31709 -38810
rect 31724 -39362 31932 -38810
rect 31952 -39362 32258 -38810
rect 32278 -39362 32486 -39010
rect 36032 -39145 36534 -38793
rect 45602 -38677 46006 -38525
rect 45530 -38810 46111 -38679
rect 36024 -39262 36525 -39149
rect -14479 -40421 -13879 -40269
rect -13642 -40421 -13042 -40269
rect -14476 -40544 -13890 -40424
rect -13639 -40544 -13053 -40424
rect -12933 -40471 -12137 -40319
rect -11779 -40421 -11179 -40269
rect -10942 -40421 -10342 -40269
rect -11776 -40544 -11190 -40424
rect -10939 -40544 -10353 -40424
rect -10233 -40471 -9437 -40319
rect 22550 -39719 25329 -39570
rect 29060 -39611 29859 -39477
rect 30965 -39625 32490 -39412
rect 37577 -39431 37883 -39079
rect 38015 -39431 38223 -39079
rect 39471 -39373 39679 -39021
rect 39941 -39373 40149 -38821
rect 40164 -39373 40372 -38821
rect 40392 -39373 40698 -38821
rect 40718 -39373 40926 -39021
rect 44895 -39184 45397 -38832
rect 54800 -38643 55204 -38491
rect 54728 -38776 55309 -38645
rect 44887 -39301 45388 -39188
rect 37500 -39622 38299 -39488
rect 39405 -39636 40930 -39423
rect 46440 -39470 46746 -39118
rect 46878 -39470 47086 -39118
rect 48334 -39412 48542 -39060
rect 48804 -39412 49012 -38860
rect 49027 -39412 49235 -38860
rect 49255 -39412 49561 -38860
rect 49581 -39412 49789 -39060
rect 54093 -39150 54595 -38798
rect 63554 -38577 63958 -38425
rect 63482 -38710 64063 -38579
rect 54085 -39267 54586 -39154
rect 55638 -39436 55944 -39084
rect 56076 -39436 56284 -39084
rect 57532 -39378 57740 -39026
rect 58002 -39378 58210 -38826
rect 58225 -39378 58433 -38826
rect 58453 -39378 58759 -38826
rect 58779 -39378 58987 -39026
rect 62847 -39084 63349 -38732
rect 72707 -38560 73111 -38408
rect 72635 -38693 73216 -38562
rect 62839 -39201 63340 -39088
rect 64392 -39370 64698 -39018
rect 64830 -39370 65038 -39018
rect 66286 -39312 66494 -38960
rect 66756 -39312 66964 -38760
rect 66979 -39312 67187 -38760
rect 67207 -39312 67513 -38760
rect 67533 -39312 67741 -38960
rect 72000 -39067 72502 -38715
rect 82071 -38522 82475 -38370
rect 81999 -38655 82580 -38524
rect 71992 -39184 72493 -39071
rect 73545 -39353 73851 -39001
rect 73983 -39353 74191 -39001
rect 75439 -39295 75647 -38943
rect 75909 -39295 76117 -38743
rect 76132 -39295 76340 -38743
rect 76360 -39295 76666 -38743
rect 76686 -39295 76894 -38943
rect 81364 -39029 81866 -38677
rect 81356 -39146 81857 -39033
rect 82909 -39315 83215 -38963
rect 83347 -39315 83555 -38963
rect 84803 -39257 85011 -38905
rect 85273 -39257 85481 -38705
rect 85496 -39257 85704 -38705
rect 85724 -39257 86030 -38705
rect 86050 -39257 86258 -38905
rect 46363 -39661 47162 -39527
rect 48268 -39675 49793 -39462
rect 55561 -39627 56360 -39493
rect 57466 -39641 58991 -39428
rect 64315 -39561 65114 -39427
rect 66220 -39575 67745 -39362
rect 73468 -39544 74267 -39410
rect 75373 -39558 76898 -39345
rect 82832 -39506 83631 -39372
rect 84737 -39520 86262 -39307
rect 18011 -40466 18660 -40325
rect 18957 -40466 19606 -40325
rect 19908 -40399 21234 -40282
rect -6605 -40688 -6005 -40536
rect -5768 -40688 -5168 -40536
rect -16975 -40953 -16176 -40819
rect -14468 -40924 -13882 -40804
rect -18451 -41292 -17950 -41179
rect -20652 -41847 -20346 -41595
rect -19747 -41848 -19441 -41596
rect -18443 -41648 -17941 -41296
rect -16898 -41362 -16592 -41010
rect -16460 -41362 -16252 -41010
rect -14479 -41079 -13879 -40927
rect -13641 -41029 -12845 -40877
rect -12725 -40924 -12139 -40804
rect -11768 -40924 -11182 -40804
rect -12736 -41079 -12136 -40927
rect -11779 -41079 -11179 -40927
rect -10941 -41029 -10145 -40877
rect -10025 -40924 -9439 -40804
rect -9143 -40924 -8557 -40804
rect -6602 -40811 -6016 -40691
rect -5765 -40811 -5179 -40691
rect -5059 -40738 -4263 -40586
rect -3905 -40688 -3305 -40536
rect -3068 -40688 -2468 -40536
rect -3902 -40811 -3316 -40691
rect -3065 -40811 -2479 -40691
rect -2359 -40738 -1563 -40586
rect -350 -40609 976 -40492
rect 4612 -40618 5938 -40501
rect -10036 -41079 -9436 -40927
rect -9154 -41079 -8554 -40927
rect -8105 -41170 -7897 -40818
rect -7765 -41170 -7459 -40818
rect -350 -41001 -142 -40749
rect -21858 -42190 -21454 -41938
rect -20773 -42043 -20124 -41902
rect -19868 -42044 -19219 -41903
rect -17808 -41801 -17227 -41670
rect -17736 -41955 -17332 -41803
rect -6594 -41191 -6008 -41071
rect -8181 -41361 -7382 -41227
rect -6605 -41346 -6005 -41194
rect -5767 -41296 -4971 -41144
rect -4851 -41191 -4265 -41071
rect -3894 -41191 -3308 -41071
rect -4862 -41346 -4262 -41194
rect -3905 -41346 -3305 -41194
rect -3067 -41296 -2271 -41144
rect -2151 -41191 -1565 -41071
rect -1269 -41191 -683 -41071
rect 63 -41101 369 -40749
rect 372 -41101 678 -40749
rect 682 -41102 988 -40750
rect 2099 -40802 2600 -40689
rect 3704 -40800 4205 -40687
rect 2090 -41158 2592 -40806
rect 3695 -41156 4197 -40804
rect 4612 -41010 4820 -40758
rect 5025 -41110 5331 -40758
rect 5334 -41110 5640 -40758
rect 5644 -41111 5950 -40759
rect 7434 -40820 8118 -40672
rect 18132 -40773 18438 -40521
rect 19078 -40773 19384 -40521
rect 6225 -41101 6433 -40849
rect 6639 -41101 6847 -40849
rect 7001 -41101 7209 -40849
rect 7295 -41101 7503 -40849
rect 7605 -41101 7813 -40849
rect 7914 -41101 8122 -40849
rect 19896 -40892 20202 -40540
rect 20206 -40891 20512 -40539
rect 20515 -40891 20821 -40539
rect 21026 -40791 21234 -40539
rect 21805 -40645 22013 -40393
rect 22015 -40645 22223 -40393
rect 22635 -40536 22843 -39784
rect 23035 -40536 23243 -39784
rect 23635 -40536 23843 -39784
rect 24035 -40536 24243 -39784
rect 24635 -40536 24843 -39784
rect 25035 -40536 25243 -39784
rect 28575 -40257 29076 -40144
rect 27636 -40437 28217 -40306
rect 21784 -40834 22315 -40701
rect 21758 -40957 22344 -40837
rect -2162 -41346 -1562 -41194
rect -1280 -41346 -680 -41194
rect 1376 -41311 1957 -41180
rect 1481 -41465 1885 -41313
rect 2981 -41309 3562 -41178
rect 3086 -41463 3490 -41311
rect 21755 -41112 22355 -40960
rect 27708 -40691 28112 -40439
rect 28583 -40613 29085 -40261
rect 32243 -40288 32744 -40175
rect 37015 -40268 37516 -40155
rect 31304 -40468 31885 -40337
rect 29218 -40766 29799 -40635
rect 31376 -40722 31780 -40470
rect 32251 -40644 32753 -40292
rect 36076 -40448 36657 -40317
rect 29290 -40920 29694 -40768
rect 32886 -40797 33467 -40666
rect 36148 -40702 36552 -40450
rect 37023 -40624 37525 -40272
rect 40683 -40299 41184 -40186
rect 39744 -40479 40325 -40348
rect 37658 -40777 38239 -40646
rect 39816 -40733 40220 -40481
rect 40691 -40655 41193 -40303
rect 45878 -40307 46379 -40194
rect 44939 -40487 45520 -40356
rect 32958 -40951 33362 -40799
rect 37730 -40931 38134 -40779
rect 41326 -40808 41907 -40677
rect 45011 -40741 45415 -40489
rect 45886 -40663 46388 -40311
rect 49546 -40338 50047 -40225
rect 55076 -40273 55577 -40160
rect 48607 -40518 49188 -40387
rect -21955 -42409 -21046 -42251
rect 28291 -42080 28695 -41928
rect 28219 -42213 28800 -42082
rect 27584 -42587 28086 -42235
rect 41398 -40962 41802 -40810
rect 46521 -40816 47102 -40685
rect 48679 -40772 49083 -40520
rect 49554 -40694 50056 -40342
rect 54137 -40453 54718 -40322
rect 54209 -40707 54613 -40455
rect 55084 -40629 55586 -40277
rect 58744 -40304 59245 -40191
rect 63830 -40207 64331 -40094
rect 57805 -40484 58386 -40353
rect 31959 -42111 32363 -41959
rect 31887 -42244 32468 -42113
rect -22195 -42944 -20869 -42827
rect 11232 -42757 11832 -42605
rect 12114 -42757 12714 -42605
rect 11235 -42880 11821 -42760
rect 12117 -42880 12703 -42760
rect 12823 -42807 13619 -42655
rect 13857 -42757 14457 -42605
rect 14814 -42757 15414 -42605
rect 13860 -42880 14446 -42760
rect 14817 -42880 15403 -42760
rect 15523 -42807 16319 -42655
rect 16557 -42757 17157 -42605
rect 27576 -42704 28077 -42591
rect 16560 -42880 17146 -42760
rect 29129 -42873 29435 -42521
rect 29567 -42873 29775 -42521
rect 31252 -42618 31754 -42266
rect 36731 -42091 37135 -41939
rect 36659 -42224 37240 -42093
rect 31244 -42735 31745 -42622
rect 32797 -42904 33103 -42552
rect 33235 -42904 33443 -42552
rect 36024 -42598 36526 -42246
rect 46593 -40970 46997 -40818
rect 50189 -40847 50770 -40716
rect 55719 -40782 56300 -40651
rect 57877 -40738 58281 -40486
rect 58752 -40660 59254 -40308
rect 62891 -40387 63472 -40256
rect 62963 -40641 63367 -40389
rect 63838 -40563 64340 -40211
rect 67498 -40238 67999 -40125
rect 72983 -40190 73484 -40077
rect 66559 -40418 67140 -40287
rect 40399 -42122 40803 -41970
rect 40327 -42255 40908 -42124
rect 36016 -42715 36517 -42602
rect 37569 -42884 37875 -42532
rect 38007 -42884 38215 -42532
rect 39692 -42629 40194 -42277
rect 50261 -41001 50665 -40849
rect 55791 -40936 56195 -40784
rect 59387 -40813 59968 -40682
rect 64473 -40716 65054 -40585
rect 66631 -40672 67035 -40420
rect 67506 -40594 68008 -40242
rect 72044 -40370 72625 -40239
rect 45594 -42130 45998 -41978
rect 45522 -42263 46103 -42132
rect 39684 -42746 40185 -42633
rect 41237 -42915 41543 -42563
rect 41675 -42915 41883 -42563
rect 44887 -42637 45389 -42285
rect 59459 -40967 59863 -40815
rect 64545 -40870 64949 -40718
rect 68141 -40747 68722 -40616
rect 72116 -40624 72520 -40372
rect 72991 -40546 73493 -40194
rect 76651 -40221 77152 -40108
rect 82347 -40152 82848 -40039
rect 75712 -40401 76293 -40270
rect 73626 -40699 74207 -40568
rect 75784 -40655 76188 -40403
rect 76659 -40577 77161 -40225
rect 81408 -40332 81989 -40201
rect 81480 -40586 81884 -40334
rect 82355 -40508 82857 -40156
rect 86015 -40183 86516 -40070
rect 85076 -40363 85657 -40232
rect 49262 -42161 49666 -42009
rect 49190 -42294 49771 -42163
rect 44879 -42754 45380 -42641
rect 46432 -42923 46738 -42571
rect 46870 -42923 47078 -42571
rect 48555 -42668 49057 -42316
rect 54792 -42096 55196 -41944
rect 54720 -42229 55301 -42098
rect 48547 -42785 49048 -42672
rect -22195 -43336 -21987 -43084
rect -21782 -43436 -21476 -43084
rect -21473 -43436 -21167 -43084
rect -21163 -43437 -20857 -43085
rect -16737 -43115 -16333 -42963
rect -5576 -43071 -4892 -42923
rect -3076 -43071 -2392 -42923
rect -576 -43071 108 -42923
rect 1924 -43071 2608 -42923
rect 4424 -43071 5108 -42923
rect 7424 -43071 8108 -42923
rect 29052 -43064 29851 -42930
rect 32720 -43095 33519 -42961
rect 37492 -43075 38291 -42941
rect 50100 -42954 50406 -42602
rect 50538 -42954 50746 -42602
rect 54085 -42603 54587 -42251
rect 68213 -40901 68617 -40749
rect 73698 -40853 74102 -40701
rect 77294 -40730 77875 -40599
rect 82990 -40661 83571 -40530
rect 85148 -40617 85552 -40365
rect 86023 -40539 86525 -40187
rect 58460 -42127 58864 -41975
rect 58388 -42260 58969 -42129
rect 54077 -42720 54578 -42607
rect 55630 -42889 55936 -42537
rect 56068 -42889 56276 -42537
rect 57753 -42634 58255 -42282
rect 63546 -42030 63950 -41878
rect 63474 -42163 64055 -42032
rect 62839 -42537 63341 -42185
rect 77366 -40884 77770 -40732
rect 83062 -40815 83466 -40663
rect 86658 -40692 87239 -40561
rect 67214 -42061 67618 -41909
rect 67142 -42194 67723 -42063
rect 57745 -42751 58246 -42638
rect 59298 -42920 59604 -42568
rect 59736 -42920 59944 -42568
rect 62831 -42654 63332 -42541
rect 64384 -42823 64690 -42471
rect 64822 -42823 65030 -42471
rect 66507 -42568 67009 -42216
rect 72699 -42013 73103 -41861
rect 72627 -42146 73208 -42015
rect 66499 -42685 67000 -42572
rect 68052 -42854 68358 -42502
rect 68490 -42854 68698 -42502
rect 71992 -42520 72494 -42168
rect 86730 -40846 87134 -40694
rect 76367 -42044 76771 -41892
rect 76295 -42177 76876 -42046
rect 71984 -42637 72485 -42524
rect 73537 -42806 73843 -42454
rect 73975 -42806 74183 -42454
rect 75660 -42551 76162 -42199
rect 82063 -41975 82467 -41823
rect 81991 -42108 82572 -41977
rect 81356 -42482 81858 -42130
rect 85731 -42006 86135 -41854
rect 85659 -42139 86240 -42008
rect 75652 -42668 76153 -42555
rect 77205 -42837 77511 -42485
rect 77643 -42837 77851 -42485
rect 81348 -42599 81849 -42486
rect 82901 -42768 83207 -42416
rect 83339 -42768 83547 -42416
rect 85024 -42513 85526 -42161
rect 85016 -42630 85517 -42517
rect 86569 -42799 86875 -42447
rect 87007 -42799 87215 -42447
rect -18319 -43444 -17915 -43192
rect -16809 -43248 -16228 -43117
rect -18391 -43577 -17810 -43446
rect -17444 -43622 -16942 -43270
rect -6785 -43352 -6577 -43100
rect -6371 -43352 -6163 -43100
rect -6009 -43352 -5801 -43100
rect -5715 -43352 -5507 -43100
rect -5405 -43352 -5197 -43100
rect -5096 -43352 -4888 -43100
rect -4285 -43352 -4077 -43100
rect -3871 -43352 -3663 -43100
rect -3509 -43352 -3301 -43100
rect -3215 -43352 -3007 -43100
rect -2905 -43352 -2697 -43100
rect -2596 -43352 -2388 -43100
rect -1785 -43352 -1577 -43100
rect -1371 -43352 -1163 -43100
rect -1009 -43352 -801 -43100
rect -715 -43352 -507 -43100
rect -405 -43352 -197 -43100
rect -96 -43352 112 -43100
rect 715 -43352 923 -43100
rect 1129 -43352 1337 -43100
rect 1491 -43352 1699 -43100
rect 1785 -43352 1993 -43100
rect 2095 -43352 2303 -43100
rect 2404 -43352 2612 -43100
rect 3215 -43352 3423 -43100
rect 3629 -43352 3837 -43100
rect 3991 -43352 4199 -43100
rect 4285 -43352 4493 -43100
rect 4595 -43352 4803 -43100
rect 4904 -43352 5112 -43100
rect 6215 -43352 6423 -43100
rect 6629 -43352 6837 -43100
rect 6991 -43352 7199 -43100
rect 7285 -43352 7493 -43100
rect 7595 -43352 7803 -43100
rect 7904 -43352 8112 -43100
rect 41160 -43106 41959 -42972
rect 46355 -43114 47154 -42980
rect 12115 -43365 12911 -43213
rect 13031 -43260 13617 -43140
rect 13868 -43260 14454 -43140
rect 13020 -43415 13620 -43263
rect 13857 -43415 14457 -43263
rect 14815 -43365 15611 -43213
rect 15731 -43260 16317 -43140
rect 16568 -43260 17154 -43140
rect 50023 -43145 50822 -43011
rect 55553 -43080 56352 -42946
rect 59221 -43111 60020 -42977
rect 64307 -43014 65106 -42880
rect 67975 -43045 68774 -42911
rect 73460 -42997 74259 -42863
rect 77128 -43028 77927 -42894
rect 82824 -42959 83623 -42825
rect 86492 -42990 87291 -42856
rect 15720 -43415 16320 -43263
rect 16557 -43415 17157 -43263
rect -17452 -43739 -16951 -43626
rect -28876 -59450 -28698 -52197
rect -28666 -59414 -28214 -52224
rect -13776 -53605 -13176 -53453
rect -12939 -53605 -12339 -53453
rect -13773 -53728 -13187 -53608
rect -12936 -53728 -12350 -53608
rect -12230 -53655 -11434 -53503
rect -11076 -53605 -10476 -53453
rect -10239 -53605 -9639 -53453
rect -11073 -53728 -10487 -53608
rect -10236 -53728 -9650 -53608
rect -9530 -53655 -8734 -53503
rect -16272 -54064 -15473 -53930
rect -13765 -54108 -13179 -53988
rect -18669 -54364 -18265 -54212
rect -21375 -54819 -21069 -54467
rect -21065 -54820 -20759 -54468
rect -20756 -54820 -20450 -54468
rect -18741 -54497 -18160 -54366
rect -17748 -54403 -17247 -54290
rect -20245 -54820 -20037 -54568
rect -19376 -54871 -18874 -54519
rect -17740 -54759 -17238 -54407
rect -16195 -54473 -15889 -54121
rect -15757 -54473 -15549 -54121
rect -13776 -54263 -13176 -54111
rect -12938 -54213 -12142 -54061
rect -12022 -54108 -11436 -53988
rect -11065 -54108 -10479 -53988
rect -12033 -54263 -11433 -54111
rect -11076 -54263 -10476 -54111
rect -10238 -54213 -9442 -54061
rect -9322 -54108 -8736 -53988
rect -8440 -54108 -7854 -53988
rect -9333 -54263 -8733 -54111
rect -8451 -54263 -7851 -54111
rect -7429 -54347 -7221 -53995
rect -7089 -54347 -6783 -53995
rect -6082 -54137 -5874 -53885
rect -5668 -54137 -5460 -53885
rect -5306 -54137 -5098 -53885
rect -5012 -54137 -4804 -53885
rect -4702 -54137 -4494 -53885
rect -4393 -54137 -4185 -53885
rect -3582 -54137 -3374 -53885
rect -3168 -54137 -2960 -53885
rect -2806 -54137 -2598 -53885
rect -2512 -54137 -2304 -53885
rect -2202 -54137 -1994 -53885
rect -1893 -54137 -1685 -53885
rect -1082 -54137 -874 -53885
rect -668 -54137 -460 -53885
rect -306 -54137 -98 -53885
rect -12 -54137 196 -53885
rect 298 -54137 506 -53885
rect 607 -54137 815 -53885
rect 1418 -54137 1626 -53885
rect 1832 -54137 2040 -53885
rect 2194 -54137 2402 -53885
rect 2488 -54137 2696 -53885
rect 2798 -54137 3006 -53885
rect 3107 -54137 3315 -53885
rect 3918 -54137 4126 -53885
rect 4332 -54137 4540 -53885
rect 4694 -54137 4902 -53885
rect 4988 -54137 5196 -53885
rect 5298 -54137 5506 -53885
rect 5607 -54137 5815 -53885
rect 6918 -54137 7126 -53885
rect 7332 -54137 7540 -53885
rect 7694 -54137 7902 -53885
rect 7988 -54137 8196 -53885
rect 8298 -54137 8506 -53885
rect 8607 -54137 8815 -53885
rect -5642 -54325 -5056 -54205
rect -4873 -54314 -4189 -54166
rect -2373 -54314 -1689 -54166
rect 127 -54314 811 -54166
rect 2627 -54314 3311 -54166
rect 5127 -54314 5811 -54166
rect 8127 -54314 8811 -54166
rect -21363 -55077 -20037 -54960
rect -19384 -54988 -18883 -54875
rect -17105 -54912 -16524 -54781
rect -17033 -55066 -16629 -54914
rect -7505 -54538 -6706 -54404
rect -5645 -54480 -5045 -54328
rect -11283 -55040 -10484 -54906
rect 29286 -54915 29787 -54802
rect 28347 -55095 28928 -54964
rect -12759 -55379 -12258 -55266
rect -12751 -55735 -12249 -55383
rect -11206 -55449 -10900 -55097
rect -10768 -55449 -10560 -55097
rect -20611 -56273 -20207 -56121
rect -16034 -56226 -15630 -56074
rect -12116 -55888 -11535 -55757
rect -12044 -56042 -11640 -55890
rect 28419 -55349 28823 -55097
rect 29294 -55271 29796 -54919
rect 37726 -54926 38227 -54813
rect 36787 -55106 37368 -54975
rect 29929 -55424 30510 -55293
rect 36859 -55360 37263 -55108
rect 37734 -55282 38236 -54930
rect 46589 -54965 47090 -54852
rect 55787 -54931 56288 -54818
rect 64541 -54865 65042 -54752
rect 73694 -54848 74195 -54735
rect 83058 -54810 83559 -54697
rect 45650 -55145 46231 -55014
rect 30001 -55578 30405 -55426
rect 38369 -55435 38950 -55304
rect 45722 -55399 46126 -55147
rect 46597 -55321 47099 -54969
rect 54848 -55111 55429 -54980
rect -5902 -56043 -5302 -55891
rect -20683 -56406 -20102 -56275
rect -21318 -56780 -20816 -56428
rect -19545 -56755 -19239 -56403
rect -19235 -56756 -18929 -56404
rect -18926 -56756 -18620 -56404
rect -18415 -56756 -18207 -56504
rect -17616 -56555 -17212 -56303
rect -16106 -56359 -15525 -56228
rect -17688 -56688 -17107 -56557
rect -16741 -56733 -16239 -56381
rect -5891 -56166 -5305 -56046
rect -5064 -56093 -4268 -55941
rect -4159 -56043 -3559 -55891
rect -3202 -56043 -2602 -55891
rect -4148 -56166 -3562 -56046
rect -3191 -56166 -2605 -56046
rect -2364 -56093 -1568 -55941
rect -1459 -56043 -859 -55891
rect -577 -56043 23 -55891
rect 2184 -55924 2588 -55772
rect -1448 -56166 -862 -56046
rect -566 -56166 20 -56046
rect 2079 -56057 2660 -55926
rect 3789 -55926 4193 -55774
rect 3684 -56059 4265 -55928
rect 18743 -55953 19652 -55795
rect -5899 -56546 -5313 -56426
rect -5062 -56546 -4476 -56426
rect -21326 -56897 -20825 -56784
rect -16749 -56850 -16248 -56737
rect -5902 -56701 -5302 -56549
rect -5065 -56701 -4465 -56549
rect -4356 -56651 -3560 -56499
rect -3199 -56546 -2613 -56426
rect -2362 -56546 -1776 -56426
rect 353 -56488 561 -56236
rect 766 -56488 1072 -56136
rect 1075 -56488 1381 -56136
rect 1385 -56487 1691 -56135
rect 2793 -56431 3295 -56079
rect 4398 -56433 4900 -56081
rect -3202 -56701 -2602 -56549
rect -2365 -56701 -1765 -56549
rect -1656 -56651 -860 -56499
rect 2802 -56548 3303 -56435
rect 4407 -56550 4908 -56437
rect 5315 -56479 5523 -56227
rect 5728 -56479 6034 -56127
rect 6037 -56479 6343 -56127
rect 6347 -56478 6653 -56126
rect 6928 -56388 7136 -56136
rect 7342 -56388 7550 -56136
rect 7704 -56388 7912 -56136
rect 7998 -56388 8206 -56136
rect 8308 -56388 8516 -56136
rect 8617 -56388 8825 -56136
rect 18840 -56266 19244 -56014
rect 38441 -55589 38845 -55437
rect 47232 -55474 47813 -55343
rect 54920 -55365 55324 -55113
rect 55795 -55287 56297 -54935
rect 63602 -55045 64183 -54914
rect 63674 -55299 64078 -55047
rect 64549 -55221 65051 -54869
rect 72755 -55028 73336 -54897
rect 56430 -55440 57011 -55309
rect 65184 -55374 65765 -55243
rect 72827 -55282 73231 -55030
rect 73702 -55204 74204 -54852
rect 82119 -54990 82700 -54859
rect 74337 -55357 74918 -55226
rect 82191 -55244 82595 -54992
rect 83066 -55166 83568 -54814
rect 83701 -55319 84282 -55188
rect 20946 -56362 21742 -56210
rect 21851 -56312 22451 -56160
rect 22688 -56312 23288 -56160
rect 8137 -56565 8821 -56417
rect 21862 -56435 22448 -56315
rect 22699 -56435 23285 -56315
rect 23646 -56362 24442 -56210
rect 24551 -56312 25151 -56160
rect 25388 -56312 25988 -56160
rect 24562 -56435 25148 -56315
rect 25399 -56435 25985 -56315
rect 353 -56745 1679 -56628
rect 5315 -56736 6641 -56619
rect -19533 -57013 -18207 -56896
rect -11045 -57202 -10641 -57050
rect -12627 -57531 -12223 -57279
rect -11117 -57335 -10536 -57204
rect 20066 -56815 20652 -56695
rect 20948 -56815 21534 -56695
rect 20063 -56970 20663 -56818
rect 20945 -56970 21545 -56818
rect 21654 -56920 22450 -56768
rect 22691 -56815 23277 -56695
rect 23648 -56815 24234 -56695
rect 22688 -56970 23288 -56818
rect 23645 -56970 24245 -56818
rect 24354 -56920 25150 -56768
rect 25391 -56815 25977 -56695
rect 29002 -56738 29406 -56586
rect 25388 -56970 25988 -56818
rect 28930 -56871 29511 -56740
rect -12699 -57664 -12118 -57533
rect -11752 -57709 -11250 -57357
rect 28295 -57245 28797 -56893
rect 47304 -55628 47708 -55476
rect 56502 -55594 56906 -55442
rect 65256 -55528 65660 -55376
rect 74409 -55511 74813 -55359
rect 83773 -55473 84177 -55321
rect 37442 -56749 37846 -56597
rect 37370 -56882 37951 -56751
rect 28287 -57362 28788 -57249
rect -11760 -57826 -11259 -57713
rect 29840 -57531 30146 -57179
rect 30278 -57531 30486 -57179
rect 31734 -57473 31942 -57121
rect 32204 -57473 32412 -56921
rect 32427 -57473 32635 -56921
rect 32655 -57473 32961 -56921
rect 32981 -57473 33189 -57121
rect 36735 -57256 37237 -56904
rect 46305 -56788 46709 -56636
rect 46233 -56921 46814 -56790
rect 36727 -57373 37228 -57260
rect -13776 -58532 -13176 -58380
rect -12939 -58532 -12339 -58380
rect -13773 -58655 -13187 -58535
rect -12936 -58655 -12350 -58535
rect -12230 -58582 -11434 -58430
rect -11076 -58532 -10476 -58380
rect -10239 -58532 -9639 -58380
rect -11073 -58655 -10487 -58535
rect -10236 -58655 -9650 -58535
rect -9530 -58582 -8734 -58430
rect 23253 -57830 26032 -57681
rect 29763 -57722 30562 -57588
rect 31668 -57736 33193 -57523
rect 38280 -57542 38586 -57190
rect 38718 -57542 38926 -57190
rect 40174 -57484 40382 -57132
rect 40644 -57484 40852 -56932
rect 40867 -57484 41075 -56932
rect 41095 -57484 41401 -56932
rect 41421 -57484 41629 -57132
rect 45598 -57295 46100 -56943
rect 55503 -56754 55907 -56602
rect 55431 -56887 56012 -56756
rect 45590 -57412 46091 -57299
rect 38203 -57733 39002 -57599
rect 40108 -57747 41633 -57534
rect 47143 -57581 47449 -57229
rect 47581 -57581 47789 -57229
rect 49037 -57523 49245 -57171
rect 49507 -57523 49715 -56971
rect 49730 -57523 49938 -56971
rect 49958 -57523 50264 -56971
rect 50284 -57523 50492 -57171
rect 54796 -57261 55298 -56909
rect 64257 -56688 64661 -56536
rect 64185 -56821 64766 -56690
rect 54788 -57378 55289 -57265
rect 56341 -57547 56647 -57195
rect 56779 -57547 56987 -57195
rect 58235 -57489 58443 -57137
rect 58705 -57489 58913 -56937
rect 58928 -57489 59136 -56937
rect 59156 -57489 59462 -56937
rect 59482 -57489 59690 -57137
rect 63550 -57195 64052 -56843
rect 73410 -56671 73814 -56519
rect 73338 -56804 73919 -56673
rect 63542 -57312 64043 -57199
rect 65095 -57481 65401 -57129
rect 65533 -57481 65741 -57129
rect 66989 -57423 67197 -57071
rect 67459 -57423 67667 -56871
rect 67682 -57423 67890 -56871
rect 67910 -57423 68216 -56871
rect 68236 -57423 68444 -57071
rect 72703 -57178 73205 -56826
rect 82774 -56633 83178 -56481
rect 82702 -56766 83283 -56635
rect 72695 -57295 73196 -57182
rect 74248 -57464 74554 -57112
rect 74686 -57464 74894 -57112
rect 76142 -57406 76350 -57054
rect 76612 -57406 76820 -56854
rect 76835 -57406 77043 -56854
rect 77063 -57406 77369 -56854
rect 77389 -57406 77597 -57054
rect 82067 -57140 82569 -56788
rect 82059 -57257 82560 -57144
rect 83612 -57426 83918 -57074
rect 84050 -57426 84258 -57074
rect 85506 -57368 85714 -57016
rect 85976 -57368 86184 -56816
rect 86199 -57368 86407 -56816
rect 86427 -57368 86733 -56816
rect 86753 -57368 86961 -57016
rect 47066 -57772 47865 -57638
rect 48971 -57786 50496 -57573
rect 56264 -57738 57063 -57604
rect 58169 -57752 59694 -57539
rect 65018 -57672 65817 -57538
rect 66923 -57686 68448 -57473
rect 74171 -57655 74970 -57521
rect 76076 -57669 77601 -57456
rect 83535 -57617 84334 -57483
rect 85440 -57631 86965 -57418
rect 18714 -58577 19363 -58436
rect 19660 -58577 20309 -58436
rect 20611 -58510 21937 -58393
rect -5902 -58799 -5302 -58647
rect -5065 -58799 -4465 -58647
rect -16272 -59064 -15473 -58930
rect -13765 -59035 -13179 -58915
rect -17748 -59403 -17247 -59290
rect -19949 -59958 -19643 -59706
rect -19044 -59959 -18738 -59707
rect -17740 -59759 -17238 -59407
rect -16195 -59473 -15889 -59121
rect -15757 -59473 -15549 -59121
rect -13776 -59190 -13176 -59038
rect -12938 -59140 -12142 -58988
rect -12022 -59035 -11436 -58915
rect -11065 -59035 -10479 -58915
rect -12033 -59190 -11433 -59038
rect -11076 -59190 -10476 -59038
rect -10238 -59140 -9442 -58988
rect -9322 -59035 -8736 -58915
rect -8440 -59035 -7854 -58915
rect -5899 -58922 -5313 -58802
rect -5062 -58922 -4476 -58802
rect -4356 -58849 -3560 -58697
rect -3202 -58799 -2602 -58647
rect -2365 -58799 -1765 -58647
rect -3199 -58922 -2613 -58802
rect -2362 -58922 -1776 -58802
rect -1656 -58849 -860 -58697
rect 353 -58720 1679 -58603
rect 5315 -58729 6641 -58612
rect -9333 -59190 -8733 -59038
rect -8451 -59190 -7851 -59038
rect -7402 -59281 -7194 -58929
rect -7062 -59281 -6756 -58929
rect 353 -59112 561 -58860
rect -21155 -60301 -20751 -60049
rect -20070 -60154 -19421 -60013
rect -19165 -60155 -18516 -60014
rect -17105 -59912 -16524 -59781
rect -17033 -60066 -16629 -59914
rect -5891 -59302 -5305 -59182
rect -7478 -59472 -6679 -59338
rect -5902 -59457 -5302 -59305
rect -5064 -59407 -4268 -59255
rect -4148 -59302 -3562 -59182
rect -3191 -59302 -2605 -59182
rect -4159 -59457 -3559 -59305
rect -3202 -59457 -2602 -59305
rect -2364 -59407 -1568 -59255
rect -1448 -59302 -862 -59182
rect -566 -59302 20 -59182
rect 766 -59212 1072 -58860
rect 1075 -59212 1381 -58860
rect 1385 -59213 1691 -58861
rect 2802 -58913 3303 -58800
rect 4407 -58911 4908 -58798
rect 2793 -59269 3295 -58917
rect 4398 -59267 4900 -58915
rect 5315 -59121 5523 -58869
rect 5728 -59221 6034 -58869
rect 6037 -59221 6343 -58869
rect 6347 -59222 6653 -58870
rect 8137 -58931 8821 -58783
rect 18835 -58884 19141 -58632
rect 19781 -58884 20087 -58632
rect 6928 -59212 7136 -58960
rect 7342 -59212 7550 -58960
rect 7704 -59212 7912 -58960
rect 7998 -59212 8206 -58960
rect 8308 -59212 8516 -58960
rect 8617 -59212 8825 -58960
rect 20599 -59003 20905 -58651
rect 20909 -59002 21215 -58650
rect 21218 -59002 21524 -58650
rect 21729 -58902 21937 -58650
rect 22508 -58756 22716 -58504
rect 22718 -58756 22926 -58504
rect 23338 -58647 23546 -57895
rect 23738 -58647 23946 -57895
rect 24338 -58647 24546 -57895
rect 24738 -58647 24946 -57895
rect 25338 -58647 25546 -57895
rect 25738 -58647 25946 -57895
rect 29278 -58368 29779 -58255
rect 28339 -58548 28920 -58417
rect 22487 -58945 23018 -58812
rect 22461 -59068 23047 -58948
rect -1459 -59457 -859 -59305
rect -577 -59457 23 -59305
rect 2079 -59422 2660 -59291
rect 2184 -59576 2588 -59424
rect 3684 -59420 4265 -59289
rect 3789 -59574 4193 -59422
rect 22458 -59223 23058 -59071
rect 28411 -58802 28815 -58550
rect 29286 -58724 29788 -58372
rect 32946 -58399 33447 -58286
rect 37718 -58379 38219 -58266
rect 32007 -58579 32588 -58448
rect 29921 -58877 30502 -58746
rect 32079 -58833 32483 -58581
rect 32954 -58755 33456 -58403
rect 36779 -58559 37360 -58428
rect 29993 -59031 30397 -58879
rect 33589 -58908 34170 -58777
rect 36851 -58813 37255 -58561
rect 37726 -58735 38228 -58383
rect 41386 -58410 41887 -58297
rect 40447 -58590 41028 -58459
rect 38361 -58888 38942 -58757
rect 40519 -58844 40923 -58592
rect 41394 -58766 41896 -58414
rect 46581 -58418 47082 -58305
rect 45642 -58598 46223 -58467
rect 33661 -59062 34065 -58910
rect 38433 -59042 38837 -58890
rect 42029 -58919 42610 -58788
rect 45714 -58852 46118 -58600
rect 46589 -58774 47091 -58422
rect 50249 -58449 50750 -58336
rect 55779 -58384 56280 -58271
rect 49310 -58629 49891 -58498
rect -21252 -60520 -20343 -60362
rect 28994 -60191 29398 -60039
rect 28922 -60324 29503 -60193
rect 28287 -60698 28789 -60346
rect 42101 -59073 42505 -58921
rect 47224 -58927 47805 -58796
rect 49382 -58883 49786 -58631
rect 50257 -58805 50759 -58453
rect 54840 -58564 55421 -58433
rect 54912 -58818 55316 -58566
rect 55787 -58740 56289 -58388
rect 59447 -58415 59948 -58302
rect 64533 -58318 65034 -58205
rect 58508 -58595 59089 -58464
rect 32662 -60222 33066 -60070
rect 32590 -60355 33171 -60224
rect -21492 -61055 -20166 -60938
rect 11935 -60868 12535 -60716
rect 12817 -60868 13417 -60716
rect 11938 -60991 12524 -60871
rect 12820 -60991 13406 -60871
rect 13526 -60918 14322 -60766
rect 14560 -60868 15160 -60716
rect 15517 -60868 16117 -60716
rect 14563 -60991 15149 -60871
rect 15520 -60991 16106 -60871
rect 16226 -60918 17022 -60766
rect 17260 -60868 17860 -60716
rect 28279 -60815 28780 -60702
rect 17263 -60991 17849 -60871
rect 29832 -60984 30138 -60632
rect 30270 -60984 30478 -60632
rect 31955 -60729 32457 -60377
rect 37434 -60202 37838 -60050
rect 37362 -60335 37943 -60204
rect 31947 -60846 32448 -60733
rect 33500 -61015 33806 -60663
rect 33938 -61015 34146 -60663
rect 36727 -60709 37229 -60357
rect 47296 -59081 47700 -58929
rect 50892 -58958 51473 -58827
rect 56422 -58893 57003 -58762
rect 58580 -58849 58984 -58597
rect 59455 -58771 59957 -58419
rect 63594 -58498 64175 -58367
rect 63666 -58752 64070 -58500
rect 64541 -58674 65043 -58322
rect 68201 -58349 68702 -58236
rect 73686 -58301 74187 -58188
rect 67262 -58529 67843 -58398
rect 41102 -60233 41506 -60081
rect 41030 -60366 41611 -60235
rect 36719 -60826 37220 -60713
rect 38272 -60995 38578 -60643
rect 38710 -60995 38918 -60643
rect 40395 -60740 40897 -60388
rect 50964 -59112 51368 -58960
rect 56494 -59047 56898 -58895
rect 60090 -58924 60671 -58793
rect 65176 -58827 65757 -58696
rect 67334 -58783 67738 -58531
rect 68209 -58705 68711 -58353
rect 72747 -58481 73328 -58350
rect 46297 -60241 46701 -60089
rect 46225 -60374 46806 -60243
rect 40387 -60857 40888 -60744
rect 41940 -61026 42246 -60674
rect 42378 -61026 42586 -60674
rect 45590 -60748 46092 -60396
rect 60162 -59078 60566 -58926
rect 65248 -58981 65652 -58829
rect 68844 -58858 69425 -58727
rect 72819 -58735 73223 -58483
rect 73694 -58657 74196 -58305
rect 77354 -58332 77855 -58219
rect 83050 -58263 83551 -58150
rect 76415 -58512 76996 -58381
rect 74329 -58810 74910 -58679
rect 76487 -58766 76891 -58514
rect 77362 -58688 77864 -58336
rect 82111 -58443 82692 -58312
rect 82183 -58697 82587 -58445
rect 83058 -58619 83560 -58267
rect 86718 -58294 87219 -58181
rect 85779 -58474 86360 -58343
rect 49965 -60272 50369 -60120
rect 49893 -60405 50474 -60274
rect 45582 -60865 46083 -60752
rect 47135 -61034 47441 -60682
rect 47573 -61034 47781 -60682
rect 49258 -60779 49760 -60427
rect 55495 -60207 55899 -60055
rect 55423 -60340 56004 -60209
rect 49250 -60896 49751 -60783
rect -21492 -61447 -21284 -61195
rect -21079 -61547 -20773 -61195
rect -20770 -61547 -20464 -61195
rect -20460 -61548 -20154 -61196
rect -16034 -61226 -15630 -61074
rect -4873 -61182 -4189 -61034
rect -2373 -61182 -1689 -61034
rect 127 -61182 811 -61034
rect 2627 -61182 3311 -61034
rect 5127 -61182 5811 -61034
rect 8127 -61182 8811 -61034
rect 29755 -61175 30554 -61041
rect 33423 -61206 34222 -61072
rect 38195 -61186 38994 -61052
rect 50803 -61065 51109 -60713
rect 51241 -61065 51449 -60713
rect 54788 -60714 55290 -60362
rect 68916 -59012 69320 -58860
rect 74401 -58964 74805 -58812
rect 77997 -58841 78578 -58710
rect 83693 -58772 84274 -58641
rect 85851 -58728 86255 -58476
rect 86726 -58650 87228 -58298
rect 59163 -60238 59567 -60086
rect 59091 -60371 59672 -60240
rect 54780 -60831 55281 -60718
rect 56333 -61000 56639 -60648
rect 56771 -61000 56979 -60648
rect 58456 -60745 58958 -60393
rect 64249 -60141 64653 -59989
rect 64177 -60274 64758 -60143
rect 63542 -60648 64044 -60296
rect 78069 -58995 78473 -58843
rect 83765 -58926 84169 -58774
rect 87361 -58803 87942 -58672
rect 67917 -60172 68321 -60020
rect 67845 -60305 68426 -60174
rect 58448 -60862 58949 -60749
rect 60001 -61031 60307 -60679
rect 60439 -61031 60647 -60679
rect 63534 -60765 64035 -60652
rect 65087 -60934 65393 -60582
rect 65525 -60934 65733 -60582
rect 67210 -60679 67712 -60327
rect 73402 -60124 73806 -59972
rect 73330 -60257 73911 -60126
rect 67202 -60796 67703 -60683
rect 68755 -60965 69061 -60613
rect 69193 -60965 69401 -60613
rect 72695 -60631 73197 -60279
rect 87433 -58957 87837 -58805
rect 77070 -60155 77474 -60003
rect 76998 -60288 77579 -60157
rect 72687 -60748 73188 -60635
rect 74240 -60917 74546 -60565
rect 74678 -60917 74886 -60565
rect 76363 -60662 76865 -60310
rect 82766 -60086 83170 -59934
rect 82694 -60219 83275 -60088
rect 82059 -60593 82561 -60241
rect 86434 -60117 86838 -59965
rect 86362 -60250 86943 -60119
rect 76355 -60779 76856 -60666
rect 77908 -60948 78214 -60596
rect 78346 -60948 78554 -60596
rect 82051 -60710 82552 -60597
rect 83604 -60879 83910 -60527
rect 84042 -60879 84250 -60527
rect 85727 -60624 86229 -60272
rect 85719 -60741 86220 -60628
rect 87272 -60910 87578 -60558
rect 87710 -60910 87918 -60558
rect -17616 -61555 -17212 -61303
rect -16106 -61359 -15525 -61228
rect -17688 -61688 -17107 -61557
rect -16741 -61733 -16239 -61381
rect -6082 -61463 -5874 -61211
rect -5668 -61463 -5460 -61211
rect -5306 -61463 -5098 -61211
rect -5012 -61463 -4804 -61211
rect -4702 -61463 -4494 -61211
rect -4393 -61463 -4185 -61211
rect -3582 -61463 -3374 -61211
rect -3168 -61463 -2960 -61211
rect -2806 -61463 -2598 -61211
rect -2512 -61463 -2304 -61211
rect -2202 -61463 -1994 -61211
rect -1893 -61463 -1685 -61211
rect -1082 -61463 -874 -61211
rect -668 -61463 -460 -61211
rect -306 -61463 -98 -61211
rect -12 -61463 196 -61211
rect 298 -61463 506 -61211
rect 607 -61463 815 -61211
rect 1418 -61463 1626 -61211
rect 1832 -61463 2040 -61211
rect 2194 -61463 2402 -61211
rect 2488 -61463 2696 -61211
rect 2798 -61463 3006 -61211
rect 3107 -61463 3315 -61211
rect 3918 -61463 4126 -61211
rect 4332 -61463 4540 -61211
rect 4694 -61463 4902 -61211
rect 4988 -61463 5196 -61211
rect 5298 -61463 5506 -61211
rect 5607 -61463 5815 -61211
rect 6918 -61463 7126 -61211
rect 7332 -61463 7540 -61211
rect 7694 -61463 7902 -61211
rect 7988 -61463 8196 -61211
rect 8298 -61463 8506 -61211
rect 8607 -61463 8815 -61211
rect 41863 -61217 42662 -61083
rect 47058 -61225 47857 -61091
rect 12818 -61476 13614 -61324
rect 13734 -61371 14320 -61251
rect 14571 -61371 15157 -61251
rect 13723 -61526 14323 -61374
rect 14560 -61526 15160 -61374
rect 15518 -61476 16314 -61324
rect 16434 -61371 17020 -61251
rect 17271 -61371 17857 -61251
rect 50726 -61256 51525 -61122
rect 56256 -61191 57055 -61057
rect 59924 -61222 60723 -61088
rect 65010 -61125 65809 -60991
rect 68678 -61156 69477 -61022
rect 74163 -61108 74962 -60974
rect 77831 -61139 78630 -61005
rect 83527 -61070 84326 -60936
rect 87195 -61101 87994 -60967
rect 16423 -61526 17023 -61374
rect 17260 -61526 17860 -61374
rect -16749 -61850 -16248 -61737
<< locali >>
rect -12872 119700 -12759 119965
rect -11318 120322 -10061 120395
rect -11346 120273 -10061 120322
rect -11346 120183 -11179 120273
rect -11333 119933 -11194 120012
rect -11308 119882 -11225 119933
rect -11327 119833 -11225 119882
rect -11090 119907 -10991 119955
rect -11090 119873 -10825 119907
rect -12872 119694 -12630 119700
rect -12872 119660 -12347 119694
rect -11327 119781 -11261 119833
rect -11451 119778 -11261 119781
rect -11451 119777 -11150 119778
rect -12043 119743 -11150 119777
rect -11451 119736 -11150 119743
rect -12872 119653 -12630 119660
rect -12872 119458 -12759 119653
rect -12872 119452 -12640 119458
rect -12872 119418 -12347 119452
rect -12872 119411 -12640 119418
rect -12872 119262 -12759 119411
rect -12872 119256 -12641 119262
rect -12872 119222 -12347 119256
rect -12872 119215 -12641 119222
rect -12872 118549 -12759 119215
rect -11327 119359 -11150 119736
rect -11450 119354 -11150 119359
rect -12043 119320 -11150 119354
rect -11450 119314 -11150 119320
rect -11327 119283 -11150 119314
rect -11090 119711 -10991 119873
rect -11090 119677 -10825 119711
rect -11090 119515 -10991 119677
rect -10546 119613 -10460 120028
rect -10183 119885 -10061 120273
rect -10183 119763 -7542 119885
rect -10702 119579 -10460 119613
rect -10546 119548 -10460 119579
rect -7664 119686 -7542 119763
rect -11090 119481 -10825 119515
rect -10546 119487 -9992 119548
rect -11090 119319 -10991 119481
rect -10546 119417 -10460 119487
rect -10702 119383 -10460 119417
rect -11090 119285 -10825 119319
rect -11327 119164 -11133 119283
rect -11453 119158 -11133 119164
rect -12043 119124 -11133 119158
rect -11453 119119 -11133 119124
rect -11327 119113 -11133 119119
rect -11303 119108 -11133 119113
rect -11090 119108 -10991 119285
rect -10546 119243 -10460 119383
rect -11303 119102 -10991 119108
rect -11303 119068 -10624 119102
rect -11996 118614 -11910 118859
rect -11465 118908 -11366 118956
rect -11631 118874 -11366 118908
rect -11465 118712 -11366 118874
rect -11631 118678 -11366 118712
rect -11996 118580 -11754 118614
rect -11996 118549 -11910 118580
rect -12872 118488 -11910 118549
rect -11465 118516 -11366 118678
rect -12464 118106 -12403 118488
rect -11996 118418 -11910 118488
rect -11631 118482 -11366 118516
rect -11996 118384 -11754 118418
rect -11996 118244 -11910 118384
rect -11465 118320 -11366 118482
rect -11631 118286 -11366 118320
rect -11303 118906 -11041 119068
rect -10053 119178 -9992 119487
rect -7664 119211 -2527 119686
rect -10053 119098 -9964 119178
rect -11303 118872 -10624 118906
rect -11303 118710 -11041 118872
rect -11303 118676 -10624 118710
rect -11303 118666 -11041 118676
rect -11303 118665 -11104 118666
rect -11303 118295 -11150 118665
rect -10050 118808 -9964 119098
rect -10395 118774 -9964 118808
rect -10087 118773 -9964 118774
rect -12482 118099 -12403 118106
rect -12482 117809 -12421 118099
rect -12482 117775 -12061 117809
rect -12482 117774 -12369 117775
rect -12482 117657 -12421 117774
rect -11465 118109 -11366 118286
rect -11465 118103 -11351 118109
rect -11317 118106 -11150 118295
rect -11832 118069 -11351 118103
rect -11310 118069 -11150 118106
rect -11415 117907 -11351 118069
rect -11832 117873 -11351 117907
rect -11929 117592 -11875 117727
rect -11415 117711 -11351 117873
rect -11832 117677 -11351 117711
rect -11415 117667 -11351 117677
rect -11303 118009 -11150 118069
rect -10960 118325 -10861 118373
rect -10960 118291 -10595 118325
rect -10960 118129 -10861 118291
rect -10050 118599 -9964 118773
rect -10217 118513 -9964 118599
rect -10960 118095 -10595 118129
rect -10960 118009 -10861 118095
rect -10217 118031 -10131 118513
rect -11303 117933 -10861 118009
rect -10473 117997 -10131 118031
rect -11303 117899 -10595 117933
rect -11303 117837 -10861 117899
rect -11303 117667 -11150 117837
rect -10960 117737 -10861 117837
rect -10217 117835 -10131 117997
rect -10473 117801 -10131 117835
rect -10960 117703 -10595 117737
rect -11921 117572 -11881 117592
rect -11919 117294 -11883 117572
rect -13051 117158 -11883 117294
rect -13051 113719 -12915 117158
rect -12841 116032 -12728 116297
rect -11250 116932 -11184 117667
rect -10960 117655 -10861 117703
rect -10217 117661 -10131 117801
rect -9372 118738 -9211 118851
rect -7664 118839 -7542 119211
rect -7825 118835 -7542 118839
rect -8117 118801 -7542 118835
rect -9372 118737 -9094 118738
rect -9372 118703 -8805 118737
rect -9372 118701 -9094 118703
rect -9372 118411 -9211 118701
rect -7825 118796 -7542 118801
rect -7665 118642 -7542 118796
rect -7827 118639 -7542 118642
rect -8117 118605 -7542 118639
rect -7827 118599 -7542 118605
rect -9372 118377 -8605 118411
rect -9372 118374 -9095 118377
rect -9372 118283 -9211 118374
rect -7665 118418 -7542 118599
rect -7842 118411 -7542 118418
rect -8317 118377 -7542 118411
rect -7842 118368 -7542 118377
rect -9372 118281 -9096 118283
rect -9372 118247 -8605 118281
rect -9372 118246 -9096 118247
rect -9372 117528 -9211 118246
rect -7665 118292 -7542 118368
rect -7845 118281 -7542 118292
rect -8317 118247 -7542 118281
rect -7845 118242 -7542 118247
rect -7665 117688 -7542 118242
rect -7822 117686 -7542 117688
rect -8317 117652 -7542 117686
rect -7822 117650 -7542 117652
rect -9372 117491 -9207 117528
rect -9372 117490 -9096 117491
rect -9372 117456 -8805 117490
rect -9372 117454 -9096 117456
rect -9372 117378 -9207 117454
rect -9320 117030 -9207 117378
rect -7665 117491 -7542 117650
rect -7824 117490 -7542 117491
rect -8317 117456 -7542 117490
rect -7824 117453 -7542 117456
rect -11250 116866 -9788 116932
rect -11268 116596 -11155 116597
rect -9854 116596 -9788 116866
rect -11268 116530 -9788 116596
rect -11268 116513 -11155 116530
rect -11059 116239 -10960 116287
rect -12841 116026 -12599 116032
rect -12841 115992 -12316 116026
rect -11296 116113 -11230 116214
rect -11420 116110 -11230 116113
rect -11059 116205 -10794 116239
rect -11420 116109 -11119 116110
rect -12012 116075 -11119 116109
rect -11420 116068 -11119 116075
rect -12841 115985 -12599 115992
rect -12841 115790 -12728 115985
rect -12841 115784 -12609 115790
rect -12841 115750 -12316 115784
rect -12841 115743 -12609 115750
rect -12841 115594 -12728 115743
rect -12841 115588 -12610 115594
rect -12841 115554 -12316 115588
rect -12841 115547 -12610 115554
rect -12841 114881 -12728 115547
rect -11296 115691 -11119 116068
rect -11419 115686 -11119 115691
rect -12012 115652 -11119 115686
rect -11419 115646 -11119 115652
rect -11296 115615 -11119 115646
rect -11059 116043 -10960 116205
rect -11059 116009 -10794 116043
rect -11059 115847 -10960 116009
rect -10515 115945 -10429 116360
rect -10671 115911 -10429 115945
rect -10515 115880 -10429 115911
rect -11059 115813 -10794 115847
rect -10515 115819 -9961 115880
rect -11059 115651 -10960 115813
rect -10515 115749 -10429 115819
rect -10671 115715 -10429 115749
rect -11059 115617 -10794 115651
rect -11296 115496 -11102 115615
rect -11422 115490 -11102 115496
rect -12012 115456 -11102 115490
rect -11422 115451 -11102 115456
rect -11296 115445 -11102 115451
rect -11272 115440 -11102 115445
rect -11059 115440 -10960 115617
rect -10515 115575 -10429 115715
rect -11272 115434 -10960 115440
rect -11272 115400 -10593 115434
rect -11965 114946 -11879 115191
rect -11434 115240 -11335 115288
rect -11600 115206 -11335 115240
rect -11434 115044 -11335 115206
rect -11600 115010 -11335 115044
rect -11965 114912 -11723 114946
rect -11965 114881 -11879 114912
rect -12841 114820 -11879 114881
rect -11434 114848 -11335 115010
rect -12433 114438 -12372 114820
rect -11965 114750 -11879 114820
rect -11600 114814 -11335 114848
rect -11965 114716 -11723 114750
rect -11965 114576 -11879 114716
rect -11434 114652 -11335 114814
rect -11600 114618 -11335 114652
rect -11272 115238 -11010 115400
rect -10022 115510 -9961 115819
rect -10022 115430 -9933 115510
rect -11272 115204 -10593 115238
rect -11272 115042 -11010 115204
rect -11272 115008 -10593 115042
rect -11272 114998 -11010 115008
rect -11272 114997 -11073 114998
rect -11272 114627 -11119 114997
rect -10019 115140 -9933 115430
rect -10364 115106 -9933 115140
rect -10056 115105 -9933 115106
rect -12451 114431 -12372 114438
rect -12451 114141 -12390 114431
rect -12451 114107 -12030 114141
rect -12451 114106 -12338 114107
rect -12451 113989 -12390 114106
rect -11434 114441 -11335 114618
rect -11434 114435 -11320 114441
rect -11286 114438 -11119 114627
rect -11801 114401 -11320 114435
rect -11279 114401 -11119 114438
rect -11384 114239 -11320 114401
rect -11801 114205 -11320 114239
rect -11898 113924 -11844 114059
rect -11384 114043 -11320 114205
rect -11801 114009 -11320 114043
rect -11384 113999 -11320 114009
rect -11272 114341 -11119 114401
rect -10929 114657 -10830 114705
rect -10929 114623 -10564 114657
rect -10929 114461 -10830 114623
rect -10019 114931 -9933 115105
rect -10186 114845 -9933 114931
rect -10929 114427 -10564 114461
rect -10929 114341 -10830 114427
rect -10186 114363 -10100 114845
rect -11272 114265 -10830 114341
rect -10442 114329 -10100 114363
rect -11272 114231 -10564 114265
rect -11272 114169 -10830 114231
rect -11272 113999 -11119 114169
rect -10929 114069 -10830 114169
rect -10186 114167 -10100 114329
rect -10442 114133 -10100 114167
rect -10929 114035 -10564 114069
rect -10929 113987 -10830 114035
rect -10186 113993 -10100 114133
rect -11890 113904 -11850 113924
rect -16160 113695 -12915 113719
rect -11888 113695 -11852 113904
rect -9388 116917 -9207 117030
rect -7729 117203 -7612 117453
rect -7856 117086 -7612 117203
rect -9388 116040 -9275 116917
rect -7856 116621 -7739 117086
rect -7862 116523 -7736 116621
rect -7850 116295 -7756 116357
rect -7836 116222 -7784 116295
rect -7606 116247 -7507 116295
rect -9388 116034 -9146 116040
rect -9388 116000 -8863 116034
rect -7843 116121 -7777 116222
rect -7967 116118 -7777 116121
rect -7606 116213 -7341 116247
rect -7967 116117 -7666 116118
rect -8559 116083 -7666 116117
rect -7967 116076 -7666 116083
rect -9388 115993 -9146 116000
rect -9388 115798 -9275 115993
rect -9388 115792 -9156 115798
rect -9388 115758 -8863 115792
rect -9388 115751 -9156 115758
rect -9388 115602 -9275 115751
rect -9388 115596 -9157 115602
rect -9388 115562 -8863 115596
rect -9388 115555 -9157 115562
rect -9388 114889 -9275 115555
rect -7843 115699 -7666 116076
rect -7966 115694 -7666 115699
rect -8559 115660 -7666 115694
rect -7966 115654 -7666 115660
rect -7843 115623 -7666 115654
rect -7606 116051 -7507 116213
rect -7606 116017 -7341 116051
rect -7606 115855 -7507 116017
rect -7062 115953 -6976 116368
rect -7218 115919 -6976 115953
rect -7062 115888 -6976 115919
rect -7606 115821 -7341 115855
rect -7062 115827 -6508 115888
rect -7606 115659 -7507 115821
rect -7062 115757 -6976 115827
rect -7218 115723 -6976 115757
rect -7606 115625 -7341 115659
rect -7843 115504 -7649 115623
rect -7969 115498 -7649 115504
rect -8559 115464 -7649 115498
rect -7969 115459 -7649 115464
rect -7843 115453 -7649 115459
rect -7819 115448 -7649 115453
rect -7606 115448 -7507 115625
rect -7062 115583 -6976 115723
rect -7819 115442 -7507 115448
rect -7819 115408 -7140 115442
rect -8512 114954 -8426 115199
rect -7981 115248 -7882 115296
rect -8147 115214 -7882 115248
rect -7981 115052 -7882 115214
rect -8147 115018 -7882 115052
rect -8512 114920 -8270 114954
rect -8512 114889 -8426 114920
rect -9388 114828 -8426 114889
rect -7981 114856 -7882 115018
rect -8980 114446 -8919 114828
rect -8512 114758 -8426 114828
rect -8147 114822 -7882 114856
rect -8512 114724 -8270 114758
rect -8512 114584 -8426 114724
rect -7981 114660 -7882 114822
rect -8147 114626 -7882 114660
rect -7819 115246 -7557 115408
rect -6569 115518 -6508 115827
rect -6569 115438 -6480 115518
rect -7819 115212 -7140 115246
rect -7819 115050 -7557 115212
rect -7819 115016 -7140 115050
rect -7819 115006 -7557 115016
rect -7819 115005 -7620 115006
rect -7819 114635 -7666 115005
rect -6566 115303 -6480 115438
rect -6124 115303 -5618 116969
rect -6566 115148 -5618 115303
rect -6911 115114 -5618 115148
rect -6603 115113 -5618 115114
rect -6566 115092 -5618 115113
rect -8998 114439 -8919 114446
rect -8998 114149 -8937 114439
rect -8998 114115 -8577 114149
rect -8998 114114 -8885 114115
rect -8998 113997 -8937 114114
rect -7981 114449 -7882 114626
rect -7981 114443 -7867 114449
rect -7833 114446 -7666 114635
rect -8348 114409 -7867 114443
rect -7826 114409 -7666 114446
rect -7931 114247 -7867 114409
rect -8348 114213 -7867 114247
rect -8445 113932 -8391 114067
rect -7931 114051 -7867 114213
rect -8348 114017 -7867 114051
rect -7931 114007 -7867 114017
rect -7819 114349 -7666 114409
rect -7476 114665 -7377 114713
rect -7476 114631 -7111 114665
rect -7476 114469 -7377 114631
rect -6566 114939 -6480 115092
rect -6733 114853 -6480 114939
rect -7476 114435 -7111 114469
rect -7476 114349 -7377 114435
rect -6733 114371 -6647 114853
rect -7819 114273 -7377 114349
rect -6989 114337 -6647 114371
rect -7819 114239 -7111 114273
rect -7819 114077 -7377 114239
rect -6733 114175 -6647 114337
rect -6989 114141 -6647 114175
rect -7819 114043 -7111 114077
rect -7819 114007 -7377 114043
rect -7763 113995 -7377 114007
rect -8437 113912 -8397 113932
rect -16160 113583 -11852 113695
rect -16404 9325 -16268 43467
rect -16414 9112 -16236 9325
rect -16404 8556 -16268 9112
rect -16160 8555 -16024 113583
rect -13051 113559 -11852 113583
rect -11888 113376 -11852 113559
rect -8435 113493 -8399 113912
rect -14192 112579 -13954 112636
rect -8510 112579 -8216 113493
rect -14192 112285 -8216 112579
rect -14192 112236 -13954 112285
rect -12910 110336 -12797 110601
rect -11356 110958 -10099 111031
rect -11384 110909 -10099 110958
rect -11384 110819 -11217 110909
rect -11371 110569 -11232 110648
rect -11346 110518 -11263 110569
rect -11365 110469 -11263 110518
rect -11128 110543 -11029 110591
rect -11128 110509 -10863 110543
rect -12910 110330 -12668 110336
rect -12910 110296 -12385 110330
rect -11365 110417 -11299 110469
rect -11489 110414 -11299 110417
rect -11489 110413 -11188 110414
rect -12081 110379 -11188 110413
rect -11489 110372 -11188 110379
rect -12910 110289 -12668 110296
rect -12910 110094 -12797 110289
rect -12910 110088 -12678 110094
rect -12910 110054 -12385 110088
rect -12910 110047 -12678 110054
rect -12910 109898 -12797 110047
rect -12910 109892 -12679 109898
rect -12910 109858 -12385 109892
rect -12910 109851 -12679 109858
rect -12910 109185 -12797 109851
rect -11365 109995 -11188 110372
rect -11488 109990 -11188 109995
rect -12081 109956 -11188 109990
rect -11488 109950 -11188 109956
rect -11365 109919 -11188 109950
rect -11128 110347 -11029 110509
rect -11128 110313 -10863 110347
rect -11128 110151 -11029 110313
rect -10584 110249 -10498 110664
rect -10221 110521 -10099 110909
rect -7763 110521 -7421 113995
rect -6733 114001 -6647 114141
rect -10221 110399 -7421 110521
rect -10740 110215 -10498 110249
rect -10584 110184 -10498 110215
rect -11128 110117 -10863 110151
rect -10584 110123 -10030 110184
rect -11128 109955 -11029 110117
rect -10584 110053 -10498 110123
rect -10740 110019 -10498 110053
rect -11128 109921 -10863 109955
rect -11365 109800 -11171 109919
rect -11491 109794 -11171 109800
rect -12081 109760 -11171 109794
rect -11491 109755 -11171 109760
rect -11365 109749 -11171 109755
rect -11341 109744 -11171 109749
rect -11128 109744 -11029 109921
rect -10584 109879 -10498 110019
rect -11341 109738 -11029 109744
rect -11341 109704 -10662 109738
rect -12034 109250 -11948 109495
rect -11503 109544 -11404 109592
rect -11669 109510 -11404 109544
rect -11503 109348 -11404 109510
rect -11669 109314 -11404 109348
rect -12034 109216 -11792 109250
rect -12034 109185 -11948 109216
rect -12910 109124 -11948 109185
rect -11503 109152 -11404 109314
rect -12502 108742 -12441 109124
rect -12034 109054 -11948 109124
rect -11669 109118 -11404 109152
rect -12034 109020 -11792 109054
rect -12034 108880 -11948 109020
rect -11503 108956 -11404 109118
rect -11669 108922 -11404 108956
rect -11341 109542 -11079 109704
rect -10091 109814 -10030 110123
rect -10091 109734 -10002 109814
rect -11341 109508 -10662 109542
rect -11341 109346 -11079 109508
rect -11341 109312 -10662 109346
rect -11341 109302 -11079 109312
rect -11341 109301 -11142 109302
rect -11341 108931 -11188 109301
rect -10088 109444 -10002 109734
rect -10433 109410 -10002 109444
rect -10125 109409 -10002 109410
rect -12520 108735 -12441 108742
rect -12520 108445 -12459 108735
rect -12520 108411 -12099 108445
rect -12520 108410 -12407 108411
rect -12520 108293 -12459 108410
rect -11503 108745 -11404 108922
rect -11503 108739 -11389 108745
rect -11355 108742 -11188 108931
rect -11870 108705 -11389 108739
rect -11348 108705 -11188 108742
rect -11453 108543 -11389 108705
rect -11870 108509 -11389 108543
rect -11967 108228 -11913 108363
rect -11453 108347 -11389 108509
rect -11870 108313 -11389 108347
rect -11453 108303 -11389 108313
rect -11341 108645 -11188 108705
rect -10998 108961 -10899 109009
rect -10998 108927 -10633 108961
rect -10998 108765 -10899 108927
rect -10088 109235 -10002 109409
rect -10255 109149 -10002 109235
rect -10998 108731 -10633 108765
rect -10998 108645 -10899 108731
rect -10255 108667 -10169 109149
rect -11341 108569 -10899 108645
rect -10511 108633 -10169 108667
rect -11341 108535 -10633 108569
rect -11341 108473 -10899 108535
rect -11341 108303 -11188 108473
rect -10998 108373 -10899 108473
rect -10255 108471 -10169 108633
rect -10511 108437 -10169 108471
rect -10998 108339 -10633 108373
rect -11959 108208 -11919 108228
rect -11957 107930 -11921 108208
rect -13089 107794 -11921 107930
rect -13089 104331 -12953 107794
rect -12879 106668 -12766 106933
rect -11288 107568 -11222 108303
rect -10998 108291 -10899 108339
rect -10255 108297 -10169 108437
rect -9410 109374 -9249 109487
rect -7763 109475 -7421 110399
rect -7863 109471 -7421 109475
rect -8155 109437 -7421 109471
rect -9410 109373 -9132 109374
rect -9410 109339 -8843 109373
rect -9410 109337 -9132 109339
rect -9410 109047 -9249 109337
rect -7863 109436 -7421 109437
rect -7863 109432 -7580 109436
rect -7703 109278 -7580 109432
rect -7865 109275 -7580 109278
rect -8155 109241 -7580 109275
rect -7865 109235 -7580 109241
rect -9410 109013 -8643 109047
rect -9410 109010 -9133 109013
rect -9410 108919 -9249 109010
rect -7703 109054 -7580 109235
rect -7880 109047 -7580 109054
rect -8355 109013 -7580 109047
rect -7880 109004 -7580 109013
rect -9410 108917 -9134 108919
rect -9410 108883 -8643 108917
rect -9410 108882 -9134 108883
rect -9410 108164 -9249 108882
rect -7703 108928 -7580 109004
rect -7883 108917 -7580 108928
rect -8355 108883 -7580 108917
rect -7883 108878 -7580 108883
rect -7703 108324 -7580 108878
rect -7860 108322 -7580 108324
rect -8355 108288 -7580 108322
rect -7860 108286 -7580 108288
rect -9410 108127 -9245 108164
rect -9410 108126 -9134 108127
rect -9410 108092 -8843 108126
rect -9410 108090 -9134 108092
rect -9410 108014 -9245 108090
rect -9358 107666 -9245 108014
rect -7703 108127 -7580 108286
rect -7862 108126 -7580 108127
rect -8355 108092 -7580 108126
rect -7862 108089 -7580 108092
rect -11288 107502 -9826 107568
rect -11306 107232 -11193 107233
rect -9892 107232 -9826 107502
rect -11306 107166 -9826 107232
rect -11306 107149 -11193 107166
rect -11097 106875 -10998 106923
rect -12879 106662 -12637 106668
rect -12879 106628 -12354 106662
rect -11334 106749 -11268 106850
rect -11458 106746 -11268 106749
rect -11097 106841 -10832 106875
rect -11458 106745 -11157 106746
rect -12050 106711 -11157 106745
rect -11458 106704 -11157 106711
rect -12879 106621 -12637 106628
rect -12879 106426 -12766 106621
rect -12879 106420 -12647 106426
rect -12879 106386 -12354 106420
rect -12879 106379 -12647 106386
rect -12879 106230 -12766 106379
rect -12879 106224 -12648 106230
rect -12879 106190 -12354 106224
rect -12879 106183 -12648 106190
rect -12879 105517 -12766 106183
rect -11334 106327 -11157 106704
rect -11457 106322 -11157 106327
rect -12050 106288 -11157 106322
rect -11457 106282 -11157 106288
rect -11334 106251 -11157 106282
rect -11097 106679 -10998 106841
rect -11097 106645 -10832 106679
rect -11097 106483 -10998 106645
rect -10553 106581 -10467 106996
rect -10709 106547 -10467 106581
rect -10553 106516 -10467 106547
rect -11097 106449 -10832 106483
rect -10553 106455 -9999 106516
rect -11097 106287 -10998 106449
rect -10553 106385 -10467 106455
rect -10709 106351 -10467 106385
rect -11097 106253 -10832 106287
rect -11334 106132 -11140 106251
rect -11460 106126 -11140 106132
rect -12050 106092 -11140 106126
rect -11460 106087 -11140 106092
rect -11334 106081 -11140 106087
rect -11310 106076 -11140 106081
rect -11097 106076 -10998 106253
rect -10553 106211 -10467 106351
rect -11310 106070 -10998 106076
rect -11310 106036 -10631 106070
rect -12003 105582 -11917 105827
rect -11472 105876 -11373 105924
rect -11638 105842 -11373 105876
rect -11472 105680 -11373 105842
rect -11638 105646 -11373 105680
rect -12003 105548 -11761 105582
rect -12003 105517 -11917 105548
rect -12879 105456 -11917 105517
rect -11472 105484 -11373 105646
rect -12471 105074 -12410 105456
rect -12003 105386 -11917 105456
rect -11638 105450 -11373 105484
rect -12003 105352 -11761 105386
rect -12003 105212 -11917 105352
rect -11472 105288 -11373 105450
rect -11638 105254 -11373 105288
rect -11310 105874 -11048 106036
rect -10060 106146 -9999 106455
rect -10060 106066 -9971 106146
rect -11310 105840 -10631 105874
rect -11310 105678 -11048 105840
rect -11310 105644 -10631 105678
rect -11310 105634 -11048 105644
rect -11310 105633 -11111 105634
rect -11310 105263 -11157 105633
rect -10057 105776 -9971 106066
rect -10402 105742 -9971 105776
rect -10094 105741 -9971 105742
rect -12489 105067 -12410 105074
rect -12489 104777 -12428 105067
rect -12489 104743 -12068 104777
rect -12489 104742 -12376 104743
rect -12489 104625 -12428 104742
rect -11472 105077 -11373 105254
rect -11472 105071 -11358 105077
rect -11324 105074 -11157 105263
rect -11839 105037 -11358 105071
rect -11317 105037 -11157 105074
rect -11422 104875 -11358 105037
rect -11839 104841 -11358 104875
rect -11936 104560 -11882 104695
rect -11422 104679 -11358 104841
rect -11839 104645 -11358 104679
rect -11422 104635 -11358 104645
rect -11310 104977 -11157 105037
rect -10967 105293 -10868 105341
rect -10967 105259 -10602 105293
rect -10967 105097 -10868 105259
rect -10057 105567 -9971 105741
rect -10224 105481 -9971 105567
rect -10967 105063 -10602 105097
rect -10967 104977 -10868 105063
rect -10224 104999 -10138 105481
rect -11310 104901 -10868 104977
rect -10480 104965 -10138 104999
rect -11310 104867 -10602 104901
rect -11310 104805 -10868 104867
rect -11310 104635 -11157 104805
rect -10967 104705 -10868 104805
rect -10224 104803 -10138 104965
rect -10480 104769 -10138 104803
rect -10967 104671 -10602 104705
rect -10967 104623 -10868 104671
rect -10224 104629 -10138 104769
rect -11928 104540 -11888 104560
rect -11926 104331 -11890 104540
rect -9426 107553 -9245 107666
rect -7767 107839 -7650 108089
rect -7894 107722 -7650 107839
rect -9426 106676 -9313 107553
rect -7894 107257 -7777 107722
rect -7900 107159 -7774 107257
rect -7888 106931 -7794 106993
rect -7874 106858 -7822 106931
rect -7644 106883 -7545 106931
rect -9426 106670 -9184 106676
rect -9426 106636 -8901 106670
rect -7881 106757 -7815 106858
rect -8005 106754 -7815 106757
rect -7644 106849 -7379 106883
rect -8005 106753 -7704 106754
rect -8597 106719 -7704 106753
rect -8005 106712 -7704 106719
rect -9426 106629 -9184 106636
rect -9426 106434 -9313 106629
rect -9426 106428 -9194 106434
rect -9426 106394 -8901 106428
rect -9426 106387 -9194 106394
rect -9426 106238 -9313 106387
rect -9426 106232 -9195 106238
rect -9426 106198 -8901 106232
rect -9426 106191 -9195 106198
rect -9426 105525 -9313 106191
rect -7881 106335 -7704 106712
rect -8004 106330 -7704 106335
rect -8597 106296 -7704 106330
rect -8004 106290 -7704 106296
rect -7881 106259 -7704 106290
rect -7644 106687 -7545 106849
rect -7644 106653 -7379 106687
rect -7644 106491 -7545 106653
rect -7100 106589 -7014 107004
rect -7256 106555 -7014 106589
rect -7100 106524 -7014 106555
rect -7644 106457 -7379 106491
rect -7100 106463 -6546 106524
rect -7644 106295 -7545 106457
rect -7100 106393 -7014 106463
rect -7256 106359 -7014 106393
rect -7644 106261 -7379 106295
rect -7881 106140 -7687 106259
rect -8007 106134 -7687 106140
rect -8597 106100 -7687 106134
rect -8007 106095 -7687 106100
rect -7881 106089 -7687 106095
rect -7857 106084 -7687 106089
rect -7644 106084 -7545 106261
rect -7100 106219 -7014 106359
rect -7857 106078 -7545 106084
rect -7857 106044 -7178 106078
rect -8550 105590 -8464 105835
rect -8019 105884 -7920 105932
rect -8185 105850 -7920 105884
rect -8019 105688 -7920 105850
rect -8185 105654 -7920 105688
rect -8550 105556 -8308 105590
rect -8550 105525 -8464 105556
rect -9426 105464 -8464 105525
rect -8019 105492 -7920 105654
rect -9018 105082 -8957 105464
rect -8550 105394 -8464 105464
rect -8185 105458 -7920 105492
rect -8550 105360 -8308 105394
rect -8550 105220 -8464 105360
rect -8019 105296 -7920 105458
rect -8185 105262 -7920 105296
rect -7857 105882 -7595 106044
rect -6607 106154 -6546 106463
rect -6607 106096 -6518 106154
rect -6124 106096 -5618 115092
rect -6607 106074 -5618 106096
rect -7857 105848 -7178 105882
rect -7857 105686 -7595 105848
rect -7857 105652 -7178 105686
rect -7857 105642 -7595 105652
rect -7857 105641 -7658 105642
rect -7857 105271 -7704 105641
rect -6604 105784 -5618 106074
rect -6949 105756 -5618 105784
rect -6949 105750 -6518 105756
rect -6641 105749 -6518 105750
rect -9036 105075 -8957 105082
rect -9036 104785 -8975 105075
rect -9036 104751 -8615 104785
rect -9036 104750 -8923 104751
rect -9036 104633 -8975 104750
rect -8019 105085 -7920 105262
rect -8019 105079 -7905 105085
rect -7871 105082 -7704 105271
rect -8386 105045 -7905 105079
rect -7864 105045 -7704 105082
rect -7969 104883 -7905 105045
rect -8386 104849 -7905 104883
rect -8483 104568 -8429 104703
rect -7969 104687 -7905 104849
rect -8386 104653 -7905 104687
rect -7969 104643 -7905 104653
rect -7857 104985 -7704 105045
rect -7514 105301 -7415 105349
rect -7514 105267 -7149 105301
rect -7514 105105 -7415 105267
rect -6604 105575 -6518 105749
rect -6771 105489 -6518 105575
rect -7514 105071 -7149 105105
rect -7514 104985 -7415 105071
rect -6771 105007 -6685 105489
rect -7857 104909 -7415 104985
rect -7027 104973 -6685 105007
rect -7857 104875 -7149 104909
rect -7857 104713 -7415 104875
rect -6771 104811 -6685 104973
rect -7027 104777 -6685 104811
rect -7857 104679 -7149 104713
rect -7857 104643 -7415 104679
rect -7754 104631 -7415 104643
rect -8475 104548 -8435 104568
rect -15790 104195 -11890 104331
rect -15790 8555 -15654 104195
rect -11926 104012 -11890 104195
rect -8473 104032 -8437 104548
rect -14196 103553 -13951 103665
rect -8543 103553 -8358 104032
rect -14196 103368 -8358 103553
rect -14196 103283 -13951 103368
rect -12927 101183 -12814 101448
rect -11373 101805 -10116 101878
rect -11401 101756 -10116 101805
rect -11401 101666 -11234 101756
rect -11388 101416 -11249 101495
rect -11363 101365 -11280 101416
rect -11382 101316 -11280 101365
rect -11145 101390 -11046 101438
rect -11145 101356 -10880 101390
rect -12927 101177 -12685 101183
rect -12927 101143 -12402 101177
rect -11382 101264 -11316 101316
rect -11506 101261 -11316 101264
rect -11506 101260 -11205 101261
rect -12098 101226 -11205 101260
rect -11506 101219 -11205 101226
rect -12927 101136 -12685 101143
rect -12927 100941 -12814 101136
rect -12927 100935 -12695 100941
rect -12927 100901 -12402 100935
rect -12927 100894 -12695 100901
rect -12927 100745 -12814 100894
rect -12927 100739 -12696 100745
rect -12927 100705 -12402 100739
rect -12927 100698 -12696 100705
rect -12927 100032 -12814 100698
rect -11382 100842 -11205 101219
rect -11505 100837 -11205 100842
rect -12098 100803 -11205 100837
rect -11505 100797 -11205 100803
rect -11382 100766 -11205 100797
rect -11145 101194 -11046 101356
rect -11145 101160 -10880 101194
rect -11145 100998 -11046 101160
rect -10601 101096 -10515 101511
rect -10238 101368 -10116 101756
rect -7754 101368 -7490 104631
rect -6771 104637 -6685 104777
rect -10238 101246 -7490 101368
rect -10757 101062 -10515 101096
rect -10601 101031 -10515 101062
rect -11145 100964 -10880 100998
rect -10601 100970 -10047 101031
rect -11145 100802 -11046 100964
rect -10601 100900 -10515 100970
rect -10757 100866 -10515 100900
rect -11145 100768 -10880 100802
rect -11382 100647 -11188 100766
rect -11508 100641 -11188 100647
rect -12098 100607 -11188 100641
rect -11508 100602 -11188 100607
rect -11382 100596 -11188 100602
rect -11358 100591 -11188 100596
rect -11145 100591 -11046 100768
rect -10601 100726 -10515 100866
rect -11358 100585 -11046 100591
rect -11358 100551 -10679 100585
rect -12051 100097 -11965 100342
rect -11520 100391 -11421 100439
rect -11686 100357 -11421 100391
rect -11520 100195 -11421 100357
rect -11686 100161 -11421 100195
rect -12051 100063 -11809 100097
rect -12051 100032 -11965 100063
rect -12927 99971 -11965 100032
rect -11520 99999 -11421 100161
rect -12519 99589 -12458 99971
rect -12051 99901 -11965 99971
rect -11686 99965 -11421 99999
rect -12051 99867 -11809 99901
rect -12051 99727 -11965 99867
rect -11520 99803 -11421 99965
rect -11686 99769 -11421 99803
rect -11358 100389 -11096 100551
rect -10108 100661 -10047 100970
rect -10108 100581 -10019 100661
rect -11358 100355 -10679 100389
rect -11358 100193 -11096 100355
rect -11358 100159 -10679 100193
rect -11358 100149 -11096 100159
rect -11358 100148 -11159 100149
rect -11358 99778 -11205 100148
rect -10105 100291 -10019 100581
rect -10450 100257 -10019 100291
rect -10142 100256 -10019 100257
rect -12537 99582 -12458 99589
rect -12537 99292 -12476 99582
rect -12537 99258 -12116 99292
rect -12537 99257 -12424 99258
rect -12537 99140 -12476 99257
rect -11520 99592 -11421 99769
rect -11520 99586 -11406 99592
rect -11372 99589 -11205 99778
rect -11887 99552 -11406 99586
rect -11365 99552 -11205 99589
rect -11470 99390 -11406 99552
rect -11887 99356 -11406 99390
rect -11984 99075 -11930 99210
rect -11470 99194 -11406 99356
rect -11887 99160 -11406 99194
rect -11470 99150 -11406 99160
rect -11358 99492 -11205 99552
rect -11015 99808 -10916 99856
rect -11015 99774 -10650 99808
rect -11015 99612 -10916 99774
rect -10105 100082 -10019 100256
rect -10272 99996 -10019 100082
rect -11015 99578 -10650 99612
rect -11015 99492 -10916 99578
rect -10272 99514 -10186 99996
rect -11358 99416 -10916 99492
rect -10528 99480 -10186 99514
rect -11358 99382 -10650 99416
rect -11358 99320 -10916 99382
rect -11358 99150 -11205 99320
rect -11015 99220 -10916 99320
rect -10272 99318 -10186 99480
rect -10528 99284 -10186 99318
rect -11015 99186 -10650 99220
rect -11976 99055 -11936 99075
rect -11974 98777 -11938 99055
rect -13106 98641 -11938 98777
rect -13106 95178 -12970 98641
rect -12896 97515 -12783 97780
rect -11305 98415 -11239 99150
rect -11015 99138 -10916 99186
rect -10272 99144 -10186 99284
rect -9427 100221 -9266 100334
rect -7754 100322 -7490 101246
rect -7880 100318 -7490 100322
rect -8172 100284 -7490 100318
rect -9427 100220 -9149 100221
rect -9427 100186 -8860 100220
rect -9427 100184 -9149 100186
rect -9427 99894 -9266 100184
rect -7880 100279 -7490 100284
rect -7754 100274 -7490 100279
rect -7720 100125 -7597 100274
rect -7882 100122 -7597 100125
rect -8172 100088 -7597 100122
rect -7882 100082 -7597 100088
rect -9427 99860 -8660 99894
rect -9427 99857 -9150 99860
rect -9427 99766 -9266 99857
rect -7720 99901 -7597 100082
rect -7897 99894 -7597 99901
rect -8372 99860 -7597 99894
rect -7897 99851 -7597 99860
rect -9427 99764 -9151 99766
rect -9427 99730 -8660 99764
rect -9427 99729 -9151 99730
rect -9427 99011 -9266 99729
rect -7720 99775 -7597 99851
rect -7900 99764 -7597 99775
rect -8372 99730 -7597 99764
rect -7900 99725 -7597 99730
rect -7720 99171 -7597 99725
rect -7877 99169 -7597 99171
rect -8372 99135 -7597 99169
rect -7877 99133 -7597 99135
rect -9427 98974 -9262 99011
rect -9427 98973 -9151 98974
rect -9427 98939 -8860 98973
rect -9427 98937 -9151 98939
rect -9427 98861 -9262 98937
rect -9375 98513 -9262 98861
rect -7720 98974 -7597 99133
rect -7879 98973 -7597 98974
rect -8372 98939 -7597 98973
rect -7879 98936 -7597 98939
rect -11305 98349 -9843 98415
rect -11323 98079 -11210 98080
rect -9909 98079 -9843 98349
rect -11323 98013 -9843 98079
rect -11323 97996 -11210 98013
rect -11114 97722 -11015 97770
rect -12896 97509 -12654 97515
rect -12896 97475 -12371 97509
rect -11351 97596 -11285 97697
rect -11475 97593 -11285 97596
rect -11114 97688 -10849 97722
rect -11475 97592 -11174 97593
rect -12067 97558 -11174 97592
rect -11475 97551 -11174 97558
rect -12896 97468 -12654 97475
rect -12896 97273 -12783 97468
rect -12896 97267 -12664 97273
rect -12896 97233 -12371 97267
rect -12896 97226 -12664 97233
rect -12896 97077 -12783 97226
rect -12896 97071 -12665 97077
rect -12896 97037 -12371 97071
rect -12896 97030 -12665 97037
rect -12896 96364 -12783 97030
rect -11351 97174 -11174 97551
rect -11474 97169 -11174 97174
rect -12067 97135 -11174 97169
rect -11474 97129 -11174 97135
rect -11351 97098 -11174 97129
rect -11114 97526 -11015 97688
rect -11114 97492 -10849 97526
rect -11114 97330 -11015 97492
rect -10570 97428 -10484 97843
rect -10726 97394 -10484 97428
rect -10570 97363 -10484 97394
rect -11114 97296 -10849 97330
rect -10570 97302 -10016 97363
rect -11114 97134 -11015 97296
rect -10570 97232 -10484 97302
rect -10726 97198 -10484 97232
rect -11114 97100 -10849 97134
rect -11351 96979 -11157 97098
rect -11477 96973 -11157 96979
rect -12067 96939 -11157 96973
rect -11477 96934 -11157 96939
rect -11351 96928 -11157 96934
rect -11327 96923 -11157 96928
rect -11114 96923 -11015 97100
rect -10570 97058 -10484 97198
rect -11327 96917 -11015 96923
rect -11327 96883 -10648 96917
rect -12020 96429 -11934 96674
rect -11489 96723 -11390 96771
rect -11655 96689 -11390 96723
rect -11489 96527 -11390 96689
rect -11655 96493 -11390 96527
rect -12020 96395 -11778 96429
rect -12020 96364 -11934 96395
rect -12896 96303 -11934 96364
rect -11489 96331 -11390 96493
rect -12488 95921 -12427 96303
rect -12020 96233 -11934 96303
rect -11655 96297 -11390 96331
rect -12020 96199 -11778 96233
rect -12020 96059 -11934 96199
rect -11489 96135 -11390 96297
rect -11655 96101 -11390 96135
rect -11327 96721 -11065 96883
rect -10077 96993 -10016 97302
rect -10077 96913 -9988 96993
rect -11327 96687 -10648 96721
rect -11327 96525 -11065 96687
rect -11327 96491 -10648 96525
rect -11327 96481 -11065 96491
rect -11327 96480 -11128 96481
rect -11327 96110 -11174 96480
rect -10074 96623 -9988 96913
rect -10419 96589 -9988 96623
rect -10111 96588 -9988 96589
rect -12506 95914 -12427 95921
rect -12506 95624 -12445 95914
rect -12506 95590 -12085 95624
rect -12506 95589 -12393 95590
rect -12506 95472 -12445 95589
rect -11489 95924 -11390 96101
rect -11489 95918 -11375 95924
rect -11341 95921 -11174 96110
rect -11856 95884 -11375 95918
rect -11334 95884 -11174 95921
rect -11439 95722 -11375 95884
rect -11856 95688 -11375 95722
rect -11953 95407 -11899 95542
rect -11439 95526 -11375 95688
rect -11856 95492 -11375 95526
rect -11439 95482 -11375 95492
rect -11327 95824 -11174 95884
rect -10984 96140 -10885 96188
rect -10984 96106 -10619 96140
rect -10984 95944 -10885 96106
rect -10074 96414 -9988 96588
rect -10241 96328 -9988 96414
rect -10984 95910 -10619 95944
rect -10984 95824 -10885 95910
rect -10241 95846 -10155 96328
rect -11327 95748 -10885 95824
rect -10497 95812 -10155 95846
rect -11327 95714 -10619 95748
rect -11327 95652 -10885 95714
rect -11327 95482 -11174 95652
rect -10984 95552 -10885 95652
rect -10241 95650 -10155 95812
rect -10497 95616 -10155 95650
rect -10984 95518 -10619 95552
rect -10984 95470 -10885 95518
rect -10241 95476 -10155 95616
rect -11945 95387 -11905 95407
rect -11943 95178 -11907 95387
rect -9443 98400 -9262 98513
rect -7784 98686 -7667 98936
rect -7911 98569 -7667 98686
rect -9443 97523 -9330 98400
rect -7911 98104 -7794 98569
rect -7917 98006 -7791 98104
rect -7905 97778 -7811 97840
rect -7891 97705 -7839 97778
rect -7661 97730 -7562 97778
rect -9443 97517 -9201 97523
rect -9443 97483 -8918 97517
rect -7898 97604 -7832 97705
rect -8022 97601 -7832 97604
rect -7661 97696 -7396 97730
rect -8022 97600 -7721 97601
rect -8614 97566 -7721 97600
rect -8022 97559 -7721 97566
rect -9443 97476 -9201 97483
rect -9443 97281 -9330 97476
rect -9443 97275 -9211 97281
rect -9443 97241 -8918 97275
rect -9443 97234 -9211 97241
rect -9443 97085 -9330 97234
rect -9443 97079 -9212 97085
rect -9443 97045 -8918 97079
rect -9443 97038 -9212 97045
rect -9443 96372 -9330 97038
rect -7898 97182 -7721 97559
rect -8021 97177 -7721 97182
rect -8614 97143 -7721 97177
rect -8021 97137 -7721 97143
rect -7898 97106 -7721 97137
rect -7661 97534 -7562 97696
rect -7661 97500 -7396 97534
rect -7661 97338 -7562 97500
rect -7117 97436 -7031 97851
rect -7273 97402 -7031 97436
rect -7117 97371 -7031 97402
rect -7661 97304 -7396 97338
rect -7117 97310 -6563 97371
rect -7661 97142 -7562 97304
rect -7117 97240 -7031 97310
rect -7273 97206 -7031 97240
rect -7661 97108 -7396 97142
rect -7898 96987 -7704 97106
rect -8024 96981 -7704 96987
rect -8614 96947 -7704 96981
rect -8024 96942 -7704 96947
rect -7898 96936 -7704 96942
rect -7874 96931 -7704 96936
rect -7661 96931 -7562 97108
rect -7117 97066 -7031 97206
rect -7874 96925 -7562 96931
rect -7874 96891 -7195 96925
rect -8567 96437 -8481 96682
rect -8036 96731 -7937 96779
rect -8202 96697 -7937 96731
rect -8036 96535 -7937 96697
rect -8202 96501 -7937 96535
rect -8567 96403 -8325 96437
rect -8567 96372 -8481 96403
rect -9443 96311 -8481 96372
rect -8036 96339 -7937 96501
rect -9035 95929 -8974 96311
rect -8567 96241 -8481 96311
rect -8202 96305 -7937 96339
rect -8567 96207 -8325 96241
rect -8567 96067 -8481 96207
rect -8036 96143 -7937 96305
rect -8202 96109 -7937 96143
rect -7874 96729 -7612 96891
rect -6624 97001 -6563 97310
rect -6624 96957 -6535 97001
rect -6124 96957 -5618 105756
rect -6624 96921 -5618 96957
rect -7874 96695 -7195 96729
rect -7874 96533 -7612 96695
rect -7874 96499 -7195 96533
rect -7874 96489 -7612 96499
rect -7874 96488 -7675 96489
rect -7874 96118 -7721 96488
rect -6621 96650 -5618 96921
rect -6621 96631 -6535 96650
rect -6966 96597 -6535 96631
rect -6658 96596 -6535 96597
rect -9053 95922 -8974 95929
rect -9053 95632 -8992 95922
rect -9053 95598 -8632 95632
rect -9053 95597 -8940 95598
rect -9053 95480 -8992 95597
rect -8036 95932 -7937 96109
rect -8036 95926 -7922 95932
rect -7888 95929 -7721 96118
rect -8403 95892 -7922 95926
rect -7881 95892 -7721 95929
rect -7986 95730 -7922 95892
rect -8403 95696 -7922 95730
rect -8500 95415 -8446 95550
rect -7986 95534 -7922 95696
rect -8403 95500 -7922 95534
rect -7986 95490 -7922 95500
rect -7874 95832 -7721 95892
rect -7531 96148 -7432 96196
rect -7531 96114 -7166 96148
rect -7531 95952 -7432 96114
rect -6621 96422 -6535 96596
rect -6788 96336 -6535 96422
rect -7531 95918 -7166 95952
rect -7531 95832 -7432 95918
rect -6788 95854 -6702 96336
rect -7874 95756 -7432 95832
rect -7044 95820 -6702 95854
rect -7874 95722 -7166 95756
rect -7874 95560 -7432 95722
rect -6788 95658 -6702 95820
rect -7044 95624 -6702 95658
rect -7874 95526 -7166 95560
rect -7874 95490 -7432 95526
rect -7848 95478 -7432 95490
rect -8492 95395 -8452 95415
rect -15491 95042 -11907 95178
rect -15491 41738 -15355 95042
rect -11943 94859 -11907 95042
rect -8490 94966 -8454 95395
rect -14186 94279 -13954 94326
rect -8569 94279 -8330 94966
rect -14186 94040 -8330 94279
rect -14186 93978 -13954 94040
rect -12993 92429 -12880 92694
rect -11439 93051 -10182 93124
rect -11467 93002 -10182 93051
rect -11467 92912 -11300 93002
rect -11454 92662 -11315 92741
rect -11429 92611 -11346 92662
rect -11448 92562 -11346 92611
rect -11211 92636 -11112 92684
rect -11211 92602 -10946 92636
rect -12993 92423 -12751 92429
rect -12993 92389 -12468 92423
rect -11448 92510 -11382 92562
rect -11572 92507 -11382 92510
rect -11572 92506 -11271 92507
rect -12164 92472 -11271 92506
rect -11572 92465 -11271 92472
rect -12993 92382 -12751 92389
rect -12993 92187 -12880 92382
rect -12993 92181 -12761 92187
rect -12993 92147 -12468 92181
rect -12993 92140 -12761 92147
rect -12993 91991 -12880 92140
rect -12993 91985 -12762 91991
rect -12993 91951 -12468 91985
rect -12993 91944 -12762 91951
rect -12993 91278 -12880 91944
rect -11448 92088 -11271 92465
rect -11571 92083 -11271 92088
rect -12164 92049 -11271 92083
rect -11571 92043 -11271 92049
rect -11448 92012 -11271 92043
rect -11211 92440 -11112 92602
rect -11211 92406 -10946 92440
rect -11211 92244 -11112 92406
rect -10667 92342 -10581 92757
rect -10304 92614 -10182 93002
rect -7848 92614 -7469 95478
rect -6788 95484 -6702 95624
rect -10304 92492 -7469 92614
rect -10823 92308 -10581 92342
rect -10667 92277 -10581 92308
rect -11211 92210 -10946 92244
rect -10667 92216 -10113 92277
rect -11211 92048 -11112 92210
rect -10667 92146 -10581 92216
rect -10823 92112 -10581 92146
rect -11211 92014 -10946 92048
rect -11448 91893 -11254 92012
rect -11574 91887 -11254 91893
rect -12164 91853 -11254 91887
rect -11574 91848 -11254 91853
rect -11448 91842 -11254 91848
rect -11424 91837 -11254 91842
rect -11211 91837 -11112 92014
rect -10667 91972 -10581 92112
rect -11424 91831 -11112 91837
rect -11424 91797 -10745 91831
rect -12117 91343 -12031 91588
rect -11586 91637 -11487 91685
rect -11752 91603 -11487 91637
rect -11586 91441 -11487 91603
rect -11752 91407 -11487 91441
rect -12117 91309 -11875 91343
rect -12117 91278 -12031 91309
rect -12993 91217 -12031 91278
rect -11586 91245 -11487 91407
rect -12585 90835 -12524 91217
rect -12117 91147 -12031 91217
rect -11752 91211 -11487 91245
rect -12117 91113 -11875 91147
rect -12117 90973 -12031 91113
rect -11586 91049 -11487 91211
rect -11752 91015 -11487 91049
rect -11424 91635 -11162 91797
rect -10174 91907 -10113 92216
rect -10174 91827 -10085 91907
rect -11424 91601 -10745 91635
rect -11424 91439 -11162 91601
rect -11424 91405 -10745 91439
rect -11424 91395 -11162 91405
rect -11424 91394 -11225 91395
rect -11424 91024 -11271 91394
rect -10171 91537 -10085 91827
rect -10516 91503 -10085 91537
rect -10208 91502 -10085 91503
rect -12603 90828 -12524 90835
rect -12603 90538 -12542 90828
rect -12603 90504 -12182 90538
rect -12603 90503 -12490 90504
rect -12603 90386 -12542 90503
rect -11586 90838 -11487 91015
rect -11586 90832 -11472 90838
rect -11438 90835 -11271 91024
rect -11953 90798 -11472 90832
rect -11431 90798 -11271 90835
rect -11536 90636 -11472 90798
rect -11953 90602 -11472 90636
rect -12050 90321 -11996 90456
rect -11536 90440 -11472 90602
rect -11953 90406 -11472 90440
rect -11536 90396 -11472 90406
rect -11424 90738 -11271 90798
rect -11081 91054 -10982 91102
rect -11081 91020 -10716 91054
rect -11081 90858 -10982 91020
rect -10171 91328 -10085 91502
rect -10338 91242 -10085 91328
rect -11081 90824 -10716 90858
rect -11081 90738 -10982 90824
rect -10338 90760 -10252 91242
rect -11424 90662 -10982 90738
rect -10594 90726 -10252 90760
rect -11424 90628 -10716 90662
rect -11424 90566 -10982 90628
rect -11424 90396 -11271 90566
rect -11081 90466 -10982 90566
rect -10338 90564 -10252 90726
rect -10594 90530 -10252 90564
rect -11081 90432 -10716 90466
rect -12042 90301 -12002 90321
rect -12040 90023 -12004 90301
rect -13172 89887 -12004 90023
rect -13172 86424 -13036 89887
rect -12962 88761 -12849 89026
rect -11371 89661 -11305 90396
rect -11081 90384 -10982 90432
rect -10338 90390 -10252 90530
rect -9493 91467 -9332 91580
rect -7848 91568 -7469 92492
rect -7946 91564 -7469 91568
rect -8238 91530 -7469 91564
rect -9493 91466 -9215 91467
rect -9493 91432 -8926 91466
rect -9493 91430 -9215 91432
rect -9493 91140 -9332 91430
rect -7946 91527 -7469 91530
rect -7946 91525 -7663 91527
rect -7786 91371 -7663 91525
rect -7948 91368 -7663 91371
rect -8238 91334 -7663 91368
rect -7948 91328 -7663 91334
rect -9493 91106 -8726 91140
rect -9493 91103 -9216 91106
rect -9493 91012 -9332 91103
rect -7786 91147 -7663 91328
rect -7963 91140 -7663 91147
rect -8438 91106 -7663 91140
rect -7963 91097 -7663 91106
rect -9493 91010 -9217 91012
rect -9493 90976 -8726 91010
rect -9493 90975 -9217 90976
rect -9493 90257 -9332 90975
rect -7786 91021 -7663 91097
rect -7966 91010 -7663 91021
rect -8438 90976 -7663 91010
rect -7966 90971 -7663 90976
rect -7786 90417 -7663 90971
rect -7943 90415 -7663 90417
rect -8438 90381 -7663 90415
rect -7943 90379 -7663 90381
rect -9493 90220 -9328 90257
rect -9493 90219 -9217 90220
rect -9493 90185 -8926 90219
rect -9493 90183 -9217 90185
rect -9493 90107 -9328 90183
rect -9441 89759 -9328 90107
rect -7786 90220 -7663 90379
rect -7945 90219 -7663 90220
rect -8438 90185 -7663 90219
rect -7945 90182 -7663 90185
rect -11371 89595 -9909 89661
rect -11389 89325 -11276 89326
rect -9975 89325 -9909 89595
rect -11389 89259 -9909 89325
rect -11389 89242 -11276 89259
rect -11180 88968 -11081 89016
rect -12962 88755 -12720 88761
rect -12962 88721 -12437 88755
rect -11417 88842 -11351 88943
rect -11541 88839 -11351 88842
rect -11180 88934 -10915 88968
rect -11541 88838 -11240 88839
rect -12133 88804 -11240 88838
rect -11541 88797 -11240 88804
rect -12962 88714 -12720 88721
rect -12962 88519 -12849 88714
rect -12962 88513 -12730 88519
rect -12962 88479 -12437 88513
rect -12962 88472 -12730 88479
rect -12962 88323 -12849 88472
rect -12962 88317 -12731 88323
rect -12962 88283 -12437 88317
rect -12962 88276 -12731 88283
rect -12962 87610 -12849 88276
rect -11417 88420 -11240 88797
rect -11540 88415 -11240 88420
rect -12133 88381 -11240 88415
rect -11540 88375 -11240 88381
rect -11417 88344 -11240 88375
rect -11180 88772 -11081 88934
rect -11180 88738 -10915 88772
rect -11180 88576 -11081 88738
rect -10636 88674 -10550 89089
rect -10792 88640 -10550 88674
rect -10636 88609 -10550 88640
rect -11180 88542 -10915 88576
rect -10636 88548 -10082 88609
rect -11180 88380 -11081 88542
rect -10636 88478 -10550 88548
rect -10792 88444 -10550 88478
rect -11180 88346 -10915 88380
rect -11417 88225 -11223 88344
rect -11543 88219 -11223 88225
rect -12133 88185 -11223 88219
rect -11543 88180 -11223 88185
rect -11417 88174 -11223 88180
rect -11393 88169 -11223 88174
rect -11180 88169 -11081 88346
rect -10636 88304 -10550 88444
rect -11393 88163 -11081 88169
rect -11393 88129 -10714 88163
rect -12086 87675 -12000 87920
rect -11555 87969 -11456 88017
rect -11721 87935 -11456 87969
rect -11555 87773 -11456 87935
rect -11721 87739 -11456 87773
rect -12086 87641 -11844 87675
rect -12086 87610 -12000 87641
rect -12962 87549 -12000 87610
rect -11555 87577 -11456 87739
rect -12554 87167 -12493 87549
rect -12086 87479 -12000 87549
rect -11721 87543 -11456 87577
rect -12086 87445 -11844 87479
rect -12086 87305 -12000 87445
rect -11555 87381 -11456 87543
rect -11721 87347 -11456 87381
rect -11393 87967 -11131 88129
rect -10143 88239 -10082 88548
rect -10143 88159 -10054 88239
rect -11393 87933 -10714 87967
rect -11393 87771 -11131 87933
rect -11393 87737 -10714 87771
rect -11393 87727 -11131 87737
rect -11393 87726 -11194 87727
rect -11393 87356 -11240 87726
rect -10140 87869 -10054 88159
rect -10485 87835 -10054 87869
rect -10177 87834 -10054 87835
rect -12572 87160 -12493 87167
rect -12572 86870 -12511 87160
rect -12572 86836 -12151 86870
rect -12572 86835 -12459 86836
rect -12572 86718 -12511 86835
rect -11555 87170 -11456 87347
rect -11555 87164 -11441 87170
rect -11407 87167 -11240 87356
rect -11922 87130 -11441 87164
rect -11400 87130 -11240 87167
rect -11505 86968 -11441 87130
rect -11922 86934 -11441 86968
rect -12019 86653 -11965 86788
rect -11505 86772 -11441 86934
rect -11922 86738 -11441 86772
rect -11505 86728 -11441 86738
rect -11393 87070 -11240 87130
rect -11050 87386 -10951 87434
rect -11050 87352 -10685 87386
rect -11050 87190 -10951 87352
rect -10140 87660 -10054 87834
rect -10307 87574 -10054 87660
rect -11050 87156 -10685 87190
rect -11050 87070 -10951 87156
rect -10307 87092 -10221 87574
rect -11393 86994 -10951 87070
rect -10563 87058 -10221 87092
rect -11393 86960 -10685 86994
rect -11393 86898 -10951 86960
rect -11393 86728 -11240 86898
rect -11050 86798 -10951 86898
rect -10307 86896 -10221 87058
rect -10563 86862 -10221 86896
rect -11050 86764 -10685 86798
rect -11050 86716 -10951 86764
rect -10307 86722 -10221 86862
rect -12011 86633 -11971 86653
rect -12009 86424 -11973 86633
rect -9509 89646 -9328 89759
rect -7850 89932 -7733 90182
rect -7977 89815 -7733 89932
rect -9509 88769 -9396 89646
rect -7977 89350 -7860 89815
rect -7983 89252 -7857 89350
rect -7971 89024 -7877 89086
rect -7957 88951 -7905 89024
rect -7727 88976 -7628 89024
rect -9509 88763 -9267 88769
rect -9509 88729 -8984 88763
rect -7964 88850 -7898 88951
rect -8088 88847 -7898 88850
rect -7727 88942 -7462 88976
rect -8088 88846 -7787 88847
rect -8680 88812 -7787 88846
rect -8088 88805 -7787 88812
rect -9509 88722 -9267 88729
rect -9509 88527 -9396 88722
rect -9509 88521 -9277 88527
rect -9509 88487 -8984 88521
rect -9509 88480 -9277 88487
rect -9509 88331 -9396 88480
rect -9509 88325 -9278 88331
rect -9509 88291 -8984 88325
rect -9509 88284 -9278 88291
rect -9509 87618 -9396 88284
rect -7964 88428 -7787 88805
rect -8087 88423 -7787 88428
rect -8680 88389 -7787 88423
rect -8087 88383 -7787 88389
rect -7964 88352 -7787 88383
rect -7727 88780 -7628 88942
rect -7727 88746 -7462 88780
rect -7727 88584 -7628 88746
rect -7183 88682 -7097 89097
rect -7339 88648 -7097 88682
rect -7183 88617 -7097 88648
rect -7727 88550 -7462 88584
rect -7183 88556 -6629 88617
rect -7727 88388 -7628 88550
rect -7183 88486 -7097 88556
rect -7339 88452 -7097 88486
rect -7727 88354 -7462 88388
rect -7964 88233 -7770 88352
rect -8090 88227 -7770 88233
rect -8680 88193 -7770 88227
rect -8090 88188 -7770 88193
rect -7964 88182 -7770 88188
rect -7940 88177 -7770 88182
rect -7727 88177 -7628 88354
rect -7183 88312 -7097 88452
rect -7940 88171 -7628 88177
rect -7940 88137 -7261 88171
rect -8633 87683 -8547 87928
rect -8102 87977 -8003 88025
rect -8268 87943 -8003 87977
rect -8102 87781 -8003 87943
rect -8268 87747 -8003 87781
rect -8633 87649 -8391 87683
rect -8633 87618 -8547 87649
rect -9509 87557 -8547 87618
rect -8102 87585 -8003 87747
rect -9101 87175 -9040 87557
rect -8633 87487 -8547 87557
rect -8268 87551 -8003 87585
rect -8633 87453 -8391 87487
rect -8633 87313 -8547 87453
rect -8102 87389 -8003 87551
rect -8268 87355 -8003 87389
rect -7940 87975 -7678 88137
rect -6690 88247 -6629 88556
rect -6690 88167 -6601 88247
rect -6687 88138 -6601 88167
rect -6124 88138 -5618 96650
rect -7940 87941 -7261 87975
rect -7940 87779 -7678 87941
rect -7940 87745 -7261 87779
rect -7940 87735 -7678 87745
rect -7940 87734 -7741 87735
rect -7940 87364 -7787 87734
rect -6687 87877 -5618 88138
rect -7032 87855 -5618 87877
rect -7032 87843 -6601 87855
rect -6724 87842 -6601 87843
rect -9119 87168 -9040 87175
rect -9119 86878 -9058 87168
rect -9119 86844 -8698 86878
rect -9119 86843 -9006 86844
rect -9119 86726 -9058 86843
rect -8102 87178 -8003 87355
rect -8102 87172 -7988 87178
rect -7954 87175 -7787 87364
rect -8469 87138 -7988 87172
rect -7947 87138 -7787 87175
rect -8052 86976 -7988 87138
rect -8469 86942 -7988 86976
rect -8566 86661 -8512 86796
rect -8052 86780 -7988 86942
rect -8469 86746 -7988 86780
rect -8052 86736 -7988 86746
rect -7940 87078 -7787 87138
rect -7597 87394 -7498 87442
rect -7597 87360 -7232 87394
rect -7597 87198 -7498 87360
rect -6687 87668 -6601 87842
rect -6854 87582 -6601 87668
rect -7597 87164 -7232 87198
rect -7597 87078 -7498 87164
rect -6854 87100 -6768 87582
rect -7940 87002 -7498 87078
rect -7110 87066 -6768 87100
rect -7940 86968 -7232 87002
rect -7940 86806 -7498 86968
rect -6854 86904 -6768 87066
rect -7110 86870 -6768 86904
rect -7940 86772 -7232 86806
rect -7940 86736 -7498 86772
rect -7880 86724 -7498 86736
rect -8558 86641 -8518 86661
rect -15205 86288 -11973 86424
rect -15491 41602 -15353 41738
rect -15491 10372 -15355 41602
rect -15496 8555 -15355 10372
rect -16182 8210 -15355 8555
rect -16182 8044 -15367 8210
rect -15205 7856 -15069 86288
rect -12009 86105 -11973 86288
rect -8556 86242 -8520 86641
rect -14174 85659 -13969 85711
rect -8601 85659 -8455 86242
rect -14174 85513 -8455 85659
rect -14174 85479 -13969 85513
rect -13027 83231 -12914 83496
rect -11473 83853 -10216 83926
rect -11501 83804 -10216 83853
rect -11501 83714 -11334 83804
rect -11488 83464 -11349 83543
rect -11463 83413 -11380 83464
rect -11482 83364 -11380 83413
rect -11245 83438 -11146 83486
rect -11245 83404 -10980 83438
rect -13027 83225 -12785 83231
rect -13027 83191 -12502 83225
rect -11482 83312 -11416 83364
rect -11606 83309 -11416 83312
rect -11606 83308 -11305 83309
rect -12198 83274 -11305 83308
rect -11606 83267 -11305 83274
rect -13027 83184 -12785 83191
rect -13027 82989 -12914 83184
rect -13027 82983 -12795 82989
rect -13027 82949 -12502 82983
rect -13027 82942 -12795 82949
rect -13027 82793 -12914 82942
rect -13027 82787 -12796 82793
rect -13027 82753 -12502 82787
rect -13027 82746 -12796 82753
rect -13027 82080 -12914 82746
rect -11482 82890 -11305 83267
rect -11605 82885 -11305 82890
rect -12198 82851 -11305 82885
rect -11605 82845 -11305 82851
rect -11482 82814 -11305 82845
rect -11245 83242 -11146 83404
rect -11245 83208 -10980 83242
rect -11245 83046 -11146 83208
rect -10701 83144 -10615 83559
rect -10338 83416 -10216 83804
rect -7880 83416 -7566 86724
rect -6854 86730 -6768 86870
rect -10338 83294 -7566 83416
rect -10857 83110 -10615 83144
rect -10701 83079 -10615 83110
rect -11245 83012 -10980 83046
rect -10701 83018 -10147 83079
rect -11245 82850 -11146 83012
rect -10701 82948 -10615 83018
rect -10857 82914 -10615 82948
rect -11245 82816 -10980 82850
rect -11482 82695 -11288 82814
rect -11608 82689 -11288 82695
rect -12198 82655 -11288 82689
rect -11608 82650 -11288 82655
rect -11482 82644 -11288 82650
rect -11458 82639 -11288 82644
rect -11245 82639 -11146 82816
rect -10701 82774 -10615 82914
rect -11458 82633 -11146 82639
rect -11458 82599 -10779 82633
rect -12151 82145 -12065 82390
rect -11620 82439 -11521 82487
rect -11786 82405 -11521 82439
rect -11620 82243 -11521 82405
rect -11786 82209 -11521 82243
rect -12151 82111 -11909 82145
rect -12151 82080 -12065 82111
rect -13027 82019 -12065 82080
rect -11620 82047 -11521 82209
rect -12619 81637 -12558 82019
rect -12151 81949 -12065 82019
rect -11786 82013 -11521 82047
rect -12151 81915 -11909 81949
rect -12151 81775 -12065 81915
rect -11620 81851 -11521 82013
rect -11786 81817 -11521 81851
rect -11458 82437 -11196 82599
rect -10208 82709 -10147 83018
rect -10208 82629 -10119 82709
rect -11458 82403 -10779 82437
rect -11458 82241 -11196 82403
rect -11458 82207 -10779 82241
rect -11458 82197 -11196 82207
rect -11458 82196 -11259 82197
rect -11458 81826 -11305 82196
rect -10205 82339 -10119 82629
rect -10550 82305 -10119 82339
rect -10242 82304 -10119 82305
rect -12637 81630 -12558 81637
rect -12637 81340 -12576 81630
rect -12637 81306 -12216 81340
rect -12637 81305 -12524 81306
rect -12637 81188 -12576 81305
rect -11620 81640 -11521 81817
rect -11620 81634 -11506 81640
rect -11472 81637 -11305 81826
rect -11987 81600 -11506 81634
rect -11465 81600 -11305 81637
rect -11570 81438 -11506 81600
rect -11987 81404 -11506 81438
rect -12084 81123 -12030 81258
rect -11570 81242 -11506 81404
rect -11987 81208 -11506 81242
rect -11570 81198 -11506 81208
rect -11458 81540 -11305 81600
rect -11115 81856 -11016 81904
rect -11115 81822 -10750 81856
rect -11115 81660 -11016 81822
rect -10205 82130 -10119 82304
rect -10372 82044 -10119 82130
rect -11115 81626 -10750 81660
rect -11115 81540 -11016 81626
rect -10372 81562 -10286 82044
rect -11458 81464 -11016 81540
rect -10628 81528 -10286 81562
rect -11458 81430 -10750 81464
rect -11458 81368 -11016 81430
rect -11458 81198 -11305 81368
rect -11115 81268 -11016 81368
rect -10372 81366 -10286 81528
rect -10628 81332 -10286 81366
rect -11115 81234 -10750 81268
rect -12076 81103 -12036 81123
rect -12074 80825 -12038 81103
rect -13206 80689 -12038 80825
rect -13206 77273 -13070 80689
rect -12996 79563 -12883 79828
rect -11405 80463 -11339 81198
rect -11115 81186 -11016 81234
rect -10372 81192 -10286 81332
rect -9527 82269 -9366 82382
rect -7880 82370 -7566 83294
rect -7980 82366 -7566 82370
rect -8272 82344 -7566 82366
rect -8272 82332 -7697 82344
rect -9527 82268 -9249 82269
rect -9527 82234 -8960 82268
rect -9527 82232 -9249 82234
rect -9527 81942 -9366 82232
rect -7980 82327 -7697 82332
rect -7820 82173 -7697 82327
rect -7982 82170 -7697 82173
rect -8272 82136 -7697 82170
rect -7982 82130 -7697 82136
rect -9527 81908 -8760 81942
rect -9527 81905 -9250 81908
rect -9527 81814 -9366 81905
rect -7820 81949 -7697 82130
rect -7997 81942 -7697 81949
rect -8472 81908 -7697 81942
rect -7997 81899 -7697 81908
rect -9527 81812 -9251 81814
rect -9527 81778 -8760 81812
rect -9527 81777 -9251 81778
rect -9527 81059 -9366 81777
rect -7820 81823 -7697 81899
rect -8000 81812 -7697 81823
rect -8472 81778 -7697 81812
rect -8000 81773 -7697 81778
rect -7820 81219 -7697 81773
rect -7977 81217 -7697 81219
rect -8472 81183 -7697 81217
rect -7977 81181 -7697 81183
rect -9527 81022 -9362 81059
rect -9527 81021 -9251 81022
rect -9527 80987 -8960 81021
rect -9527 80985 -9251 80987
rect -9527 80909 -9362 80985
rect -9475 80561 -9362 80909
rect -7820 81022 -7697 81181
rect -7979 81021 -7697 81022
rect -8472 80987 -7697 81021
rect -7979 80984 -7697 80987
rect -11405 80397 -9943 80463
rect -11423 80127 -11310 80128
rect -10009 80127 -9943 80397
rect -11423 80061 -9943 80127
rect -11423 80044 -11310 80061
rect -11214 79770 -11115 79818
rect -12996 79557 -12754 79563
rect -12996 79523 -12471 79557
rect -11451 79644 -11385 79745
rect -11575 79641 -11385 79644
rect -11214 79736 -10949 79770
rect -11575 79640 -11274 79641
rect -12167 79606 -11274 79640
rect -11575 79599 -11274 79606
rect -12996 79516 -12754 79523
rect -12996 79321 -12883 79516
rect -12996 79315 -12764 79321
rect -12996 79281 -12471 79315
rect -12996 79274 -12764 79281
rect -12996 79125 -12883 79274
rect -12996 79119 -12765 79125
rect -12996 79085 -12471 79119
rect -12996 79078 -12765 79085
rect -12996 78412 -12883 79078
rect -11451 79222 -11274 79599
rect -11574 79217 -11274 79222
rect -12167 79183 -11274 79217
rect -11574 79177 -11274 79183
rect -11451 79146 -11274 79177
rect -11214 79574 -11115 79736
rect -11214 79540 -10949 79574
rect -11214 79378 -11115 79540
rect -10670 79476 -10584 79891
rect -10826 79442 -10584 79476
rect -10670 79411 -10584 79442
rect -11214 79344 -10949 79378
rect -10670 79350 -10116 79411
rect -11214 79182 -11115 79344
rect -10670 79280 -10584 79350
rect -10826 79246 -10584 79280
rect -11214 79148 -10949 79182
rect -11451 79027 -11257 79146
rect -11577 79021 -11257 79027
rect -12167 78987 -11257 79021
rect -11577 78982 -11257 78987
rect -11451 78976 -11257 78982
rect -11427 78971 -11257 78976
rect -11214 78971 -11115 79148
rect -10670 79106 -10584 79246
rect -11427 78965 -11115 78971
rect -11427 78931 -10748 78965
rect -12120 78477 -12034 78722
rect -11589 78771 -11490 78819
rect -11755 78737 -11490 78771
rect -11589 78575 -11490 78737
rect -11755 78541 -11490 78575
rect -12120 78443 -11878 78477
rect -12120 78412 -12034 78443
rect -12996 78351 -12034 78412
rect -11589 78379 -11490 78541
rect -12588 77969 -12527 78351
rect -12120 78281 -12034 78351
rect -11755 78345 -11490 78379
rect -12120 78247 -11878 78281
rect -12120 78107 -12034 78247
rect -11589 78183 -11490 78345
rect -11755 78149 -11490 78183
rect -11427 78769 -11165 78931
rect -10177 79041 -10116 79350
rect -10177 78961 -10088 79041
rect -11427 78735 -10748 78769
rect -11427 78573 -11165 78735
rect -11427 78539 -10748 78573
rect -11427 78529 -11165 78539
rect -11427 78528 -11228 78529
rect -11427 78158 -11274 78528
rect -10174 78671 -10088 78961
rect -10519 78637 -10088 78671
rect -10211 78636 -10088 78637
rect -12606 77962 -12527 77969
rect -12606 77672 -12545 77962
rect -12606 77638 -12185 77672
rect -12606 77637 -12493 77638
rect -12606 77520 -12545 77637
rect -11589 77972 -11490 78149
rect -11589 77966 -11475 77972
rect -11441 77969 -11274 78158
rect -11956 77932 -11475 77966
rect -11434 77932 -11274 77969
rect -11539 77770 -11475 77932
rect -11956 77736 -11475 77770
rect -12053 77455 -11999 77590
rect -11539 77574 -11475 77736
rect -11956 77540 -11475 77574
rect -11539 77530 -11475 77540
rect -11427 77872 -11274 77932
rect -11084 78188 -10985 78236
rect -11084 78154 -10719 78188
rect -11084 77992 -10985 78154
rect -10174 78462 -10088 78636
rect -10341 78376 -10088 78462
rect -11084 77958 -10719 77992
rect -11084 77872 -10985 77958
rect -10341 77894 -10255 78376
rect -11427 77796 -10985 77872
rect -10597 77860 -10255 77894
rect -11427 77762 -10719 77796
rect -11427 77700 -10985 77762
rect -11427 77530 -11274 77700
rect -11084 77600 -10985 77700
rect -10341 77698 -10255 77860
rect -10597 77664 -10255 77698
rect -11084 77566 -10719 77600
rect -11084 77518 -10985 77566
rect -10341 77524 -10255 77664
rect -12045 77435 -12005 77455
rect -19000 7720 -15069 7856
rect -14950 77226 -13056 77273
rect -12043 77226 -12007 77435
rect -9543 80448 -9362 80561
rect -7884 80734 -7767 80984
rect -8011 80617 -7767 80734
rect -9543 79571 -9430 80448
rect -8011 80152 -7894 80617
rect -8017 80054 -7891 80152
rect -8005 79826 -7911 79888
rect -7991 79753 -7939 79826
rect -7761 79778 -7662 79826
rect -9543 79565 -9301 79571
rect -9543 79531 -9018 79565
rect -7998 79652 -7932 79753
rect -8122 79649 -7932 79652
rect -7761 79744 -7496 79778
rect -8122 79648 -7821 79649
rect -8714 79614 -7821 79648
rect -8122 79607 -7821 79614
rect -9543 79524 -9301 79531
rect -9543 79329 -9430 79524
rect -9543 79323 -9311 79329
rect -9543 79289 -9018 79323
rect -9543 79282 -9311 79289
rect -9543 79133 -9430 79282
rect -9543 79127 -9312 79133
rect -9543 79093 -9018 79127
rect -9543 79086 -9312 79093
rect -9543 78420 -9430 79086
rect -7998 79230 -7821 79607
rect -8121 79225 -7821 79230
rect -8714 79191 -7821 79225
rect -8121 79185 -7821 79191
rect -7998 79154 -7821 79185
rect -7761 79582 -7662 79744
rect -7761 79548 -7496 79582
rect -7761 79386 -7662 79548
rect -7217 79484 -7131 79899
rect -7373 79450 -7131 79484
rect -7217 79419 -7131 79450
rect -7761 79352 -7496 79386
rect -7217 79358 -6663 79419
rect -7761 79190 -7662 79352
rect -7217 79288 -7131 79358
rect -7373 79254 -7131 79288
rect -7761 79156 -7496 79190
rect -7998 79035 -7804 79154
rect -8124 79029 -7804 79035
rect -8714 78995 -7804 79029
rect -8124 78990 -7804 78995
rect -7998 78984 -7804 78990
rect -7974 78979 -7804 78984
rect -7761 78979 -7662 79156
rect -7217 79114 -7131 79254
rect -7974 78973 -7662 78979
rect -7974 78939 -7295 78973
rect -8667 78485 -8581 78730
rect -8136 78779 -8037 78827
rect -8302 78745 -8037 78779
rect -8136 78583 -8037 78745
rect -8302 78549 -8037 78583
rect -8667 78451 -8425 78485
rect -8667 78420 -8581 78451
rect -9543 78359 -8581 78420
rect -8136 78387 -8037 78549
rect -9135 77977 -9074 78359
rect -8667 78289 -8581 78359
rect -8302 78353 -8037 78387
rect -8667 78255 -8425 78289
rect -8667 78115 -8581 78255
rect -8136 78191 -8037 78353
rect -8302 78157 -8037 78191
rect -7974 78777 -7712 78939
rect -6724 79049 -6663 79358
rect -6724 78969 -6635 79049
rect -7974 78743 -7295 78777
rect -7974 78581 -7712 78743
rect -7974 78547 -7295 78581
rect -7974 78537 -7712 78547
rect -7974 78536 -7775 78537
rect -7974 78166 -7821 78536
rect -6721 78919 -6635 78969
rect -6124 78919 -5618 87855
rect -6721 78679 -5618 78919
rect -7066 78645 -5618 78679
rect -6758 78644 -5618 78645
rect -6721 78636 -5618 78644
rect -9153 77970 -9074 77977
rect -9153 77680 -9092 77970
rect -9153 77646 -8732 77680
rect -9153 77645 -9040 77646
rect -9153 77528 -9092 77645
rect -8136 77980 -8037 78157
rect -8136 77974 -8022 77980
rect -7988 77977 -7821 78166
rect -8503 77940 -8022 77974
rect -7981 77940 -7821 77977
rect -8086 77778 -8022 77940
rect -8503 77744 -8022 77778
rect -8600 77463 -8546 77598
rect -8086 77582 -8022 77744
rect -8503 77548 -8022 77582
rect -8086 77538 -8022 77548
rect -7974 77880 -7821 77940
rect -7631 78196 -7532 78244
rect -7631 78162 -7266 78196
rect -7631 78000 -7532 78162
rect -6721 78470 -6635 78636
rect -6888 78384 -6635 78470
rect -7631 77966 -7266 78000
rect -7631 77880 -7532 77966
rect -6888 77902 -6802 78384
rect -7974 77804 -7532 77880
rect -7144 77868 -6802 77902
rect -7974 77770 -7266 77804
rect -7974 77608 -7532 77770
rect -6888 77706 -6802 77868
rect -7144 77672 -6802 77706
rect -7974 77574 -7266 77608
rect -7974 77538 -7532 77574
rect -7870 77526 -7532 77538
rect -8592 77443 -8552 77463
rect -14950 77137 -12007 77226
rect -14950 7153 -14814 77137
rect -13206 77090 -12007 77137
rect -12043 76907 -12007 77090
rect -8590 76961 -8554 77443
rect -14147 76340 -14008 76392
rect -8693 76340 -8547 76961
rect -14147 76194 -8547 76340
rect -14147 76140 -14008 76194
rect -12988 74368 -12875 74633
rect -11434 74990 -10177 75063
rect -11462 74941 -10177 74990
rect -11462 74851 -11295 74941
rect -11449 74601 -11310 74680
rect -11424 74550 -11341 74601
rect -11443 74501 -11341 74550
rect -11206 74575 -11107 74623
rect -11206 74541 -10941 74575
rect -12988 74362 -12746 74368
rect -12988 74328 -12463 74362
rect -11443 74449 -11377 74501
rect -11567 74446 -11377 74449
rect -11567 74445 -11266 74446
rect -12159 74411 -11266 74445
rect -11567 74404 -11266 74411
rect -12988 74321 -12746 74328
rect -12988 74126 -12875 74321
rect -12988 74120 -12756 74126
rect -12988 74086 -12463 74120
rect -12988 74079 -12756 74086
rect -12988 73930 -12875 74079
rect -12988 73924 -12757 73930
rect -12988 73890 -12463 73924
rect -12988 73883 -12757 73890
rect -12988 73217 -12875 73883
rect -11443 74027 -11266 74404
rect -11566 74022 -11266 74027
rect -12159 73988 -11266 74022
rect -11566 73982 -11266 73988
rect -11443 73951 -11266 73982
rect -11206 74379 -11107 74541
rect -11206 74345 -10941 74379
rect -11206 74183 -11107 74345
rect -10662 74281 -10576 74696
rect -10299 74553 -10177 74941
rect -7870 74553 -7616 77526
rect -6888 77532 -6802 77672
rect -10299 74431 -7616 74553
rect -10818 74247 -10576 74281
rect -10662 74216 -10576 74247
rect -11206 74149 -10941 74183
rect -10662 74155 -10108 74216
rect -11206 73987 -11107 74149
rect -10662 74085 -10576 74155
rect -10818 74051 -10576 74085
rect -11206 73953 -10941 73987
rect -11443 73832 -11249 73951
rect -11569 73826 -11249 73832
rect -12159 73792 -11249 73826
rect -11569 73787 -11249 73792
rect -11443 73781 -11249 73787
rect -11419 73776 -11249 73781
rect -11206 73776 -11107 73953
rect -10662 73911 -10576 74051
rect -11419 73770 -11107 73776
rect -11419 73736 -10740 73770
rect -12112 73282 -12026 73527
rect -11581 73576 -11482 73624
rect -11747 73542 -11482 73576
rect -11581 73380 -11482 73542
rect -11747 73346 -11482 73380
rect -12112 73248 -11870 73282
rect -12112 73217 -12026 73248
rect -12988 73156 -12026 73217
rect -11581 73184 -11482 73346
rect -12580 72774 -12519 73156
rect -12112 73086 -12026 73156
rect -11747 73150 -11482 73184
rect -12112 73052 -11870 73086
rect -12112 72912 -12026 73052
rect -11581 72988 -11482 73150
rect -11747 72954 -11482 72988
rect -11419 73574 -11157 73736
rect -10169 73846 -10108 74155
rect -10169 73766 -10080 73846
rect -11419 73540 -10740 73574
rect -11419 73378 -11157 73540
rect -11419 73344 -10740 73378
rect -11419 73334 -11157 73344
rect -11419 73333 -11220 73334
rect -11419 72963 -11266 73333
rect -10166 73476 -10080 73766
rect -10511 73442 -10080 73476
rect -10203 73441 -10080 73442
rect -12598 72767 -12519 72774
rect -12598 72477 -12537 72767
rect -12598 72443 -12177 72477
rect -12598 72442 -12485 72443
rect -12598 72325 -12537 72442
rect -11581 72777 -11482 72954
rect -11581 72771 -11467 72777
rect -11433 72774 -11266 72963
rect -11948 72737 -11467 72771
rect -11426 72737 -11266 72774
rect -11531 72575 -11467 72737
rect -11948 72541 -11467 72575
rect -12045 72260 -11991 72395
rect -11531 72379 -11467 72541
rect -11948 72345 -11467 72379
rect -11531 72335 -11467 72345
rect -11419 72677 -11266 72737
rect -11076 72993 -10977 73041
rect -11076 72959 -10711 72993
rect -11076 72797 -10977 72959
rect -10166 73267 -10080 73441
rect -10333 73181 -10080 73267
rect -11076 72763 -10711 72797
rect -11076 72677 -10977 72763
rect -10333 72699 -10247 73181
rect -11419 72601 -10977 72677
rect -10589 72665 -10247 72699
rect -11419 72567 -10711 72601
rect -11419 72505 -10977 72567
rect -11419 72335 -11266 72505
rect -11076 72405 -10977 72505
rect -10333 72503 -10247 72665
rect -10589 72469 -10247 72503
rect -11076 72371 -10711 72405
rect -12037 72240 -11997 72260
rect -12035 71962 -11999 72240
rect -13167 71826 -11999 71962
rect -13167 68363 -13031 71826
rect -12957 70700 -12844 70965
rect -11366 71600 -11300 72335
rect -11076 72323 -10977 72371
rect -10333 72329 -10247 72469
rect -9488 73406 -9327 73519
rect -7870 73507 -7616 74431
rect -7941 73503 -7616 73507
rect -8233 73493 -7616 73503
rect -8233 73469 -7658 73493
rect -9488 73405 -9210 73406
rect -9488 73371 -8921 73405
rect -9488 73369 -9210 73371
rect -9488 73079 -9327 73369
rect -7941 73464 -7658 73469
rect -7781 73310 -7658 73464
rect -7943 73307 -7658 73310
rect -8233 73273 -7658 73307
rect -7943 73267 -7658 73273
rect -9488 73045 -8721 73079
rect -9488 73042 -9211 73045
rect -9488 72951 -9327 73042
rect -7781 73086 -7658 73267
rect -7958 73079 -7658 73086
rect -8433 73045 -7658 73079
rect -7958 73036 -7658 73045
rect -9488 72949 -9212 72951
rect -9488 72915 -8721 72949
rect -9488 72914 -9212 72915
rect -9488 72196 -9327 72914
rect -7781 72960 -7658 73036
rect -7961 72949 -7658 72960
rect -8433 72915 -7658 72949
rect -7961 72910 -7658 72915
rect -7781 72356 -7658 72910
rect -7938 72354 -7658 72356
rect -8433 72320 -7658 72354
rect -7938 72318 -7658 72320
rect -9488 72159 -9323 72196
rect -9488 72158 -9212 72159
rect -9488 72124 -8921 72158
rect -9488 72122 -9212 72124
rect -9488 72046 -9323 72122
rect -9436 71698 -9323 72046
rect -7781 72159 -7658 72318
rect -7940 72158 -7658 72159
rect -8433 72124 -7658 72158
rect -7940 72121 -7658 72124
rect -11366 71534 -9904 71600
rect -11384 71264 -11271 71265
rect -9970 71264 -9904 71534
rect -11384 71198 -9904 71264
rect -11384 71181 -11271 71198
rect -11175 70907 -11076 70955
rect -12957 70694 -12715 70700
rect -12957 70660 -12432 70694
rect -11412 70781 -11346 70882
rect -11536 70778 -11346 70781
rect -11175 70873 -10910 70907
rect -11536 70777 -11235 70778
rect -12128 70743 -11235 70777
rect -11536 70736 -11235 70743
rect -12957 70653 -12715 70660
rect -12957 70458 -12844 70653
rect -12957 70452 -12725 70458
rect -12957 70418 -12432 70452
rect -12957 70411 -12725 70418
rect -12957 70262 -12844 70411
rect -12957 70256 -12726 70262
rect -12957 70222 -12432 70256
rect -12957 70215 -12726 70222
rect -12957 69549 -12844 70215
rect -11412 70359 -11235 70736
rect -11535 70354 -11235 70359
rect -12128 70320 -11235 70354
rect -11535 70314 -11235 70320
rect -11412 70283 -11235 70314
rect -11175 70711 -11076 70873
rect -11175 70677 -10910 70711
rect -11175 70515 -11076 70677
rect -10631 70613 -10545 71028
rect -10787 70579 -10545 70613
rect -10631 70548 -10545 70579
rect -11175 70481 -10910 70515
rect -10631 70487 -10077 70548
rect -11175 70319 -11076 70481
rect -10631 70417 -10545 70487
rect -10787 70383 -10545 70417
rect -11175 70285 -10910 70319
rect -11412 70164 -11218 70283
rect -11538 70158 -11218 70164
rect -12128 70124 -11218 70158
rect -11538 70119 -11218 70124
rect -11412 70113 -11218 70119
rect -11388 70108 -11218 70113
rect -11175 70108 -11076 70285
rect -10631 70243 -10545 70383
rect -11388 70102 -11076 70108
rect -11388 70068 -10709 70102
rect -12081 69614 -11995 69859
rect -11550 69908 -11451 69956
rect -11716 69874 -11451 69908
rect -11550 69712 -11451 69874
rect -11716 69678 -11451 69712
rect -12081 69580 -11839 69614
rect -12081 69549 -11995 69580
rect -12957 69488 -11995 69549
rect -11550 69516 -11451 69678
rect -12549 69106 -12488 69488
rect -12081 69418 -11995 69488
rect -11716 69482 -11451 69516
rect -12081 69384 -11839 69418
rect -12081 69244 -11995 69384
rect -11550 69320 -11451 69482
rect -11716 69286 -11451 69320
rect -11388 69906 -11126 70068
rect -10138 70178 -10077 70487
rect -10138 70098 -10049 70178
rect -11388 69872 -10709 69906
rect -11388 69710 -11126 69872
rect -11388 69676 -10709 69710
rect -11388 69666 -11126 69676
rect -11388 69665 -11189 69666
rect -11388 69295 -11235 69665
rect -10135 69808 -10049 70098
rect -10480 69774 -10049 69808
rect -10172 69773 -10049 69774
rect -12567 69099 -12488 69106
rect -12567 68809 -12506 69099
rect -12567 68775 -12146 68809
rect -12567 68774 -12454 68775
rect -12567 68657 -12506 68774
rect -11550 69109 -11451 69286
rect -11550 69103 -11436 69109
rect -11402 69106 -11235 69295
rect -11917 69069 -11436 69103
rect -11395 69069 -11235 69106
rect -11500 68907 -11436 69069
rect -11917 68873 -11436 68907
rect -12014 68592 -11960 68727
rect -11500 68711 -11436 68873
rect -11917 68677 -11436 68711
rect -11500 68667 -11436 68677
rect -11388 69009 -11235 69069
rect -11045 69325 -10946 69373
rect -11045 69291 -10680 69325
rect -11045 69129 -10946 69291
rect -10135 69599 -10049 69773
rect -10302 69513 -10049 69599
rect -11045 69095 -10680 69129
rect -11045 69009 -10946 69095
rect -10302 69031 -10216 69513
rect -11388 68933 -10946 69009
rect -10558 68997 -10216 69031
rect -11388 68899 -10680 68933
rect -11388 68837 -10946 68899
rect -11388 68667 -11235 68837
rect -11045 68737 -10946 68837
rect -10302 68835 -10216 68997
rect -10558 68801 -10216 68835
rect -11045 68703 -10680 68737
rect -11045 68655 -10946 68703
rect -10302 68661 -10216 68801
rect -12006 68572 -11966 68592
rect -12004 68363 -11968 68572
rect -9504 71585 -9323 71698
rect -7845 71871 -7728 72121
rect -7972 71754 -7728 71871
rect -9504 70708 -9391 71585
rect -7972 71289 -7855 71754
rect -7978 71191 -7852 71289
rect -7966 70963 -7872 71025
rect -7952 70890 -7900 70963
rect -7722 70915 -7623 70963
rect -9504 70702 -9262 70708
rect -9504 70668 -8979 70702
rect -7959 70789 -7893 70890
rect -8083 70786 -7893 70789
rect -7722 70881 -7457 70915
rect -8083 70785 -7782 70786
rect -8675 70751 -7782 70785
rect -8083 70744 -7782 70751
rect -9504 70661 -9262 70668
rect -9504 70466 -9391 70661
rect -9504 70460 -9272 70466
rect -9504 70426 -8979 70460
rect -9504 70419 -9272 70426
rect -9504 70270 -9391 70419
rect -9504 70264 -9273 70270
rect -9504 70230 -8979 70264
rect -9504 70223 -9273 70230
rect -9504 69557 -9391 70223
rect -7959 70367 -7782 70744
rect -8082 70362 -7782 70367
rect -8675 70328 -7782 70362
rect -8082 70322 -7782 70328
rect -7959 70291 -7782 70322
rect -7722 70719 -7623 70881
rect -7722 70685 -7457 70719
rect -7722 70523 -7623 70685
rect -7178 70621 -7092 71036
rect -7334 70587 -7092 70621
rect -7178 70556 -7092 70587
rect -7722 70489 -7457 70523
rect -7178 70495 -6624 70556
rect -7722 70327 -7623 70489
rect -7178 70425 -7092 70495
rect -7334 70391 -7092 70425
rect -7722 70293 -7457 70327
rect -7959 70172 -7765 70291
rect -8085 70166 -7765 70172
rect -8675 70132 -7765 70166
rect -8085 70127 -7765 70132
rect -7959 70121 -7765 70127
rect -7935 70116 -7765 70121
rect -7722 70116 -7623 70293
rect -7178 70251 -7092 70391
rect -7935 70110 -7623 70116
rect -7935 70076 -7256 70110
rect -8628 69622 -8542 69867
rect -8097 69916 -7998 69964
rect -8263 69882 -7998 69916
rect -8097 69720 -7998 69882
rect -8263 69686 -7998 69720
rect -8628 69588 -8386 69622
rect -8628 69557 -8542 69588
rect -9504 69496 -8542 69557
rect -8097 69524 -7998 69686
rect -9096 69114 -9035 69496
rect -8628 69426 -8542 69496
rect -8263 69490 -7998 69524
rect -8628 69392 -8386 69426
rect -8628 69252 -8542 69392
rect -8097 69328 -7998 69490
rect -8263 69294 -7998 69328
rect -7935 69914 -7673 70076
rect -6685 70186 -6624 70495
rect -6685 70106 -6596 70186
rect -7935 69880 -7256 69914
rect -7935 69718 -7673 69880
rect -7935 69684 -7256 69718
rect -7935 69674 -7673 69684
rect -7935 69673 -7736 69674
rect -7935 69303 -7782 69673
rect -6682 70007 -6596 70106
rect -6124 70007 -5618 78636
rect -6682 69816 -5618 70007
rect -7027 69782 -5618 69816
rect -6719 69781 -5618 69782
rect -6682 69724 -5618 69781
rect -9114 69107 -9035 69114
rect -9114 68817 -9053 69107
rect -9114 68783 -8693 68817
rect -9114 68782 -9001 68783
rect -9114 68665 -9053 68782
rect -8097 69117 -7998 69294
rect -8097 69111 -7983 69117
rect -7949 69114 -7782 69303
rect -8464 69077 -7983 69111
rect -7942 69077 -7782 69114
rect -8047 68915 -7983 69077
rect -8464 68881 -7983 68915
rect -8561 68600 -8507 68735
rect -8047 68719 -7983 68881
rect -8464 68685 -7983 68719
rect -8047 68675 -7983 68685
rect -7935 69017 -7782 69077
rect -7592 69333 -7493 69381
rect -7592 69299 -7227 69333
rect -7592 69137 -7493 69299
rect -6682 69607 -6596 69724
rect -6849 69521 -6596 69607
rect -7592 69103 -7227 69137
rect -7592 69017 -7493 69103
rect -6849 69039 -6763 69521
rect -7935 68941 -7493 69017
rect -7105 69005 -6763 69039
rect -7935 68907 -7227 68941
rect -7935 68845 -7493 68907
rect -8553 68580 -8513 68600
rect -19851 7017 -14814 7153
rect -14717 68227 -11968 68363
rect -14717 5489 -14581 68227
rect -12004 68044 -11968 68227
rect -8551 68160 -8515 68580
rect -14193 67658 -13990 67717
rect -8607 67658 -8461 68160
rect -14193 67512 -8461 67658
rect -14193 67443 -13990 67512
rect -12977 65928 -12864 66193
rect -11423 66550 -10166 66623
rect -11451 66501 -10166 66550
rect -11451 66411 -11284 66501
rect -11438 66161 -11299 66240
rect -11413 66110 -11330 66161
rect -11432 66061 -11330 66110
rect -11195 66135 -11096 66183
rect -11195 66101 -10930 66135
rect -12977 65922 -12735 65928
rect -12977 65888 -12452 65922
rect -11432 66009 -11366 66061
rect -11556 66006 -11366 66009
rect -11556 66005 -11255 66006
rect -12148 65971 -11255 66005
rect -11556 65964 -11255 65971
rect -12977 65881 -12735 65888
rect -12977 65686 -12864 65881
rect -12977 65680 -12745 65686
rect -12977 65646 -12452 65680
rect -12977 65639 -12745 65646
rect -12977 65490 -12864 65639
rect -12977 65484 -12746 65490
rect -12977 65450 -12452 65484
rect -12977 65443 -12746 65450
rect -12977 64777 -12864 65443
rect -11432 65587 -11255 65964
rect -11555 65582 -11255 65587
rect -12148 65548 -11255 65582
rect -11555 65542 -11255 65548
rect -11432 65511 -11255 65542
rect -11195 65939 -11096 66101
rect -11195 65905 -10930 65939
rect -11195 65743 -11096 65905
rect -10651 65841 -10565 66256
rect -10288 66113 -10166 66501
rect -7935 66113 -7782 68845
rect -7592 68745 -7493 68845
rect -6849 68843 -6763 69005
rect -7105 68809 -6763 68843
rect -7592 68711 -7227 68745
rect -7592 68663 -7493 68711
rect -6849 68669 -6763 68809
rect -10288 65991 -7647 66113
rect -10807 65807 -10565 65841
rect -10651 65776 -10565 65807
rect -11195 65709 -10930 65743
rect -10651 65715 -10097 65776
rect -11195 65547 -11096 65709
rect -10651 65645 -10565 65715
rect -10807 65611 -10565 65645
rect -11195 65513 -10930 65547
rect -11432 65392 -11238 65511
rect -11558 65386 -11238 65392
rect -12148 65352 -11238 65386
rect -11558 65347 -11238 65352
rect -11432 65341 -11238 65347
rect -11408 65336 -11238 65341
rect -11195 65336 -11096 65513
rect -10651 65471 -10565 65611
rect -11408 65330 -11096 65336
rect -11408 65296 -10729 65330
rect -12101 64842 -12015 65087
rect -11570 65136 -11471 65184
rect -11736 65102 -11471 65136
rect -11570 64940 -11471 65102
rect -11736 64906 -11471 64940
rect -12101 64808 -11859 64842
rect -12101 64777 -12015 64808
rect -12977 64716 -12015 64777
rect -11570 64744 -11471 64906
rect -12569 64334 -12508 64716
rect -12101 64646 -12015 64716
rect -11736 64710 -11471 64744
rect -12101 64612 -11859 64646
rect -12101 64472 -12015 64612
rect -11570 64548 -11471 64710
rect -11736 64514 -11471 64548
rect -11408 65134 -11146 65296
rect -10158 65406 -10097 65715
rect -10158 65326 -10069 65406
rect -11408 65100 -10729 65134
rect -11408 64938 -11146 65100
rect -11408 64904 -10729 64938
rect -11408 64894 -11146 64904
rect -11408 64893 -11209 64894
rect -11408 64523 -11255 64893
rect -10155 65036 -10069 65326
rect -10500 65002 -10069 65036
rect -10192 65001 -10069 65002
rect -12587 64327 -12508 64334
rect -12587 64037 -12526 64327
rect -12587 64003 -12166 64037
rect -12587 64002 -12474 64003
rect -12587 63885 -12526 64002
rect -11570 64337 -11471 64514
rect -11570 64331 -11456 64337
rect -11422 64334 -11255 64523
rect -11937 64297 -11456 64331
rect -11415 64297 -11255 64334
rect -11520 64135 -11456 64297
rect -11937 64101 -11456 64135
rect -12034 63820 -11980 63955
rect -11520 63939 -11456 64101
rect -11937 63905 -11456 63939
rect -11520 63895 -11456 63905
rect -11408 64237 -11255 64297
rect -11065 64553 -10966 64601
rect -11065 64519 -10700 64553
rect -11065 64357 -10966 64519
rect -10155 64827 -10069 65001
rect -10322 64741 -10069 64827
rect -11065 64323 -10700 64357
rect -11065 64237 -10966 64323
rect -10322 64259 -10236 64741
rect -11408 64161 -10966 64237
rect -10578 64225 -10236 64259
rect -11408 64127 -10700 64161
rect -11408 64065 -10966 64127
rect -11408 63895 -11255 64065
rect -11065 63965 -10966 64065
rect -10322 64063 -10236 64225
rect -10578 64029 -10236 64063
rect -11065 63931 -10700 63965
rect -12026 63800 -11986 63820
rect -12024 63522 -11988 63800
rect -13156 63386 -11988 63522
rect -13156 59923 -13020 63386
rect -12946 62260 -12833 62525
rect -11355 63160 -11289 63895
rect -11065 63883 -10966 63931
rect -10322 63889 -10236 64029
rect -9477 64966 -9316 65079
rect -7769 65067 -7647 65991
rect -7930 65063 -7647 65067
rect -8222 65029 -7647 65063
rect -9477 64965 -9199 64966
rect -9477 64931 -8910 64965
rect -9477 64929 -9199 64931
rect -9477 64639 -9316 64929
rect -7930 65024 -7647 65029
rect -7770 64870 -7647 65024
rect -7932 64867 -7647 64870
rect -8222 64833 -7647 64867
rect -7932 64827 -7647 64833
rect -9477 64605 -8710 64639
rect -9477 64602 -9200 64605
rect -9477 64511 -9316 64602
rect -7770 64646 -7647 64827
rect -7947 64639 -7647 64646
rect -8422 64605 -7647 64639
rect -7947 64596 -7647 64605
rect -9477 64509 -9201 64511
rect -9477 64475 -8710 64509
rect -9477 64474 -9201 64475
rect -9477 63756 -9316 64474
rect -7770 64520 -7647 64596
rect -7950 64509 -7647 64520
rect -8422 64475 -7647 64509
rect -7950 64470 -7647 64475
rect -7770 63916 -7647 64470
rect -7927 63914 -7647 63916
rect -8422 63880 -7647 63914
rect -7927 63878 -7647 63880
rect -9477 63719 -9312 63756
rect -9477 63718 -9201 63719
rect -9477 63684 -8910 63718
rect -9477 63682 -9201 63684
rect -9477 63606 -9312 63682
rect -9425 63258 -9312 63606
rect -7770 63719 -7647 63878
rect -7929 63718 -7647 63719
rect -8422 63684 -7647 63718
rect -7929 63681 -7647 63684
rect -11355 63094 -9893 63160
rect -11373 62824 -11260 62825
rect -9959 62824 -9893 63094
rect -11373 62758 -9893 62824
rect -11373 62741 -11260 62758
rect -11164 62467 -11065 62515
rect -12946 62254 -12704 62260
rect -12946 62220 -12421 62254
rect -11401 62341 -11335 62442
rect -11525 62338 -11335 62341
rect -11164 62433 -10899 62467
rect -11525 62337 -11224 62338
rect -12117 62303 -11224 62337
rect -11525 62296 -11224 62303
rect -12946 62213 -12704 62220
rect -12946 62018 -12833 62213
rect -12946 62012 -12714 62018
rect -12946 61978 -12421 62012
rect -12946 61971 -12714 61978
rect -12946 61822 -12833 61971
rect -12946 61816 -12715 61822
rect -12946 61782 -12421 61816
rect -12946 61775 -12715 61782
rect -12946 61109 -12833 61775
rect -11401 61919 -11224 62296
rect -11524 61914 -11224 61919
rect -12117 61880 -11224 61914
rect -11524 61874 -11224 61880
rect -11401 61843 -11224 61874
rect -11164 62271 -11065 62433
rect -11164 62237 -10899 62271
rect -11164 62075 -11065 62237
rect -10620 62173 -10534 62588
rect -10776 62139 -10534 62173
rect -10620 62108 -10534 62139
rect -11164 62041 -10899 62075
rect -10620 62047 -10066 62108
rect -11164 61879 -11065 62041
rect -10620 61977 -10534 62047
rect -10776 61943 -10534 61977
rect -11164 61845 -10899 61879
rect -11401 61724 -11207 61843
rect -11527 61718 -11207 61724
rect -12117 61684 -11207 61718
rect -11527 61679 -11207 61684
rect -11401 61673 -11207 61679
rect -11377 61668 -11207 61673
rect -11164 61668 -11065 61845
rect -10620 61803 -10534 61943
rect -11377 61662 -11065 61668
rect -11377 61628 -10698 61662
rect -12070 61174 -11984 61419
rect -11539 61468 -11440 61516
rect -11705 61434 -11440 61468
rect -11539 61272 -11440 61434
rect -11705 61238 -11440 61272
rect -12070 61140 -11828 61174
rect -12070 61109 -11984 61140
rect -12946 61048 -11984 61109
rect -11539 61076 -11440 61238
rect -12538 60666 -12477 61048
rect -12070 60978 -11984 61048
rect -11705 61042 -11440 61076
rect -12070 60944 -11828 60978
rect -12070 60804 -11984 60944
rect -11539 60880 -11440 61042
rect -11705 60846 -11440 60880
rect -11377 61466 -11115 61628
rect -10127 61738 -10066 62047
rect -10127 61658 -10038 61738
rect -11377 61432 -10698 61466
rect -11377 61270 -11115 61432
rect -11377 61236 -10698 61270
rect -11377 61226 -11115 61236
rect -11377 61225 -11178 61226
rect -11377 60855 -11224 61225
rect -10124 61368 -10038 61658
rect -10469 61334 -10038 61368
rect -10161 61333 -10038 61334
rect -12556 60659 -12477 60666
rect -12556 60369 -12495 60659
rect -12556 60335 -12135 60369
rect -12556 60334 -12443 60335
rect -12556 60217 -12495 60334
rect -11539 60669 -11440 60846
rect -11539 60663 -11425 60669
rect -11391 60666 -11224 60855
rect -11906 60629 -11425 60663
rect -11384 60629 -11224 60666
rect -11489 60467 -11425 60629
rect -11906 60433 -11425 60467
rect -12003 60152 -11949 60287
rect -11489 60271 -11425 60433
rect -11906 60237 -11425 60271
rect -11489 60227 -11425 60237
rect -11377 60569 -11224 60629
rect -11034 60885 -10935 60933
rect -11034 60851 -10669 60885
rect -11034 60689 -10935 60851
rect -10124 61159 -10038 61333
rect -10291 61073 -10038 61159
rect -11034 60655 -10669 60689
rect -11034 60569 -10935 60655
rect -10291 60591 -10205 61073
rect -11377 60493 -10935 60569
rect -10547 60557 -10205 60591
rect -11377 60459 -10669 60493
rect -11377 60397 -10935 60459
rect -11377 60227 -11224 60397
rect -11034 60297 -10935 60397
rect -10291 60395 -10205 60557
rect -10547 60361 -10205 60395
rect -11034 60263 -10669 60297
rect -11034 60215 -10935 60263
rect -10291 60221 -10205 60361
rect -11995 60132 -11955 60152
rect -11993 59923 -11957 60132
rect -9493 63145 -9312 63258
rect -7834 63431 -7717 63681
rect -7961 63314 -7717 63431
rect -9493 62268 -9380 63145
rect -7961 62849 -7844 63314
rect -7967 62751 -7841 62849
rect -7955 62523 -7861 62585
rect -7941 62450 -7889 62523
rect -7711 62475 -7612 62523
rect -9493 62262 -9251 62268
rect -9493 62228 -8968 62262
rect -7948 62349 -7882 62450
rect -8072 62346 -7882 62349
rect -7711 62441 -7446 62475
rect -8072 62345 -7771 62346
rect -8664 62311 -7771 62345
rect -8072 62304 -7771 62311
rect -9493 62221 -9251 62228
rect -9493 62026 -9380 62221
rect -9493 62020 -9261 62026
rect -9493 61986 -8968 62020
rect -9493 61979 -9261 61986
rect -9493 61830 -9380 61979
rect -9493 61824 -9262 61830
rect -9493 61790 -8968 61824
rect -9493 61783 -9262 61790
rect -9493 61117 -9380 61783
rect -7948 61927 -7771 62304
rect -8071 61922 -7771 61927
rect -8664 61888 -7771 61922
rect -8071 61882 -7771 61888
rect -7948 61851 -7771 61882
rect -7711 62279 -7612 62441
rect -7711 62245 -7446 62279
rect -7711 62083 -7612 62245
rect -7167 62181 -7081 62596
rect -7323 62147 -7081 62181
rect -7167 62116 -7081 62147
rect -7711 62049 -7446 62083
rect -7167 62055 -6613 62116
rect -7711 61887 -7612 62049
rect -7167 61985 -7081 62055
rect -7323 61951 -7081 61985
rect -7711 61853 -7446 61887
rect -7948 61732 -7754 61851
rect -8074 61726 -7754 61732
rect -8664 61692 -7754 61726
rect -8074 61687 -7754 61692
rect -7948 61681 -7754 61687
rect -7924 61676 -7754 61681
rect -7711 61676 -7612 61853
rect -7167 61811 -7081 61951
rect -7924 61670 -7612 61676
rect -7924 61636 -7245 61670
rect -8617 61182 -8531 61427
rect -8086 61476 -7987 61524
rect -8252 61442 -7987 61476
rect -8086 61280 -7987 61442
rect -8252 61246 -7987 61280
rect -8617 61148 -8375 61182
rect -8617 61117 -8531 61148
rect -9493 61056 -8531 61117
rect -8086 61084 -7987 61246
rect -9085 60674 -9024 61056
rect -8617 60986 -8531 61056
rect -8252 61050 -7987 61084
rect -8617 60952 -8375 60986
rect -8617 60812 -8531 60952
rect -8086 60888 -7987 61050
rect -8252 60854 -7987 60888
rect -7924 61474 -7662 61636
rect -6674 61746 -6613 62055
rect -6674 61666 -6585 61746
rect -7924 61440 -7245 61474
rect -7924 61278 -7662 61440
rect -7924 61244 -7245 61278
rect -7924 61234 -7662 61244
rect -7924 61233 -7725 61234
rect -7924 60863 -7771 61233
rect -7202 61159 -7148 61294
rect -6671 61608 -6585 61666
rect -6124 61608 -5618 69724
rect -6671 61376 -5618 61608
rect -7016 61342 -5618 61376
rect -6708 61341 -5618 61342
rect -6671 61325 -5618 61341
rect -7196 61139 -7156 61159
rect -9103 60667 -9024 60674
rect -9103 60377 -9042 60667
rect -9103 60343 -8682 60377
rect -9103 60342 -8990 60343
rect -9103 60225 -9042 60342
rect -8086 60677 -7987 60854
rect -8086 60671 -7972 60677
rect -7938 60674 -7771 60863
rect -8453 60637 -7972 60671
rect -7931 60637 -7771 60674
rect -8036 60475 -7972 60637
rect -8453 60441 -7972 60475
rect -8550 60160 -8496 60295
rect -8036 60279 -7972 60441
rect -8453 60245 -7972 60279
rect -8036 60235 -7972 60245
rect -7924 60577 -7771 60637
rect -7581 60893 -7482 60941
rect -7194 60932 -7158 61139
rect -7581 60859 -7216 60893
rect -7581 60697 -7482 60859
rect -6671 61167 -6585 61325
rect -6838 61081 -6585 61167
rect -7581 60663 -7216 60697
rect -7581 60577 -7482 60663
rect -6838 60599 -6752 61081
rect -7924 60501 -7482 60577
rect -7094 60565 -6752 60599
rect -7924 60467 -7216 60501
rect -7924 60305 -7482 60467
rect -6838 60403 -6752 60565
rect -7094 60369 -6752 60403
rect -7924 60271 -7216 60305
rect -7924 60235 -7482 60271
rect -7840 60223 -7482 60235
rect -8542 60140 -8502 60160
rect -19980 5353 -14581 5489
rect -14717 5310 -14581 5353
rect -14518 59787 -11957 59923
rect -14518 41221 -14382 59787
rect -11993 59604 -11957 59787
rect -14170 59217 -13975 59438
rect -8540 59770 -8504 60140
rect -8613 59511 -8350 59770
rect -8598 58645 -8393 59511
rect -7840 58111 -7546 60223
rect -6838 60229 -6752 60369
rect -6802 58922 -6623 59771
rect -6834 58592 -6540 58922
rect -11507 58022 -7418 58111
rect -11507 57918 -11404 58022
rect -11507 57884 -10569 57918
rect -11507 57722 -11404 57884
rect -11507 57688 -10569 57722
rect -11507 57518 -11404 57688
rect -9571 57722 -9474 57918
rect -10392 57688 -9474 57722
rect -11507 57484 -10569 57518
rect -11507 57322 -11404 57484
rect -11507 57288 -10569 57322
rect -11507 56918 -11404 57288
rect -9571 57322 -9474 57688
rect -10392 57288 -9474 57322
rect -11507 56884 -10569 56918
rect -11507 56722 -11404 56884
rect -11507 56688 -10569 56722
rect -11507 56518 -11404 56688
rect -9571 56722 -9474 57288
rect -9249 57824 -9181 58022
rect -9249 57764 -9178 57824
rect -9249 57730 -8887 57764
rect -9249 57568 -9178 57730
rect -8556 57764 -8488 57863
rect -8715 57730 -8488 57764
rect -9249 57534 -8887 57568
rect -9249 57372 -9178 57534
rect -8556 57568 -8488 57730
rect -8176 57862 -8108 57871
rect -8176 57828 -7949 57862
rect -8176 57666 -8108 57828
rect -7486 57862 -7418 58022
rect -7777 57828 -7418 57862
rect -8715 57534 -8488 57568
rect -9249 57338 -8887 57372
rect -9249 57329 -9178 57338
rect -9249 57007 -9181 57329
rect -8556 57372 -8488 57534
rect -8715 57338 -8488 57372
rect -8556 57329 -8488 57338
rect -10392 56688 -9474 56722
rect -11507 56484 -10569 56518
rect -11507 56322 -11404 56484
rect -11507 56288 -10569 56322
rect -11507 55918 -11404 56288
rect -9571 56322 -9474 56688
rect -10392 56288 -9474 56322
rect -11507 55884 -10569 55918
rect -11507 55722 -11404 55884
rect -11507 55688 -10569 55722
rect -11507 55518 -11404 55688
rect -9571 55722 -9474 56288
rect -10392 55688 -9474 55722
rect -11507 55484 -10569 55518
rect -11507 55322 -11404 55484
rect -11507 55288 -10569 55322
rect -11507 54834 -11404 55288
rect -9571 55322 -9474 55688
rect -10392 55288 -9474 55322
rect -9571 55064 -9474 55288
rect -10809 54994 -9474 55064
rect -9246 56082 -9183 57007
rect -9246 56021 -9178 56082
rect -9246 55987 -8887 56021
rect -9246 55825 -9178 55987
rect -8556 56021 -8488 56120
rect -8715 55987 -8488 56021
rect -9246 55791 -8887 55825
rect -9246 55629 -9178 55791
rect -8556 55825 -8488 55987
rect -8715 55791 -8488 55825
rect -9246 55595 -8887 55629
rect -9246 55064 -9178 55595
rect -8823 55483 -8749 55651
rect -8556 55629 -8488 55791
rect -8715 55595 -8488 55629
rect -8812 55423 -8754 55483
rect -8813 55363 -8681 55423
rect -9246 55030 -8887 55064
rect -10809 54904 -10608 54994
rect -11507 54822 -11140 54834
rect -11499 54800 -11140 54822
rect -11499 54638 -11431 54800
rect -10809 54834 -10605 54904
rect -10968 54800 -10605 54834
rect -9530 54884 -9466 54890
rect -10047 54850 -9466 54884
rect -11499 54604 -11140 54638
rect -11499 54442 -11431 54604
rect -10809 54638 -10605 54800
rect -10968 54604 -10605 54638
rect -10809 54492 -10605 54604
rect -9530 54738 -9466 54850
rect -9246 54868 -9178 55030
rect -8556 55064 -8488 55595
rect -8715 55030 -8488 55064
rect -9246 54834 -8887 54868
rect -9246 54789 -9178 54834
rect -9247 54738 -9178 54789
rect -8556 54868 -8488 55030
rect -8715 54834 -8488 54868
rect -9530 54688 -9178 54738
rect -10047 54672 -9178 54688
rect -10047 54654 -8887 54672
rect -9530 54638 -8887 54654
rect -9530 54629 -9178 54638
rect -11499 54408 -11140 54442
rect -11499 54179 -11431 54408
rect -10809 54458 -10293 54492
rect -10809 54442 -10605 54458
rect -10968 54425 -10605 54442
rect -10968 54408 -10608 54425
rect -10809 54399 -10608 54408
rect -11512 54105 -11425 54179
rect -11506 53909 -11439 54105
rect -10766 54096 -10608 54399
rect -9530 54506 -9179 54629
rect -8556 54672 -8488 54834
rect -8715 54638 -8488 54672
rect -8556 54629 -8488 54638
rect -9530 54492 -9466 54506
rect -10047 54458 -9466 54492
rect -9530 54448 -9466 54458
rect -10267 54096 -10186 54097
rect -10766 54015 -10186 54096
rect -9247 54316 -9179 54506
rect -11506 53875 -11147 53909
rect -11506 53713 -11439 53875
rect -10302 53781 -10186 54015
rect -11506 53679 -11147 53713
rect -11506 53487 -11439 53679
rect -10251 53713 -10186 53781
rect -10647 53679 -10186 53713
rect -11523 53424 -11425 53487
rect -11512 53171 -11443 53424
rect -11512 53137 -11147 53171
rect -11512 52975 -11443 53137
rect -11512 52941 -11147 52975
rect -11512 52779 -11443 52941
rect -11512 52745 -11147 52779
rect -11512 52583 -11443 52745
rect -11512 52549 -11147 52583
rect -11512 52390 -11443 52549
rect -11516 52304 -11423 52390
rect -11500 51871 -11431 52304
rect -10251 52681 -10186 53679
rect -10748 52647 -10186 52681
rect -10318 52501 -10186 52647
rect -9246 53382 -9183 54316
rect -9246 53321 -9178 53382
rect -9246 53287 -8887 53321
rect -9246 53125 -9178 53287
rect -8556 53321 -8488 53420
rect -8715 53287 -8488 53321
rect -9246 53091 -8887 53125
rect -9246 52929 -9178 53091
rect -8556 53125 -8488 53287
rect -8715 53091 -8488 53125
rect -9246 52895 -8887 52929
rect -11500 51863 -11298 51871
rect -11500 51829 -10913 51863
rect -11500 51823 -11298 51829
rect -11500 51674 -11431 51823
rect -10318 51965 -10229 52501
rect -9246 52439 -9178 52895
rect -8556 52929 -8488 53091
rect -8715 52895 -8488 52929
rect -9246 52405 -8887 52439
rect -9246 52243 -9178 52405
rect -8556 52439 -8488 52895
rect -8355 55472 -8316 57651
rect -8263 57634 -8224 57651
rect -8276 57623 -8216 57634
rect -8176 57632 -7949 57666
rect -8176 57623 -8108 57632
rect -8276 57512 -8108 57623
rect -7486 57666 -7418 57828
rect -7777 57632 -7418 57666
rect -8276 57497 -8216 57512
rect -8263 56812 -8224 57497
rect -8176 57470 -8108 57512
rect -8176 57436 -7949 57470
rect -8176 57025 -8108 57436
rect -7486 57470 -7418 57632
rect -7777 57436 -7418 57470
rect -8176 56991 -7949 57025
rect -8176 56829 -8108 56991
rect -7486 57025 -7418 57436
rect -7777 56991 -7418 57025
rect -8176 56812 -7949 56829
rect -8263 56795 -7949 56812
rect -8263 56701 -8108 56795
rect -7486 56829 -7418 56991
rect -7777 56795 -7418 56829
rect -8365 55335 -8305 55472
rect -8355 54526 -8316 55335
rect -8263 55037 -8224 56701
rect -8176 56633 -8108 56701
rect -8176 56599 -7949 56633
rect -8176 56500 -8108 56599
rect -7486 56633 -7418 56795
rect -7777 56599 -7418 56633
rect -7486 56538 -7418 56599
rect -7481 55640 -7418 56538
rect -8176 55162 -8108 55171
rect -8176 55128 -7949 55162
rect -8282 55014 -8222 55037
rect -8176 55014 -8108 55128
rect -7486 55162 -7418 55640
rect -7777 55128 -7418 55162
rect -8282 54966 -8108 55014
rect -8282 54932 -7949 54966
rect -8282 54903 -8108 54932
rect -8282 54900 -8222 54903
rect -8366 54394 -8306 54526
rect -8715 52405 -8488 52439
rect -9246 52209 -8887 52243
rect -9246 52047 -9178 52209
rect -8556 52243 -8488 52405
rect -8715 52209 -8488 52243
rect -9246 52013 -8887 52047
rect -9246 52004 -9178 52013
rect -10469 51961 -10229 51965
rect -10629 51927 -10229 51961
rect -10469 51921 -10229 51927
rect -11500 51667 -11304 51674
rect -11500 51633 -10913 51667
rect -11500 51626 -11304 51633
rect -11500 50925 -11431 51626
rect -10318 51855 -10229 51921
rect -8823 51960 -8749 52069
rect -8556 52047 -8488 52209
rect -8715 52013 -8488 52047
rect -8556 52004 -8488 52013
rect -8355 52027 -8316 54394
rect -8263 54136 -8224 54900
rect -8176 54831 -8108 54903
rect -7486 54966 -7418 55128
rect -7777 54932 -7418 54966
rect -8178 54770 -8108 54831
rect -8178 54736 -7949 54770
rect -8178 54637 -8108 54736
rect -7486 54770 -7418 54932
rect -7777 54736 -7418 54770
rect -8178 54334 -8110 54637
rect -8074 54437 -7852 54497
rect -8178 54325 -8108 54334
rect -8178 54311 -7949 54325
rect -8176 54291 -7949 54311
rect -8176 54136 -8108 54291
rect -7915 54269 -7841 54437
rect -7486 54325 -7418 54736
rect -7777 54291 -7418 54325
rect -8263 54129 -8108 54136
rect -8263 54095 -7949 54129
rect -8263 54025 -8108 54095
rect -7486 54129 -7418 54291
rect -7777 54095 -7418 54129
rect -8263 52451 -8224 54025
rect -8176 53933 -8108 54025
rect -8176 53899 -7949 53933
rect -8176 53800 -8108 53899
rect -7486 53933 -7418 54095
rect -7777 53899 -7418 53933
rect -7486 53838 -7418 53899
rect -7481 52886 -7418 53838
rect -8263 52399 -7588 52451
rect -8282 52267 -7588 52399
rect -8263 52266 -8224 52267
rect -7694 52124 -7588 52267
rect -6124 52124 -5618 61325
rect -3630 59641 -2527 119211
rect -5019 58538 -2527 59641
rect -7981 52027 -7846 52053
rect -8355 51960 -7846 52027
rect -8823 51921 -7846 51960
rect -8823 51901 -8749 51921
rect -7694 51855 -3747 52124
rect -10318 51771 -3747 51855
rect -10470 51765 -3747 51771
rect -10629 51731 -3747 51765
rect -10470 51727 -3747 51731
rect -10318 51706 -3747 51727
rect -11500 50917 -11298 50925
rect -11500 50883 -10913 50917
rect -11500 50877 -11298 50883
rect -11500 50728 -11431 50877
rect -10318 51019 -10229 51706
rect -10469 51015 -10229 51019
rect -10629 50981 -10229 51015
rect -10469 50975 -10229 50981
rect -11500 50721 -11304 50728
rect -11500 50687 -10913 50721
rect -11500 50680 -11304 50687
rect -11500 49983 -11431 50680
rect -10318 50825 -10229 50975
rect -10470 50819 -10229 50825
rect -10629 50785 -10229 50819
rect -10470 50781 -10229 50785
rect -13802 49894 -11431 49983
rect -13802 49734 -13734 49894
rect -12039 49857 -11431 49894
rect -13802 49700 -13443 49734
rect -13802 49538 -13734 49700
rect -13112 49734 -13044 49743
rect -13271 49700 -13044 49734
rect -13802 49504 -13443 49538
rect -13802 49342 -13734 49504
rect -13112 49538 -13044 49700
rect -13271 49504 -13044 49538
rect -12732 49636 -12664 49735
rect -12039 49696 -11971 49857
rect -12732 49602 -12505 49636
rect -12996 49506 -12957 49523
rect -13112 49495 -13044 49504
rect -13004 49495 -12944 49506
rect -13802 49308 -13443 49342
rect -13802 48897 -13734 49308
rect -13112 49384 -12944 49495
rect -13112 49342 -13044 49384
rect -13004 49369 -12944 49384
rect -13271 49308 -13044 49342
rect -13802 48863 -13443 48897
rect -13802 48701 -13734 48863
rect -13112 48897 -13044 49308
rect -13271 48863 -13044 48897
rect -13802 48667 -13443 48701
rect -13802 48505 -13734 48667
rect -13112 48701 -13044 48863
rect -13271 48684 -13044 48701
rect -12996 48684 -12957 49369
rect -13271 48667 -12957 48684
rect -13112 48573 -12957 48667
rect -13802 48471 -13443 48505
rect -13802 48410 -13734 48471
rect -13112 48505 -13044 48573
rect -13271 48471 -13044 48505
rect -13802 47512 -13739 48410
rect -13112 48372 -13044 48471
rect -13802 47034 -13734 47512
rect -13802 47000 -13443 47034
rect -13802 46838 -13734 47000
rect -13112 47034 -13044 47043
rect -13271 47000 -13044 47034
rect -13802 46804 -13443 46838
rect -13802 46642 -13734 46804
rect -13112 46886 -13044 47000
rect -12996 46909 -12957 48573
rect -12904 47344 -12865 49523
rect -12732 49440 -12664 49602
rect -12042 49636 -11971 49696
rect -12333 49602 -11971 49636
rect -12732 49406 -12505 49440
rect -12732 49244 -12664 49406
rect -12042 49440 -11971 49602
rect -12333 49406 -11971 49440
rect -12732 49210 -12505 49244
rect -12732 49201 -12664 49210
rect -12042 49244 -11971 49406
rect -12333 49210 -11971 49244
rect -12042 49201 -11971 49210
rect -12915 47207 -12855 47344
rect -12998 46886 -12938 46909
rect -13112 46838 -12938 46886
rect -13271 46804 -12938 46838
rect -13112 46775 -12938 46804
rect -13112 46703 -13044 46775
rect -12998 46772 -12938 46775
rect -13802 46608 -13443 46642
rect -13802 46197 -13734 46608
rect -13112 46642 -13042 46703
rect -13271 46608 -13042 46642
rect -13112 46509 -13042 46608
rect -13368 46309 -13146 46369
rect -13802 46163 -13443 46197
rect -13802 46001 -13734 46163
rect -13379 46141 -13305 46309
rect -13110 46206 -13042 46509
rect -13112 46197 -13042 46206
rect -13271 46183 -13042 46197
rect -13271 46163 -13044 46183
rect -13802 45967 -13443 46001
rect -13802 45805 -13734 45967
rect -13112 46008 -13044 46163
rect -12996 46008 -12957 46772
rect -12904 46398 -12865 47207
rect -12914 46266 -12854 46398
rect -13112 46001 -12957 46008
rect -13271 45967 -12957 46001
rect -13112 45897 -12957 45967
rect -13802 45771 -13443 45805
rect -13802 45710 -13734 45771
rect -13112 45805 -13044 45897
rect -13271 45771 -13044 45805
rect -13802 44758 -13739 45710
rect -13112 45672 -13044 45771
rect -12996 44504 -12957 45897
rect -13915 44271 -12957 44504
rect -13915 44243 -12938 44271
rect -13915 42720 -13654 44243
rect -12998 44139 -12938 44243
rect -12996 44138 -12957 44139
rect -12904 43832 -12865 46266
rect -12039 48879 -11971 49201
rect -12732 47893 -12664 47992
rect -12037 47954 -11974 48879
rect -12732 47859 -12505 47893
rect -12732 47697 -12664 47859
rect -12042 47893 -11974 47954
rect -12333 47859 -11974 47893
rect -12732 47663 -12505 47697
rect -12732 47501 -12664 47663
rect -12042 47697 -11974 47859
rect -12333 47663 -11974 47697
rect -12732 47467 -12505 47501
rect -12732 46936 -12664 47467
rect -12471 47355 -12397 47523
rect -12042 47501 -11974 47663
rect -10318 50652 -10229 50781
rect -9212 50932 -9079 51551
rect -9212 50922 -8951 50932
rect -9212 50888 -8367 50922
rect -9212 50879 -8951 50888
rect -9212 50736 -9079 50879
rect -9212 50726 -8967 50736
rect -9212 50692 -8367 50726
rect -9212 50683 -8967 50692
rect -12333 47467 -11974 47501
rect -12466 47295 -12408 47355
rect -12539 47235 -12407 47295
rect -12732 46902 -12505 46936
rect -12732 46740 -12664 46902
rect -12042 46936 -11974 47467
rect -12333 46902 -11974 46936
rect -12732 46706 -12505 46740
rect -12732 46544 -12664 46706
rect -12042 46740 -11974 46902
rect -12333 46706 -11974 46740
rect -12042 46661 -11974 46706
rect -12732 46510 -12505 46544
rect -12732 46501 -12664 46510
rect -12042 46544 -11973 46661
rect -12333 46510 -11973 46544
rect -12042 46501 -11973 46510
rect -12041 46188 -11973 46501
rect -12732 45193 -12664 45292
rect -12037 45254 -11974 46188
rect -12732 45159 -12505 45193
rect -12732 44997 -12664 45159
rect -12042 45193 -11974 45254
rect -12333 45159 -11974 45193
rect -12732 44963 -12505 44997
rect -12732 44801 -12664 44963
rect -12042 44997 -11974 45159
rect -12333 44963 -11974 44997
rect -12732 44767 -12505 44801
rect -12732 44311 -12664 44767
rect -12042 44801 -11974 44963
rect -12333 44767 -11974 44801
rect -12732 44277 -12505 44311
rect -12732 44115 -12664 44277
rect -12042 44311 -11974 44767
rect -12333 44277 -11974 44311
rect -12732 44081 -12505 44115
rect -12732 43919 -12664 44081
rect -12042 44115 -11974 44277
rect -12333 44081 -11974 44115
rect -12732 43885 -12505 43919
rect -12732 43876 -12664 43885
rect -12471 43832 -12397 43941
rect -12042 43919 -11974 44081
rect -12333 43885 -11974 43919
rect -12042 43876 -11974 43885
rect -12904 43793 -12397 43832
rect -12904 43467 -12865 43793
rect -12471 43773 -12397 43793
rect -12970 43172 -12767 43467
rect -13915 42459 -11613 42720
rect -14114 42305 -13935 42326
rect -14114 42222 -11987 42305
rect -14114 42198 -13935 42222
rect -12317 41994 -12269 42046
rect -14069 41940 -12269 41994
rect -14069 41896 -14015 41940
rect -12317 41898 -12269 41940
rect -12070 41933 -11987 42222
rect -11874 42011 -11613 42459
rect -7694 51579 -3747 51706
rect -7694 51027 -7588 51579
rect -7843 51020 -7588 51027
rect -8011 50986 -7588 51020
rect -6124 50996 -5618 51579
rect -7843 50979 -7588 50986
rect -7694 50833 -7588 50979
rect -7840 50824 -7588 50833
rect -8011 50790 -7588 50824
rect -7840 50785 -7588 50790
rect -7694 50681 -7588 50785
rect -6763 50532 -6517 50569
rect -7809 50390 -6517 50532
rect -7809 50353 -7620 50390
rect -6763 50351 -6517 50390
rect -14110 41842 -13985 41896
rect -12452 41851 -12408 41865
rect -12937 41797 -12408 41851
rect -12937 41752 -12883 41797
rect -14110 41698 -12883 41752
rect -12452 41742 -12408 41797
rect -12088 41742 -11981 41933
rect -11874 41750 -10558 42011
rect -6828 48691 -6560 48815
rect -6830 48580 -6560 48691
rect -6830 43172 -6583 48580
rect -12579 41637 -12539 41740
rect -14110 41583 -12539 41637
rect -11106 41527 -10971 41593
rect -14327 41471 -10971 41527
rect -11106 41448 -10971 41471
rect -12722 41426 -12678 41431
rect -14110 41372 -12678 41426
rect -13350 41321 -13213 41329
rect -14110 41267 -13213 41321
rect -12722 41308 -12678 41372
rect -13350 41264 -13213 41267
rect -12164 41222 -12120 41288
rect -12972 41221 -12120 41222
rect -14518 41165 -12120 41221
rect -14518 4472 -14382 41165
rect -12972 41164 -12121 41165
rect -10819 41117 -10558 41750
rect -4080 44102 -3747 51579
rect -4820 42470 -3747 44102
rect -4080 41117 -3747 42470
rect -12941 40856 -3747 41117
rect -14218 40696 -14025 40741
rect -14218 40689 -13796 40696
rect -14218 40655 -13606 40689
rect -14218 40650 -13796 40655
rect -14218 40499 -13918 40650
rect -12941 40693 -12814 40856
rect -13009 40689 -12814 40693
rect -13208 40655 -12814 40689
rect -13009 40650 -12814 40655
rect -14218 40493 -13784 40499
rect -14218 40459 -13606 40493
rect -14218 40453 -13784 40459
rect -14218 40386 -13918 40453
rect -14218 40380 -13794 40386
rect -14218 40346 -13606 40380
rect -14218 40340 -13794 40346
rect -14218 40190 -13918 40340
rect -13346 40327 -13292 40466
rect -12941 40384 -12814 40650
rect -13007 40380 -12814 40384
rect -13208 40346 -12814 40380
rect -13007 40341 -12814 40346
rect -14218 40184 -13789 40190
rect -14218 40150 -13606 40184
rect -14218 40144 -13789 40150
rect -14218 40077 -13918 40144
rect -14218 40070 -13793 40077
rect -14218 40036 -13606 40070
rect -14218 40031 -13793 40036
rect -14218 39879 -13918 40031
rect -12941 40049 -12814 40341
rect -11736 40699 -11545 40706
rect -11736 40665 -11355 40699
rect -11736 40660 -11545 40665
rect -11736 40509 -11667 40660
rect -10672 40703 -10576 40707
rect -10758 40699 -10576 40703
rect -10957 40665 -10576 40699
rect -10758 40660 -10576 40665
rect -10672 40658 -10576 40660
rect -10131 40658 -9870 40856
rect -11736 40503 -11533 40509
rect -11736 40469 -11355 40503
rect -11736 40463 -11533 40469
rect -11736 40396 -11667 40463
rect -11736 40390 -11543 40396
rect -11736 40356 -11355 40390
rect -11736 40350 -11543 40356
rect -11736 40200 -11667 40350
rect -11095 40337 -11041 40476
rect -10672 40461 -9870 40658
rect -10672 40394 -10576 40461
rect -10756 40390 -10576 40394
rect -10957 40356 -10576 40390
rect -10756 40351 -10576 40356
rect -11736 40194 -11538 40200
rect -11736 40160 -11355 40194
rect -11736 40154 -11538 40160
rect -11736 40087 -11667 40154
rect -11736 40080 -11542 40087
rect -14218 39874 -13789 39879
rect -14218 39840 -13606 39874
rect -14218 39833 -13789 39840
rect -14218 39684 -13918 39833
rect -14218 39678 -13789 39684
rect -14218 39644 -13606 39678
rect -14218 37514 -14025 39644
rect -13352 39249 -13298 39388
rect -13260 39282 -13000 39316
rect -13260 39279 -13202 39282
rect -13260 39197 -13223 39279
rect -13321 39160 -13223 39197
rect -13321 38903 -13284 39160
rect -12889 38903 -12836 40049
rect -11736 40046 -11355 40080
rect -11736 40041 -11542 40046
rect -11736 39889 -11667 40041
rect -10672 40155 -10576 40351
rect -10131 40155 -9870 40461
rect -10672 40075 -9870 40155
rect -11736 39884 -11538 39889
rect -11736 39850 -11355 39884
rect -11736 39843 -11538 39850
rect -11736 39776 -11667 39843
rect -11763 39694 -11627 39776
rect -11763 39688 -11538 39694
rect -11763 39654 -11355 39688
rect -11763 39653 -11627 39654
rect -13321 38902 -13201 38903
rect -13012 38902 -12836 38903
rect -13321 38868 -12836 38902
rect -11101 39259 -11047 39398
rect -11009 39292 -10749 39326
rect -11009 39289 -10951 39292
rect -11009 39207 -10972 39289
rect -11070 39170 -10972 39207
rect -13321 38866 -13201 38868
rect -13012 38864 -12836 38868
rect -13987 37689 -13796 37696
rect -13987 37655 -13606 37689
rect -13987 37650 -13796 37655
rect -13987 37514 -13918 37650
rect -12889 37697 -12836 38864
rect -11070 38913 -11033 39170
rect -10638 39958 -9870 40075
rect -10638 39642 -10585 39958
rect -10131 39642 -9870 39958
rect -10638 39623 -9870 39642
rect -9012 40658 -8751 40856
rect -8306 40703 -8210 40707
rect -8306 40699 -8124 40703
rect -8306 40665 -7925 40699
rect -8306 40660 -8124 40665
rect -8306 40658 -8210 40660
rect -9012 40461 -8210 40658
rect -7337 40699 -7146 40706
rect -7527 40665 -7146 40699
rect -7337 40660 -7146 40665
rect -9012 40155 -8751 40461
rect -8306 40394 -8210 40461
rect -8306 40390 -8126 40394
rect -8306 40356 -7925 40390
rect -8306 40351 -8126 40356
rect -8306 40155 -8210 40351
rect -7841 40337 -7787 40476
rect -7215 40509 -7146 40660
rect -7349 40503 -7146 40509
rect -7527 40469 -7146 40503
rect -7349 40463 -7146 40469
rect -7215 40396 -7146 40463
rect -7339 40390 -7146 40396
rect -7527 40356 -7146 40390
rect -7339 40350 -7146 40356
rect -7215 40200 -7146 40350
rect -7344 40194 -7146 40200
rect -9012 40075 -8210 40155
rect -9012 39958 -8244 40075
rect -9012 39642 -8751 39958
rect -8297 39642 -8244 39958
rect -9012 39623 -8244 39642
rect -10638 39445 -8244 39623
rect -10638 39109 -10585 39445
rect -10131 39362 -8751 39445
rect -10131 39109 -9870 39362
rect -10638 38913 -9870 39109
rect -11070 38912 -10950 38913
rect -10761 38912 -9870 38913
rect -11070 38878 -10585 38912
rect -11070 38876 -10950 38878
rect -10761 38874 -10585 38878
rect -11764 38527 -11628 38560
rect -11764 38493 -11366 38527
rect -11764 38437 -11628 38493
rect -12923 37693 -12827 37697
rect -13009 37689 -12827 37693
rect -13208 37655 -12827 37689
rect -13009 37650 -12827 37655
rect -14218 37499 -13918 37514
rect -14218 37493 -13784 37499
rect -14218 37459 -13606 37493
rect -14218 37453 -13784 37459
rect -14218 37386 -13918 37453
rect -14218 37380 -13794 37386
rect -14218 37346 -13606 37380
rect -14218 37340 -13794 37346
rect -14218 37190 -13918 37340
rect -13346 37327 -13292 37466
rect -12923 37384 -12827 37650
rect -13007 37380 -12827 37384
rect -13208 37346 -12827 37380
rect -13007 37341 -12827 37346
rect -14218 37184 -13789 37190
rect -14218 37150 -13606 37184
rect -14218 37144 -13789 37150
rect -14218 37077 -13918 37144
rect -14218 37070 -13793 37077
rect -14218 37036 -13606 37070
rect -14218 37031 -13793 37036
rect -14218 36921 -13918 37031
rect -12923 37065 -12827 37341
rect -14218 35101 -14025 36921
rect -13987 36879 -13918 36921
rect -13987 36874 -13789 36879
rect -13987 36840 -13606 36874
rect -13987 36833 -13789 36840
rect -13987 36684 -13918 36833
rect -13987 36678 -13789 36684
rect -13987 36644 -13606 36678
rect -13352 36249 -13298 36388
rect -13260 36282 -13000 36316
rect -13260 36279 -13202 36282
rect -13260 36197 -13223 36279
rect -13321 36160 -13223 36197
rect -13321 35903 -13284 36160
rect -12889 35903 -12836 37065
rect -13321 35902 -13201 35903
rect -13012 35902 -12836 35903
rect -13321 35868 -12836 35902
rect -13321 35866 -13201 35868
rect -13012 35864 -12836 35868
rect -13987 35189 -13796 35196
rect -13987 35155 -13606 35189
rect -13987 35150 -13796 35155
rect -13987 35101 -13918 35150
rect -12889 35197 -12836 35864
rect -11731 38331 -11662 38437
rect -11731 38297 -11366 38331
rect -11731 38135 -11662 38297
rect -11731 38101 -11366 38135
rect -11731 37977 -11662 38101
rect -10470 38494 -10405 38527
rect -10131 38494 -9870 38912
rect -10470 38429 -9870 38494
rect -10967 38395 -9870 38429
rect -10470 38348 -9870 38395
rect -11736 37939 -11662 37977
rect -11736 37905 -11366 37939
rect -11736 37402 -11663 37905
rect -10470 38134 -10405 38348
rect -10131 38134 -9870 38348
rect -10470 37988 -9870 38134
rect -10470 37868 -10405 37988
rect -10131 37868 -9870 37988
rect -10470 37722 -9870 37868
rect -11736 37397 -11658 37402
rect -11736 37363 -11366 37397
rect -11736 37204 -11658 37363
rect -10470 37423 -10405 37722
rect -10131 37677 -9870 37722
rect -9012 39109 -8751 39362
rect -8297 39109 -8244 39445
rect -9012 38913 -8244 39109
rect -7527 40160 -7146 40194
rect -7344 40154 -7146 40160
rect -7215 40087 -7146 40154
rect -7340 40080 -7146 40087
rect -7527 40046 -7146 40080
rect -6068 40693 -5941 40856
rect -6068 40689 -5873 40693
rect -6068 40655 -5674 40689
rect -6068 40650 -5873 40655
rect -6068 40384 -5941 40650
rect -4857 40696 -4664 40741
rect -5086 40689 -4664 40696
rect -5276 40655 -4664 40689
rect -5086 40650 -4664 40655
rect -6068 40380 -5875 40384
rect -6068 40346 -5674 40380
rect -6068 40341 -5875 40346
rect -6068 40049 -5941 40341
rect -5590 40327 -5536 40466
rect -4964 40499 -4664 40650
rect -3510 40571 -2748 58538
rect -5098 40493 -4664 40499
rect -5276 40459 -4664 40493
rect -5098 40453 -4664 40459
rect -4964 40386 -4664 40453
rect -5088 40380 -4664 40386
rect -5276 40346 -4664 40380
rect -5088 40340 -4664 40346
rect -4964 40272 -4664 40340
rect -3742 40272 -2527 40571
rect -4964 40190 -2527 40272
rect -5093 40184 -2527 40190
rect -7340 40041 -7146 40046
rect -7215 39889 -7146 40041
rect -7344 39884 -7146 39889
rect -7527 39850 -7146 39884
rect -7344 39843 -7146 39850
rect -7215 39776 -7146 39843
rect -7255 39694 -7119 39776
rect -7344 39688 -7119 39694
rect -7527 39654 -7119 39688
rect -7255 39653 -7119 39654
rect -8133 39292 -7873 39326
rect -7931 39289 -7873 39292
rect -7910 39207 -7873 39289
rect -7835 39259 -7781 39398
rect -7910 39170 -7812 39207
rect -7849 38913 -7812 39170
rect -9012 38912 -8121 38913
rect -7932 38912 -7812 38913
rect -9012 38494 -8751 38912
rect -8297 38878 -7812 38912
rect -8297 38874 -8121 38878
rect -7932 38876 -7812 38878
rect -6046 38903 -5993 40049
rect -5276 40150 -2527 40184
rect -5093 40144 -2527 40150
rect -4964 40077 -2527 40144
rect -5089 40070 -2527 40077
rect -5276 40036 -2527 40070
rect -5089 40031 -2527 40036
rect -4964 39879 -2527 40031
rect -5093 39874 -2527 39879
rect -5276 39840 -2527 39874
rect -5093 39833 -2527 39840
rect -4964 39684 -2527 39833
rect -5093 39678 -2527 39684
rect -5276 39644 -2527 39678
rect -5882 39282 -5622 39316
rect -5680 39279 -5622 39282
rect -5659 39197 -5622 39279
rect -5584 39249 -5530 39388
rect -5659 39160 -5561 39197
rect -5598 38903 -5561 39160
rect -6046 38902 -5870 38903
rect -5681 38902 -5561 38903
rect -6046 38868 -5561 38902
rect -6046 38864 -5870 38868
rect -5681 38866 -5561 38868
rect -8477 38494 -8412 38527
rect -9012 38429 -8412 38494
rect -9012 38395 -7915 38429
rect -9012 38348 -8412 38395
rect -9012 38134 -8751 38348
rect -8477 38134 -8412 38348
rect -9012 37988 -8412 38134
rect -9012 37868 -8751 37988
rect -8477 37868 -8412 37988
rect -9012 37722 -8412 37868
rect -7254 38527 -7118 38560
rect -7516 38493 -7118 38527
rect -7254 38437 -7118 38493
rect -7220 38331 -7151 38437
rect -7516 38297 -7151 38331
rect -7220 38135 -7151 38297
rect -7516 38101 -7151 38135
rect -7220 37977 -7151 38101
rect -7220 37939 -7146 37977
rect -7516 37905 -7146 37939
rect -9012 37677 -8751 37722
rect -10131 37423 -8751 37677
rect -8477 37423 -8412 37722
rect -10470 37416 -8412 37423
rect -10470 37397 -9870 37416
rect -10866 37363 -9870 37397
rect -10470 37277 -9870 37363
rect -11769 37201 -11633 37204
rect -11769 37167 -11366 37201
rect -11769 37081 -11633 37167
rect -10470 37253 -10405 37277
rect -12923 35193 -12827 35197
rect -13009 35189 -12827 35193
rect -13208 35155 -12827 35189
rect -13009 35150 -12827 35155
rect -14218 34999 -13918 35101
rect -14218 34993 -13784 34999
rect -14218 34959 -13606 34993
rect -14218 34953 -13784 34959
rect -14218 34886 -13918 34953
rect -14218 34880 -13794 34886
rect -14218 34846 -13606 34880
rect -14218 34840 -13794 34846
rect -14218 34690 -13918 34840
rect -13346 34827 -13292 34966
rect -12923 34884 -12827 35150
rect -13007 34880 -12827 34884
rect -13208 34846 -12827 34880
rect -13007 34841 -12827 34846
rect -14218 34684 -13789 34690
rect -14218 34650 -13606 34684
rect -14218 34644 -13789 34650
rect -14218 34577 -13918 34644
rect -14218 34570 -13793 34577
rect -14218 34536 -13606 34570
rect -14218 34531 -13793 34536
rect -14218 34508 -13918 34531
rect -12923 34565 -12827 34841
rect -14218 33136 -14025 34508
rect -13987 34379 -13918 34508
rect -13987 34374 -13789 34379
rect -13987 34340 -13606 34374
rect -13987 34333 -13789 34340
rect -13987 34184 -13918 34333
rect -13987 34178 -13789 34184
rect -13987 34144 -13606 34178
rect -13352 33749 -13298 33888
rect -13260 33782 -13000 33816
rect -13260 33779 -13202 33782
rect -13260 33697 -13223 33779
rect -13321 33660 -13223 33697
rect -13321 33403 -13284 33660
rect -12889 33403 -12836 34565
rect -11767 36774 -11631 36803
rect -11767 36740 -11241 36774
rect -11767 36680 -11631 36740
rect -10652 36788 -10591 36794
rect -10131 36788 -9870 37277
rect -11722 36578 -11658 36680
rect -11722 36544 -11241 36578
rect -11722 36382 -11658 36544
rect -11722 36348 -11241 36382
rect -11722 36342 -11608 36348
rect -11707 36165 -11608 36342
rect -10652 36677 -9870 36788
rect -10704 36676 -9870 36677
rect -11012 36642 -9870 36676
rect -10652 36637 -9870 36642
rect -10652 36495 -10591 36637
rect -10131 36495 -9870 36637
rect -10652 36463 -9870 36495
rect -9012 37397 -8412 37416
rect -9012 37363 -8016 37397
rect -9012 37277 -8412 37363
rect -7219 37402 -7146 37905
rect -7224 37397 -7146 37402
rect -7516 37363 -7146 37397
rect -9012 36788 -8751 37277
rect -8477 37253 -8412 37277
rect -7224 37204 -7146 37363
rect -7249 37201 -7113 37204
rect -7516 37167 -7113 37201
rect -7249 37081 -7113 37167
rect -8291 36788 -8230 36794
rect -9012 36677 -8230 36788
rect -9012 36676 -8178 36677
rect -9012 36642 -7870 36676
rect -9012 36637 -8230 36642
rect -9012 36495 -8751 36637
rect -8291 36495 -8230 36637
rect -9012 36463 -8230 36495
rect -10652 36352 -8230 36463
rect -7251 36774 -7115 36803
rect -7641 36740 -7115 36774
rect -7251 36680 -7115 36740
rect -7224 36578 -7160 36680
rect -7641 36544 -7160 36578
rect -10670 36344 -8212 36352
rect -11707 36131 -11442 36165
rect -11707 35969 -11608 36131
rect -11163 36067 -11077 36207
rect -11319 36033 -11077 36067
rect -11707 35935 -11442 35969
rect -11163 35963 -11077 36033
rect -10670 36053 -10609 36344
rect -10131 36202 -8751 36344
rect -10131 36053 -9870 36202
rect -10670 35963 -9870 36053
rect -11707 35773 -11608 35935
rect -11163 35902 -9870 35963
rect -11163 35871 -11077 35902
rect -11319 35837 -11077 35871
rect -11707 35739 -11442 35773
rect -11707 35577 -11608 35739
rect -11707 35575 -11442 35577
rect -11744 35543 -11442 35575
rect -11163 35592 -11077 35837
rect -11744 35452 -11608 35543
rect -13321 33402 -13201 33403
rect -13012 33402 -12836 33403
rect -13321 33368 -12836 33402
rect -13321 33366 -13201 33368
rect -13012 33364 -12836 33368
rect -13153 33136 -13017 33139
rect -14218 33021 -13017 33136
rect -14218 32567 -14025 33021
rect -13153 33016 -13017 33021
rect -13987 32689 -13796 32696
rect -13987 32655 -13606 32689
rect -13987 32650 -13796 32655
rect -13987 32567 -13918 32650
rect -12889 32697 -12836 33364
rect -12923 32693 -12827 32697
rect -13009 32689 -12827 32693
rect -13208 32655 -12827 32689
rect -13009 32650 -12827 32655
rect -14218 32499 -13918 32567
rect -14218 32493 -13784 32499
rect -14218 32459 -13606 32493
rect -14218 32453 -13784 32459
rect -14218 32386 -13918 32453
rect -14218 32380 -13794 32386
rect -14218 32346 -13606 32380
rect -14218 32340 -13794 32346
rect -14218 32190 -13918 32340
rect -13346 32327 -13292 32466
rect -12923 32384 -12827 32650
rect -13007 32380 -12827 32384
rect -13208 32346 -12827 32380
rect -13007 32341 -12827 32346
rect -14218 32184 -13789 32190
rect -14218 32150 -13606 32184
rect -14218 32144 -13789 32150
rect -14218 32077 -13918 32144
rect -14218 32070 -13793 32077
rect -14218 32036 -13606 32070
rect -14218 32031 -13793 32036
rect -14218 31974 -13918 32031
rect -12923 32065 -12827 32341
rect -14218 30653 -14025 31974
rect -13987 31879 -13918 31974
rect -13987 31874 -13789 31879
rect -13987 31840 -13606 31874
rect -13987 31833 -13789 31840
rect -13987 31684 -13918 31833
rect -13987 31678 -13789 31684
rect -13987 31644 -13606 31678
rect -13352 31249 -13298 31388
rect -13260 31282 -13000 31316
rect -13260 31279 -13202 31282
rect -13260 31197 -13223 31279
rect -13321 31160 -13223 31197
rect -13321 30903 -13284 31160
rect -12889 30903 -12836 32065
rect -11743 35169 -11607 35186
rect -11743 35135 -11243 35169
rect -11743 35063 -11607 35135
rect -11729 34973 -11650 35063
rect -11729 34939 -11243 34973
rect -11729 34777 -11650 34939
rect -11729 34743 -11243 34777
rect -11729 34560 -11610 34743
rect -10654 35128 -10593 35189
rect -10131 35128 -9870 35902
rect -10654 35072 -9870 35128
rect -10706 35071 -9870 35072
rect -11014 35037 -9870 35071
rect -10654 35005 -9870 35037
rect -9012 36053 -8751 36202
rect -8273 36053 -8212 36344
rect -7224 36382 -7160 36544
rect -7641 36348 -7160 36382
rect -7274 36342 -7160 36348
rect -9012 35963 -8212 36053
rect -7805 36067 -7719 36207
rect -7274 36165 -7175 36342
rect -7440 36131 -7175 36165
rect -7805 36033 -7563 36067
rect -7805 35963 -7719 36033
rect -7274 35969 -7175 36131
rect -9012 35902 -7719 35963
rect -7440 35935 -7175 35969
rect -9012 35128 -8751 35902
rect -7805 35871 -7719 35902
rect -7805 35837 -7563 35871
rect -7805 35592 -7719 35837
rect -7274 35773 -7175 35935
rect -7440 35739 -7175 35773
rect -7274 35577 -7175 35739
rect -7440 35575 -7175 35577
rect -7440 35543 -7138 35575
rect -7274 35452 -7138 35543
rect -6046 37697 -5993 38864
rect -4857 39510 -2527 39644
rect -6055 37693 -5959 37697
rect -6055 37689 -5873 37693
rect -6055 37655 -5674 37689
rect -6055 37650 -5873 37655
rect -6055 37384 -5959 37650
rect -5086 37689 -4895 37696
rect -5276 37655 -4895 37689
rect -5086 37650 -4895 37655
rect -6055 37380 -5875 37384
rect -6055 37346 -5674 37380
rect -6055 37341 -5875 37346
rect -6055 37065 -5959 37341
rect -5590 37327 -5536 37466
rect -4964 37514 -4895 37650
rect -4857 37514 -4664 39510
rect -3742 39356 -2527 39510
rect -4964 37499 -4664 37514
rect -5098 37493 -4664 37499
rect -5276 37459 -4664 37493
rect -5098 37453 -4664 37459
rect -4964 37386 -4664 37453
rect -5088 37380 -4664 37386
rect -5276 37346 -4664 37380
rect -5088 37340 -4664 37346
rect -4964 37190 -4664 37340
rect -5093 37184 -4664 37190
rect -6046 35903 -5993 37065
rect -5276 37150 -4664 37184
rect -5093 37144 -4664 37150
rect -4964 37077 -4664 37144
rect -5089 37070 -4664 37077
rect -5276 37036 -4664 37070
rect -5089 37031 -4664 37036
rect -4964 36921 -4664 37031
rect -4964 36879 -4895 36921
rect -5093 36874 -4895 36879
rect -5276 36840 -4895 36874
rect -5093 36833 -4895 36840
rect -4964 36684 -4895 36833
rect -5093 36678 -4895 36684
rect -5276 36644 -4895 36678
rect -5882 36282 -5622 36316
rect -5680 36279 -5622 36282
rect -5659 36197 -5622 36279
rect -5584 36249 -5530 36388
rect -5659 36160 -5561 36197
rect -5598 35903 -5561 36160
rect -6046 35902 -5870 35903
rect -5681 35902 -5561 35903
rect -6046 35868 -5561 35902
rect -6046 35864 -5870 35868
rect -5681 35866 -5561 35868
rect -8289 35128 -8228 35189
rect -9012 35072 -8228 35128
rect -9012 35071 -8176 35072
rect -9012 35037 -7868 35071
rect -9012 35005 -8228 35037
rect -10654 35004 -8228 35005
rect -10654 34798 -10593 35004
rect -10131 34798 -8751 35004
rect -8289 34798 -8228 35004
rect -10654 34747 -8228 34798
rect -7275 35169 -7139 35186
rect -7639 35135 -7139 35169
rect -7275 35063 -7139 35135
rect -7232 34973 -7153 35063
rect -7639 34939 -7153 34973
rect -10672 34744 -8210 34747
rect -10672 34674 -9870 34744
rect -11729 34526 -11444 34560
rect -11729 34364 -11610 34526
rect -11165 34462 -11079 34602
rect -11321 34428 -11079 34462
rect -11729 34330 -11444 34364
rect -11165 34358 -11079 34428
rect -10672 34448 -10611 34674
rect -10131 34448 -9870 34674
rect -10672 34358 -9870 34448
rect -11729 34168 -11610 34330
rect -11165 34297 -9870 34358
rect -11165 34266 -11079 34297
rect -11321 34232 -11079 34266
rect -11729 34134 -11444 34168
rect -11729 33972 -11610 34134
rect -11729 33938 -11444 33972
rect -11165 33987 -11079 34232
rect -10131 33965 -9870 34297
rect -9012 34674 -8210 34744
rect -9012 34448 -8751 34674
rect -8271 34448 -8210 34674
rect -7232 34777 -7153 34939
rect -7639 34743 -7153 34777
rect -9012 34358 -8210 34448
rect -7803 34462 -7717 34602
rect -7272 34560 -7153 34743
rect -7438 34526 -7153 34560
rect -7803 34428 -7561 34462
rect -7803 34358 -7717 34428
rect -7272 34364 -7153 34526
rect -9012 34297 -7717 34358
rect -7438 34330 -7153 34364
rect -9012 33965 -8751 34297
rect -7803 34266 -7717 34297
rect -7803 34232 -7561 34266
rect -7803 33987 -7717 34232
rect -7272 34168 -7153 34330
rect -7438 34134 -7153 34168
rect -11729 33890 -11610 33938
rect -11729 33565 -11650 33890
rect -11729 33531 -11357 33565
rect -11729 33369 -11650 33531
rect -11729 33335 -11357 33369
rect -12599 33138 -12537 33321
rect -12600 33135 -12537 33138
rect -11729 33173 -11650 33335
rect -11729 33139 -11357 33173
rect -11729 33135 -11650 33139
rect -12600 33020 -11650 33135
rect -10131 33704 -8751 33965
rect -7272 33972 -7153 34134
rect -10461 33503 -10396 33565
rect -10131 33503 -9870 33704
rect -10461 33467 -9870 33503
rect -10958 33433 -9870 33467
rect -10461 33373 -9870 33433
rect -12600 33015 -12537 33020
rect -11729 32977 -11650 33020
rect -11729 32943 -11357 32977
rect -11729 32440 -11650 32943
rect -10461 33057 -10396 33373
rect -10131 33128 -9870 33373
rect -9012 33503 -8751 33704
rect -7438 33938 -7153 33972
rect -8486 33503 -8421 33565
rect -9012 33467 -8421 33503
rect -9012 33433 -7924 33467
rect -9012 33373 -8421 33433
rect -9012 33128 -8751 33373
rect -10131 33057 -8751 33128
rect -8486 33057 -8421 33373
rect -10461 32927 -8421 33057
rect -10461 32740 -10396 32927
rect -10131 32867 -8751 32927
rect -10131 32740 -9870 32867
rect -10461 32610 -9870 32740
rect -11729 32435 -11649 32440
rect -11729 32401 -11357 32435
rect -11729 32239 -11649 32401
rect -10461 32435 -10396 32610
rect -10857 32434 -10396 32435
rect -10131 32434 -9870 32610
rect -10857 32401 -9870 32434
rect -10461 32304 -9870 32401
rect -11729 32208 -11357 32239
rect -11756 32205 -11357 32208
rect -11910 31989 -11859 32087
rect -11756 32085 -11620 32205
rect -10461 32291 -10396 32304
rect -11310 31989 -11236 32009
rect -11910 31950 -10803 31989
rect -11755 31897 -11619 31914
rect -11755 31863 -11374 31897
rect -11755 31791 -11619 31863
rect -11310 31841 -11236 31950
rect -11043 31897 -10975 31906
rect -11202 31863 -10975 31897
rect -11733 31701 -11665 31791
rect -11733 31667 -11374 31701
rect -11733 31505 -11665 31667
rect -11043 31701 -10975 31863
rect -11202 31667 -10975 31701
rect -11733 31471 -11374 31505
rect -11733 31015 -11665 31471
rect -11043 31505 -10975 31667
rect -11202 31471 -10975 31505
rect -11733 30981 -11374 31015
rect -13321 30902 -13201 30903
rect -13012 30902 -12836 30903
rect -13321 30868 -12836 30902
rect -13321 30866 -13201 30868
rect -13012 30864 -12836 30868
rect -13153 30653 -13017 30656
rect -14218 30539 -13017 30653
rect -14218 30051 -14025 30539
rect -13153 30533 -13017 30539
rect -13987 30189 -13796 30196
rect -13987 30155 -13606 30189
rect -13987 30150 -13796 30155
rect -13987 30051 -13918 30150
rect -12889 30197 -12836 30864
rect -11733 30819 -11665 30981
rect -11043 31015 -10975 31471
rect -11202 30981 -10975 31015
rect -11733 30785 -11374 30819
rect -12565 30651 -12429 30655
rect -11733 30651 -11665 30785
rect -11043 30819 -10975 30981
rect -11202 30785 -10975 30819
rect -12565 30623 -11665 30651
rect -12565 30589 -11374 30623
rect -12565 30536 -11665 30589
rect -12565 30532 -12429 30536
rect -11733 30528 -11665 30536
rect -11043 30623 -10975 30785
rect -11202 30589 -10975 30623
rect -12923 30193 -12827 30197
rect -13009 30189 -12827 30193
rect -13208 30155 -12827 30189
rect -13009 30150 -12827 30155
rect -14218 29999 -13918 30051
rect -14218 29993 -13784 29999
rect -14218 29959 -13606 29993
rect -14218 29953 -13784 29959
rect -14218 29886 -13918 29953
rect -14218 29880 -13794 29886
rect -14218 29846 -13606 29880
rect -14218 29840 -13794 29846
rect -14218 29690 -13918 29840
rect -13346 29827 -13292 29966
rect -12923 29884 -12827 30150
rect -13007 29880 -12827 29884
rect -13208 29846 -12827 29880
rect -13007 29841 -12827 29846
rect -14218 29684 -13789 29690
rect -14218 29650 -13606 29684
rect -14218 29644 -13789 29650
rect -14218 29577 -13918 29644
rect -14218 29570 -13793 29577
rect -14218 29536 -13606 29570
rect -14218 29531 -13793 29536
rect -14218 29458 -13918 29531
rect -12923 29565 -12827 29841
rect -11733 29594 -11670 30528
rect -11043 30490 -10975 30589
rect -14218 28086 -14025 29458
rect -13987 29379 -13918 29458
rect -13987 29374 -13789 29379
rect -13987 29340 -13606 29374
rect -13987 29333 -13789 29340
rect -13987 29184 -13918 29333
rect -13987 29178 -13789 29184
rect -13987 29144 -13606 29178
rect -13352 28749 -13298 28888
rect -13260 28782 -13000 28816
rect -13260 28779 -13202 28782
rect -13260 28697 -13223 28779
rect -13321 28660 -13223 28697
rect -13321 28403 -13284 28660
rect -12889 28403 -12836 29565
rect -11734 29281 -11666 29594
rect -11734 29272 -11665 29281
rect -11734 29238 -11374 29272
rect -11734 29121 -11665 29238
rect -11043 29272 -10975 29281
rect -11202 29238 -10975 29272
rect -13321 28402 -13201 28403
rect -13012 28402 -12836 28403
rect -13321 28368 -12836 28402
rect -13321 28366 -13201 28368
rect -13012 28364 -12836 28368
rect -11733 29076 -11665 29121
rect -11733 29042 -11374 29076
rect -11733 28880 -11665 29042
rect -11043 29076 -10975 29238
rect -11202 29042 -10975 29076
rect -11733 28846 -11374 28880
rect -13188 28086 -13052 28089
rect -14218 27971 -13052 28086
rect -14218 27696 -14025 27971
rect -13188 27966 -13052 27971
rect -14218 27689 -13796 27696
rect -14218 27655 -13606 27689
rect -14218 27650 -13796 27655
rect -14218 27499 -13918 27650
rect -12924 27697 -12837 28364
rect -11733 28315 -11665 28846
rect -11043 28880 -10975 29042
rect -11202 28846 -10975 28880
rect -11300 28487 -11168 28547
rect -11299 28427 -11241 28487
rect -11733 28281 -11374 28315
rect -11733 28119 -11665 28281
rect -11310 28259 -11236 28427
rect -11043 28315 -10975 28846
rect -11202 28281 -10975 28315
rect -12421 28085 -12285 28088
rect -11733 28085 -11374 28119
rect -12421 27970 -11665 28085
rect -11043 28119 -10975 28281
rect -11202 28085 -10975 28119
rect -12421 27965 -12285 27970
rect -11733 27923 -11665 27970
rect -11733 27889 -11374 27923
rect -11733 27828 -11665 27889
rect -11043 27923 -10975 28085
rect -11202 27889 -10975 27923
rect -12924 27693 -12827 27697
rect -13009 27689 -12827 27693
rect -13208 27655 -12827 27689
rect -13009 27650 -12827 27655
rect -12924 27576 -12827 27650
rect -14218 27493 -13784 27499
rect -14218 27459 -13606 27493
rect -14218 27453 -13784 27459
rect -14218 27386 -13918 27453
rect -14218 27380 -13794 27386
rect -14218 27346 -13606 27380
rect -14218 27340 -13794 27346
rect -14218 27190 -13918 27340
rect -13346 27327 -13292 27466
rect -12923 27384 -12827 27576
rect -13007 27380 -12827 27384
rect -13208 27346 -12827 27380
rect -13007 27341 -12827 27346
rect -14218 27184 -13789 27190
rect -14218 27150 -13606 27184
rect -14218 27144 -13789 27150
rect -14218 27077 -13918 27144
rect -14218 27070 -13793 27077
rect -14218 27036 -13606 27070
rect -14218 27031 -13793 27036
rect -14218 26879 -13918 27031
rect -12923 27065 -12827 27341
rect -14218 26874 -13789 26879
rect -14218 26840 -13606 26874
rect -14218 26833 -13789 26840
rect -14218 26684 -13918 26833
rect -14218 26678 -13789 26684
rect -14218 26644 -13606 26678
rect -14218 25779 -14025 26644
rect -13352 26249 -13298 26388
rect -13260 26282 -13000 26316
rect -13260 26279 -13202 26282
rect -13260 26197 -13223 26279
rect -13321 26160 -13223 26197
rect -13321 25903 -13284 26160
rect -12889 25903 -12836 27065
rect -11733 26903 -11670 27828
rect -11043 27790 -10975 27889
rect -13321 25902 -13201 25903
rect -13012 25902 -12836 25903
rect -13321 25868 -12836 25902
rect -13321 25866 -13201 25868
rect -13012 25864 -12836 25868
rect -11736 26581 -11668 26903
rect -10842 29516 -10803 31950
rect -10750 31643 -10711 31644
rect -10769 31556 -10709 31643
rect -10131 31556 -9870 32304
rect -9012 32740 -8751 32867
rect -8486 32740 -8421 32927
rect -7272 33890 -7153 33938
rect -7232 33565 -7153 33890
rect -7525 33531 -7153 33565
rect -7232 33369 -7153 33531
rect -7525 33335 -7153 33369
rect -7232 33173 -7153 33335
rect -7525 33139 -7153 33173
rect -7232 33135 -7153 33139
rect -6345 33138 -6283 33321
rect -6345 33135 -6282 33138
rect -7232 33020 -6282 33135
rect -7232 32977 -7153 33020
rect -6345 33015 -6282 33020
rect -7525 32943 -7153 32977
rect -9012 32610 -8421 32740
rect -9012 32434 -8751 32610
rect -8486 32435 -8421 32610
rect -8486 32434 -8025 32435
rect -9012 32401 -8025 32434
rect -9012 32304 -8421 32401
rect -7232 32440 -7153 32943
rect -7233 32435 -7153 32440
rect -7525 32401 -7153 32435
rect -9012 31556 -8751 32304
rect -8486 32291 -8421 32304
rect -7233 32239 -7153 32401
rect -7525 32208 -7153 32239
rect -7525 32205 -7126 32208
rect -7262 32085 -7126 32205
rect -7646 31989 -7572 32009
rect -7023 31989 -6972 32087
rect -7993 31950 -6972 31989
rect -8171 31773 -8132 31774
rect -8173 31641 -8113 31773
rect -8171 31556 -8132 31641
rect -10769 31511 -8132 31556
rect -10750 31258 -8132 31511
rect -10750 29885 -10711 31258
rect -9968 30575 -9905 31024
rect -8977 30575 -8914 31024
rect -9968 30306 -8914 30575
rect -10663 30011 -10595 30110
rect -9968 30072 -9905 30306
rect -10663 29977 -10436 30011
rect -10663 29885 -10595 29977
rect -9973 30011 -9905 30072
rect -10264 29977 -9905 30011
rect -10750 29815 -10595 29885
rect -10750 29781 -10436 29815
rect -10750 29774 -10595 29781
rect -10853 29384 -10793 29516
rect -10842 28575 -10803 29384
rect -10750 29010 -10711 29774
rect -10663 29619 -10595 29774
rect -9973 29815 -9905 29977
rect -10264 29781 -9905 29815
rect -10663 29599 -10436 29619
rect -10665 29585 -10436 29599
rect -10665 29576 -10595 29585
rect -10665 29273 -10597 29576
rect -10402 29473 -10328 29641
rect -9973 29619 -9905 29781
rect -10264 29585 -9905 29619
rect -9973 29544 -9905 29585
rect -8977 30072 -8914 30306
rect -8977 30011 -8909 30072
rect -8977 29977 -8618 30011
rect -8977 29815 -8909 29977
rect -8287 30011 -8219 30110
rect -8446 29977 -8219 30011
rect -8287 29885 -8219 29977
rect -8171 29885 -8132 31258
rect -8977 29781 -8618 29815
rect -8977 29619 -8909 29781
rect -8287 29815 -8132 29885
rect -8446 29781 -8132 29815
rect -8287 29774 -8132 29781
rect -8977 29585 -8618 29619
rect -8977 29544 -8909 29585
rect -10561 29413 -10339 29473
rect -10665 29174 -10595 29273
rect -9973 29275 -8909 29544
rect -8287 29619 -8219 29774
rect -8446 29599 -8219 29619
rect -8446 29585 -8217 29599
rect -8287 29576 -8217 29585
rect -10665 29140 -10436 29174
rect -10665 29079 -10595 29140
rect -9973 29174 -9905 29275
rect -10264 29140 -9905 29174
rect -10769 29007 -10709 29010
rect -10663 29007 -10595 29079
rect -10769 28978 -10595 29007
rect -10769 28944 -10436 28978
rect -10769 28896 -10595 28944
rect -10769 28873 -10709 28896
rect -10852 28438 -10792 28575
rect -11736 26572 -11665 26581
rect -11736 26538 -11374 26572
rect -11736 26376 -11665 26538
rect -11043 26572 -10975 26581
rect -11202 26538 -10975 26572
rect -11736 26342 -11374 26376
rect -11736 26180 -11665 26342
rect -11043 26376 -10975 26538
rect -11202 26342 -10975 26376
rect -11736 26146 -11374 26180
rect -11736 26086 -11665 26146
rect -11043 26180 -10975 26342
rect -10842 26259 -10803 28438
rect -10750 27209 -10711 28873
rect -10663 28782 -10595 28896
rect -9973 28978 -9905 29140
rect -10264 28944 -9905 28978
rect -10663 28748 -10436 28782
rect -10663 28739 -10595 28748
rect -9973 28782 -9905 28944
rect -10264 28748 -9905 28782
rect -9973 28641 -9905 28748
rect -8977 29174 -8909 29275
rect -8285 29273 -8217 29576
rect -8977 29140 -8618 29174
rect -8977 28978 -8909 29140
rect -8287 29174 -8217 29273
rect -8446 29140 -8217 29174
rect -8287 29079 -8217 29140
rect -8977 28944 -8618 28978
rect -8977 28782 -8909 28944
rect -8287 29007 -8219 29079
rect -8171 29010 -8132 29774
rect -7993 30431 -7954 31950
rect -7907 31897 -7839 31906
rect -7907 31863 -7680 31897
rect -7907 31701 -7839 31863
rect -7646 31841 -7572 31950
rect -7263 31897 -7127 31914
rect -7508 31863 -7127 31897
rect -7263 31791 -7127 31863
rect -7907 31667 -7680 31701
rect -7907 31505 -7839 31667
rect -7217 31701 -7149 31791
rect -7508 31667 -7149 31701
rect -7907 31471 -7680 31505
rect -7907 31015 -7839 31471
rect -7217 31505 -7149 31667
rect -7508 31471 -7149 31505
rect -7641 31127 -7583 31162
rect -7907 30981 -7680 31015
rect -7907 30819 -7839 30981
rect -7646 30959 -7572 31127
rect -7217 31015 -7149 31471
rect -7508 30981 -7149 31015
rect -6046 35197 -5993 35864
rect -6055 35193 -5959 35197
rect -6055 35189 -5873 35193
rect -6055 35155 -5674 35189
rect -6055 35150 -5873 35155
rect -6055 34884 -5959 35150
rect -5086 35189 -4895 35196
rect -5276 35155 -4895 35189
rect -5086 35150 -4895 35155
rect -4964 35101 -4895 35150
rect -4857 35101 -4664 36921
rect -6055 34880 -5875 34884
rect -6055 34846 -5674 34880
rect -6055 34841 -5875 34846
rect -6055 34565 -5959 34841
rect -5590 34827 -5536 34966
rect -4964 34999 -4664 35101
rect -5098 34993 -4664 34999
rect -5276 34959 -4664 34993
rect -5098 34953 -4664 34959
rect -4964 34886 -4664 34953
rect -5088 34880 -4664 34886
rect -5276 34846 -4664 34880
rect -5088 34840 -4664 34846
rect -4964 34690 -4664 34840
rect -5093 34684 -4664 34690
rect -6046 33403 -5993 34565
rect -5276 34650 -4664 34684
rect -5093 34644 -4664 34650
rect -4964 34577 -4664 34644
rect -5089 34570 -4664 34577
rect -5276 34536 -4664 34570
rect -5089 34531 -4664 34536
rect -4964 34508 -4664 34531
rect -4964 34379 -4895 34508
rect -5093 34374 -4895 34379
rect -5276 34340 -4895 34374
rect -5093 34333 -4895 34340
rect -4964 34184 -4895 34333
rect -5093 34178 -4895 34184
rect -5276 34144 -4895 34178
rect -5882 33782 -5622 33816
rect -5680 33779 -5622 33782
rect -5659 33697 -5622 33779
rect -5584 33749 -5530 33888
rect -5659 33660 -5561 33697
rect -5598 33403 -5561 33660
rect -6046 33402 -5870 33403
rect -5681 33402 -5561 33403
rect -6046 33368 -5561 33402
rect -6046 33364 -5870 33368
rect -5681 33366 -5561 33368
rect -6046 32697 -5993 33364
rect -5865 33136 -5729 33139
rect -4857 33136 -4664 34508
rect -5865 33021 -4664 33136
rect -5865 33016 -5729 33021
rect -6055 32693 -5959 32697
rect -6055 32689 -5873 32693
rect -6055 32655 -5674 32689
rect -6055 32650 -5873 32655
rect -6055 32384 -5959 32650
rect -5086 32689 -4895 32696
rect -5276 32655 -4895 32689
rect -5086 32650 -4895 32655
rect -4964 32567 -4895 32650
rect -4857 32567 -4664 33021
rect -6055 32380 -5875 32384
rect -6055 32346 -5674 32380
rect -6055 32341 -5875 32346
rect -6055 32065 -5959 32341
rect -5590 32327 -5536 32466
rect -4964 32499 -4664 32567
rect -5098 32493 -4664 32499
rect -5276 32459 -4664 32493
rect -5098 32453 -4664 32459
rect -4964 32386 -4664 32453
rect -5088 32380 -4664 32386
rect -5276 32346 -4664 32380
rect -5088 32340 -4664 32346
rect -4964 32190 -4664 32340
rect -5093 32184 -4664 32190
rect -7907 30785 -7680 30819
rect -7907 30623 -7839 30785
rect -7217 30819 -7149 30981
rect -7508 30785 -7149 30819
rect -7907 30589 -7680 30623
rect -7907 30490 -7839 30589
rect -7217 30651 -7149 30785
rect -6046 30903 -5993 32065
rect -5276 32150 -4664 32184
rect -5093 32144 -4664 32150
rect -4964 32077 -4664 32144
rect -5089 32070 -4664 32077
rect -5276 32036 -4664 32070
rect -5089 32031 -4664 32036
rect -4964 31974 -4664 32031
rect -4964 31879 -4895 31974
rect -5093 31874 -4895 31879
rect -5276 31840 -4895 31874
rect -5093 31833 -4895 31840
rect -4964 31684 -4895 31833
rect -5093 31678 -4895 31684
rect -5276 31644 -4895 31678
rect -5882 31282 -5622 31316
rect -5680 31279 -5622 31282
rect -5659 31197 -5622 31279
rect -5584 31249 -5530 31388
rect -5659 31160 -5561 31197
rect -5598 30903 -5561 31160
rect -6046 30902 -5870 30903
rect -5681 30902 -5561 30903
rect -6046 30868 -5561 30902
rect -6046 30864 -5870 30868
rect -5681 30866 -5561 30868
rect -6453 30651 -6317 30655
rect -7217 30623 -6317 30651
rect -7508 30589 -6317 30623
rect -7217 30536 -6317 30589
rect -7217 30528 -7149 30536
rect -6453 30532 -6317 30536
rect -7993 30430 -7831 30431
rect -7993 30356 -7672 30430
rect -8173 29007 -8113 29010
rect -8287 28978 -8113 29007
rect -8446 28944 -8113 28978
rect -8287 28896 -8113 28944
rect -8977 28748 -8618 28782
rect -8977 28641 -8909 28748
rect -9973 28372 -8909 28641
rect -8287 28782 -8219 28896
rect -8173 28873 -8113 28896
rect -8446 28748 -8219 28782
rect -8287 28739 -8219 28748
rect -9973 28270 -9905 28372
rect -9968 27779 -9905 28270
rect -8977 28270 -8909 28372
rect -8977 27779 -8914 28270
rect -9968 27510 -8914 27779
rect -10663 27311 -10595 27410
rect -9968 27372 -9905 27510
rect -10663 27277 -10436 27311
rect -10663 27209 -10595 27277
rect -9973 27311 -9905 27372
rect -10264 27277 -9905 27311
rect -10750 27115 -10595 27209
rect -10750 27098 -10436 27115
rect -10750 26413 -10711 27098
rect -10663 27081 -10436 27098
rect -10663 26919 -10595 27081
rect -9973 27115 -9905 27277
rect -10264 27081 -9905 27115
rect -10663 26885 -10436 26919
rect -10663 26474 -10595 26885
rect -9973 26919 -9905 27081
rect -10264 26902 -9905 26919
rect -8977 27372 -8914 27510
rect -8977 27311 -8909 27372
rect -8977 27277 -8618 27311
rect -8977 27115 -8909 27277
rect -8287 27311 -8219 27410
rect -8446 27277 -8219 27311
rect -8287 27209 -8219 27277
rect -8171 27209 -8132 28873
rect -8977 27081 -8618 27115
rect -8977 26919 -8909 27081
rect -8287 27115 -8132 27209
rect -8446 27098 -8132 27115
rect -8446 27081 -8219 27098
rect -8977 26902 -8618 26919
rect -10264 26885 -8618 26902
rect -9973 26633 -8909 26885
rect -8554 26773 -8480 26941
rect -8287 26919 -8219 27081
rect -8446 26885 -8219 26919
rect -10663 26440 -10436 26474
rect -10763 26398 -10703 26413
rect -10663 26398 -10595 26440
rect -10763 26287 -10595 26398
rect -9973 26474 -9905 26633
rect -10264 26440 -9905 26474
rect -9973 26356 -9905 26440
rect -8977 26474 -8909 26633
rect -8543 26761 -8480 26773
rect -8543 26738 -8336 26761
rect -8542 26701 -8336 26738
rect -8977 26440 -8618 26474
rect -8977 26356 -8909 26440
rect -8287 26474 -8219 26885
rect -8446 26440 -8219 26474
rect -8287 26398 -8219 26440
rect -8171 26413 -8132 27098
rect -8179 26398 -8119 26413
rect -10763 26276 -10703 26287
rect -10663 26278 -10595 26287
rect -10750 26259 -10711 26276
rect -11202 26146 -10975 26180
rect -11736 25888 -11668 26086
rect -11043 26047 -10975 26146
rect -10663 26244 -10436 26278
rect -10663 26082 -10595 26244
rect -9973 26278 -8909 26356
rect -10264 26244 -8618 26278
rect -10663 26048 -10436 26082
rect -10663 26039 -10595 26048
rect -9973 26087 -8909 26244
rect -8287 26287 -8119 26398
rect -8287 26278 -8219 26287
rect -8446 26244 -8219 26278
rect -8179 26276 -8119 26287
rect -8171 26259 -8132 26276
rect -7993 26797 -7954 30356
rect -7212 29594 -7149 30528
rect -6046 30197 -5993 30864
rect -5865 30653 -5729 30656
rect -4857 30653 -4664 31974
rect -5865 30539 -4664 30653
rect -5865 30533 -5729 30539
rect -6055 30193 -5959 30197
rect -6055 30189 -5873 30193
rect -6055 30155 -5674 30189
rect -6055 30150 -5873 30155
rect -6055 29884 -5959 30150
rect -5086 30189 -4895 30196
rect -5276 30155 -4895 30189
rect -5086 30150 -4895 30155
rect -6055 29880 -5875 29884
rect -6055 29846 -5674 29880
rect -6055 29841 -5875 29846
rect -7907 29272 -7839 29281
rect -7907 29238 -7680 29272
rect -7907 29076 -7839 29238
rect -7216 29281 -7148 29594
rect -6055 29565 -5959 29841
rect -5590 29827 -5536 29966
rect -4964 30051 -4895 30150
rect -4857 30051 -4664 30539
rect -4964 29999 -4664 30051
rect -5098 29993 -4664 29999
rect -5276 29959 -4664 29993
rect -5098 29953 -4664 29959
rect -4964 29886 -4664 29953
rect -5088 29880 -4664 29886
rect -5276 29846 -4664 29880
rect -5088 29840 -4664 29846
rect -4964 29690 -4664 29840
rect -5093 29684 -4664 29690
rect -7217 29272 -7148 29281
rect -7508 29238 -7148 29272
rect -7907 29042 -7680 29076
rect -7907 28880 -7839 29042
rect -7217 29121 -7148 29238
rect -7217 29076 -7149 29121
rect -7508 29042 -7149 29076
rect -7907 28846 -7680 28880
rect -7907 28315 -7839 28846
rect -7217 28880 -7149 29042
rect -7508 28846 -7149 28880
rect -7907 28281 -7680 28315
rect -7907 28119 -7839 28281
rect -7217 28315 -7149 28846
rect -6046 28403 -5993 29565
rect -5276 29650 -4664 29684
rect -5093 29644 -4664 29650
rect -4964 29577 -4664 29644
rect -5089 29570 -4664 29577
rect -5276 29536 -4664 29570
rect -5089 29531 -4664 29536
rect -4964 29458 -4664 29531
rect -4964 29379 -4895 29458
rect -5093 29374 -4895 29379
rect -5276 29340 -4895 29374
rect -5093 29333 -4895 29340
rect -4964 29184 -4895 29333
rect -5093 29178 -4895 29184
rect -5276 29144 -4895 29178
rect -5882 28782 -5622 28816
rect -5680 28779 -5622 28782
rect -5659 28697 -5622 28779
rect -5584 28749 -5530 28888
rect -5659 28660 -5561 28697
rect -5598 28403 -5561 28660
rect -6046 28402 -5870 28403
rect -5681 28402 -5561 28403
rect -6046 28368 -5561 28402
rect -6046 28364 -5870 28368
rect -5681 28366 -5561 28368
rect -7508 28281 -7149 28315
rect -7907 28085 -7680 28119
rect -7907 27923 -7839 28085
rect -7217 28119 -7149 28281
rect -7508 28085 -7149 28119
rect -6597 28085 -6461 28088
rect -7907 27889 -7680 27923
rect -7907 27790 -7839 27889
rect -7217 27970 -6461 28085
rect -7217 27923 -7149 27970
rect -6597 27965 -6461 27970
rect -7508 27889 -7149 27923
rect -7217 27828 -7149 27889
rect -7212 26903 -7149 27828
rect -8001 26665 -7941 26797
rect -7214 26765 -7146 26903
rect -6045 27697 -5958 28364
rect -5830 28086 -5694 28089
rect -4857 28086 -4664 29458
rect -5830 27971 -4664 28086
rect -5830 27966 -5694 27971
rect -6055 27693 -5958 27697
rect -6055 27689 -5873 27693
rect -6055 27655 -5674 27689
rect -6055 27650 -5873 27655
rect -6055 27576 -5958 27650
rect -4857 27696 -4664 27971
rect -5086 27689 -4664 27696
rect -5276 27655 -4664 27689
rect -5086 27650 -4664 27655
rect -6055 27384 -5959 27576
rect -6055 27380 -5875 27384
rect -6055 27346 -5674 27380
rect -6055 27341 -5875 27346
rect -6055 27065 -5959 27341
rect -4964 27499 -4664 27650
rect -5098 27493 -4664 27499
rect -5276 27459 -4664 27493
rect -5098 27453 -4664 27459
rect -4964 27386 -4664 27453
rect -5088 27380 -4664 27386
rect -5276 27346 -4664 27380
rect -5088 27340 -4664 27346
rect -4964 27190 -4664 27340
rect -5093 27184 -4664 27190
rect -6046 26830 -5993 27065
rect -6756 26765 -6688 26791
rect -7214 26731 -6688 26765
rect -7214 26697 -6397 26731
rect -7993 26259 -7954 26665
rect -7907 26572 -7839 26581
rect -7907 26538 -7680 26572
rect -7907 26376 -7839 26538
rect -7214 26677 -6688 26697
rect -7214 26583 -7146 26677
rect -6756 26583 -6688 26677
rect -6066 26731 -5993 26830
rect -6225 26697 -5993 26731
rect -7214 26581 -6688 26583
rect -7217 26572 -6688 26581
rect -7508 26538 -6688 26572
rect -7217 26535 -6688 26538
rect -7217 26501 -6397 26535
rect -7217 26495 -6688 26501
rect -7907 26342 -7680 26376
rect -9973 26082 -9905 26087
rect -10264 26048 -9905 26082
rect -9973 25889 -9905 26048
rect -8977 26082 -8909 26087
rect -8977 26048 -8618 26082
rect -9973 25888 -9816 25889
rect -8977 25888 -8909 26048
rect -8287 26082 -8219 26244
rect -8446 26048 -8219 26082
rect -8287 26039 -8219 26048
rect -7907 26180 -7839 26342
rect -7217 26400 -7146 26495
rect -6756 26400 -6688 26495
rect -6066 26535 -5993 26697
rect -6225 26501 -5993 26535
rect -7217 26376 -6688 26400
rect -7508 26342 -6688 26376
rect -7217 26339 -6688 26342
rect -7217 26312 -6397 26339
rect -7907 26146 -7680 26180
rect -7907 26047 -7839 26146
rect -7217 26180 -7146 26312
rect -6756 26305 -6397 26312
rect -6756 26296 -6688 26305
rect -7508 26146 -7146 26180
rect -6333 26173 -6259 26361
rect -6066 26339 -5993 26501
rect -6225 26305 -5993 26339
rect -6066 26296 -5993 26305
rect -7217 26086 -7146 26146
rect -7214 25888 -7146 26086
rect -11736 25799 -7146 25888
rect -6046 25903 -5993 26296
rect -5276 27150 -4664 27184
rect -5093 27144 -4664 27150
rect -4964 27077 -4664 27144
rect -5089 27070 -4664 27077
rect -5276 27036 -4664 27070
rect -5089 27031 -4664 27036
rect -4964 26879 -4664 27031
rect -5093 26874 -4664 26879
rect -5276 26840 -4664 26874
rect -5093 26833 -4664 26840
rect -4964 26684 -4664 26833
rect -5093 26678 -4664 26684
rect -5276 26644 -4664 26678
rect -5882 26282 -5622 26316
rect -5680 26279 -5622 26282
rect -5659 26197 -5622 26279
rect -5659 26160 -5561 26197
rect -5598 25903 -5561 26160
rect -6046 25902 -5870 25903
rect -5681 25902 -5561 25903
rect -6046 25868 -5561 25902
rect -6046 25864 -5870 25868
rect -5681 25866 -5561 25868
rect -11220 25589 -11125 25694
rect -11213 25125 -11131 25589
rect -11213 25118 -11012 25125
rect -11213 25084 -10718 25118
rect -11213 25078 -11012 25084
rect -11213 24929 -11131 25078
rect -11213 24922 -11011 24929
rect -11213 24888 -10718 24922
rect -11213 24882 -11011 24888
rect -11213 24687 -11131 24882
rect -9701 25221 -9616 25799
rect -9824 25216 -9616 25221
rect -10414 25182 -9616 25216
rect -9824 25176 -9616 25182
rect -9701 25026 -9616 25176
rect -9821 25020 -9616 25026
rect -10414 24986 -9616 25020
rect -9821 24981 -9616 24986
rect -11213 24680 -11001 24687
rect -11213 24646 -10718 24680
rect -11213 24640 -11001 24646
rect -11213 24460 -11131 24640
rect -9701 24604 -9616 24981
rect -9822 24597 -9616 24604
rect -10414 24563 -9616 24597
rect -9822 24559 -9616 24563
rect -11466 24023 -11398 24032
rect -11466 23989 -11107 24023
rect -11466 23827 -11398 23989
rect -10776 24023 -10708 24032
rect -10935 23989 -10708 24023
rect -11466 23793 -11107 23827
rect -11466 23631 -11398 23793
rect -10776 23827 -10708 23989
rect -10935 23793 -10708 23827
rect -11466 23597 -11107 23631
rect -11466 23141 -11398 23597
rect -10776 23631 -10708 23793
rect -10935 23597 -10708 23631
rect -11466 23107 -11107 23141
rect -11466 22945 -11398 23107
rect -10776 23141 -10708 23597
rect -10935 23107 -10708 23141
rect -11466 22911 -11107 22945
rect -11466 22749 -11398 22911
rect -10776 22945 -10708 23107
rect -10935 22911 -10708 22945
rect -11466 22715 -11107 22749
rect -11466 22654 -11398 22715
rect -10776 22749 -10708 22911
rect -10935 22715 -10708 22749
rect -11466 21720 -11403 22654
rect -10776 22616 -10708 22715
rect -11467 21407 -11399 21720
rect -11467 21398 -11398 21407
rect -11467 21364 -11107 21398
rect -11467 21247 -11398 21364
rect -10776 21398 -10708 21407
rect -10935 21364 -10708 21398
rect -11466 21202 -11398 21247
rect -11466 21168 -11107 21202
rect -11466 21006 -11398 21168
rect -10776 21202 -10708 21364
rect -10935 21168 -10708 21202
rect -11466 20972 -11107 21006
rect -11466 20441 -11398 20972
rect -10776 21006 -10708 21168
rect -10935 20972 -10708 21006
rect -11466 20407 -11107 20441
rect -11466 20245 -11398 20407
rect -10776 20441 -10708 20972
rect -10935 20407 -10708 20441
rect -11466 20211 -11107 20245
rect -11466 20049 -11398 20211
rect -10776 20245 -10708 20407
rect -10935 20211 -10708 20245
rect -11466 20015 -11107 20049
rect -11466 19954 -11398 20015
rect -10776 20049 -10708 20211
rect -10935 20015 -10708 20049
rect -11466 19029 -11403 19954
rect -10776 19916 -10708 20015
rect -11469 18707 -11401 19029
rect -10483 23769 -10444 23770
rect -10502 23637 -10442 23769
rect -10483 22011 -10444 23637
rect -10396 22137 -10328 22236
rect -9701 22198 -9616 24559
rect -6279 25098 -6197 25180
rect -6279 25091 -6078 25098
rect -6279 25057 -5784 25091
rect -6279 25051 -6078 25057
rect -6279 24902 -6197 25051
rect -6279 24895 -6077 24902
rect -6279 24861 -5784 24895
rect -6279 24855 -6077 24861
rect -6279 24660 -6197 24855
rect -4857 25281 -4664 26644
rect -4857 25279 -4675 25281
rect -4764 25194 -4675 25279
rect -4890 25189 -4675 25194
rect -5480 25155 -4675 25189
rect -4890 25149 -4675 25155
rect -4764 24999 -4675 25149
rect -4887 24993 -4675 24999
rect -5480 24959 -4675 24993
rect -4887 24954 -4675 24959
rect -6279 24653 -6067 24660
rect -6279 24619 -5784 24653
rect -6279 24613 -6067 24619
rect -6279 24467 -6197 24613
rect -4764 24577 -4675 24954
rect -4888 24570 -4675 24577
rect -5480 24536 -4675 24570
rect -4888 24532 -4675 24536
rect -6279 24189 -6196 24467
rect -10396 22103 -10169 22137
rect -10396 22011 -10328 22103
rect -9706 22137 -9616 22198
rect -9997 22103 -9616 22137
rect -10483 21941 -10328 22011
rect -9706 22003 -9616 22103
rect -10483 21907 -10169 21941
rect -10483 21900 -10328 21907
rect -10483 21136 -10444 21900
rect -10396 21745 -10328 21900
rect -9706 21941 -9638 22003
rect -9997 21907 -9638 21941
rect -10396 21725 -10169 21745
rect -10398 21711 -10169 21725
rect -10398 21702 -10328 21711
rect -10398 21399 -10330 21702
rect -9706 21745 -9638 21907
rect -9997 21711 -9638 21745
rect -10398 21300 -10328 21399
rect -10398 21266 -10169 21300
rect -10398 21205 -10328 21266
rect -9706 21300 -9638 21711
rect -9997 21266 -9638 21300
rect -10502 21133 -10442 21136
rect -10396 21133 -10328 21205
rect -10502 21104 -10328 21133
rect -10502 21070 -10169 21104
rect -10502 21022 -10328 21070
rect -10502 20999 -10442 21022
rect -11469 18698 -11398 18707
rect -11469 18664 -11107 18698
rect -11469 18502 -11398 18664
rect -10776 18698 -10708 18707
rect -10935 18664 -10708 18698
rect -11469 18468 -11107 18502
rect -11469 18306 -11398 18468
rect -10776 18502 -10708 18664
rect -10935 18468 -10708 18502
rect -11469 18272 -11107 18306
rect -11469 18212 -11398 18272
rect -10776 18306 -10708 18468
rect -10483 19335 -10444 20999
rect -10396 20908 -10328 21022
rect -9706 21104 -9638 21266
rect -9997 21070 -9638 21104
rect -9081 21135 -8995 21550
rect -8550 21429 -8451 21477
rect -8716 21395 -8451 21429
rect -6539 24023 -6471 24032
rect -6539 23989 -6180 24023
rect -6539 23827 -6471 23989
rect -5849 24023 -5781 24032
rect -6008 23989 -5781 24023
rect -6539 23793 -6180 23827
rect -6539 23631 -6471 23793
rect -5849 23827 -5781 23989
rect -6008 23793 -5781 23827
rect -6539 23597 -6180 23631
rect -6539 23141 -6471 23597
rect -5849 23631 -5781 23793
rect -6008 23597 -5781 23631
rect -6539 23107 -6180 23141
rect -6539 22945 -6471 23107
rect -5849 23141 -5781 23597
rect -6008 23107 -5781 23141
rect -6539 22911 -6180 22945
rect -6539 22749 -6471 22911
rect -5849 22945 -5781 23107
rect -6008 22911 -5781 22945
rect -6539 22715 -6180 22749
rect -6539 22654 -6471 22715
rect -5849 22749 -5781 22911
rect -6008 22715 -5781 22749
rect -6539 21720 -6476 22654
rect -5849 22616 -5781 22715
rect -8550 21233 -8451 21395
rect -8280 21303 -8214 21404
rect -8280 21300 -8090 21303
rect -8716 21199 -8451 21233
rect -9081 21101 -8839 21135
rect -9081 21070 -8995 21101
rect -10396 20874 -10169 20908
rect -10396 20865 -10328 20874
rect -9706 20908 -9638 21070
rect -9997 20874 -9638 20908
rect -9706 20396 -9638 20874
rect -9549 21009 -8995 21070
rect -8550 21037 -8451 21199
rect -9549 20700 -9488 21009
rect -9081 20939 -8995 21009
rect -8716 21003 -8451 21037
rect -9081 20905 -8839 20939
rect -9081 20765 -8995 20905
rect -8550 20841 -8451 21003
rect -8716 20807 -8451 20841
rect -10396 19437 -10328 19536
rect -9701 19498 -9638 20396
rect -9577 20620 -9488 20700
rect -9577 20330 -9491 20620
rect -9577 20296 -9146 20330
rect -9577 20295 -9454 20296
rect -9577 20121 -9491 20295
rect -8550 20630 -8451 20807
rect -8391 21299 -8090 21300
rect -8391 21265 -7498 21299
rect -8391 21258 -8090 21265
rect -8391 20881 -8214 21258
rect -6782 21222 -6669 21487
rect -6540 21407 -6472 21720
rect -6540 21398 -6471 21407
rect -6540 21364 -6180 21398
rect -6540 21247 -6471 21364
rect -5849 21398 -5781 21407
rect -6008 21364 -5781 21398
rect -6911 21216 -6669 21222
rect -7194 21182 -6669 21216
rect -6911 21175 -6669 21182
rect -8391 20876 -8091 20881
rect -8391 20842 -7498 20876
rect -8391 20836 -8091 20842
rect -8391 20805 -8214 20836
rect -8408 20686 -8214 20805
rect -8408 20680 -8088 20686
rect -8408 20646 -7498 20680
rect -8408 20641 -8088 20646
rect -8408 20635 -8214 20641
rect -8408 20630 -8238 20635
rect -8550 20624 -8238 20630
rect -8917 20590 -8238 20624
rect -8500 20428 -8238 20590
rect -6782 20980 -6669 21175
rect -6901 20974 -6669 20980
rect -7194 20940 -6669 20974
rect -6901 20933 -6669 20940
rect -6782 20784 -6669 20933
rect -6900 20778 -6669 20784
rect -7194 20744 -6669 20778
rect -6900 20737 -6669 20744
rect -8917 20394 -8238 20428
rect -9577 20035 -9324 20121
rect -10396 19403 -10169 19437
rect -10396 19335 -10328 19403
rect -9706 19437 -9638 19498
rect -9997 19403 -9638 19437
rect -10483 19241 -10328 19335
rect -10483 19224 -10169 19241
rect -10483 18539 -10444 19224
rect -10396 19207 -10169 19224
rect -10396 19045 -10328 19207
rect -9706 19241 -9638 19403
rect -9997 19207 -9638 19241
rect -10396 19011 -10169 19045
rect -10396 18600 -10328 19011
rect -9706 19045 -9638 19207
rect -9410 19553 -9324 20035
rect -8500 20232 -8238 20394
rect -8917 20198 -8238 20232
rect -8500 20188 -8238 20198
rect -8437 20187 -8238 20188
rect -8680 19847 -8581 19895
rect -8946 19813 -8581 19847
rect -8680 19651 -8581 19813
rect -8946 19617 -8581 19651
rect -9410 19519 -9068 19553
rect -8680 19531 -8581 19617
rect -8391 19817 -8238 20187
rect -8175 20430 -8076 20478
rect -8175 20396 -7910 20430
rect -8175 20234 -8076 20396
rect -8175 20200 -7910 20234
rect -8175 20038 -8076 20200
rect -7631 20136 -7545 20381
rect -7787 20102 -7545 20136
rect -7631 20071 -7545 20102
rect -6782 20071 -6669 20737
rect -8175 20004 -7910 20038
rect -7631 20010 -6669 20071
rect -6539 21202 -6471 21247
rect -6539 21168 -6180 21202
rect -6539 21006 -6471 21168
rect -5849 21202 -5781 21364
rect -6008 21168 -5781 21202
rect -6539 20972 -6180 21006
rect -6539 20441 -6471 20972
rect -5849 21006 -5781 21168
rect -6008 20972 -5781 21006
rect -6539 20407 -6180 20441
rect -6539 20245 -6471 20407
rect -5849 20441 -5781 20972
rect -6008 20407 -5781 20441
rect -6539 20211 -6180 20245
rect -6539 20049 -6471 20211
rect -5849 20245 -5781 20407
rect -6008 20211 -5781 20245
rect -6539 20015 -6180 20049
rect -8175 19842 -8076 20004
rect -7631 19940 -7545 20010
rect -7787 19906 -7545 19940
rect -8391 19628 -8224 19817
rect -8175 19808 -7910 19842
rect -8175 19631 -8076 19808
rect -7631 19766 -7545 19906
rect -8391 19591 -8231 19628
rect -8190 19625 -8076 19631
rect -8190 19591 -7709 19625
rect -8391 19531 -8238 19591
rect -9410 19357 -9324 19519
rect -8680 19455 -8238 19531
rect -8946 19421 -8238 19455
rect -8680 19359 -8238 19421
rect -9410 19323 -9068 19357
rect -9410 19183 -9324 19323
rect -9040 19205 -8980 19278
rect -8680 19259 -8581 19359
rect -8946 19225 -8581 19259
rect -9034 19161 -8993 19205
rect -8680 19177 -8581 19225
rect -9997 19011 -9638 19045
rect -9126 19031 -8976 19161
rect -10396 18566 -10169 18600
rect -10496 18524 -10436 18539
rect -10396 18524 -10328 18566
rect -10496 18413 -10328 18524
rect -9706 18600 -9638 19011
rect -9997 18566 -9638 18600
rect -9706 18540 -9638 18566
rect -8391 18540 -8238 19359
rect -8190 19429 -8126 19591
rect -7588 19579 -7517 19653
rect -7138 19628 -7077 20010
rect -6539 19954 -6471 20015
rect -5849 20049 -5781 20211
rect -6008 20015 -5781 20049
rect -7138 19621 -7059 19628
rect -8190 19395 -7709 19429
rect -8190 19233 -8126 19395
rect -8190 19199 -7709 19233
rect -8190 19189 -8126 19199
rect -7562 19238 -7523 19579
rect -7120 19331 -7059 19621
rect -7480 19297 -7059 19331
rect -7172 19296 -7059 19297
rect -7562 19168 -7522 19238
rect -7120 19179 -7059 19296
rect -7564 19167 -7522 19168
rect -7564 18941 -7524 19167
rect -6539 19029 -6476 19954
rect -5849 19916 -5781 20015
rect -6542 18707 -6474 19029
rect -5556 23769 -5517 23770
rect -5575 23637 -5515 23769
rect -5556 22011 -5517 23637
rect -4764 23150 -4675 24532
rect -4774 22950 -4675 23150
rect -5469 22137 -5401 22236
rect -4774 22198 -4711 22950
rect -5469 22103 -5242 22137
rect -5469 22011 -5401 22103
rect -4779 22137 -4711 22198
rect -5070 22103 -4711 22137
rect -5556 21941 -5401 22011
rect -5556 21907 -5242 21941
rect -5556 21900 -5401 21907
rect -5556 21136 -5517 21900
rect -5469 21745 -5401 21900
rect -4779 21941 -4711 22103
rect -5070 21907 -4711 21941
rect -5469 21725 -5242 21745
rect -5471 21711 -5242 21725
rect -5471 21702 -5401 21711
rect -5471 21399 -5403 21702
rect -4779 21745 -4711 21907
rect -5070 21711 -4711 21745
rect -5471 21300 -5401 21399
rect -5471 21266 -5242 21300
rect -5471 21205 -5401 21266
rect -4779 21300 -4711 21711
rect -5070 21266 -4711 21300
rect -5575 21133 -5515 21136
rect -5469 21133 -5401 21205
rect -5575 21104 -5401 21133
rect -5575 21070 -5242 21104
rect -5575 21022 -5401 21070
rect -5575 20999 -5515 21022
rect -6542 18698 -6471 18707
rect -6542 18664 -6180 18698
rect -6542 18540 -6471 18664
rect -5849 18698 -5781 18707
rect -6008 18664 -5781 18698
rect -9706 18502 -6471 18540
rect -9706 18468 -6180 18502
rect -10496 18402 -10436 18413
rect -10396 18404 -10328 18413
rect -10483 18385 -10444 18402
rect -10935 18272 -10708 18306
rect -11469 18014 -11401 18212
rect -10776 18173 -10708 18272
rect -10396 18370 -10169 18404
rect -10396 18208 -10328 18370
rect -9706 18404 -6471 18468
rect -5849 18502 -5781 18664
rect -6008 18468 -5781 18502
rect -9997 18387 -6471 18404
rect -9997 18370 -9638 18387
rect -10396 18174 -10169 18208
rect -10396 18165 -10328 18174
rect -9706 18208 -9638 18370
rect -9997 18174 -9638 18208
rect -10498 18014 -10331 18015
rect -9706 18014 -9638 18174
rect -11469 17925 -9638 18014
rect -6542 18306 -6471 18387
rect -6542 18272 -6180 18306
rect -6542 18212 -6471 18272
rect -5849 18306 -5781 18468
rect -5556 19335 -5517 20999
rect -5469 20908 -5401 21022
rect -4779 21104 -4711 21266
rect -5070 21070 -4711 21104
rect -5469 20874 -5242 20908
rect -5469 20865 -5401 20874
rect -4779 20908 -4711 21070
rect -5070 20874 -4711 20908
rect -4779 20396 -4711 20874
rect -5469 19437 -5401 19536
rect -4774 19498 -4711 20396
rect -5469 19403 -5242 19437
rect -5469 19335 -5401 19403
rect -4779 19437 -4711 19498
rect -5070 19403 -4711 19437
rect -5556 19241 -5401 19335
rect -5556 19224 -5242 19241
rect -5556 18539 -5517 19224
rect -5469 19207 -5242 19224
rect -5469 19045 -5401 19207
rect -4779 19241 -4711 19403
rect -5070 19207 -4711 19241
rect -5469 19011 -5242 19045
rect -5469 18600 -5401 19011
rect -4779 19045 -4711 19207
rect -5070 19011 -4711 19045
rect -5469 18566 -5242 18600
rect -5569 18524 -5509 18539
rect -5469 18524 -5401 18566
rect -5569 18413 -5401 18524
rect -4779 18600 -4711 19011
rect -5070 18566 -4711 18600
rect -5569 18402 -5509 18413
rect -5469 18404 -5401 18413
rect -5556 18385 -5517 18402
rect -6008 18272 -5781 18306
rect -6542 18014 -6474 18212
rect -5849 18173 -5781 18272
rect -5469 18370 -5242 18404
rect -5469 18208 -5401 18370
rect -4779 18404 -4711 18566
rect -5070 18370 -4711 18404
rect -5469 18174 -5242 18208
rect -5469 18165 -5401 18174
rect -4779 18208 -4711 18370
rect -5070 18174 -4711 18208
rect -4779 18014 -4711 18174
rect -6542 17925 -4711 18014
rect -13105 16146 -13019 16561
rect -12574 16440 -12475 16488
rect -12740 16406 -12475 16440
rect -12574 16244 -12475 16406
rect -12304 16314 -12238 16415
rect -12304 16311 -12114 16314
rect -12740 16210 -12475 16244
rect -13105 16112 -12863 16146
rect -13105 16081 -13019 16112
rect -13573 16020 -13019 16081
rect -12574 16048 -12475 16210
rect -13573 15711 -13512 16020
rect -13105 15950 -13019 16020
rect -12740 16014 -12475 16048
rect -13105 15916 -12863 15950
rect -13105 15776 -13019 15916
rect -12574 15852 -12475 16014
rect -12740 15818 -12475 15852
rect -13601 15631 -13512 15711
rect -13601 15341 -13515 15631
rect -13601 15307 -13170 15341
rect -13601 15306 -13478 15307
rect -13601 15132 -13515 15306
rect -12574 15641 -12475 15818
rect -12415 16310 -12114 16311
rect -12415 16276 -11522 16310
rect -12415 16269 -12114 16276
rect -12415 15892 -12238 16269
rect -10806 16233 -10693 16498
rect -10935 16227 -10693 16233
rect -11218 16193 -10693 16227
rect -10935 16186 -10693 16193
rect -12415 15887 -12115 15892
rect -12415 15853 -11522 15887
rect -12415 15847 -12115 15853
rect -12415 15816 -12238 15847
rect -12432 15697 -12238 15816
rect -12432 15691 -12112 15697
rect -12432 15657 -11522 15691
rect -12432 15652 -12112 15657
rect -12432 15646 -12238 15652
rect -12432 15641 -12262 15646
rect -12574 15635 -12262 15641
rect -12941 15601 -12262 15635
rect -12524 15439 -12262 15601
rect -10806 15991 -10693 16186
rect -10925 15985 -10693 15991
rect -11218 15951 -10693 15985
rect -10925 15944 -10693 15951
rect -10806 15795 -10693 15944
rect -10924 15789 -10693 15795
rect -11218 15755 -10693 15789
rect -10924 15748 -10693 15755
rect -12941 15405 -12262 15439
rect -13601 15046 -13348 15132
rect -13434 14564 -13348 15046
rect -12524 15243 -12262 15405
rect -12941 15209 -12262 15243
rect -12524 15199 -12262 15209
rect -12461 15198 -12262 15199
rect -12704 14858 -12605 14906
rect -12970 14824 -12605 14858
rect -12704 14662 -12605 14824
rect -12970 14628 -12605 14662
rect -13434 14530 -13092 14564
rect -12704 14542 -12605 14628
rect -12415 14828 -12262 15198
rect -12199 15441 -12100 15489
rect -12199 15407 -11934 15441
rect -12199 15245 -12100 15407
rect -12199 15211 -11934 15245
rect -12199 15049 -12100 15211
rect -11655 15147 -11569 15392
rect -11811 15113 -11569 15147
rect -11655 15082 -11569 15113
rect -10806 15082 -10693 15748
rect -12199 15015 -11934 15049
rect -11655 15021 -10693 15082
rect -12199 14853 -12100 15015
rect -11655 14951 -11569 15021
rect -11811 14917 -11569 14951
rect -12415 14639 -12248 14828
rect -12199 14819 -11934 14853
rect -12199 14642 -12100 14819
rect -11655 14777 -11569 14917
rect -12415 14602 -12255 14639
rect -12214 14636 -12100 14642
rect -12214 14602 -11733 14636
rect -12415 14542 -12262 14602
rect -13434 14368 -13348 14530
rect -12704 14466 -12262 14542
rect -12970 14432 -12262 14466
rect -12704 14370 -12262 14432
rect -13434 14334 -13092 14368
rect -13434 14194 -13348 14334
rect -12704 14270 -12605 14370
rect -12970 14236 -12605 14270
rect -12704 14188 -12605 14236
rect -14060 11720 -13968 13140
rect -13516 13138 -13429 13140
rect -12434 13138 -12262 14370
rect -12214 14440 -12150 14602
rect -11162 14639 -11101 15021
rect -12214 14406 -11733 14440
rect -12214 14244 -12150 14406
rect -12214 14210 -11733 14244
rect -12214 14200 -12150 14210
rect -11162 14342 -11083 14639
rect -11504 14308 -11083 14342
rect -11196 14307 -11083 14308
rect -11162 14190 -11083 14307
rect -11162 13739 -11101 14190
rect -11581 13678 -11101 13739
rect -11896 13352 -11807 13370
rect -11581 13352 -11520 13678
rect -11896 13291 -11520 13352
rect -11896 13154 -11807 13291
rect -13516 12966 -12262 13138
rect -11957 13140 -11807 13154
rect -11957 13136 -11656 13140
rect -11957 13102 -11496 13136
rect -11957 13096 -11656 13102
rect -13516 12964 -13429 12966
rect -11957 12946 -11807 13096
rect -11381 13035 -11321 13178
rect -11957 12940 -11655 12946
rect -11957 12906 -11496 12940
rect -11957 12902 -11655 12906
rect -11957 12773 -11807 12902
rect -11461 12812 -11401 12958
rect -11453 12774 -11417 12812
rect -12650 12710 -12513 12768
rect -14060 11686 -13692 11720
rect -14060 11524 -13968 11686
rect -14060 11490 -13692 11524
rect -14060 11328 -13968 11490
rect -14060 11294 -13692 11328
rect -14060 11132 -13968 11294
rect -12796 11622 -12731 11720
rect -13293 11588 -12731 11622
rect -12796 11425 -12731 11588
rect -14060 11098 -13692 11132
rect -14060 10590 -13968 11098
rect -14060 10556 -13692 10590
rect -14060 10538 -13968 10556
rect -14051 10394 -13984 10538
rect -12815 10590 -12700 11425
rect -13192 10556 -12700 10590
rect -12815 10442 -12700 10556
rect -14051 10360 -13692 10394
rect -14051 10350 -13984 10360
rect -12650 10258 -12609 12710
rect -12746 10200 -12609 10258
rect -12573 12617 -12436 12675
rect -12573 10113 -12532 12617
rect -11957 12465 -11841 12773
rect -11542 12716 -11405 12774
rect -11364 12697 -11328 13035
rect -10694 13348 -10625 13350
rect -10498 13348 -10331 17925
rect -10694 13046 -10331 13348
rect -10827 13038 -10331 13046
rect -11212 13004 -10331 13038
rect -10827 12998 -10331 13004
rect -10694 12849 -10331 12998
rect -10821 12842 -10331 12849
rect -11212 12808 -10331 12842
rect -10821 12801 -10331 12808
rect -10694 12796 -10331 12801
rect -10666 12795 -10331 12796
rect -11370 12639 -11233 12697
rect -11957 12235 -11806 12465
rect -11957 12231 -11655 12235
rect -11957 12197 -11495 12231
rect -11957 12191 -11655 12197
rect -11957 12041 -11806 12191
rect -11380 12130 -11320 12273
rect -11957 12035 -11654 12041
rect -11957 12001 -11495 12035
rect -11957 11997 -11654 12001
rect -11957 11868 -11806 11997
rect -11460 11907 -11400 12053
rect -12494 11796 -12357 11854
rect -12668 10055 -12531 10113
rect -12494 9999 -12453 11796
rect -12415 11703 -12278 11761
rect -12587 9941 -12450 9999
rect -12415 9886 -12374 11703
rect -12261 11459 -12155 11543
rect -12288 11429 -12138 11459
rect -11957 11429 -11841 11868
rect -11452 11856 -11416 11907
rect -11540 11798 -11403 11856
rect -11363 11781 -11327 12130
rect -10693 12424 -10624 12445
rect -10498 12424 -10331 12795
rect -10693 12141 -10331 12424
rect -10826 12133 -10331 12141
rect -11211 12099 -10331 12133
rect -10826 12093 -10331 12099
rect -10693 11944 -10331 12093
rect -10820 11937 -10331 11944
rect -11211 11906 -10331 11937
rect -11211 11903 -10624 11906
rect -10820 11896 -10624 11903
rect -10693 11891 -10624 11896
rect -11369 11723 -11232 11781
rect -12288 11313 -11841 11429
rect -12288 11032 -12138 11313
rect -11691 11318 -11635 11403
rect -11691 11258 -11589 11318
rect -12288 11025 -12006 11032
rect -12288 10991 -11838 11025
rect -12288 10984 -12006 10991
rect -12288 10838 -12138 10984
rect -11723 10938 -11667 11083
rect -12288 10829 -12009 10838
rect -12288 10795 -11838 10829
rect -12288 10790 -12009 10795
rect -12288 10655 -12138 10790
rect -11818 10609 -11762 10754
rect -12415 9828 -12278 9886
rect -11811 9790 -11770 10609
rect -12005 9730 -11768 9790
rect -11719 9680 -11678 10938
rect -11902 9620 -11665 9680
rect -11630 9489 -11589 11258
rect -10770 11530 -10637 11556
rect -10498 11530 -10331 11906
rect -10770 10937 -10331 11530
rect -10898 10927 -10331 10937
rect -11482 10893 -10331 10927
rect -10898 10884 -10331 10893
rect -10770 10748 -10331 10884
rect -10770 10741 -10637 10748
rect -10882 10731 -10637 10741
rect -11482 10697 -10637 10731
rect -10882 10688 -10637 10697
rect -10498 10378 -10331 10748
rect -11645 9429 -11408 9489
rect -8105 16146 -8019 16561
rect -7574 16440 -7475 16488
rect -7740 16406 -7475 16440
rect -7574 16244 -7475 16406
rect -7304 16314 -7238 16415
rect -7304 16311 -7114 16314
rect -7740 16210 -7475 16244
rect -8105 16112 -7863 16146
rect -8105 16081 -8019 16112
rect -8573 16020 -8019 16081
rect -7574 16048 -7475 16210
rect -8573 15711 -8512 16020
rect -8105 15950 -8019 16020
rect -7740 16014 -7475 16048
rect -8105 15916 -7863 15950
rect -8105 15776 -8019 15916
rect -7574 15852 -7475 16014
rect -7740 15818 -7475 15852
rect -8601 15631 -8512 15711
rect -8601 15341 -8515 15631
rect -8601 15307 -8170 15341
rect -8601 15306 -8478 15307
rect -8601 15292 -8515 15306
rect -8817 15132 -8515 15292
rect -7574 15641 -7475 15818
rect -7415 16310 -7114 16311
rect -7415 16276 -6522 16310
rect -7415 16269 -7114 16276
rect -7415 15892 -7238 16269
rect -5806 16233 -5693 16498
rect -5935 16227 -5693 16233
rect -6218 16193 -5693 16227
rect -5935 16186 -5693 16193
rect -7415 15887 -7115 15892
rect -7415 15853 -6522 15887
rect -7415 15847 -7115 15853
rect -7415 15816 -7238 15847
rect -7432 15697 -7238 15816
rect -7432 15691 -7112 15697
rect -7432 15657 -6522 15691
rect -7432 15652 -7112 15657
rect -7432 15646 -7238 15652
rect -7432 15641 -7262 15646
rect -7574 15635 -7262 15641
rect -7941 15601 -7262 15635
rect -7524 15439 -7262 15601
rect -5806 15991 -5693 16186
rect -5925 15985 -5693 15991
rect -6218 15951 -5693 15985
rect -5925 15944 -5693 15951
rect -5806 15795 -5693 15944
rect -5924 15789 -5693 15795
rect -6218 15755 -5693 15789
rect -5924 15748 -5693 15755
rect -7941 15405 -7262 15439
rect -8817 15082 -8348 15132
rect -8817 13569 -8662 15082
rect -8601 15046 -8348 15082
rect -8434 14564 -8348 15046
rect -7524 15243 -7262 15405
rect -7941 15209 -7262 15243
rect -7524 15199 -7262 15209
rect -7461 15198 -7262 15199
rect -7704 14858 -7605 14906
rect -7970 14824 -7605 14858
rect -7704 14662 -7605 14824
rect -7970 14628 -7605 14662
rect -8434 14530 -8092 14564
rect -7704 14542 -7605 14628
rect -7415 14828 -7262 15198
rect -7199 15441 -7100 15489
rect -7199 15407 -6934 15441
rect -7199 15245 -7100 15407
rect -7199 15211 -6934 15245
rect -7199 15049 -7100 15211
rect -6655 15147 -6569 15392
rect -6811 15113 -6569 15147
rect -6655 15082 -6569 15113
rect -5806 15082 -5693 15748
rect -7199 15015 -6934 15049
rect -6655 15021 -5693 15082
rect -7199 14853 -7100 15015
rect -6655 14951 -6569 15021
rect -6811 14917 -6569 14951
rect -7415 14639 -7248 14828
rect -7199 14819 -6934 14853
rect -7199 14642 -7100 14819
rect -6655 14777 -6569 14917
rect -7415 14602 -7255 14639
rect -7214 14636 -7100 14642
rect -7214 14602 -6733 14636
rect -7415 14542 -7262 14602
rect -8434 14368 -8348 14530
rect -7704 14466 -7262 14542
rect -7970 14432 -7262 14466
rect -7704 14370 -7262 14432
rect -8434 14334 -8092 14368
rect -8434 14194 -8348 14334
rect -7704 14270 -7605 14370
rect -7970 14236 -7605 14270
rect -7704 14188 -7605 14236
rect -7415 14200 -7262 14370
rect -7214 14440 -7150 14602
rect -6162 14639 -6101 15021
rect -7214 14406 -6733 14440
rect -7214 14244 -7150 14406
rect -7214 14210 -6733 14244
rect -7214 14200 -7150 14210
rect -7415 13775 -7302 14200
rect -6690 14125 -6636 14260
rect -6162 14342 -6083 14639
rect -6504 14308 -6083 14342
rect -6196 14307 -6083 14308
rect -6162 14190 -6083 14307
rect -6684 14105 -6644 14125
rect -6682 13848 -6646 14105
rect -7501 13765 -7302 13775
rect -7793 13731 -7302 13765
rect -8817 13535 -8293 13569
rect -8817 13334 -8662 13535
rect -7534 13569 -7302 13731
rect -7793 13535 -7302 13569
rect -8817 12537 -8689 13334
rect -7534 13027 -7302 13535
rect -7793 12993 -7302 13027
rect -8817 12503 -8192 12537
rect -8817 12405 -8689 12503
rect -8817 12223 -8692 12405
rect -7534 12831 -7302 12993
rect -7793 12797 -7302 12831
rect -8817 12108 -8559 12223
rect -7534 12635 -7302 12797
rect -7793 12601 -7302 12635
rect -7534 12439 -7302 12601
rect -7793 12405 -7302 12439
rect -8674 11504 -8559 12108
rect -8152 11569 -8066 11814
rect -7534 11911 -7302 12405
rect -7621 11863 -7302 11911
rect -7787 11829 -7302 11863
rect -7621 11667 -7302 11829
rect -7787 11633 -7302 11667
rect -8152 11535 -7910 11569
rect -8152 11504 -8066 11535
rect -8674 11443 -8066 11504
rect -7621 11471 -7302 11633
rect -8674 11054 -8559 11443
rect -8152 11373 -8066 11443
rect -7787 11437 -7302 11471
rect -8152 11339 -7910 11373
rect -8152 11199 -8066 11339
rect -7621 11275 -7302 11437
rect -7787 11241 -7302 11275
rect -8674 11053 -8577 11054
rect -8638 10764 -8577 11053
rect -8180 11012 -8109 11086
rect -8638 10730 -8217 10764
rect -8638 10729 -8525 10730
rect -8638 10612 -8577 10729
rect -8174 10671 -8135 11012
rect -7621 11058 -7302 11241
rect -7988 11024 -7302 11058
rect -7571 10862 -7302 11024
rect -7988 10828 -7302 10862
rect -8175 10601 -8135 10671
rect -8175 10600 -8133 10601
rect -8515 10114 -8278 10117
rect -8173 10114 -8133 10600
rect -8085 10547 -8031 10682
rect -7571 10666 -7302 10828
rect -7988 10632 -7302 10666
rect -7571 10622 -7302 10632
rect -8077 10527 -8037 10547
rect -8075 10260 -8039 10527
rect -8077 10200 -7840 10260
rect -8515 10074 -8133 10114
rect -8515 10057 -8278 10074
rect -7534 9234 -7302 10622
rect -7261 13791 -6646 13848
rect -7261 9382 -7198 13791
rect -6682 13714 -6646 13791
rect -6162 13775 -6101 14190
rect -6245 13714 -6101 13775
rect -6243 13511 -6157 13714
rect -5712 13849 -5613 13853
rect -5551 13849 -5338 17925
rect -5712 13805 -5338 13849
rect -5878 13771 -5338 13805
rect -5712 13609 -5338 13771
rect -5878 13575 -5338 13609
rect -6243 13477 -6001 13511
rect -6816 13446 -6664 13476
rect -6243 13446 -6157 13477
rect -6816 13385 -6157 13446
rect -5712 13413 -5338 13575
rect -6816 12996 -6650 13385
rect -6243 13315 -6157 13385
rect -5878 13379 -5338 13413
rect -6243 13281 -6001 13315
rect -6243 13141 -6157 13281
rect -5712 13217 -5338 13379
rect -5878 13183 -5338 13217
rect -6816 12706 -6664 12996
rect -6271 12954 -6200 13028
rect -6816 12672 -6308 12706
rect -6816 12671 -6616 12672
rect -7104 12245 -7051 12377
rect -7100 9888 -7060 12245
rect -7013 12229 -6881 12282
rect -7013 10002 -6977 12229
rect -6816 11849 -6664 12671
rect -6265 12613 -6226 12954
rect -5712 13000 -5338 13183
rect -6079 12966 -5338 13000
rect -5668 12804 -5338 12966
rect -6079 12770 -5338 12804
rect -6266 12543 -6226 12613
rect -6266 12542 -6224 12543
rect -6264 12491 -6224 12542
rect -6278 12354 -6220 12491
rect -6176 12489 -6122 12624
rect -5668 12608 -5338 12770
rect -6079 12574 -5338 12608
rect -5668 12522 -5338 12574
rect -6168 12469 -6128 12489
rect -6166 12396 -6130 12469
rect -6264 12316 -6224 12354
rect -6171 12259 -6113 12396
rect -5551 11945 -5338 12522
rect -5565 11935 -5338 11945
rect -5857 11901 -5338 11935
rect -6818 11739 -6664 11849
rect -6818 11705 -6357 11739
rect -6818 11520 -6664 11705
rect -5565 11739 -5338 11901
rect -5857 11705 -5338 11739
rect -5565 11700 -5338 11705
rect -6818 10707 -6753 11520
rect -5551 11197 -5338 11700
rect -6110 11022 -6056 11157
rect -5857 11163 -5338 11197
rect -6818 10673 -6256 10707
rect -6818 10575 -6753 10673
rect -7015 9941 -6799 10002
rect -6983 9888 -6943 9896
rect -7104 9828 -6867 9888
rect -6103 9490 -6069 11022
rect -6032 10834 -5978 10969
rect -5561 11001 -5338 11163
rect -5857 10967 -5338 11001
rect -6025 9681 -5987 10834
rect -5561 10805 -5338 10967
rect -5857 10771 -5338 10805
rect -5950 10498 -5896 10633
rect -5561 10609 -5338 10771
rect -5857 10575 -5338 10609
rect -5941 10479 -5904 10498
rect -5939 9790 -5904 10479
rect -5939 9729 -5701 9790
rect -6025 9620 -5787 9681
rect -6104 9429 -5866 9490
rect -7268 9281 -7025 9382
rect -5561 9234 -5338 10575
rect -7534 8962 -5338 9234
rect -2105 8544 -746 44258
rect 16949 13005 17282 16839
rect 16949 11350 17315 13005
rect 14597 10257 15867 10291
rect 14597 10215 14631 10257
rect 14469 9909 14662 10215
rect 15833 10167 15867 10257
rect 17125 10250 17315 11350
rect 17118 10172 17337 10250
rect 15584 10133 15867 10167
rect 16014 10138 16222 10172
rect 16814 10138 17337 10172
rect 14469 9875 14989 9909
rect 14469 9807 14662 9875
rect 3428 9393 14662 9807
rect 15833 9651 15867 10133
rect 15584 9617 15867 9651
rect 3428 9359 14989 9393
rect 3428 9172 14662 9359
rect -20516 4336 -14382 4472
rect -6647 7185 -745 8544
rect 3428 8200 4063 9172
rect 14469 9053 14662 9172
rect 15833 9135 15867 9617
rect 16014 9622 16222 9656
rect 17118 9656 17337 10138
rect 69244 10012 92336 10046
rect 69244 9682 69278 10012
rect 92302 9682 92336 10012
rect 69244 9668 92336 9682
rect 16814 9622 17337 9656
rect 15584 9101 15867 9135
rect 16014 9106 16222 9140
rect 15833 9006 15867 9101
rect 15722 8972 15890 9006
rect 16029 8972 16121 9006
rect 17118 9140 17337 9622
rect 16814 9106 17337 9140
rect 17118 8908 17337 9106
rect 69243 9648 92336 9668
rect 17125 8341 17315 8908
rect 69243 8878 92311 9648
rect 17671 8341 92311 8878
rect 3375 7918 4103 8200
rect 17125 8151 92311 8341
rect 3375 7840 8854 7918
rect 3375 7659 12714 7840
rect 3375 7565 4103 7659
rect 8144 7658 12714 7659
rect 14552 7821 14795 7846
rect 16664 7821 16961 7884
rect 14552 7685 16961 7821
rect -12975 6803 -11404 6943
rect -12975 5558 -2388 6803
rect -12975 5372 -11404 5558
rect -2105 4551 -746 7185
rect 8144 6692 8178 7658
rect 9860 6692 9894 7658
rect 11576 6692 11740 7658
rect 12622 6692 12656 7658
rect 14552 7642 14795 7685
rect 16664 7621 16961 7685
rect 17671 7646 92311 8151
rect 26753 7623 38073 7646
rect 2866 4551 3250 4560
rect 8180 4551 8214 6447
rect 9012 5496 9098 5582
rect 9038 4639 9072 5496
rect 9896 4551 9930 6447
rect 10711 5501 10837 5592
rect 10754 4639 10788 5501
rect 11612 4643 11646 6447
rect 14443 6151 14691 6213
rect 12023 6038 14691 6151
rect 12023 5710 12136 6038
rect 14443 6016 14691 6038
rect 11815 5565 12295 5710
rect 11612 4551 11647 4643
rect -2197 4085 12654 4551
rect 23929 4367 61121 4741
rect 23929 4290 98798 4367
rect 15817 4168 16331 4171
rect 23929 4168 24380 4290
rect 14819 3717 24380 4168
rect 25573 3778 26392 3779
rect 26583 3778 38866 3886
rect 14819 3692 15270 3717
rect -13207 3241 15270 3692
rect 21388 3591 21612 3717
rect 21003 3539 22224 3591
rect 20268 3533 20657 3534
rect 21003 3533 21130 3539
rect 19785 3465 21130 3533
rect 21567 3527 22102 3539
rect -13326 2204 -9322 2305
rect -2198 2250 -1747 3241
rect -13347 2138 -5909 2204
rect -2375 2198 -1154 2250
rect -3110 2192 -2721 2193
rect -2375 2192 -2248 2198
rect -12359 2066 -12300 2138
rect -11882 2066 -11823 2138
rect -11651 2066 -11592 2138
rect -11415 2066 -11356 2138
rect -11177 2066 -11118 2138
rect -10937 2066 -10878 2138
rect -10707 2066 -10648 2138
rect -10470 2066 -10411 2138
rect -10236 2066 -10177 2138
rect -10002 2066 -9943 2138
rect -9277 2066 -9218 2138
rect -9046 2066 -8987 2138
rect -8810 2066 -8751 2138
rect -8575 2066 -8516 2138
rect -8336 2066 -8277 2138
rect -8107 2066 -8048 2138
rect -7501 2066 -7442 2138
rect -7269 2066 -7210 2138
rect -7028 2066 -6969 2138
rect -6757 2066 -6698 2138
rect -6169 2066 -6110 2138
rect -3593 2124 -2248 2192
rect -1811 2186 -1276 2198
rect -13457 2018 -5905 2066
rect -13409 1425 -13375 1979
rect -13291 1571 -13257 2018
rect -13173 1571 -13139 1979
rect -13055 1571 -13021 2018
rect -12937 1571 -12903 1979
rect -12819 1571 -12785 2018
rect -12701 1571 -12667 1979
rect -12583 1571 -12549 2018
rect -12465 1571 -12431 1979
rect -12347 1571 -12313 2018
rect -12229 1571 -12195 1979
rect -12111 1571 -12077 2018
rect -11993 1571 -11959 1979
rect -11875 1571 -11841 2018
rect -11757 1571 -11723 1979
rect -11639 1571 -11605 2018
rect -11521 1571 -11487 1979
rect -11403 1571 -11369 2018
rect -11285 1571 -11251 1979
rect -11167 1571 -11133 2018
rect -11049 1571 -11015 1979
rect -10931 1571 -10897 2018
rect -10813 1571 -10779 1979
rect -10695 1571 -10661 2018
rect -10577 1571 -10543 1979
rect -10459 1571 -10425 2018
rect -10341 1571 -10307 1979
rect -10223 1571 -10189 2018
rect -10105 1571 -10071 1979
rect -9987 1571 -9953 2018
rect -9869 1571 -9835 1979
rect -9751 1571 -9717 2018
rect -9633 1571 -9599 1979
rect -9503 1571 -9469 2018
rect -22664 1391 -13375 1425
rect -9267 1571 -9233 2018
rect -9031 1571 -8997 2018
rect -8795 1571 -8761 2018
rect -8559 1571 -8525 2018
rect -8323 1571 -8289 2018
rect -8087 1571 -8053 2018
rect -7851 1571 -7817 2018
rect -7615 1571 -7581 2018
rect -7485 1571 -7451 2018
rect -7249 1571 -7215 2018
rect -7013 1571 -6979 2018
rect -6777 1571 -6743 2018
rect -6541 1571 -6507 2018
rect -6411 1571 -6377 2018
rect -6175 1571 -6141 2018
rect -5939 1571 -5905 2018
rect -3584 1833 -3550 2124
rect -3388 1833 -3354 2124
rect -3192 1833 -3158 2124
rect -2734 1833 -2700 2124
rect -2538 1833 -2504 2124
rect -2342 1833 -2308 2124
rect -3827 1695 -3528 1769
rect -9653 763 -9619 1171
rect -9417 763 -9383 1171
rect -9181 763 -9147 1171
rect -8945 763 -8911 1171
rect -8709 763 -8675 1171
rect -8473 763 -8439 1171
rect -8237 763 -8203 1171
rect -8001 763 -7967 1171
rect -3699 1090 -3647 1695
rect -2846 1090 -2678 1104
rect -3699 1038 -2678 1090
rect -18039 457 -17604 565
rect -6543 457 -5591 465
rect -22512 320 -5591 457
rect -6543 299 -5591 320
rect -3695 212 -3643 1038
rect -2846 1030 -2678 1038
rect -2734 675 -2700 966
rect -2538 675 -2504 966
rect -2342 675 -2308 966
rect -2088 1049 -2054 1312
rect -1892 1049 -1858 1312
rect -1696 1049 -1662 1312
rect -1500 1049 -1466 1312
rect -1304 1049 -1270 1312
rect -2088 1015 -1270 1049
rect -2088 758 -2054 1015
rect -1892 758 -1858 1015
rect -1696 758 -1662 1015
rect -1500 758 -1466 1015
rect -1304 758 -1270 1015
rect -2743 607 -2248 675
rect -2404 601 -2248 607
rect -1811 601 -1276 613
rect -1206 601 -1154 2198
rect 2820 2367 3099 2508
rect 6011 2426 6354 3241
rect 11748 2486 12550 3241
rect 18156 3110 18330 3181
rect 19794 3174 19828 3465
rect 19990 3174 20024 3465
rect 20186 3174 20220 3465
rect 20644 3174 20678 3465
rect 20840 3174 20874 3465
rect 21036 3174 21070 3465
rect 18156 3036 19850 3110
rect 18156 2985 18330 3036
rect 19567 2877 19632 2878
rect 19563 2800 19636 2877
rect 18629 2540 18739 2549
rect 19341 2540 19481 2579
rect 5724 2374 6945 2426
rect 7622 2420 15060 2486
rect 18629 2447 19481 2540
rect 18629 2441 18739 2447
rect 19341 2444 19481 2447
rect 4989 2368 5378 2369
rect 5724 2368 5851 2374
rect 565 2274 3099 2367
rect 4506 2300 5851 2368
rect 6288 2362 6823 2374
rect 565 2272 2965 2274
rect 591 2172 792 2272
rect 713 1997 747 2172
rect 1225 1986 1259 2272
rect 1515 1991 1549 2272
rect 2455 2172 2965 2272
rect 1947 1998 1981 2126
rect 713 1591 747 1825
rect 577 1576 795 1591
rect 1049 1576 1083 1823
rect 577 1539 1083 1576
rect 1225 1539 1259 1823
rect 2183 1998 2217 2126
rect 2500 1997 2534 2172
rect 1401 1576 1435 1823
rect 1690 1576 1724 1823
rect 1836 1576 1870 1823
rect 2809 1997 2843 2172
rect 2500 1591 2534 1825
rect 4515 2009 4549 2300
rect 4711 2009 4745 2300
rect 4907 2009 4941 2300
rect 5365 2009 5399 2300
rect 5561 2009 5595 2300
rect 5757 2009 5791 2300
rect 2809 1591 2843 1825
rect 2452 1576 2979 1591
rect 1401 1574 2979 1576
rect 3500 1574 3875 1654
rect 4272 1871 4571 1945
rect 1401 1539 3875 1574
rect 577 1323 3875 1539
rect 577 1286 1083 1323
rect 577 1271 795 1286
rect 713 1037 747 1271
rect 1049 1039 1083 1286
rect -2404 549 -1154 601
rect -2404 364 -2075 549
rect 1225 1039 1259 1323
rect 1401 1319 3875 1323
rect 1401 1286 2979 1319
rect 1401 1039 1435 1286
rect 1690 1039 1724 1286
rect 1836 1039 1870 1286
rect 2452 1271 2979 1286
rect 3500 1279 3875 1319
rect 713 690 747 865
rect 591 590 792 690
rect 1225 590 1259 876
rect 1515 590 1549 871
rect 2500 1037 2534 1271
rect 1947 736 1981 864
rect 2183 736 2217 864
rect 2809 1037 2843 1271
rect 2500 690 2534 865
rect 2809 690 2843 865
rect 2455 593 2965 690
rect 4196 595 4326 1504
rect 4400 1266 4452 1871
rect 4515 1678 4549 1837
rect 4711 1678 4745 1837
rect 4907 1678 4941 1837
rect 5365 1678 5399 1837
rect 5561 1678 5595 1837
rect 5757 1678 5791 1837
rect 4506 1610 5890 1678
rect 4626 1517 4768 1610
rect 4600 1392 4817 1517
rect 5356 1473 5890 1610
rect 5365 1314 5399 1473
rect 5253 1266 5421 1280
rect 4400 1243 5421 1266
rect 4388 1214 5421 1243
rect 4388 1066 4549 1214
rect 5253 1206 5421 1214
rect 5561 1314 5595 1473
rect 5757 1314 5791 1473
rect 5365 851 5399 1142
rect 5561 851 5595 1142
rect 5757 851 5791 1142
rect 6011 1225 6045 1488
rect 6207 1225 6241 1488
rect 6403 1225 6437 1488
rect 6599 1225 6633 1488
rect 6795 1225 6829 1488
rect 6011 1191 6829 1225
rect 6011 934 6045 1191
rect 6207 934 6241 1191
rect 6403 934 6437 1191
rect 6599 934 6633 1191
rect 6795 934 6829 1191
rect 5356 783 5851 851
rect 5724 777 5851 783
rect 6288 777 6823 789
rect 6893 777 6945 2374
rect 7823 2348 7882 2420
rect 8411 2348 8470 2420
rect 8682 2348 8741 2420
rect 8923 2348 8982 2420
rect 9155 2348 9214 2420
rect 9761 2348 9820 2420
rect 9990 2348 10049 2420
rect 10229 2348 10288 2420
rect 10464 2348 10523 2420
rect 10700 2348 10759 2420
rect 10931 2348 10990 2420
rect 11656 2348 11715 2420
rect 11890 2348 11949 2420
rect 12124 2348 12183 2420
rect 12361 2348 12420 2420
rect 12591 2348 12650 2420
rect 12831 2348 12890 2420
rect 13069 2348 13128 2420
rect 13305 2348 13364 2420
rect 13536 2348 13595 2420
rect 14013 2348 14072 2420
rect 7618 2300 15170 2348
rect 7618 1853 7652 2300
rect 7854 1853 7888 2300
rect 8090 1853 8124 2300
rect 8220 1853 8254 2300
rect 8456 1853 8490 2300
rect 8692 1853 8726 2300
rect 8928 1853 8962 2300
rect 9164 1853 9198 2300
rect 9294 1853 9328 2300
rect 9530 1853 9564 2300
rect 9766 1853 9800 2300
rect 10002 1853 10036 2300
rect 10238 1853 10272 2300
rect 10474 1853 10508 2300
rect 10710 1853 10744 2300
rect 10946 1853 10980 2300
rect 11182 1853 11216 2300
rect 11312 1853 11346 2261
rect 11430 1853 11464 2300
rect 11548 1853 11582 2261
rect 11666 1853 11700 2300
rect 11784 1853 11818 2261
rect 11902 1853 11936 2300
rect 12020 1853 12054 2261
rect 12138 1853 12172 2300
rect 12256 1853 12290 2261
rect 12374 1853 12408 2300
rect 12492 1853 12526 2261
rect 12610 1853 12644 2300
rect 12728 1853 12762 2261
rect 12846 1853 12880 2300
rect 12964 1853 12998 2261
rect 13082 1853 13116 2300
rect 13200 1853 13234 2261
rect 13318 1853 13352 2300
rect 13436 1853 13470 2261
rect 13554 1853 13588 2300
rect 13672 1853 13706 2261
rect 13790 1853 13824 2300
rect 13908 1853 13942 2261
rect 14026 1853 14060 2300
rect 14144 1853 14178 2261
rect 14262 1853 14296 2300
rect 14380 1853 14414 2261
rect 14498 1853 14532 2300
rect 14616 1853 14650 2261
rect 14734 1853 14768 2300
rect 14852 1853 14886 2261
rect 14970 1853 15004 2300
rect 15088 1707 15122 2261
rect 15522 1707 15742 1833
rect 15088 1673 15742 1707
rect 15522 1597 15742 1673
rect 11568 1517 15050 1545
rect 11420 1453 15050 1517
rect 7910 960 7944 1453
rect 8146 960 8180 1453
rect 8382 960 8416 1453
rect 8618 960 8652 1453
rect 8854 960 8888 1453
rect 9090 960 9124 1453
rect 9326 960 9360 1453
rect 9562 971 9596 1453
rect 9680 1045 9714 1453
rect 9394 960 9762 971
rect 9798 960 9832 1453
rect 9916 1045 9950 1453
rect 10034 960 10068 1453
rect 10152 1045 10186 1453
rect 10270 960 10304 1453
rect 10388 1045 10422 1453
rect 10506 960 10540 1453
rect 10624 1045 10658 1453
rect 10742 960 10776 1453
rect 10860 1045 10894 1453
rect 10978 960 11012 1453
rect 11096 1045 11130 1453
rect 11214 960 11248 1453
rect 11332 1045 11366 1453
rect 11450 960 11484 1453
rect 11568 1045 11602 1453
rect 11686 1045 11720 1453
rect 11804 1045 11838 1453
rect 11922 1045 11956 1453
rect 12040 1045 12074 1453
rect 12158 1045 12192 1453
rect 12276 1045 12310 1453
rect 12394 1045 12428 1453
rect 12512 1045 12546 1453
rect 12630 1045 12664 1453
rect 12748 1045 12782 1453
rect 12866 1045 12900 1453
rect 12984 1045 13018 1453
rect 13102 1045 13136 1453
rect 13220 1045 13254 1453
rect 13338 1045 13372 1453
rect 13456 1045 13490 1453
rect 13574 1045 13608 1453
rect 13692 1045 13726 1453
rect 13810 1045 13844 1453
rect 13928 1045 13962 1453
rect 14046 1045 14080 1453
rect 14164 1045 14198 1453
rect 14282 1045 14316 1453
rect 14400 1045 14434 1453
rect 14518 1045 14552 1453
rect 14636 1045 14670 1453
rect 14754 1045 14788 1453
rect 14872 1045 14906 1453
rect 14990 1045 15024 1453
rect 19567 1242 19632 2800
rect 19679 2431 19731 3036
rect 19794 2844 19828 3002
rect 19990 2844 20024 3002
rect 20186 2844 20220 3002
rect 19794 2843 20301 2844
rect 20644 2843 20678 3002
rect 20840 2843 20874 3002
rect 21036 2843 21070 3002
rect 19785 2775 21169 2843
rect 20635 2638 21169 2775
rect 20644 2479 20678 2638
rect 20532 2431 20700 2445
rect 19679 2379 20700 2431
rect 20532 2371 20700 2379
rect 20840 2479 20874 2638
rect 21036 2479 21070 2638
rect 20644 2016 20678 2307
rect 20840 2016 20874 2307
rect 21036 2016 21070 2307
rect 21290 2390 21324 2653
rect 21486 2390 21520 2653
rect 21682 2390 21716 2653
rect 21878 2390 21912 2653
rect 22074 2390 22108 2653
rect 21290 2356 22108 2390
rect 21290 2099 21324 2356
rect 21486 2099 21520 2356
rect 21682 2099 21716 2356
rect 21878 2099 21912 2356
rect 22074 2099 22108 2356
rect 20635 1948 21130 2016
rect 21003 1942 21130 1948
rect 21567 1942 22102 1954
rect 22172 1942 22224 3539
rect 25573 3484 47674 3778
rect 21003 1890 22224 1942
rect 19404 1241 19736 1242
rect 7868 840 15055 960
rect 19404 943 19770 1241
rect 5724 725 6945 777
rect 8203 744 8571 840
rect 9394 744 9762 840
rect 10640 744 11008 840
rect 12204 744 12572 840
rect 13329 744 13697 840
rect 14498 744 14866 840
rect 19404 744 19742 943
rect 5730 686 6208 725
rect 8089 595 19742 744
rect 3030 593 19742 595
rect 2455 590 19742 593
rect 565 495 19742 590
rect -22962 160 -3643 212
rect -3192 35 -2075 364
rect 2764 382 19742 495
rect 2764 336 3099 382
rect 15818 275 16268 345
rect 3985 213 4186 265
rect -1806 100 4186 213
rect -3192 -122 -2863 35
rect -3843 -174 -2622 -122
rect -4578 -180 -4189 -179
rect -3843 -180 -3716 -174
rect -5061 -248 -3716 -180
rect -3279 -186 -2744 -174
rect -5052 -539 -5018 -248
rect -4856 -539 -4822 -248
rect -4660 -539 -4626 -248
rect -4202 -539 -4168 -248
rect -4006 -539 -3972 -248
rect -3810 -539 -3776 -248
rect -22114 -677 -4996 -603
rect -5167 -1282 -5115 -677
rect -4314 -1282 -4146 -1268
rect -5167 -1334 -4146 -1282
rect -4314 -1342 -4146 -1334
rect -4202 -1697 -4168 -1406
rect -4006 -1697 -3972 -1406
rect -3810 -1697 -3776 -1406
rect -4211 -1765 -3716 -1697
rect -3843 -1771 -3716 -1765
rect -3279 -1771 -2744 -1759
rect -2674 -1771 -2622 -174
rect -3843 -1823 -2622 -1771
rect -1806 -1962 -1693 100
rect 3985 76 4186 100
rect 4383 -36 4585 -15
rect -1577 -85 4585 -36
rect -1581 -175 4585 -85
rect -1581 -342 -1323 -175
rect 4383 -213 4585 -175
rect 5857 -176 16268 275
rect 21288 241 21541 1890
rect 21915 241 22067 1890
rect 25573 1356 25868 3484
rect 26289 3483 47674 3484
rect 26688 2858 26963 2876
rect 26688 2669 28014 2858
rect 26688 2653 26963 2669
rect 27825 2314 28014 2669
rect 30305 2689 31641 2779
rect 33299 2689 33705 3483
rect 41815 3093 44205 3238
rect 41815 3091 45284 3093
rect 41489 3090 45284 3091
rect 39177 3027 45284 3090
rect 39177 3022 40555 3027
rect 41489 3023 43255 3027
rect 44180 3025 45284 3027
rect 41802 3022 43255 3023
rect 44502 3022 44997 3025
rect 35040 2689 36376 2801
rect 30305 2676 36376 2689
rect 30305 2654 35099 2676
rect 28132 2314 29133 2327
rect 27721 2309 29133 2314
rect 27721 2280 29505 2309
rect 27721 2106 27755 2280
rect 28132 2275 29505 2280
rect 28132 2262 29133 2275
rect 28336 2183 28377 2262
rect 28732 2183 28773 2262
rect 29471 2196 29505 2275
rect 28267 2149 29063 2183
rect 27721 2037 27914 2106
rect 27721 1464 27755 2037
rect 27879 1464 27913 2037
rect 28267 1853 28301 2149
rect 28583 1853 28617 2149
rect 29029 1858 29063 2149
rect 29359 2123 29505 2196
rect 29313 1858 29347 2066
rect 29471 1858 29505 2123
rect 30330 2092 30364 2654
rect 30646 2092 30680 2654
rect 30962 2092 30996 2654
rect 31120 2074 31154 2500
rect 31278 2074 31312 2654
rect 31594 2564 35099 2654
rect 31436 2074 31470 2500
rect 31594 2074 31628 2564
rect 32987 2307 33988 2320
rect 31120 2040 31628 2074
rect 32576 2302 33988 2307
rect 32576 2273 34360 2302
rect 32576 2099 32610 2273
rect 32987 2268 34360 2273
rect 32987 2255 33988 2268
rect 33191 2176 33232 2255
rect 33587 2176 33628 2255
rect 34326 2189 34360 2268
rect 33122 2142 33918 2176
rect 31169 1987 31572 2040
rect 32576 2030 32769 2099
rect 22419 876 25868 1356
rect 28267 1464 28301 1672
rect 28583 1464 28617 1672
rect 29029 1464 29063 1672
rect 29317 1463 29351 1671
rect 29475 1463 29509 1671
rect 30330 1286 30364 1844
rect 30646 1286 30680 1844
rect 30962 1286 30996 1844
rect 31278 1286 31312 1844
rect 31594 1286 31628 1844
rect 21175 189 22396 241
rect 20440 183 20829 184
rect 21175 183 21302 189
rect 19957 115 21302 183
rect 21739 177 22274 189
rect 19966 -176 20000 115
rect 5877 -264 6211 -176
rect 5739 -316 6960 -264
rect 8303 -270 8754 -176
rect 9891 -270 10342 -176
rect 11432 -270 11883 -176
rect 12650 -270 13101 -176
rect 13848 -270 14299 -176
rect 15818 -209 16268 -176
rect 20162 -176 20196 115
rect 20358 -176 20392 115
rect 20816 -176 20850 115
rect 21012 -176 21046 115
rect 21208 -176 21242 115
rect 5004 -322 5393 -321
rect 5739 -322 5866 -316
rect 4521 -390 5866 -322
rect 6303 -328 6838 -316
rect 3281 -745 3574 -645
rect 4530 -681 4564 -390
rect 4726 -681 4760 -390
rect 4922 -681 4956 -390
rect 5380 -681 5414 -390
rect 5576 -681 5610 -390
rect 5772 -681 5806 -390
rect 3281 -819 4586 -745
rect 3281 -911 3574 -819
rect 4415 -1424 4467 -819
rect 4530 -1012 4564 -853
rect 4726 -1012 4760 -853
rect 4922 -1012 4956 -853
rect 5380 -1012 5414 -853
rect 5576 -1012 5610 -853
rect 5772 -1012 5806 -853
rect 4521 -1080 5905 -1012
rect 5371 -1217 5905 -1080
rect 5380 -1376 5414 -1217
rect 5268 -1424 5436 -1410
rect 4415 -1476 5436 -1424
rect 5268 -1484 5436 -1476
rect 5576 -1376 5610 -1217
rect 5772 -1376 5806 -1217
rect 5380 -1839 5414 -1548
rect 5576 -1839 5610 -1548
rect 5772 -1839 5806 -1548
rect 6026 -1465 6060 -1202
rect 6222 -1465 6256 -1202
rect 6418 -1465 6452 -1202
rect 6614 -1465 6648 -1202
rect 6810 -1465 6844 -1202
rect 6026 -1499 6844 -1465
rect 6026 -1756 6060 -1499
rect 6222 -1756 6256 -1499
rect 6418 -1756 6452 -1499
rect 6614 -1756 6648 -1499
rect 6810 -1756 6844 -1499
rect 5371 -1907 5866 -1839
rect -26391 -2075 -1693 -1962
rect 5739 -1913 5866 -1907
rect 6303 -1913 6838 -1901
rect 6908 -1913 6960 -316
rect 7581 -336 15019 -270
rect 19723 -314 20022 -240
rect 7782 -408 7841 -336
rect 8370 -408 8429 -336
rect 8641 -408 8700 -336
rect 8882 -408 8941 -336
rect 9114 -408 9173 -336
rect 9720 -408 9779 -336
rect 9949 -408 10008 -336
rect 10188 -408 10247 -336
rect 10423 -408 10482 -336
rect 10659 -408 10718 -336
rect 10890 -408 10949 -336
rect 11615 -408 11674 -336
rect 11849 -408 11908 -336
rect 12083 -408 12142 -336
rect 12320 -408 12379 -336
rect 12550 -408 12609 -336
rect 12790 -408 12849 -336
rect 13028 -408 13087 -336
rect 13264 -408 13323 -336
rect 13495 -408 13554 -336
rect 13972 -408 14031 -336
rect 7577 -456 15129 -408
rect 7577 -903 7611 -456
rect 7813 -903 7847 -456
rect 8049 -903 8083 -456
rect 8179 -903 8213 -456
rect 8415 -903 8449 -456
rect 8651 -903 8685 -456
rect 8887 -903 8921 -456
rect 9123 -903 9157 -456
rect 9253 -903 9287 -456
rect 9489 -903 9523 -456
rect 9725 -903 9759 -456
rect 9961 -903 9995 -456
rect 10197 -903 10231 -456
rect 10433 -903 10467 -456
rect 10669 -903 10703 -456
rect 10905 -903 10939 -456
rect 11141 -903 11175 -456
rect 11271 -903 11305 -495
rect 11389 -903 11423 -456
rect 11507 -903 11541 -495
rect 11625 -903 11659 -456
rect 11743 -903 11777 -495
rect 11861 -903 11895 -456
rect 11979 -903 12013 -495
rect 12097 -903 12131 -456
rect 12215 -903 12249 -495
rect 12333 -903 12367 -456
rect 12451 -903 12485 -495
rect 12569 -903 12603 -456
rect 12687 -903 12721 -495
rect 12805 -903 12839 -456
rect 12923 -903 12957 -495
rect 13041 -903 13075 -456
rect 13159 -903 13193 -495
rect 13277 -903 13311 -456
rect 13395 -903 13429 -495
rect 13513 -903 13547 -456
rect 13631 -903 13665 -495
rect 13749 -903 13783 -456
rect 13867 -903 13901 -495
rect 13985 -903 14019 -456
rect 14103 -903 14137 -495
rect 14221 -903 14255 -456
rect 14339 -903 14373 -495
rect 14457 -903 14491 -456
rect 14575 -903 14609 -495
rect 14693 -903 14727 -456
rect 14811 -903 14845 -495
rect 14929 -903 14963 -456
rect 15047 -1021 15081 -495
rect 16101 -1021 16445 -871
rect 19851 -916 19903 -314
rect 19966 -507 20000 -348
rect 20162 -507 20196 -348
rect 20358 -507 20392 -348
rect 20816 -507 20850 -348
rect 21012 -507 21046 -348
rect 21208 -507 21242 -348
rect 19957 -575 21341 -507
rect 20807 -712 21341 -575
rect 20816 -871 20850 -712
rect 15047 -1127 16445 -1021
rect 11527 -1239 15009 -1211
rect 16101 -1228 16445 -1127
rect 19836 -919 20098 -916
rect 20704 -919 20872 -905
rect 19836 -971 20872 -919
rect 19836 -1129 20098 -971
rect 20704 -979 20872 -971
rect 21012 -871 21046 -712
rect 21208 -871 21242 -712
rect 11379 -1303 15009 -1239
rect 19836 -1279 20093 -1129
rect 7869 -1796 7903 -1303
rect 8105 -1796 8139 -1303
rect 8341 -1796 8375 -1303
rect 8577 -1796 8611 -1303
rect 8813 -1796 8847 -1303
rect 9049 -1796 9083 -1303
rect 9285 -1796 9319 -1303
rect 9521 -1796 9555 -1303
rect 9639 -1711 9673 -1303
rect 9757 -1796 9791 -1303
rect 9875 -1711 9909 -1303
rect 9993 -1796 10027 -1303
rect 10111 -1711 10145 -1303
rect 10229 -1796 10263 -1303
rect 10347 -1711 10381 -1303
rect 10465 -1796 10499 -1303
rect 10583 -1711 10617 -1303
rect 10701 -1796 10735 -1303
rect 10819 -1711 10853 -1303
rect 10937 -1796 10971 -1303
rect 11055 -1711 11089 -1303
rect 11173 -1796 11207 -1303
rect 11291 -1711 11325 -1303
rect 11409 -1796 11443 -1303
rect 11527 -1711 11561 -1303
rect 11645 -1711 11679 -1303
rect 11763 -1711 11797 -1303
rect 11881 -1711 11915 -1303
rect 11999 -1711 12033 -1303
rect 12117 -1711 12151 -1303
rect 12235 -1711 12269 -1303
rect 12353 -1711 12387 -1303
rect 12471 -1711 12505 -1303
rect 12589 -1711 12623 -1303
rect 12707 -1711 12741 -1303
rect 12825 -1711 12859 -1303
rect 12943 -1711 12977 -1303
rect 13061 -1711 13095 -1303
rect 13179 -1711 13213 -1303
rect 13297 -1711 13331 -1303
rect 13415 -1711 13449 -1303
rect 13533 -1711 13567 -1303
rect 13651 -1711 13685 -1303
rect 13769 -1711 13803 -1303
rect 13887 -1711 13921 -1303
rect 14005 -1711 14039 -1303
rect 14123 -1711 14157 -1303
rect 14241 -1711 14275 -1303
rect 14359 -1711 14393 -1303
rect 14477 -1711 14511 -1303
rect 14595 -1711 14629 -1303
rect 14713 -1711 14747 -1303
rect 14831 -1711 14865 -1303
rect 14949 -1711 14983 -1303
rect 20816 -1334 20850 -1043
rect 21012 -1334 21046 -1043
rect 21208 -1334 21242 -1043
rect 21462 -960 21496 -697
rect 21658 -960 21692 -697
rect 21854 -960 21888 -697
rect 22050 -960 22084 -697
rect 22246 -960 22280 -697
rect 21462 -994 22280 -960
rect 21462 -1251 21496 -994
rect 21658 -1251 21692 -994
rect 21854 -1251 21888 -994
rect 22050 -1251 22084 -994
rect 22246 -1251 22280 -994
rect 20807 -1402 21302 -1334
rect 21175 -1408 21302 -1402
rect 21739 -1408 22274 -1396
rect 22344 -1408 22396 189
rect 21175 -1460 22396 -1408
rect 25573 -1155 25868 876
rect 27816 937 27850 1145
rect 27974 937 28008 1145
rect 30321 1179 31628 1286
rect 29122 858 29156 1141
rect 29280 858 29314 1141
rect 30321 994 31628 1101
rect 27816 486 27850 693
rect 27974 486 28008 693
rect 27816 403 28008 486
rect 29101 777 29336 858
rect 29121 485 29155 777
rect 29279 485 29313 777
rect 30330 436 30364 994
rect 30646 436 30680 994
rect 30962 436 30996 994
rect 31278 436 31312 994
rect 31594 436 31628 994
rect 32576 1457 32610 2030
rect 32734 1457 32768 2030
rect 33122 1846 33156 2142
rect 33438 1846 33472 2142
rect 33884 1851 33918 2142
rect 34214 2116 34360 2189
rect 34168 1851 34202 2059
rect 34326 1851 34360 2116
rect 35065 2114 35099 2564
rect 35381 2114 35415 2676
rect 35697 2114 35731 2676
rect 35855 2096 35889 2522
rect 36013 2096 36047 2676
rect 36329 2641 36363 2676
rect 36761 2644 38097 2758
rect 39186 2731 39220 3022
rect 39382 2731 39416 3022
rect 39578 2731 39612 3022
rect 40068 2731 40102 3022
rect 40264 2731 40298 3022
rect 40460 2731 40494 3022
rect 36761 2641 38938 2644
rect 36329 2633 38938 2641
rect 36329 2548 36820 2633
rect 36171 2096 36205 2522
rect 36329 2096 36363 2548
rect 35855 2062 36363 2096
rect 36786 2071 36820 2548
rect 35904 2009 36307 2062
rect 33122 1457 33156 1665
rect 33438 1457 33472 1665
rect 33884 1457 33918 1665
rect 34172 1456 34206 1664
rect 34330 1456 34364 1664
rect 35065 1308 35099 1866
rect 37102 2071 37136 2633
rect 37418 2071 37452 2633
rect 37576 2053 37610 2479
rect 37734 2053 37768 2633
rect 38050 2548 38938 2633
rect 37892 2053 37926 2479
rect 38050 2053 38084 2548
rect 38874 2407 38938 2548
rect 38780 2149 38972 2407
rect 39186 2400 39220 2559
rect 39382 2400 39416 2559
rect 39578 2400 39612 2559
rect 40068 2400 40102 2559
rect 40264 2400 40298 2559
rect 41811 2731 41845 3022
rect 42007 2731 42041 3022
rect 42203 2731 42237 3022
rect 40460 2400 40494 2559
rect 42768 2731 42802 3022
rect 42964 2731 42998 3022
rect 43160 2731 43194 3022
rect 39177 2332 40593 2400
rect 41811 2400 41845 2559
rect 42007 2400 42041 2559
rect 42203 2400 42237 2559
rect 42768 2400 42802 2559
rect 42964 2400 42998 2559
rect 44511 2731 44545 3022
rect 44707 2731 44741 3022
rect 44903 2731 44937 3022
rect 43160 2400 43194 2559
rect 41802 2332 43293 2400
rect 44511 2400 44545 2559
rect 44707 2400 44741 2559
rect 44903 2400 44937 2559
rect 44502 2332 45036 2400
rect 37576 2019 38084 2053
rect 35381 1308 35415 1866
rect 35697 1308 35731 1866
rect 36013 1308 36047 1866
rect 37625 1966 38028 2019
rect 36329 1363 36363 1866
rect 36786 1363 36820 1823
rect 39440 2107 39572 2126
rect 42073 2107 42210 2126
rect 44670 2107 44807 2120
rect 39439 2068 44824 2107
rect 39440 2066 39572 2068
rect 41198 2020 41309 2068
rect 42073 2066 42210 2068
rect 41484 2020 42004 2022
rect 42076 2020 42187 2066
rect 36329 1308 36820 1363
rect 35056 1299 36820 1308
rect 32671 930 32705 1138
rect 32829 930 32863 1138
rect 35056 1201 36363 1299
rect 36786 1265 36820 1299
rect 37102 1265 37136 1823
rect 37418 1265 37452 1823
rect 37734 1265 37768 1823
rect 38050 1326 38084 1823
rect 40973 1954 42344 2020
rect 40973 1952 41507 1954
rect 41810 1952 42344 1954
rect 43874 2020 43985 2068
rect 44670 2060 44807 2068
rect 44685 2020 44796 2060
rect 41072 1793 41106 1952
rect 41268 1793 41302 1952
rect 41464 1793 41498 1952
rect 41909 1793 41943 1952
rect 42105 1793 42139 1952
rect 42301 1793 42335 1952
rect 43673 1952 45044 2020
rect 41072 1330 41106 1621
rect 41268 1330 41302 1621
rect 43772 1793 43806 1952
rect 41464 1330 41498 1621
rect 41909 1330 41943 1621
rect 42105 1330 42139 1621
rect 42301 1330 42335 1621
rect 43968 1793 44002 1952
rect 44164 1793 44198 1952
rect 44609 1793 44643 1952
rect 44805 1793 44839 1952
rect 45001 1793 45035 1952
rect 43772 1330 43806 1621
rect 43968 1330 44002 1621
rect 44164 1330 44198 1621
rect 44609 1330 44643 1621
rect 44805 1330 44839 1621
rect 45001 1330 45035 1621
rect 45195 1472 45284 3025
rect 45804 2255 45950 2441
rect 45853 2110 45897 2255
rect 45570 2042 46104 2110
rect 45579 1883 45613 2042
rect 45775 1883 45809 2042
rect 45971 1883 46005 2042
rect 45579 1472 45613 1711
rect 45195 1420 45613 1472
rect 45775 1420 45809 1711
rect 45971 1420 46005 1711
rect 45195 1415 46065 1420
rect 45195 1330 45284 1415
rect 45570 1352 46065 1415
rect 38049 1325 40098 1326
rect 41011 1325 42813 1330
rect 43711 1325 45284 1330
rect 38049 1265 45284 1325
rect 33977 851 34011 1134
rect 34135 851 34169 1134
rect 35065 1124 35099 1201
rect 35381 1124 35415 1201
rect 35697 1124 35731 1201
rect 36013 1124 36047 1201
rect 36329 1124 36363 1201
rect 35056 1017 36363 1124
rect 36777 1262 45284 1265
rect 36777 1242 40098 1262
rect 36777 1060 38084 1242
rect 32671 479 32705 686
rect 32829 479 32863 686
rect 32671 396 32863 479
rect 33956 770 34191 851
rect 33976 478 34010 770
rect 34134 478 34168 770
rect 35065 459 35099 1017
rect 35381 459 35415 1017
rect 35697 459 35731 1017
rect 36013 459 36047 1017
rect 36329 1011 36363 1017
rect 36786 1011 36820 1060
rect 36329 947 36820 1011
rect 36329 459 36363 947
rect 36786 502 36820 947
rect 37102 502 37136 1060
rect 37418 502 37452 1060
rect 37734 502 37768 1060
rect 38050 502 38084 1060
rect 47379 824 47674 3483
rect 51135 3263 51730 4290
rect 53312 3263 53907 4290
rect 55261 3263 55856 4290
rect 57618 3263 58213 4290
rect 50900 3197 58338 3263
rect 51101 3125 51160 3197
rect 51689 3125 51748 3197
rect 51960 3125 52019 3197
rect 52201 3125 52260 3197
rect 52433 3125 52492 3197
rect 53039 3125 53098 3197
rect 53268 3125 53327 3197
rect 53507 3125 53566 3197
rect 53742 3125 53801 3197
rect 53978 3125 54037 3197
rect 54209 3125 54268 3197
rect 54934 3125 54993 3197
rect 55168 3125 55227 3197
rect 55402 3125 55461 3197
rect 55639 3125 55698 3197
rect 55869 3125 55928 3197
rect 56109 3125 56168 3197
rect 56347 3125 56406 3197
rect 56583 3125 56642 3197
rect 56814 3125 56873 3197
rect 57291 3125 57350 3197
rect 50896 3077 58448 3125
rect 50896 2630 50930 3077
rect 51132 2630 51166 3077
rect 51368 2630 51402 3077
rect 51498 2630 51532 3077
rect 51734 2630 51768 3077
rect 51970 2630 52004 3077
rect 52206 2630 52240 3077
rect 52442 2630 52476 3077
rect 52572 2630 52606 3077
rect 52808 2630 52842 3077
rect 53044 2630 53078 3077
rect 53280 2630 53314 3077
rect 53516 2630 53550 3077
rect 53752 2630 53786 3077
rect 53988 2630 54022 3077
rect 54224 2630 54258 3077
rect 54460 2630 54494 3077
rect 54590 2630 54624 3038
rect 54708 2630 54742 3077
rect 54826 2630 54860 3038
rect 54944 2630 54978 3077
rect 55062 2630 55096 3038
rect 55180 2630 55214 3077
rect 55298 2630 55332 3038
rect 55416 2630 55450 3077
rect 55534 2630 55568 3038
rect 55652 2630 55686 3077
rect 55770 2630 55804 3038
rect 55888 2630 55922 3077
rect 56006 2630 56040 3038
rect 56124 2630 56158 3077
rect 56242 2630 56276 3038
rect 56360 2630 56394 3077
rect 56478 2630 56512 3038
rect 56596 2630 56630 3077
rect 56714 2630 56748 3038
rect 56832 2630 56866 3077
rect 56950 2630 56984 3038
rect 57068 2630 57102 3077
rect 57186 2630 57220 3038
rect 57304 2630 57338 3077
rect 57422 2630 57456 3038
rect 57540 2630 57574 3077
rect 57658 2630 57692 3038
rect 57776 2630 57810 3077
rect 57894 2630 57928 3038
rect 58012 2630 58046 3077
rect 58130 2630 58164 3038
rect 58248 2630 58282 3077
rect 58366 2484 58400 3038
rect 58711 2484 58930 2597
rect 58366 2450 58930 2484
rect 58711 2334 58930 2450
rect 54846 2294 58328 2322
rect 54698 2230 58328 2294
rect 51188 1737 51222 2230
rect 51424 1737 51458 2230
rect 51660 1737 51694 2230
rect 51896 1737 51930 2230
rect 52132 1737 52166 2230
rect 52368 1737 52402 2230
rect 52604 1737 52638 2230
rect 52840 1737 52874 2230
rect 52958 1822 52992 2230
rect 53076 1737 53110 2230
rect 53194 1822 53228 2230
rect 53312 1737 53346 2230
rect 53430 1822 53464 2230
rect 53548 1737 53582 2230
rect 53666 1822 53700 2230
rect 53784 1737 53818 2230
rect 53902 1822 53936 2230
rect 54020 1737 54054 2230
rect 54138 1822 54172 2230
rect 54256 1737 54290 2230
rect 54374 1822 54408 2230
rect 54492 1737 54526 2230
rect 54610 1822 54644 2230
rect 54728 1737 54762 2230
rect 54846 1822 54880 2230
rect 54964 1822 54998 2230
rect 55082 1822 55116 2230
rect 55200 1822 55234 2230
rect 55318 1822 55352 2230
rect 55436 1822 55470 2230
rect 55554 1822 55588 2230
rect 55672 1822 55706 2230
rect 55790 1822 55824 2230
rect 55908 1822 55942 2230
rect 56026 1822 56060 2230
rect 56144 1822 56178 2230
rect 56262 1822 56296 2230
rect 56380 1822 56414 2230
rect 56498 1822 56532 2230
rect 56616 1822 56650 2230
rect 56734 1822 56768 2230
rect 56852 1822 56886 2230
rect 56970 1822 57004 2230
rect 57088 1822 57122 2230
rect 57206 1822 57240 2230
rect 57324 1822 57358 2230
rect 57442 1822 57476 2230
rect 57560 1822 57594 2230
rect 57678 1822 57712 2230
rect 57796 1822 57830 2230
rect 57914 1822 57948 2230
rect 58032 1822 58066 2230
rect 58150 1822 58184 2230
rect 58268 1822 58302 2230
rect 51146 1617 58333 1737
rect 51870 824 52157 1617
rect 60670 1398 98798 4290
rect 60670 1310 61121 1398
rect 47379 537 52157 824
rect 53362 859 64533 1310
rect 27537 202 27729 274
rect 26988 -69 27304 -38
rect 26885 -149 27304 -69
rect 26988 -166 27304 -149
rect 27537 -191 27571 202
rect 27695 -27 27729 202
rect 27767 -69 27920 -59
rect 27605 -133 27920 -69
rect 27605 -149 27767 -133
rect 27967 -182 28001 183
rect 28283 -182 28317 183
rect 28599 -182 28633 183
rect 28915 -182 28949 183
rect 29231 -182 29265 183
rect 29506 -41 29540 183
rect 29664 -41 29698 183
rect 29506 -132 29698 -41
rect 29589 -182 29647 -132
rect 30330 -182 30364 188
rect 27781 -191 30364 -182
rect 27537 -225 30364 -191
rect 27537 -1155 27726 -225
rect 27781 -240 30364 -225
rect 29583 -291 30364 -240
rect 30330 -374 30364 -291
rect 30646 -374 30680 188
rect 31169 240 31572 293
rect 31120 206 31628 240
rect 30962 -374 30996 188
rect 31120 -220 31154 206
rect 31278 -374 31312 206
rect 31436 -220 31470 206
rect 31594 -217 31628 206
rect 32392 195 32584 267
rect 32392 -198 32426 195
rect 32550 -34 32584 195
rect 32622 -72 32775 -66
rect 32461 -140 32775 -72
rect 32461 -152 32623 -140
rect 32822 -189 32856 176
rect 33138 -189 33172 176
rect 33454 -189 33488 176
rect 33770 -189 33804 176
rect 34086 -189 34120 176
rect 34361 -48 34395 176
rect 34519 -48 34553 176
rect 34361 -139 34553 -48
rect 34444 -189 34502 -139
rect 32636 -198 34502 -189
rect 32392 -217 34502 -198
rect 31594 -232 34502 -217
rect 31594 -307 32499 -232
rect 32636 -247 34502 -232
rect 34420 -260 34502 -247
rect 35065 -260 35099 211
rect 34420 -294 35099 -260
rect 31594 -374 31628 -307
rect 35065 -351 35099 -294
rect 35381 -351 35415 211
rect 35904 263 36307 316
rect 35855 229 36363 263
rect 35697 -351 35731 211
rect 35855 -197 35889 229
rect 36013 -351 36047 229
rect 36171 -197 36205 229
rect 36329 -210 36363 229
rect 36786 -210 36820 254
rect 36329 -265 36820 -210
rect 36329 -351 36363 -265
rect 36786 -308 36820 -265
rect 37102 -308 37136 254
rect 37625 306 38028 359
rect 37576 272 38084 306
rect 37418 -308 37452 254
rect 37576 -154 37610 272
rect 37734 -308 37768 272
rect 37892 -154 37926 272
rect 38050 -308 38084 272
rect 30305 -499 31641 -374
rect 35040 -476 36376 -351
rect 36761 -433 38097 -308
rect 47379 -1155 47674 537
rect 53362 352 54000 859
rect 54759 352 55397 859
rect 56173 352 56811 859
rect 57259 352 57897 859
rect 50697 286 58135 352
rect 50898 214 50957 286
rect 51486 214 51545 286
rect 51757 214 51816 286
rect 51998 214 52057 286
rect 52230 214 52289 286
rect 52836 214 52895 286
rect 53065 214 53124 286
rect 53304 214 53363 286
rect 53539 214 53598 286
rect 53775 214 53834 286
rect 54006 214 54065 286
rect 54731 214 54790 286
rect 54965 214 55024 286
rect 55199 214 55258 286
rect 55436 214 55495 286
rect 55666 214 55725 286
rect 55906 214 55965 286
rect 56144 214 56203 286
rect 56380 214 56439 286
rect 56611 214 56670 286
rect 57088 214 57147 286
rect 50693 166 58245 214
rect 50693 -281 50727 166
rect 50929 -281 50963 166
rect 51165 -281 51199 166
rect 51295 -281 51329 166
rect 51531 -281 51565 166
rect 51767 -281 51801 166
rect 52003 -281 52037 166
rect 52239 -281 52273 166
rect 52369 -281 52403 166
rect 52605 -281 52639 166
rect 52841 -281 52875 166
rect 53077 -281 53111 166
rect 53313 -281 53347 166
rect 53549 -281 53583 166
rect 53785 -281 53819 166
rect 54021 -281 54055 166
rect 54257 -281 54291 166
rect 54387 -281 54421 127
rect 54505 -281 54539 166
rect 54623 -281 54657 127
rect 54741 -281 54775 166
rect 54859 -281 54893 127
rect 54977 -281 55011 166
rect 55095 -281 55129 127
rect 55213 -281 55247 166
rect 55331 -281 55365 127
rect 55449 -281 55483 166
rect 55567 -281 55601 127
rect 55685 -281 55719 166
rect 55803 -281 55837 127
rect 55921 -281 55955 166
rect 56039 -281 56073 127
rect 56157 -281 56191 166
rect 56275 -281 56309 127
rect 56393 -281 56427 166
rect 56511 -281 56545 127
rect 56629 -281 56663 166
rect 56747 -281 56781 127
rect 56865 -281 56899 166
rect 56983 -281 57017 127
rect 57101 -281 57135 166
rect 57219 -281 57253 127
rect 57337 -281 57371 166
rect 57455 -281 57489 127
rect 57573 -281 57607 166
rect 57691 -281 57725 127
rect 57809 -281 57843 166
rect 57927 -281 57961 127
rect 58045 -281 58079 166
rect 58163 -427 58197 127
rect 60613 -427 61078 -338
rect 58163 -461 61078 -427
rect 54643 -617 58125 -589
rect 54495 -681 58125 -617
rect 58324 -618 61078 -461
rect 60613 -669 61078 -618
rect 25573 -1450 47674 -1155
rect 50985 -1174 51019 -681
rect 51221 -1174 51255 -681
rect 51457 -1174 51491 -681
rect 51693 -1174 51727 -681
rect 51929 -1174 51963 -681
rect 52165 -1174 52199 -681
rect 52401 -1174 52435 -681
rect 52637 -1174 52671 -681
rect 52755 -1089 52789 -681
rect 52873 -1174 52907 -681
rect 52991 -1089 53025 -681
rect 53109 -1174 53143 -681
rect 53227 -1089 53261 -681
rect 53345 -1174 53379 -681
rect 53463 -1089 53497 -681
rect 53581 -1174 53615 -681
rect 53699 -1089 53733 -681
rect 53817 -1174 53851 -681
rect 53935 -1089 53969 -681
rect 54053 -1174 54087 -681
rect 54171 -1089 54205 -681
rect 54289 -1174 54323 -681
rect 54407 -1089 54441 -681
rect 54525 -1174 54559 -681
rect 54643 -1089 54677 -681
rect 54761 -1089 54795 -681
rect 54879 -1089 54913 -681
rect 54997 -1089 55031 -681
rect 55115 -1089 55149 -681
rect 55233 -1089 55267 -681
rect 55351 -1089 55385 -681
rect 55469 -1089 55503 -681
rect 55587 -1089 55621 -681
rect 55705 -1089 55739 -681
rect 55823 -1089 55857 -681
rect 55941 -1089 55975 -681
rect 56059 -1089 56093 -681
rect 56177 -1089 56211 -681
rect 56295 -1089 56329 -681
rect 56413 -1089 56447 -681
rect 56531 -1089 56565 -681
rect 56649 -1089 56683 -681
rect 56767 -1089 56801 -681
rect 56885 -1089 56919 -681
rect 57003 -1089 57037 -681
rect 57121 -1089 57155 -681
rect 57239 -1089 57273 -681
rect 57357 -1089 57391 -681
rect 57475 -1089 57509 -681
rect 57593 -1089 57627 -681
rect 57711 -1089 57745 -681
rect 57829 -1089 57863 -681
rect 57947 -1089 57981 -681
rect 58065 -1089 58099 -681
rect 50943 -1294 58130 -1174
rect 5739 -1965 6960 -1913
rect 7827 -1916 15014 -1796
rect 8336 -1966 8557 -1916
rect 9274 -1966 9547 -1916
rect 10255 -1966 10528 -1916
rect 11457 -1966 11730 -1916
rect 12412 -1966 12685 -1916
rect 13206 -1966 13479 -1916
rect 13931 -1966 14204 -1916
rect 26281 -1966 26638 -1450
rect 4310 -2204 4465 -2171
rect -26307 -2300 4465 -2204
rect 4310 -2309 4465 -2300
rect 8168 -2323 26638 -1966
rect 46864 -1737 47369 -1450
rect 52463 -1737 52968 -1294
rect 55332 -1517 55783 -1516
rect 56669 -1517 57120 -1516
rect 57856 -1517 58307 -1516
rect 64082 -1517 64533 859
rect 46864 -2242 52968 -1737
rect 53892 -1968 64533 -1517
rect -1585 -2393 -1283 -2369
rect -26253 -2533 -1283 -2393
rect 46864 -2515 47369 -2242
rect -1585 -2584 -1283 -2533
rect 3196 -2628 3624 -2539
rect -26211 -2873 3624 -2628
rect 53892 -2695 54343 -1968
rect 55332 -2695 55783 -1968
rect 56669 -2695 57120 -1968
rect 57856 -2695 58307 -1968
rect 64082 -2625 64533 -1968
rect 63602 -2677 64823 -2625
rect 62867 -2683 63256 -2682
rect 63602 -2683 63729 -2677
rect 50697 -2731 58307 -2695
rect 50697 -2761 58135 -2731
rect 62384 -2751 63729 -2683
rect 64166 -2689 64701 -2677
rect 50898 -2833 50957 -2761
rect 51486 -2833 51545 -2761
rect 51757 -2833 51816 -2761
rect 51998 -2833 52057 -2761
rect 52230 -2833 52289 -2761
rect 52836 -2833 52895 -2761
rect 53065 -2833 53124 -2761
rect 53304 -2833 53363 -2761
rect 53539 -2833 53598 -2761
rect 53775 -2833 53834 -2761
rect 54006 -2833 54065 -2761
rect 54731 -2833 54790 -2761
rect 54965 -2833 55024 -2761
rect 55199 -2833 55258 -2761
rect 55436 -2833 55495 -2761
rect 55666 -2833 55725 -2761
rect 55906 -2833 55965 -2761
rect 56144 -2833 56203 -2761
rect 56380 -2833 56439 -2761
rect 56611 -2833 56670 -2761
rect 57088 -2833 57147 -2761
rect 3196 -2900 3624 -2873
rect 15440 -2934 15853 -2842
rect -26114 -3188 15853 -2934
rect 15440 -3211 15853 -3188
rect 50693 -2881 58245 -2833
rect 16088 -3296 16483 -3292
rect -26140 -3586 16483 -3296
rect 50693 -3328 50727 -2881
rect 50929 -3328 50963 -2881
rect 16088 -3623 16483 -3586
rect 51165 -3328 51199 -2881
rect 51295 -3328 51329 -2881
rect 51531 -3328 51565 -2881
rect 51767 -3328 51801 -2881
rect 52003 -3328 52037 -2881
rect 52239 -3328 52273 -2881
rect 52369 -3328 52403 -2881
rect 52605 -3328 52639 -2881
rect 52841 -3328 52875 -2881
rect 53077 -3328 53111 -2881
rect 53313 -3328 53347 -2881
rect 53549 -3328 53583 -2881
rect 53785 -3328 53819 -2881
rect 54021 -3328 54055 -2881
rect 54257 -3328 54291 -2881
rect 54505 -3328 54539 -2881
rect 54741 -3328 54775 -2881
rect 54977 -3328 55011 -2881
rect 55213 -3328 55247 -2881
rect 55449 -3328 55483 -2881
rect 55685 -3328 55719 -2881
rect 55921 -3328 55955 -2881
rect 56157 -3328 56191 -2881
rect 56393 -3328 56427 -2881
rect 56629 -3328 56663 -2881
rect 56865 -3328 56899 -2881
rect 57101 -3328 57135 -2881
rect 57337 -3328 57371 -2881
rect 57573 -3328 57607 -2881
rect 57809 -3328 57843 -2881
rect 58045 -3328 58079 -2881
rect 62393 -3042 62427 -2751
rect 62589 -3042 62623 -2751
rect 62785 -3042 62819 -2751
rect 63243 -3042 63277 -2751
rect 63439 -3042 63473 -2751
rect 63635 -3042 63669 -2751
rect 62150 -3180 62449 -3106
rect 54643 -3664 58125 -3636
rect 54495 -3728 58125 -3664
rect 50985 -4221 51019 -3728
rect 51221 -4221 51255 -3728
rect 51457 -4221 51491 -3728
rect 51693 -4221 51727 -3728
rect 51929 -4221 51963 -3728
rect 52165 -4221 52199 -3728
rect 52401 -4221 52435 -3728
rect 52637 -4221 52671 -3728
rect 52873 -4221 52907 -3728
rect 53109 -4221 53143 -3728
rect 53345 -4221 53379 -3728
rect 53581 -4221 53615 -3728
rect 53817 -4221 53851 -3728
rect 54053 -4221 54087 -3728
rect 54289 -4221 54323 -3728
rect 54525 -4221 54559 -3728
rect 54643 -4136 54677 -3728
rect 54761 -4136 54795 -3728
rect 54879 -4136 54913 -3728
rect 54997 -4136 55031 -3728
rect 55115 -4136 55149 -3728
rect 55233 -4136 55267 -3728
rect 55351 -4136 55385 -3728
rect 55469 -4136 55503 -3728
rect 55587 -4136 55621 -3728
rect 55705 -4136 55739 -3728
rect 55823 -4136 55857 -3728
rect 55941 -4136 55975 -3728
rect 56059 -4136 56093 -3728
rect 56177 -4136 56211 -3728
rect 56295 -4136 56329 -3728
rect 56413 -4136 56447 -3728
rect 56531 -4136 56565 -3728
rect 56649 -4136 56683 -3728
rect 56767 -4136 56801 -3728
rect 56885 -4136 56919 -3728
rect 57003 -4136 57037 -3728
rect 57121 -4136 57155 -3728
rect 57239 -4136 57273 -3728
rect 57357 -4136 57391 -3728
rect 57475 -4136 57509 -3728
rect 57593 -4136 57627 -3728
rect 57711 -4136 57745 -3728
rect 57829 -4136 57863 -3728
rect 57947 -4136 57981 -3728
rect 58065 -4136 58099 -3728
rect 62278 -3785 62330 -3180
rect 62393 -3373 62427 -3214
rect 62589 -3373 62623 -3214
rect 62785 -3373 62819 -3214
rect 63243 -3373 63277 -3214
rect 63439 -3373 63473 -3214
rect 63635 -3373 63669 -3214
rect 62384 -3441 63768 -3373
rect 63234 -3578 63768 -3441
rect 63243 -3737 63277 -3578
rect 63131 -3785 63299 -3771
rect 62278 -3837 63299 -3785
rect 62432 -4139 62779 -3837
rect 63131 -3845 63299 -3837
rect 63439 -3737 63473 -3578
rect 63635 -3737 63669 -3578
rect 63243 -4200 63277 -3909
rect 63439 -4200 63473 -3909
rect 63635 -4200 63669 -3909
rect 63889 -3826 63923 -3563
rect 64085 -3826 64119 -3563
rect 64281 -3826 64315 -3563
rect 64477 -3826 64511 -3563
rect 64673 -3826 64707 -3563
rect 63889 -3860 64707 -3826
rect 63889 -4117 63923 -3860
rect 64085 -4117 64119 -3860
rect 64281 -4117 64315 -3860
rect 64477 -4117 64511 -3860
rect 64673 -4117 64707 -3860
rect 17293 -4336 17906 -4235
rect 16975 -4354 17906 -4336
rect 50943 -4341 58130 -4221
rect 63234 -4268 63729 -4200
rect 63602 -4274 63729 -4268
rect 64166 -4274 64701 -4262
rect 64771 -4274 64823 -2677
rect 63602 -4326 64823 -4274
rect -26205 -4766 17906 -4354
rect 17293 -4848 17906 -4766
rect 46778 -4698 47398 -4670
rect 52571 -4698 53148 -4341
rect 95829 -4698 98798 1398
rect 17978 -5013 18468 -4849
rect -26311 -5399 18468 -5013
rect 46778 -5275 92959 -4698
rect 46778 -5304 47412 -5275
rect 17978 -5437 18468 -5399
rect 18534 -5664 18990 -5587
rect -26321 -6062 18990 -5664
rect -26321 -6098 18704 -6062
rect 18949 -6346 19611 -6293
rect -26653 -6787 19611 -6346
rect 18949 -6850 19611 -6787
rect 19665 -7100 20295 -7025
rect -26746 -7593 20295 -7100
rect 19665 -7634 20295 -7593
rect 70077 -7667 92959 -5275
rect 95743 -7667 98798 -4698
rect 70077 -7803 73046 -7667
rect 81551 -7803 84520 -7667
rect -31467 -9060 -30570 -8797
rect 58913 -9060 59860 -8831
rect -34283 -9713 59860 -9060
rect -31467 -10014 -30570 -9713
rect 58913 -9909 59860 -9713
rect -29173 -9983 -28472 -9982
rect 60423 -9983 61454 -9617
rect -29347 -10522 61454 -9983
rect -29564 -10681 61454 -10522
rect -29564 -11751 -28286 -10681
rect 60423 -10731 61454 -10681
rect -29173 -12595 -28472 -11751
rect -6611 -11274 -5937 -11153
rect 61366 -11274 62272 -11116
rect -6611 -11839 62272 -11274
rect -6611 -11894 -5937 -11839
rect 61366 -11971 62272 -11839
rect 62246 -12546 63072 -12441
rect -34369 -13296 -28472 -12595
rect -26996 -13121 63072 -12546
rect 95829 -12668 98798 -7667
rect -26996 -13991 -26421 -13121
rect 62246 -13180 63072 -13121
rect -34505 -14566 -26421 -13991
rect -11293 -15732 -11259 -15324
rect -11057 -15732 -11023 -15324
rect -10821 -15732 -10787 -15324
rect -10585 -15732 -10551 -15324
rect -10349 -15732 -10315 -15324
rect -10113 -15732 -10079 -15324
rect -9877 -15732 -9843 -15324
rect -9641 -15732 -9607 -15324
rect -34293 -15952 -15114 -15892
rect -34293 -15986 -15015 -15952
rect -34293 -16022 -15114 -15986
rect -15049 -16540 -15015 -15986
rect -14931 -16579 -14897 -16132
rect -14813 -16540 -14779 -16132
rect -14695 -16579 -14661 -16132
rect -14577 -16540 -14543 -16132
rect -14459 -16579 -14425 -16132
rect -14341 -16540 -14307 -16132
rect -14223 -16579 -14189 -16132
rect -14105 -16540 -14071 -16132
rect -13987 -16579 -13953 -16132
rect -13869 -16540 -13835 -16132
rect -13751 -16579 -13717 -16132
rect -13633 -16540 -13599 -16132
rect -13515 -16579 -13481 -16132
rect -13397 -16540 -13363 -16132
rect -13279 -16579 -13245 -16132
rect -13161 -16540 -13127 -16132
rect -13043 -16579 -13009 -16132
rect -12925 -16540 -12891 -16132
rect -12807 -16579 -12773 -16132
rect -12689 -16540 -12655 -16132
rect -12571 -16579 -12537 -16132
rect -12453 -16540 -12419 -16132
rect -12335 -16579 -12301 -16132
rect -12217 -16540 -12183 -16132
rect -12099 -16579 -12065 -16132
rect -11981 -16540 -11947 -16132
rect -11863 -16579 -11829 -16132
rect -11745 -16540 -11711 -16132
rect -11627 -16579 -11593 -16132
rect -11509 -16540 -11475 -16132
rect -11391 -16579 -11357 -16132
rect -11273 -16540 -11239 -16132
rect -11143 -16579 -11109 -16132
rect -10907 -16579 -10873 -16132
rect -10671 -16579 -10637 -16132
rect -10435 -16579 -10401 -16132
rect -10199 -16579 -10165 -16132
rect -9963 -16579 -9929 -16132
rect -9727 -16579 -9693 -16132
rect -9491 -16579 -9457 -16132
rect -9255 -16579 -9221 -16132
rect -9125 -16579 -9091 -16132
rect 81378 -15816 98798 -12668
rect 81378 -16058 84526 -15816
rect -8889 -16579 -8855 -16132
rect -8653 -16579 -8619 -16132
rect -8417 -16579 -8383 -16132
rect -8181 -16579 -8147 -16132
rect -8051 -16579 -8017 -16132
rect -7815 -16579 -7781 -16132
rect -7579 -16579 -7545 -16132
rect 25225 -16279 86373 -16058
rect -15097 -16627 -7545 -16579
rect -13999 -16699 -13940 -16627
rect -13522 -16699 -13463 -16627
rect -13291 -16699 -13232 -16627
rect -13055 -16699 -12996 -16627
rect -12817 -16699 -12758 -16627
rect -12577 -16699 -12518 -16627
rect -12347 -16699 -12288 -16627
rect -12110 -16699 -12051 -16627
rect -11876 -16699 -11817 -16627
rect -11642 -16699 -11583 -16627
rect -10917 -16699 -10858 -16627
rect -10686 -16699 -10627 -16627
rect -10450 -16699 -10391 -16627
rect -10215 -16699 -10156 -16627
rect -9976 -16699 -9917 -16627
rect -9747 -16699 -9688 -16627
rect -9141 -16699 -9082 -16627
rect -8909 -16699 -8850 -16627
rect -8668 -16699 -8609 -16627
rect -8397 -16699 -8338 -16627
rect -7809 -16699 -7750 -16627
rect -14987 -16765 -7549 -16699
rect -14106 -18242 -13756 -16765
rect -11883 -18242 -11533 -16765
rect -9810 -18206 -9410 -16765
rect 6197 -17041 86373 -16279
rect 6197 -18195 6959 -17041
rect 25225 -17161 86373 -17041
rect -8032 -18206 7428 -18195
rect -10363 -18242 7428 -18206
rect -15388 -18295 7428 -18242
rect -15388 -18305 -10163 -18295
rect -15388 -18310 -13815 -18305
rect -12917 -18310 -11115 -18305
rect -15388 -18869 -15299 -18310
rect -15139 -18601 -15105 -18310
rect -14943 -18601 -14909 -18310
rect -14747 -18601 -14713 -18310
rect -14302 -18601 -14268 -18310
rect -24351 -19082 -15299 -18869
rect -24351 -19092 -22116 -19082
rect -24351 -20833 -24079 -19092
rect -23884 -19600 -23823 -19397
rect -23693 -19518 -23632 -19318
rect -23584 -19435 -23523 -19232
rect -22738 -19388 -22704 -19092
rect -22542 -19388 -22508 -19092
rect -22346 -19388 -22312 -19092
rect -22150 -19388 -22116 -19092
rect -21613 -19096 -21368 -19082
rect -21608 -19388 -21574 -19096
rect -22815 -19435 -22680 -19427
rect -23584 -19470 -22680 -19435
rect -22834 -19472 -22680 -19470
rect -22815 -19481 -22680 -19472
rect -22479 -19518 -22344 -19509
rect -23693 -19556 -22344 -19518
rect -22479 -19563 -22344 -19556
rect -22291 -19600 -22156 -19587
rect -23884 -19634 -22156 -19600
rect -23884 -19635 -23823 -19634
rect -22291 -19641 -22156 -19634
rect -21412 -19388 -21378 -19096
rect -20791 -19144 -19464 -19082
rect -20791 -19199 -19460 -19144
rect -20739 -19610 -20705 -19199
rect -21054 -19661 -20917 -19644
rect -20543 -19610 -20509 -19199
rect -20347 -19243 -19460 -19199
rect -20347 -19610 -20313 -19243
rect -20130 -19409 -20096 -19243
rect -19934 -19409 -19900 -19243
rect -19738 -19409 -19704 -19243
rect -19542 -19409 -19508 -19243
rect -20824 -19659 -20689 -19653
rect -20844 -19661 -20689 -19659
rect -21054 -19697 -20689 -19661
rect -21054 -19702 -20917 -19697
rect -20844 -19699 -20689 -19697
rect -20824 -19707 -20689 -19699
rect -20959 -19755 -20822 -19751
rect -20997 -19757 -20770 -19755
rect -20359 -19757 -20285 -19731
rect -20997 -19795 -20285 -19757
rect -20959 -19809 -20822 -19795
rect -20771 -19796 -20285 -19795
rect -20771 -19797 -20700 -19796
rect -20359 -19802 -20285 -19796
rect -23485 -20474 -23425 -20398
rect -23485 -20514 -23417 -20474
rect -23372 -20508 -23311 -20330
rect -21084 -20508 -21031 -20412
rect -23485 -20591 -23425 -20514
rect -23372 -20544 -21031 -20508
rect -23372 -20546 -23311 -20544
rect -21068 -20591 -20936 -20582
rect -23485 -20631 -20936 -20591
rect -23485 -20635 -23425 -20631
rect -21068 -20635 -20936 -20631
rect -19103 -20681 -19069 -20264
rect -18907 -20681 -18873 -20264
rect -18711 -20631 -18677 -20264
rect -18494 -20631 -18460 -20465
rect -18298 -20631 -18264 -20465
rect -18102 -20631 -18068 -20465
rect -17906 -20631 -17872 -20465
rect -18711 -20681 -17824 -20631
rect -17656 -20643 -17622 -20053
rect -19113 -20730 -17824 -20681
rect -19113 -20745 -18671 -20730
rect -17661 -20769 -17616 -20643
rect -17460 -20646 -17426 -20053
rect -17466 -20769 -17421 -20646
rect -17037 -20645 -17003 -20053
rect -17044 -20769 -16999 -20645
rect -18674 -20786 -18485 -20779
rect -18711 -20793 -18485 -20786
rect -17667 -20793 -16898 -20769
rect -19113 -20833 -16898 -20793
rect -24351 -20835 -16898 -20833
rect -24351 -20946 -17002 -20835
rect -24351 -21032 -19538 -20946
rect -24351 -21065 -19548 -21032
rect -22691 -21102 -21402 -21065
rect -23113 -21570 -23053 -21371
rect -22681 -21519 -22647 -21102
rect -22485 -21519 -22451 -21102
rect -22289 -21152 -21402 -21102
rect -22289 -21519 -22255 -21152
rect -22072 -21318 -22038 -21152
rect -21876 -21318 -21842 -21152
rect -21680 -21318 -21646 -21152
rect -21484 -21318 -21450 -21152
rect -20908 -21324 -20874 -21065
rect -20712 -21324 -20678 -21065
rect -20516 -21324 -20482 -21065
rect -20320 -21324 -20286 -21065
rect -19778 -21324 -19744 -21065
rect -22766 -21568 -22631 -21562
rect -22786 -21570 -22631 -21568
rect -23113 -21606 -22631 -21570
rect -23113 -21608 -23053 -21606
rect -22786 -21608 -22631 -21606
rect -22766 -21616 -22631 -21608
rect -23239 -21666 -22712 -21664
rect -22301 -21666 -22227 -21640
rect -23239 -21704 -22227 -21666
rect -23239 -21809 -23199 -21704
rect -22713 -21705 -22227 -21704
rect -22713 -21706 -22642 -21705
rect -22301 -21711 -22227 -21705
rect -23256 -22046 -23196 -21809
rect -19582 -21324 -19548 -21065
rect -18943 -21136 -18771 -20946
rect -18115 -20963 -17497 -20946
rect -18115 -20992 -17672 -20963
rect -18114 -21006 -17672 -20992
rect -18114 -21055 -16825 -21006
rect -19125 -21235 -18407 -21136
rect -19077 -21501 -19043 -21235
rect -18881 -21501 -18847 -21235
rect -18685 -21501 -18651 -21235
rect -18489 -21501 -18455 -21235
rect -18104 -21472 -18070 -21055
rect -17908 -21472 -17874 -21055
rect -17712 -21105 -16825 -21055
rect -17712 -21472 -17678 -21105
rect -17495 -21271 -17461 -21105
rect -17299 -21271 -17265 -21105
rect -17103 -21271 -17069 -21105
rect -16907 -21271 -16873 -21105
rect -15388 -20005 -15299 -19082
rect -14106 -18601 -14072 -18310
rect -13910 -18601 -13876 -18310
rect -12439 -18601 -12405 -18310
rect -12243 -18601 -12209 -18310
rect -12047 -18601 -12013 -18310
rect -11602 -18601 -11568 -18310
rect -11406 -18601 -11372 -18310
rect -11210 -18601 -11176 -18310
rect -8781 -18419 -8736 -18295
rect -8777 -19011 -8743 -18419
rect -8359 -18418 -8314 -18295
rect -8354 -19011 -8320 -18418
rect -8164 -18421 -8119 -18295
rect -8034 -18388 7428 -18295
rect -8158 -19011 -8124 -18421
rect -15041 -20002 -15007 -19711
rect -14845 -20002 -14811 -19711
rect -14649 -20002 -14615 -19711
rect -13298 -20002 -13264 -19711
rect -13102 -20002 -13068 -19711
rect -12906 -20002 -12872 -19711
rect -12341 -20002 -12307 -19711
rect -12145 -20002 -12111 -19711
rect -11949 -20002 -11915 -19711
rect -10598 -20002 -10564 -19711
rect -10402 -20002 -10368 -19711
rect -10206 -20002 -10172 -19711
rect -9716 -20002 -9682 -19711
rect -9520 -20002 -9486 -19711
rect -9324 -20002 -9290 -19711
rect -15101 -20005 -14606 -20002
rect -13359 -20003 -11906 -20002
rect -15388 -20007 -14284 -20005
rect -13359 -20007 -11593 -20003
rect -10659 -20007 -9281 -20002
rect -15388 -20070 -9281 -20007
rect -15388 -20073 -14284 -20070
rect -12066 -20071 -11593 -20070
rect -14926 -21769 -14773 -20073
rect -14146 -21054 -14075 -21053
rect -13734 -21054 -13660 -21048
rect -14146 -21055 -13660 -21054
rect -14372 -21093 -13660 -21055
rect -14372 -21095 -14145 -21093
rect -13734 -21119 -13660 -21093
rect -14114 -21657 -14080 -21240
rect -13918 -21657 -13884 -21240
rect -13722 -21607 -13688 -21240
rect -13505 -21607 -13471 -21441
rect -13309 -21607 -13275 -21441
rect -13113 -21607 -13079 -21441
rect -12917 -21607 -12883 -21441
rect -13722 -21657 -12835 -21607
rect -12667 -21619 -12633 -21029
rect -14124 -21706 -12835 -21657
rect -14124 -21721 -13682 -21706
rect -12672 -21745 -12627 -21619
rect -12471 -21622 -12437 -21029
rect -12477 -21745 -12432 -21622
rect -12048 -21621 -12014 -21029
rect -12055 -21745 -12010 -21621
rect -13685 -21762 -13496 -21755
rect -13722 -21769 -13496 -21762
rect -12678 -21769 -11909 -21745
rect -14926 -21811 -11909 -21769
rect -14926 -21922 -12013 -21811
rect -14926 -23169 -14773 -21922
rect -13954 -22112 -13782 -21922
rect -13126 -21939 -12508 -21922
rect -13126 -21968 -12683 -21939
rect -13125 -21982 -12683 -21968
rect -13125 -22031 -11836 -21982
rect -14136 -22211 -13418 -22112
rect -14088 -22477 -14054 -22211
rect -13892 -22477 -13858 -22211
rect -13696 -22477 -13662 -22211
rect -13500 -22477 -13466 -22211
rect -13115 -22448 -13081 -22031
rect -12919 -22448 -12885 -22031
rect -12723 -22081 -11836 -22031
rect -12723 -22448 -12689 -22081
rect -12506 -22247 -12472 -22081
rect -12310 -22247 -12276 -22081
rect -12114 -22247 -12080 -22081
rect -11918 -22247 -11884 -22081
rect -6669 -18495 -5617 -18388
rect -6669 -18624 -6629 -18495
rect -6669 -18807 -6635 -18624
rect -6480 -18624 -6434 -18495
rect -6473 -18807 -6439 -18624
rect -6282 -18620 -6236 -18495
rect -6277 -18807 -6243 -18620
rect -6169 -18624 -6123 -18495
rect -6163 -18807 -6129 -18624
rect -5973 -18619 -5927 -18495
rect -5967 -18807 -5933 -18619
rect -5860 -18629 -5814 -18495
rect -5854 -18807 -5820 -18629
rect -5663 -18617 -5617 -18495
rect -5658 -18807 -5624 -18617
rect -5342 -19225 -5227 -18388
rect -3855 -18426 -3262 -18388
rect -5347 -19361 -5224 -19225
rect -4169 -18495 -3117 -18426
rect -4169 -18624 -4129 -18495
rect -4169 -18807 -4135 -18624
rect -3980 -18624 -3934 -18495
rect -3973 -18807 -3939 -18624
rect -3782 -18620 -3736 -18495
rect -3777 -18807 -3743 -18620
rect -3669 -18624 -3623 -18495
rect -3663 -18807 -3629 -18624
rect -3473 -18619 -3427 -18495
rect -4564 -19115 -4425 -19061
rect -3467 -18807 -3433 -18619
rect -3360 -18629 -3314 -18495
rect -3354 -18807 -3320 -18629
rect -3163 -18617 -3117 -18495
rect -3158 -18807 -3124 -18617
rect -3486 -19121 -3347 -19067
rect -2774 -19260 -2660 -18388
rect -1339 -18426 -746 -18388
rect -1669 -18495 -617 -18426
rect -1669 -18624 -1629 -18495
rect -1669 -18807 -1635 -18624
rect -1480 -18624 -1434 -18495
rect -1473 -18807 -1439 -18624
rect -1282 -18620 -1236 -18495
rect -1277 -18807 -1243 -18620
rect -1169 -18624 -1123 -18495
rect -1163 -18807 -1129 -18624
rect -973 -18619 -927 -18495
rect -2064 -19115 -1925 -19061
rect -2780 -19396 -2657 -19260
rect -967 -18807 -933 -18619
rect -860 -18629 -814 -18495
rect -854 -18807 -820 -18629
rect -663 -18617 -617 -18495
rect -658 -18807 -624 -18617
rect -986 -19121 -847 -19067
rect -292 -19260 -177 -18388
rect 1195 -18426 1788 -18388
rect 3608 -18426 4201 -18388
rect 831 -18495 1883 -18426
rect 831 -18624 871 -18495
rect 831 -18807 865 -18624
rect 1020 -18624 1066 -18495
rect 1027 -18807 1061 -18624
rect 1218 -18620 1264 -18495
rect 1223 -18807 1257 -18620
rect 1331 -18624 1377 -18495
rect 1337 -18807 1371 -18624
rect 1527 -18619 1573 -18495
rect 436 -19115 575 -19061
rect -297 -19396 -174 -19260
rect 1533 -18807 1567 -18619
rect 1640 -18629 1686 -18495
rect 1646 -18807 1680 -18629
rect 1837 -18617 1883 -18495
rect 1842 -18807 1876 -18617
rect 1514 -19121 1653 -19067
rect 3331 -18495 4383 -18426
rect 3331 -18624 3371 -18495
rect 3331 -18807 3365 -18624
rect 3520 -18624 3566 -18495
rect 3527 -18807 3561 -18624
rect 3718 -18620 3764 -18495
rect 3723 -18807 3757 -18620
rect 3831 -18624 3877 -18495
rect 3837 -18807 3871 -18624
rect 4027 -18619 4073 -18495
rect 2936 -19115 3075 -19061
rect 4033 -18807 4067 -18619
rect 4140 -18629 4186 -18495
rect 4146 -18807 4180 -18629
rect 4337 -18617 4383 -18495
rect 4342 -18807 4376 -18617
rect 4014 -19121 4153 -19067
rect 6331 -18495 7383 -18388
rect 6331 -18624 6371 -18495
rect 6331 -18807 6365 -18624
rect 6520 -18624 6566 -18495
rect 6527 -18807 6561 -18624
rect 6718 -18620 6764 -18495
rect 6723 -18807 6757 -18620
rect 6831 -18624 6877 -18495
rect 6837 -18807 6871 -18624
rect 7027 -18619 7073 -18495
rect 5936 -19115 6075 -19061
rect 7033 -18807 7067 -18619
rect 7140 -18629 7186 -18495
rect 7146 -18807 7180 -18629
rect 7337 -18617 7383 -18495
rect 7342 -18807 7376 -18617
rect 7014 -19121 7153 -19067
rect -7140 -19864 -6952 -19790
rect -298 -19814 -175 -19813
rect -7008 -20219 -6974 -19928
rect -6812 -20219 -6778 -19928
rect -6616 -20219 -6582 -19928
rect -5348 -20128 -5225 -19992
rect -2781 -19984 -2658 -19848
rect -298 -19876 8 -19814
rect -7017 -20287 -6522 -20219
rect -7001 -20677 -6913 -20287
rect -6818 -20677 -6730 -20287
rect -6636 -20677 -6548 -20287
rect -7514 -20680 -6410 -20677
rect -5343 -20680 -5228 -20128
rect -4192 -20680 -3719 -20679
rect -2777 -20680 -2662 -19984
rect -1522 -20680 -1399 -20658
rect -7514 -20743 -1399 -20680
rect -7514 -20745 -6410 -20743
rect -14282 -22524 -14152 -22507
rect -14108 -22524 -14035 -22511
rect -14282 -22565 -14035 -22524
rect -7514 -22440 -7425 -20745
rect -7227 -20748 -6732 -20745
rect -5485 -20747 -3719 -20743
rect -5485 -20748 -4032 -20747
rect -2785 -20748 -1399 -20743
rect -7167 -21039 -7133 -20748
rect -6971 -21039 -6937 -20748
rect -6775 -21039 -6741 -20748
rect -5424 -21039 -5390 -20748
rect -5228 -21039 -5194 -20748
rect -5032 -21039 -4998 -20748
rect -4467 -21039 -4433 -20748
rect -4271 -21039 -4237 -20748
rect -4075 -21039 -4041 -20748
rect -2724 -21039 -2690 -20748
rect -2528 -21039 -2494 -20748
rect -2332 -21039 -2298 -20748
rect -1842 -21039 -1808 -20748
rect -1646 -21039 -1612 -20748
rect -1522 -20794 -1399 -20748
rect -1450 -21039 -1416 -20794
rect -1228 -20684 -1105 -20657
rect -293 -20684 -178 -19876
rect 1750 -20684 1873 -20670
rect -1228 -20763 1873 -20684
rect -1228 -20764 -873 -20763
rect -1228 -20793 -1074 -20764
rect -1108 -21056 -1074 -20793
rect -912 -21056 -878 -20764
rect -370 -21056 -336 -20763
rect -174 -21056 -140 -20763
rect 22 -21056 56 -20763
rect 218 -21056 252 -20763
rect 577 -20803 1464 -20763
rect 625 -20969 659 -20803
rect 821 -20969 855 -20803
rect 1017 -20969 1051 -20803
rect 1213 -20969 1247 -20803
rect -7265 -22440 -7231 -22149
rect -7069 -22440 -7035 -22149
rect -6873 -22440 -6839 -22149
rect -6428 -22440 -6394 -22149
rect -6232 -22440 -6198 -22149
rect -6036 -22440 -6002 -22149
rect -4565 -22440 -4531 -22149
rect -4369 -22440 -4335 -22149
rect -4173 -22440 -4139 -22149
rect -3728 -22440 -3694 -22149
rect -3532 -22440 -3498 -22149
rect -3336 -22440 -3302 -22149
rect 1430 -21170 1464 -20803
rect 1626 -21170 1660 -20763
rect 1750 -20806 1873 -20763
rect 1822 -21170 1856 -20806
rect 2139 -20706 2262 -20669
rect 3367 -20691 3490 -20646
rect 3029 -20706 3490 -20691
rect 2139 -20755 3490 -20706
rect 2139 -20805 3069 -20755
rect 2230 -20971 2264 -20805
rect 2426 -20971 2460 -20805
rect 2622 -20971 2656 -20805
rect 2818 -20971 2852 -20805
rect 3035 -21172 3069 -20805
rect 3231 -21172 3265 -20755
rect 3367 -20782 3490 -20755
rect 3427 -21172 3461 -20782
rect 3768 -20677 3891 -20644
rect 3768 -20682 4664 -20677
rect 5124 -20682 5247 -20649
rect 3768 -20750 5247 -20682
rect 3768 -20755 4089 -20750
rect 4592 -20751 5247 -20750
rect 3768 -20780 3891 -20755
rect 3854 -21047 3888 -20780
rect 4050 -21047 4084 -20755
rect 4592 -21047 4626 -20751
rect 4788 -21047 4822 -20751
rect 4984 -21047 5018 -20751
rect 5124 -20785 5247 -20751
rect 5180 -21047 5214 -20785
rect 6340 -20677 6463 -20650
rect 6340 -20746 7393 -20677
rect 6340 -20786 6463 -20746
rect 6341 -20875 6381 -20786
rect 6341 -21058 6375 -20875
rect 6530 -20875 6576 -20746
rect 6537 -21058 6571 -20875
rect 6728 -20871 6774 -20746
rect 6733 -21058 6767 -20871
rect 6841 -20875 6887 -20746
rect 6847 -21058 6881 -20875
rect 7037 -20870 7083 -20746
rect 5946 -21366 6085 -21312
rect 7043 -21058 7077 -20870
rect 7150 -20880 7196 -20746
rect 7156 -21058 7190 -20880
rect 7347 -20868 7393 -20746
rect 7352 -21058 7386 -20868
rect 7024 -21372 7163 -21318
rect 25225 -18550 26328 -17161
rect 19573 -21012 24798 -20949
rect 20525 -21017 22327 -21012
rect 23225 -21017 24798 -21012
rect 26958 -21013 26992 -20747
rect 27154 -21013 27188 -20747
rect 27350 -21013 27384 -20747
rect 27546 -21013 27580 -20747
rect -7514 -22445 -5941 -22440
rect -5043 -22445 -3241 -22440
rect -7514 -22508 -2289 -22445
rect -14282 -22657 -14152 -22565
rect -14108 -22571 -14035 -22565
rect -7514 -23147 -7425 -22508
rect -11310 -23169 -7425 -23147
rect -15388 -23232 -7425 -23169
rect -15388 -23237 -13815 -23232
rect -12917 -23237 -11115 -23232
rect -15388 -23862 -15299 -23237
rect -15139 -23528 -15105 -23237
rect -14943 -23528 -14909 -23237
rect -14747 -23528 -14713 -23237
rect -14302 -23528 -14268 -23237
rect -14106 -23528 -14072 -23237
rect -13910 -23528 -13876 -23237
rect -22935 -24029 -15298 -23862
rect -22565 -24168 -21783 -24029
rect -21407 -24155 -20889 -24029
rect -22625 -24301 -21757 -24168
rect -21422 -24224 -20868 -24155
rect -20518 -24156 -19965 -24029
rect -20518 -24197 -19963 -24156
rect -22625 -24413 -22572 -24301
rect -23884 -25120 -23824 -24939
rect -22616 -25013 -22582 -24413
rect -22429 -24429 -22376 -24301
rect -21417 -24351 -21369 -24224
rect -22420 -25013 -22386 -24429
rect -21410 -24742 -21376 -24351
rect -21220 -24357 -21172 -24224
rect -20517 -24225 -19963 -24197
rect -21590 -24858 -21532 -24763
rect -21214 -24742 -21180 -24357
rect -20512 -24352 -20464 -24225
rect -21183 -24858 -21040 -24851
rect -21590 -24894 -21040 -24858
rect -21590 -24900 -21532 -24894
rect -21183 -24911 -21040 -24894
rect -20505 -24743 -20471 -24352
rect -20315 -24358 -20267 -24225
rect -20674 -24859 -20616 -24764
rect -20309 -24743 -20275 -24358
rect -20278 -24859 -20135 -24852
rect -20674 -24895 -20135 -24859
rect -20674 -24901 -20616 -24895
rect -20278 -24912 -20135 -24895
rect -21515 -24947 -21457 -24934
rect -21406 -24947 -21260 -24931
rect -21515 -24983 -21260 -24947
rect -21515 -25071 -21457 -24983
rect -21406 -24991 -21260 -24983
rect -20597 -24948 -20539 -24936
rect -20501 -24948 -20355 -24932
rect -20597 -24984 -20355 -24948
rect -23884 -25161 -21995 -25120
rect -23884 -25176 -23824 -25161
rect -22055 -25166 -21995 -25161
rect -23693 -25209 -23633 -25196
rect -22375 -25209 -22230 -25198
rect -23693 -25250 -22230 -25209
rect -22055 -25222 -21910 -25166
rect -23693 -25433 -23633 -25250
rect -22375 -25254 -22230 -25250
rect -23583 -25301 -23523 -25299
rect -22704 -25301 -22559 -25293
rect -23583 -25342 -22559 -25301
rect -23583 -25536 -23523 -25342
rect -22704 -25349 -22559 -25342
rect -20597 -25073 -20539 -24984
rect -20501 -24992 -20355 -24984
rect -19103 -25681 -19069 -25264
rect -18907 -25681 -18873 -25264
rect -18711 -25631 -18677 -25264
rect -18494 -25631 -18460 -25465
rect -18298 -25631 -18264 -25465
rect -18102 -25631 -18068 -25465
rect -17906 -25631 -17872 -25465
rect -18711 -25681 -17824 -25631
rect -17656 -25643 -17622 -25053
rect -19113 -25730 -17824 -25681
rect -19113 -25745 -18671 -25730
rect -17661 -25769 -17616 -25643
rect -17460 -25646 -17426 -25053
rect -17466 -25769 -17421 -25646
rect -17037 -25645 -17003 -25053
rect -15388 -24932 -15299 -24029
rect -12439 -23528 -12405 -23237
rect -12243 -23528 -12209 -23237
rect -12047 -23528 -12013 -23237
rect -11602 -23528 -11568 -23237
rect -11406 -23528 -11372 -23237
rect -11210 -23528 -11176 -23237
rect -8754 -23353 -8709 -23232
rect -8750 -23945 -8716 -23353
rect -8332 -23352 -8287 -23232
rect -8327 -23945 -8293 -23352
rect -8137 -23355 -8092 -23232
rect -7514 -23347 -7425 -23232
rect -8131 -23945 -8097 -23355
rect -7514 -23436 -7424 -23347
rect -7226 -23436 -6957 -22508
rect -6680 -23436 -6411 -22508
rect -5803 -23436 -5534 -22508
rect -4941 -23436 -4672 -22508
rect -4038 -23436 -3769 -22508
rect -3007 -23436 -2738 -22508
rect 17379 -22498 17413 -21898
rect 17370 -22610 17423 -22498
rect 17575 -22482 17609 -21898
rect 17566 -22610 17619 -22482
rect 17370 -22743 18238 -22610
rect -7514 -23499 -2289 -23436
rect -7514 -23504 -5941 -23499
rect -5043 -23504 -3241 -23499
rect -15041 -24929 -15007 -24638
rect -14845 -24929 -14811 -24638
rect -14649 -24929 -14615 -24638
rect -13298 -24929 -13264 -24638
rect -13102 -24929 -13068 -24638
rect -12906 -24929 -12872 -24638
rect -12341 -24929 -12307 -24638
rect -12145 -24929 -12111 -24638
rect -11949 -24929 -11915 -24638
rect -10598 -24929 -10564 -24638
rect -10402 -24929 -10368 -24638
rect -10206 -24929 -10172 -24638
rect -9716 -24929 -9682 -24638
rect -9520 -24929 -9486 -24638
rect -9324 -24929 -9290 -24638
rect -15101 -24932 -14606 -24929
rect -13359 -24930 -11906 -24929
rect -15388 -24934 -14284 -24932
rect -13359 -24934 -11593 -24930
rect -10659 -24934 -9281 -24929
rect -15388 -24997 -9281 -24934
rect -17044 -25769 -16999 -25645
rect -18674 -25786 -18485 -25779
rect -23485 -25905 -23427 -25809
rect -18711 -25793 -18485 -25786
rect -17667 -25793 -16898 -25769
rect -21610 -25905 -21552 -25809
rect -20347 -25835 -16898 -25793
rect -23485 -25946 -21552 -25905
rect -23372 -25984 -23314 -25981
rect -21517 -25984 -21459 -25888
rect -20347 -25946 -17002 -25835
rect -20347 -25965 -18771 -25946
rect -23372 -26025 -21459 -25984
rect -23372 -26118 -23314 -26025
rect -23258 -26063 -23200 -26062
rect -20696 -26063 -20638 -25967
rect -23258 -26104 -20638 -26063
rect -23258 -26199 -23200 -26104
rect -20603 -26140 -20545 -26044
rect -23113 -26181 -20545 -26140
rect -23113 -26277 -23055 -26181
rect -22953 -27515 -22919 -27223
rect -20347 -26960 -20175 -25965
rect -18943 -26136 -18771 -25965
rect -18115 -25963 -17497 -25946
rect -18115 -25992 -17672 -25963
rect -18114 -26006 -17672 -25992
rect -18114 -26055 -16825 -26006
rect -19125 -26235 -18407 -26136
rect -19077 -26501 -19043 -26235
rect -18881 -26501 -18847 -26235
rect -18685 -26501 -18651 -26235
rect -18489 -26501 -18455 -26235
rect -18104 -26472 -18070 -26055
rect -17908 -26472 -17874 -26055
rect -17712 -26105 -16825 -26055
rect -17712 -26472 -17678 -26105
rect -17495 -26271 -17461 -26105
rect -17299 -26271 -17265 -26105
rect -17103 -26271 -17069 -26105
rect -16907 -26271 -16873 -26105
rect -15388 -25000 -14284 -24997
rect -12066 -24998 -11593 -24997
rect -7514 -25199 -7425 -23504
rect -7265 -23795 -7231 -23504
rect -7069 -23795 -7035 -23504
rect -6873 -23795 -6839 -23504
rect -6428 -23795 -6394 -23504
rect -6232 -23795 -6198 -23504
rect -6036 -23795 -6002 -23504
rect -4565 -23795 -4531 -23504
rect -4369 -23795 -4335 -23504
rect -4173 -23795 -4139 -23504
rect -3728 -23795 -3694 -23504
rect -3532 -23795 -3498 -23504
rect -3336 -23795 -3302 -23504
rect -7167 -25196 -7133 -24905
rect -6971 -25196 -6937 -24905
rect -6775 -25196 -6741 -24905
rect -5424 -25196 -5390 -24905
rect -5228 -25196 -5194 -24905
rect -5032 -25196 -4998 -24905
rect -4467 -25196 -4433 -24905
rect -4271 -25196 -4237 -24905
rect -4075 -25196 -4041 -24905
rect -2724 -25196 -2690 -24905
rect -2528 -25196 -2494 -24905
rect -2332 -25196 -2298 -24905
rect -1842 -25196 -1808 -24905
rect -1646 -25196 -1612 -24905
rect -1450 -25150 -1416 -24905
rect -1522 -25196 -1399 -25150
rect -7227 -25199 -6732 -25196
rect -5485 -25197 -4032 -25196
rect -7514 -25201 -6410 -25199
rect -5485 -25201 -3719 -25197
rect -2785 -25201 -1399 -25196
rect -7514 -25264 -1399 -25201
rect -7514 -25267 -6410 -25264
rect -20349 -27047 -20173 -26960
rect -5343 -25816 -5228 -25264
rect -4192 -25265 -3719 -25264
rect -5348 -25952 -5225 -25816
rect -2777 -25960 -2662 -25264
rect -1522 -25286 -1399 -25264
rect -1108 -25151 -1074 -24888
rect -1228 -25180 -1074 -25151
rect -912 -25180 -878 -24888
rect -1228 -25181 -873 -25180
rect -370 -25181 -336 -24888
rect -174 -25181 -140 -24888
rect 22 -25181 56 -24888
rect 218 -25181 252 -24888
rect 625 -25141 659 -24975
rect 821 -25141 855 -24975
rect 1017 -25141 1051 -24975
rect 1213 -25141 1247 -24975
rect 1430 -25141 1464 -24774
rect 577 -25181 1464 -25141
rect 1626 -25181 1660 -24774
rect 1822 -25138 1856 -24774
rect 1750 -25181 1873 -25138
rect -1228 -25260 1873 -25181
rect -1228 -25287 -1105 -25260
rect -2781 -26096 -2658 -25960
rect -293 -26068 -178 -25260
rect 1750 -25274 1873 -25260
rect 2230 -25139 2264 -24973
rect 2426 -25139 2460 -24973
rect 2622 -25139 2656 -24973
rect 2818 -25139 2852 -24973
rect 3035 -25139 3069 -24772
rect 2139 -25189 3069 -25139
rect 3231 -25189 3265 -24772
rect 3427 -25162 3461 -24772
rect 3367 -25189 3490 -25162
rect 2139 -25238 3490 -25189
rect 2139 -25275 2262 -25238
rect 3029 -25253 3490 -25238
rect 3367 -25298 3490 -25253
rect -298 -26130 8 -26068
rect -298 -26131 -175 -26130
rect 3854 -25164 3888 -24897
rect 20586 -21308 20620 -21017
rect 20782 -21308 20816 -21017
rect 20978 -21308 21012 -21017
rect 21423 -21308 21457 -21017
rect 21619 -21308 21653 -21017
rect 21815 -21308 21849 -21017
rect 23286 -21308 23320 -21017
rect 23482 -21308 23516 -21017
rect 23678 -21308 23712 -21017
rect 24123 -21308 24157 -21017
rect 24319 -21308 24353 -21017
rect 24515 -21308 24549 -21017
rect 24709 -21077 24798 -21017
rect 26910 -21077 27628 -21013
rect 24709 -21112 27628 -21077
rect 24709 -21302 27264 -21112
rect 27931 -21193 27965 -20776
rect 28127 -21193 28161 -20776
rect 28323 -21143 28357 -20776
rect 28540 -21143 28574 -20977
rect 28736 -21143 28770 -20977
rect 28932 -21143 28966 -20977
rect 29128 -21143 29162 -20977
rect 28323 -21193 29210 -21143
rect 27921 -21242 29210 -21193
rect 27921 -21256 28363 -21242
rect 27920 -21285 28363 -21256
rect 27920 -21302 28538 -21285
rect 24709 -21371 29033 -21302
rect 18700 -22709 18734 -22418
rect 18896 -22709 18930 -22418
rect 19092 -22709 19126 -22418
rect 19582 -22709 19616 -22418
rect 19778 -22709 19812 -22418
rect 19974 -22709 20008 -22418
rect 21325 -22709 21359 -22418
rect 21521 -22709 21555 -22418
rect 21717 -22709 21751 -22418
rect 22282 -22709 22316 -22418
rect 22478 -22709 22512 -22418
rect 22674 -22709 22708 -22418
rect 24025 -22709 24059 -22418
rect 24221 -22709 24255 -22418
rect 24417 -22709 24451 -22418
rect 18691 -22714 20069 -22709
rect 21316 -22710 22769 -22709
rect 21003 -22714 22769 -22710
rect 24016 -22712 24511 -22709
rect 24709 -22712 24798 -21371
rect 26922 -21413 29033 -21371
rect 26922 -21420 29137 -21413
rect 29210 -21420 29272 -21392
rect 26922 -21455 29272 -21420
rect 27324 -21462 27550 -21455
rect 27361 -21469 27550 -21462
rect 28368 -21472 29272 -21455
rect 28368 -21479 29137 -21472
rect 26922 -21518 27364 -21503
rect 26922 -21567 28211 -21518
rect 26932 -21984 26966 -21567
rect 27128 -21984 27162 -21567
rect 27324 -21617 28211 -21567
rect 28374 -21605 28419 -21479
rect 27324 -21984 27358 -21617
rect 27541 -21783 27575 -21617
rect 27737 -21783 27771 -21617
rect 27933 -21783 27967 -21617
rect 28129 -21783 28163 -21617
rect 23694 -22714 24798 -22712
rect 18691 -22777 24798 -22714
rect 21003 -22778 21476 -22777
rect 21193 -22997 21425 -22778
rect 23694 -22780 24798 -22777
rect 21135 -23061 21577 -22997
rect 21145 -23578 21179 -23061
rect 21341 -23578 21375 -23061
rect 21537 -23578 21571 -23061
rect 5946 -24632 6085 -24578
rect 3768 -25189 3891 -25164
rect 4050 -25189 4084 -24897
rect 3768 -25194 4089 -25189
rect 4592 -25193 4626 -24897
rect 4788 -25193 4822 -24897
rect 4984 -25193 5018 -24897
rect 5180 -25159 5214 -24897
rect 5124 -25193 5247 -25159
rect 4592 -25194 5247 -25193
rect 3768 -25262 5247 -25194
rect 3768 -25267 4664 -25262
rect 3768 -25300 3891 -25267
rect 5124 -25295 5247 -25262
rect 6341 -25069 6375 -24886
rect 6341 -25158 6381 -25069
rect 6537 -25069 6571 -24886
rect 6340 -25198 6463 -25158
rect 6530 -25198 6576 -25069
rect 6733 -25073 6767 -24886
rect 6847 -25069 6881 -24886
rect 7024 -24626 7163 -24572
rect 6728 -25198 6774 -25073
rect 6841 -25198 6887 -25069
rect 7043 -25074 7077 -24886
rect 7156 -25064 7190 -24886
rect 7037 -25198 7083 -25074
rect 7150 -25198 7196 -25064
rect 7352 -25076 7386 -24886
rect 7347 -25198 7393 -25076
rect 6340 -25267 7393 -25198
rect 6340 -25294 6463 -25267
rect 8135 -24637 8280 -24502
rect 7852 -25652 7975 -25651
rect -7064 -26883 -6925 -26829
rect -22757 -27499 -22723 -27223
rect -22215 -27499 -22181 -27223
rect -22019 -27499 -21985 -27223
rect -21823 -27499 -21789 -27223
rect -21627 -27499 -21593 -27223
rect -6669 -27320 -6635 -27137
rect -6669 -27449 -6629 -27320
rect -6473 -27320 -6439 -27137
rect -6480 -27449 -6434 -27320
rect -6277 -27324 -6243 -27137
rect -6163 -27320 -6129 -27137
rect -5986 -26877 -5847 -26823
rect -5347 -26719 -5224 -26583
rect -6282 -27449 -6236 -27324
rect -6169 -27449 -6123 -27320
rect -5967 -27325 -5933 -27137
rect -5854 -27315 -5820 -27137
rect -5973 -27449 -5927 -27325
rect -5860 -27449 -5814 -27315
rect -5658 -27327 -5624 -27137
rect -5663 -27449 -5617 -27327
rect -22775 -27515 -20173 -27499
rect -22963 -27582 -20173 -27515
rect -22775 -27591 -20173 -27582
rect -6669 -27556 -5617 -27449
rect -5342 -27556 -5227 -26719
rect -4564 -26883 -4425 -26829
rect -4169 -27320 -4135 -27137
rect -4169 -27449 -4129 -27320
rect -3973 -27320 -3939 -27137
rect -3980 -27449 -3934 -27320
rect -3777 -27324 -3743 -27137
rect -3663 -27320 -3629 -27137
rect -3486 -26877 -3347 -26823
rect -2780 -26684 -2657 -26548
rect -3782 -27449 -3736 -27324
rect -3669 -27449 -3623 -27320
rect -3467 -27325 -3433 -27137
rect -3354 -27315 -3320 -27137
rect -3473 -27449 -3427 -27325
rect -3360 -27449 -3314 -27315
rect -3158 -27327 -3124 -27137
rect -3163 -27449 -3117 -27327
rect -4169 -27518 -3117 -27449
rect -3855 -27556 -3262 -27518
rect -2774 -27556 -2660 -26684
rect -2064 -26883 -1925 -26829
rect -1669 -27320 -1635 -27137
rect -1669 -27449 -1629 -27320
rect -1473 -27320 -1439 -27137
rect -1480 -27449 -1434 -27320
rect -1277 -27324 -1243 -27137
rect -1163 -27320 -1129 -27137
rect -986 -26877 -847 -26823
rect -297 -26684 -174 -26548
rect -1282 -27449 -1236 -27324
rect -1169 -27449 -1123 -27320
rect -967 -27325 -933 -27137
rect -854 -27315 -820 -27137
rect -973 -27449 -927 -27325
rect -860 -27449 -814 -27315
rect -658 -27327 -624 -27137
rect -663 -27449 -617 -27327
rect -1669 -27518 -617 -27449
rect -1339 -27556 -746 -27518
rect -292 -27556 -177 -26684
rect 436 -26883 575 -26829
rect 831 -27320 865 -27137
rect 831 -27449 871 -27320
rect 1027 -27320 1061 -27137
rect 1020 -27449 1066 -27320
rect 1223 -27324 1257 -27137
rect 1337 -27320 1371 -27137
rect 1514 -26877 1653 -26823
rect 1218 -27449 1264 -27324
rect 1331 -27449 1377 -27320
rect 1533 -27325 1567 -27137
rect 1646 -27315 1680 -27137
rect 2936 -26883 3075 -26829
rect 1527 -27449 1573 -27325
rect 1640 -27449 1686 -27315
rect 1842 -27327 1876 -27137
rect 1837 -27449 1883 -27327
rect 831 -27518 1883 -27449
rect 3331 -27320 3365 -27137
rect 3331 -27449 3371 -27320
rect 3527 -27320 3561 -27137
rect 3520 -27449 3566 -27320
rect 3723 -27324 3757 -27137
rect 3837 -27320 3871 -27137
rect 4014 -26877 4153 -26823
rect 7851 -25695 7975 -25652
rect 3718 -27449 3764 -27324
rect 3831 -27449 3877 -27320
rect 4033 -27325 4067 -27137
rect 4146 -27315 4180 -27137
rect 7851 -26503 7909 -25695
rect 7995 -26253 8118 -26209
rect 5936 -26883 6075 -26829
rect 4027 -27449 4073 -27325
rect 4140 -27449 4186 -27315
rect 4342 -27327 4376 -27137
rect 4337 -27449 4383 -27327
rect 3331 -27518 4383 -27449
rect 6331 -27320 6365 -27137
rect 6331 -27449 6371 -27320
rect 6527 -27320 6561 -27137
rect 6520 -27449 6566 -27320
rect 6723 -27324 6757 -27137
rect 6837 -27320 6871 -27137
rect 7014 -26877 7153 -26823
rect 6718 -27449 6764 -27324
rect 6831 -27449 6877 -27320
rect 7033 -27325 7067 -27137
rect 7146 -27315 7180 -27137
rect 7027 -27449 7073 -27325
rect 7140 -27449 7186 -27315
rect 7342 -27327 7376 -27137
rect 7337 -27449 7383 -27327
rect 1195 -27556 1788 -27518
rect 3608 -27556 4201 -27518
rect 6331 -27556 7383 -27449
rect -7534 -27749 7428 -27556
rect 7852 -27913 7908 -26503
rect 7951 -26881 8016 -26744
rect 7954 -27641 8008 -26881
rect 8059 -27641 8113 -26253
rect 8158 -27858 8214 -24637
rect 17374 -24835 17408 -24444
rect 17367 -24962 17415 -24835
rect 17570 -24829 17604 -24444
rect 17564 -24962 17612 -24829
rect 18320 -24835 18354 -24444
rect 18313 -24962 18361 -24835
rect 18516 -24829 18550 -24444
rect 18510 -24962 18558 -24829
rect 18991 -24962 19077 -24954
rect 16544 -24974 19077 -24962
rect 19236 -24974 19270 -24678
rect 19432 -24974 19466 -24678
rect 19628 -24974 19662 -24678
rect 19824 -24974 19858 -24678
rect 20111 -24970 20174 -24956
rect 20366 -24970 20400 -24678
rect 20562 -24970 20596 -24678
rect 20792 -24962 20866 -24956
rect 21095 -24962 21129 -24671
rect 21291 -24962 21325 -24671
rect 21487 -24935 21521 -24671
rect 21975 -24935 22009 -24100
rect 22171 -24935 22205 -24100
rect 22375 -24935 22409 -24100
rect 22571 -24935 22605 -24100
rect 22975 -24935 23009 -24100
rect 23171 -24935 23205 -24100
rect 23375 -24935 23409 -24100
rect 23571 -24935 23605 -24100
rect 23975 -24935 24009 -24100
rect 24171 -24935 24205 -24100
rect 24375 -24935 24409 -24100
rect 24571 -24935 24605 -24100
rect 24709 -24935 24798 -22780
rect 28379 -22195 28413 -21605
rect 28569 -21602 28614 -21479
rect 28575 -22195 28609 -21602
rect 28991 -21603 29036 -21479
rect 29210 -21486 29272 -21472
rect 28998 -22195 29032 -21603
rect 35398 -21024 35432 -20758
rect 35594 -21024 35628 -20758
rect 35790 -21024 35824 -20758
rect 35986 -21024 36020 -20758
rect 35350 -21123 36068 -21024
rect 30368 -21248 32800 -21178
rect 30001 -21300 32800 -21248
rect 30001 -21301 31754 -21300
rect 30001 -21365 30406 -21301
rect 29438 -21375 29536 -21372
rect 30001 -21375 30118 -21365
rect 29438 -21492 30118 -21375
rect 30368 -21460 30406 -21365
rect 29438 -21498 29536 -21492
rect 30371 -21953 30405 -21460
rect 30565 -21458 30603 -21301
rect 30567 -21953 30601 -21458
rect 31157 -21481 31207 -21301
rect 31283 -21478 31333 -21301
rect 31162 -21953 31196 -21481
rect 31292 -21953 31326 -21478
rect 31514 -21463 31557 -21301
rect 31520 -21753 31554 -21463
rect 31711 -21461 31754 -21301
rect 32678 -21313 32800 -21300
rect 35532 -21313 35704 -21123
rect 36371 -21204 36405 -20787
rect 36567 -21204 36601 -20787
rect 36763 -21154 36797 -20787
rect 36980 -21154 37014 -20988
rect 37176 -21154 37210 -20988
rect 37372 -21154 37406 -20988
rect 37568 -21154 37602 -20988
rect 36763 -21204 37650 -21154
rect 36361 -21253 37650 -21204
rect 36361 -21267 36803 -21253
rect 36360 -21296 36803 -21267
rect 36360 -21313 36978 -21296
rect 32678 -21424 37473 -21313
rect 32678 -21431 37577 -21424
rect 37650 -21431 37712 -21403
rect 31716 -21753 31750 -21461
rect 32678 -21466 37712 -21431
rect 21487 -24962 24798 -24935
rect 20792 -24970 24798 -24962
rect 20111 -24974 24798 -24970
rect 16544 -25030 24798 -24974
rect 16544 -25031 20866 -25030
rect 8585 -25848 8733 -25800
rect 8429 -25983 8552 -25939
rect 8270 -26110 8427 -26070
rect 8270 -27641 8324 -26110
rect 8484 -26414 8538 -25983
rect 8385 -26468 8538 -26414
rect 8385 -27641 8439 -26468
rect 8529 -27546 8583 -27516
rect 8627 -27546 8681 -25848
rect 16544 -25502 16670 -25031
rect 18991 -25037 20866 -25031
rect 18991 -25043 20174 -25037
rect 20792 -25043 20866 -25037
rect 21509 -25038 24798 -25030
rect 18991 -25047 19077 -25043
rect 20111 -25054 20174 -25043
rect 12875 -25505 13348 -25504
rect 15566 -25505 16670 -25502
rect 10563 -25568 16670 -25505
rect 10563 -25573 11941 -25568
rect 12875 -25572 14641 -25568
rect 15566 -25570 16670 -25568
rect 13188 -25573 14641 -25572
rect 15888 -25573 16383 -25570
rect 10572 -25864 10606 -25573
rect 10768 -25864 10802 -25573
rect 10964 -25864 10998 -25573
rect 11454 -25864 11488 -25573
rect 11650 -25864 11684 -25573
rect 11846 -25864 11880 -25573
rect 13197 -25864 13231 -25573
rect 13393 -25864 13427 -25573
rect 13589 -25864 13623 -25573
rect 14154 -25864 14188 -25573
rect 14350 -25864 14384 -25573
rect 14546 -25864 14580 -25573
rect 15897 -25864 15931 -25573
rect 16093 -25864 16127 -25573
rect 16289 -25864 16323 -25573
rect 12458 -27265 12492 -26974
rect 12654 -27265 12688 -26974
rect 12850 -27265 12884 -26974
rect 13295 -27265 13329 -26974
rect 13491 -27265 13525 -26974
rect 13687 -27265 13721 -26974
rect 15158 -27265 15192 -26974
rect 15354 -27265 15388 -26974
rect 15550 -27265 15584 -26974
rect 15995 -27265 16029 -26974
rect 16191 -27265 16225 -26974
rect 16387 -27265 16421 -26974
rect 16581 -27265 16670 -25570
rect 29445 -23490 29847 -23424
rect 26950 -24466 26984 -24200
rect 27146 -24466 27180 -24200
rect 27342 -24466 27376 -24200
rect 27538 -24466 27572 -24200
rect 26902 -24565 27620 -24466
rect 27084 -24755 27256 -24565
rect 27923 -24646 27957 -24229
rect 28119 -24646 28153 -24229
rect 28315 -24596 28349 -24229
rect 28532 -24596 28566 -24430
rect 28728 -24596 28762 -24430
rect 28924 -24596 28958 -24430
rect 29120 -24596 29154 -24430
rect 28315 -24646 29202 -24596
rect 27913 -24695 29202 -24646
rect 27913 -24709 28355 -24695
rect 27912 -24738 28355 -24709
rect 27912 -24755 28530 -24738
rect 26914 -24866 29025 -24755
rect 26914 -24908 29129 -24866
rect 27316 -24915 27542 -24908
rect 27353 -24922 27542 -24915
rect 28360 -24932 29129 -24908
rect 26914 -24971 27356 -24956
rect 26914 -25020 28203 -24971
rect 26924 -25437 26958 -25020
rect 27120 -25437 27154 -25020
rect 27316 -25070 28203 -25020
rect 28366 -25058 28411 -24932
rect 27316 -25437 27350 -25070
rect 27533 -25236 27567 -25070
rect 27729 -25236 27763 -25070
rect 27925 -25236 27959 -25070
rect 28121 -25236 28155 -25070
rect 26839 -25486 26974 -25480
rect 26819 -25488 26974 -25486
rect 26291 -25524 26974 -25488
rect 12397 -27270 14199 -27265
rect 15097 -27270 16670 -27265
rect 11445 -27333 16670 -27270
rect 26474 -26551 26610 -25524
rect 26819 -25526 26974 -25524
rect 26839 -25534 26974 -25526
rect 28371 -25648 28405 -25058
rect 28561 -25055 28606 -24932
rect 28567 -25648 28601 -25055
rect 28983 -25056 29028 -24932
rect 28990 -25648 29024 -25056
rect 29445 -24791 29511 -23490
rect 29428 -24904 29512 -24791
rect 29781 -24820 29847 -23490
rect 32678 -23697 32800 -21466
rect 35764 -21473 35990 -21466
rect 35801 -21480 35990 -21473
rect 36808 -21483 37712 -21466
rect 36808 -21490 37577 -21483
rect 35362 -21529 35804 -21514
rect 35362 -21578 36651 -21529
rect 35372 -21995 35406 -21578
rect 35568 -21995 35602 -21578
rect 35764 -21628 36651 -21578
rect 36814 -21616 36859 -21490
rect 35764 -21995 35798 -21628
rect 35981 -21794 36015 -21628
rect 36177 -21794 36211 -21628
rect 36373 -21794 36407 -21628
rect 36569 -21794 36603 -21628
rect 32678 -23819 33310 -23697
rect 30618 -24497 30652 -24231
rect 30814 -24497 30848 -24231
rect 31010 -24497 31044 -24231
rect 31206 -24497 31240 -24231
rect 30570 -24596 31288 -24497
rect 30752 -24786 30924 -24596
rect 31591 -24677 31625 -24260
rect 31787 -24677 31821 -24260
rect 31983 -24627 32017 -24260
rect 32200 -24627 32234 -24461
rect 32396 -24627 32430 -24461
rect 32592 -24627 32626 -24461
rect 32788 -24627 32822 -24461
rect 31983 -24677 32870 -24627
rect 31581 -24726 32870 -24677
rect 31581 -24740 32023 -24726
rect 31580 -24769 32023 -24740
rect 31580 -24786 32198 -24769
rect 30582 -24820 32693 -24786
rect 29781 -24886 32693 -24820
rect 32848 -24861 32927 -24830
rect 30582 -24897 32693 -24886
rect 32748 -24897 32927 -24861
rect 30582 -24939 32927 -24897
rect 30984 -24946 31210 -24939
rect 31021 -24953 31210 -24946
rect 32028 -24944 32927 -24939
rect 32028 -24963 32797 -24944
rect 30582 -25002 31024 -24987
rect 30582 -25051 31871 -25002
rect 30592 -25468 30626 -25051
rect 30788 -25468 30822 -25051
rect 30984 -25101 31871 -25051
rect 32034 -25089 32079 -24963
rect 30984 -25468 31018 -25101
rect 31201 -25267 31235 -25101
rect 31397 -25267 31431 -25101
rect 31593 -25267 31627 -25101
rect 31789 -25267 31823 -25101
rect 30507 -25517 30642 -25511
rect 30487 -25519 30642 -25517
rect 30073 -25555 30642 -25519
rect 30073 -26551 30209 -25555
rect 30487 -25557 30642 -25555
rect 30507 -25565 30642 -25557
rect 32039 -25679 32073 -25089
rect 32229 -25086 32274 -24963
rect 32235 -25679 32269 -25086
rect 32651 -25087 32696 -24963
rect 32848 -24969 32927 -24944
rect 32658 -25679 32692 -25087
rect 33188 -24815 33310 -23819
rect 33098 -24954 33310 -24815
rect 33098 -24982 33237 -24954
rect 26474 -26687 30209 -26551
rect 8529 -27600 8681 -27546
rect 8529 -27641 8583 -27600
rect 26474 -27913 26610 -26687
rect 36819 -22206 36853 -21616
rect 37009 -21613 37054 -21490
rect 37015 -22206 37049 -21613
rect 37431 -21614 37476 -21490
rect 37650 -21497 37712 -21483
rect 37438 -22206 37472 -21614
rect 44261 -21063 44295 -20797
rect 44457 -21063 44491 -20797
rect 44653 -21063 44687 -20797
rect 44849 -21063 44883 -20797
rect 44213 -21147 44931 -21063
rect 40180 -21162 44931 -21147
rect 40180 -21189 44567 -21162
rect 38808 -21259 44567 -21189
rect 45234 -21243 45268 -20826
rect 45430 -21243 45464 -20826
rect 45626 -21193 45660 -20826
rect 45843 -21193 45877 -21027
rect 46039 -21193 46073 -21027
rect 46235 -21193 46269 -21027
rect 46431 -21193 46465 -21027
rect 45626 -21243 46513 -21193
rect 38441 -21312 44567 -21259
rect 45224 -21292 46513 -21243
rect 45224 -21306 45666 -21292
rect 38441 -21376 38846 -21312
rect 37878 -21386 37976 -21383
rect 38441 -21386 38558 -21376
rect 37878 -21503 38558 -21386
rect 38808 -21471 38846 -21376
rect 37878 -21509 37976 -21503
rect 38811 -21964 38845 -21471
rect 39005 -21469 39043 -21312
rect 39007 -21964 39041 -21469
rect 39597 -21492 39647 -21312
rect 39723 -21489 39773 -21312
rect 39602 -21964 39636 -21492
rect 39732 -21964 39766 -21489
rect 39954 -21474 39997 -21312
rect 40151 -21352 44567 -21312
rect 45223 -21335 45666 -21306
rect 45223 -21352 45841 -21335
rect 40151 -21401 46336 -21352
rect 39960 -21764 39994 -21474
rect 40151 -21472 40194 -21401
rect 40156 -21764 40190 -21472
rect 37885 -23501 38287 -23435
rect 35390 -24477 35424 -24211
rect 35586 -24477 35620 -24211
rect 35782 -24477 35816 -24211
rect 35978 -24477 36012 -24211
rect 35342 -24576 36060 -24477
rect 35524 -24766 35696 -24576
rect 36363 -24657 36397 -24240
rect 36559 -24657 36593 -24240
rect 36755 -24607 36789 -24240
rect 36972 -24607 37006 -24441
rect 37168 -24607 37202 -24441
rect 37364 -24607 37398 -24441
rect 37560 -24607 37594 -24441
rect 36755 -24657 37642 -24607
rect 36353 -24706 37642 -24657
rect 36353 -24720 36795 -24706
rect 36352 -24749 36795 -24720
rect 36352 -24766 36970 -24749
rect 35354 -24877 37465 -24766
rect 35354 -24919 37569 -24877
rect 35756 -24926 35982 -24919
rect 35793 -24933 35982 -24926
rect 36800 -24943 37569 -24919
rect 35354 -24982 35796 -24967
rect 35354 -25031 36643 -24982
rect 35364 -25448 35398 -25031
rect 35560 -25448 35594 -25031
rect 35756 -25081 36643 -25031
rect 36806 -25069 36851 -24943
rect 35756 -25448 35790 -25081
rect 35973 -25247 36007 -25081
rect 36169 -25247 36203 -25081
rect 36365 -25247 36399 -25081
rect 36561 -25247 36595 -25081
rect 35279 -25497 35414 -25491
rect 35259 -25499 35414 -25497
rect 34731 -25535 35414 -25499
rect 34914 -26562 35050 -25535
rect 35259 -25537 35414 -25535
rect 35279 -25545 35414 -25537
rect 36811 -25659 36845 -25069
rect 37001 -25066 37046 -24943
rect 37007 -25659 37041 -25066
rect 37423 -25067 37468 -24943
rect 37430 -25659 37464 -25067
rect 37885 -24802 37951 -23501
rect 37868 -24915 37952 -24802
rect 38221 -24831 38287 -23501
rect 41118 -23708 41240 -21401
rect 44225 -21463 46336 -21401
rect 44225 -21470 46440 -21463
rect 46513 -21470 46575 -21442
rect 44225 -21505 46575 -21470
rect 44627 -21512 44853 -21505
rect 44664 -21519 44853 -21512
rect 45671 -21522 46575 -21505
rect 45671 -21529 46440 -21522
rect 44225 -21568 44667 -21553
rect 44225 -21617 45514 -21568
rect 44235 -22034 44269 -21617
rect 44431 -22034 44465 -21617
rect 44627 -21667 45514 -21617
rect 45677 -21655 45722 -21529
rect 44627 -22034 44661 -21667
rect 44844 -21833 44878 -21667
rect 45040 -21833 45074 -21667
rect 45236 -21833 45270 -21667
rect 45432 -21833 45466 -21667
rect 41118 -23830 41750 -23708
rect 39058 -24508 39092 -24242
rect 39254 -24508 39288 -24242
rect 39450 -24508 39484 -24242
rect 39646 -24508 39680 -24242
rect 39010 -24607 39728 -24508
rect 39192 -24797 39364 -24607
rect 40031 -24688 40065 -24271
rect 40227 -24688 40261 -24271
rect 40423 -24638 40457 -24271
rect 40640 -24638 40674 -24472
rect 40836 -24638 40870 -24472
rect 41032 -24638 41066 -24472
rect 41228 -24638 41262 -24472
rect 40423 -24688 41310 -24638
rect 40021 -24737 41310 -24688
rect 40021 -24751 40463 -24737
rect 40020 -24780 40463 -24751
rect 40020 -24797 40638 -24780
rect 39022 -24831 41133 -24797
rect 38221 -24897 41133 -24831
rect 41288 -24872 41367 -24841
rect 39022 -24908 41133 -24897
rect 41188 -24908 41367 -24872
rect 39022 -24950 41367 -24908
rect 39424 -24957 39650 -24950
rect 39461 -24964 39650 -24957
rect 40468 -24955 41367 -24950
rect 40468 -24974 41237 -24955
rect 39022 -25013 39464 -24998
rect 39022 -25062 40311 -25013
rect 39032 -25479 39066 -25062
rect 39228 -25479 39262 -25062
rect 39424 -25112 40311 -25062
rect 40474 -25100 40519 -24974
rect 39424 -25479 39458 -25112
rect 39641 -25278 39675 -25112
rect 39837 -25278 39871 -25112
rect 40033 -25278 40067 -25112
rect 40229 -25278 40263 -25112
rect 38947 -25528 39082 -25522
rect 38927 -25530 39082 -25528
rect 38513 -25566 39082 -25530
rect 38513 -26562 38649 -25566
rect 38927 -25568 39082 -25566
rect 38947 -25576 39082 -25568
rect 40479 -25690 40513 -25100
rect 40669 -25097 40714 -24974
rect 40675 -25690 40709 -25097
rect 41091 -25098 41136 -24974
rect 41288 -24980 41367 -24955
rect 41098 -25690 41132 -25098
rect 41628 -24826 41750 -23830
rect 41538 -24965 41750 -24826
rect 41538 -24993 41677 -24965
rect 34914 -26698 38649 -26562
rect -32565 -28049 26610 -27913
rect 34914 -28112 35050 -26698
rect -32538 -28248 35050 -28112
rect 45682 -22245 45716 -21655
rect 45872 -21652 45917 -21529
rect 45878 -22245 45912 -21652
rect 46294 -21653 46339 -21529
rect 46513 -21536 46575 -21522
rect 46301 -22245 46335 -21653
rect 53459 -21029 53493 -20763
rect 53655 -21029 53689 -20763
rect 53851 -21029 53885 -20763
rect 54047 -21029 54081 -20763
rect 53411 -21097 54129 -21029
rect 49031 -21128 54129 -21097
rect 49031 -21228 53765 -21128
rect 54432 -21209 54466 -20792
rect 54628 -21209 54662 -20792
rect 54824 -21159 54858 -20792
rect 55041 -21159 55075 -20993
rect 55237 -21159 55271 -20993
rect 55433 -21159 55467 -20993
rect 55629 -21159 55663 -20993
rect 54824 -21209 55711 -21159
rect 47671 -21298 53765 -21228
rect 54422 -21258 55711 -21209
rect 54422 -21272 54864 -21258
rect 47304 -21318 53765 -21298
rect 54421 -21301 54864 -21272
rect 54421 -21318 55039 -21301
rect 47304 -21351 55534 -21318
rect 47304 -21415 47709 -21351
rect 46741 -21425 46839 -21422
rect 47304 -21425 47421 -21415
rect 46741 -21542 47421 -21425
rect 47671 -21510 47709 -21415
rect 46741 -21548 46839 -21542
rect 47674 -22003 47708 -21510
rect 47868 -21508 47906 -21351
rect 47870 -22003 47904 -21508
rect 48460 -21531 48510 -21351
rect 48586 -21528 48636 -21351
rect 48465 -22003 48499 -21531
rect 48595 -22003 48629 -21528
rect 48817 -21513 48860 -21351
rect 49014 -21411 55534 -21351
rect 48823 -21803 48857 -21513
rect 49014 -21511 49057 -21411
rect 49019 -21803 49053 -21511
rect 46748 -23540 47150 -23474
rect 44253 -24516 44287 -24250
rect 44449 -24516 44483 -24250
rect 44645 -24516 44679 -24250
rect 44841 -24516 44875 -24250
rect 44205 -24615 44923 -24516
rect 44387 -24805 44559 -24615
rect 45226 -24696 45260 -24279
rect 45422 -24696 45456 -24279
rect 45618 -24646 45652 -24279
rect 45835 -24646 45869 -24480
rect 46031 -24646 46065 -24480
rect 46227 -24646 46261 -24480
rect 46423 -24646 46457 -24480
rect 45618 -24696 46505 -24646
rect 45216 -24745 46505 -24696
rect 45216 -24759 45658 -24745
rect 45215 -24788 45658 -24759
rect 45215 -24805 45833 -24788
rect 44217 -24916 46328 -24805
rect 44217 -24958 46432 -24916
rect 44619 -24965 44845 -24958
rect 44656 -24972 44845 -24965
rect 45663 -24982 46432 -24958
rect 44217 -25021 44659 -25006
rect 44217 -25070 45506 -25021
rect 44227 -25487 44261 -25070
rect 44423 -25487 44457 -25070
rect 44619 -25120 45506 -25070
rect 45669 -25108 45714 -24982
rect 44619 -25487 44653 -25120
rect 44836 -25286 44870 -25120
rect 45032 -25286 45066 -25120
rect 45228 -25286 45262 -25120
rect 45424 -25286 45458 -25120
rect 44142 -25536 44277 -25530
rect 44122 -25538 44277 -25536
rect 43594 -25574 44277 -25538
rect 43777 -26587 43913 -25574
rect 44122 -25576 44277 -25574
rect 44142 -25584 44277 -25576
rect 45674 -25698 45708 -25108
rect 45864 -25105 45909 -24982
rect 45870 -25698 45904 -25105
rect 46286 -25106 46331 -24982
rect 46293 -25698 46327 -25106
rect 46748 -24841 46814 -23540
rect 46731 -24954 46815 -24841
rect 47084 -24870 47150 -23540
rect 49981 -23747 50103 -21411
rect 53423 -21429 55534 -21411
rect 53423 -21436 55638 -21429
rect 55711 -21436 55773 -21408
rect 53423 -21471 55773 -21436
rect 53825 -21478 54051 -21471
rect 53862 -21485 54051 -21478
rect 54869 -21488 55773 -21471
rect 54869 -21495 55638 -21488
rect 53423 -21534 53865 -21519
rect 53423 -21583 54712 -21534
rect 53433 -22000 53467 -21583
rect 53629 -22000 53663 -21583
rect 53825 -21633 54712 -21583
rect 54875 -21621 54920 -21495
rect 53825 -22000 53859 -21633
rect 54042 -21799 54076 -21633
rect 54238 -21799 54272 -21633
rect 54434 -21799 54468 -21633
rect 54630 -21799 54664 -21633
rect 49981 -23869 50613 -23747
rect 47921 -24547 47955 -24281
rect 48117 -24547 48151 -24281
rect 48313 -24547 48347 -24281
rect 48509 -24547 48543 -24281
rect 47873 -24646 48591 -24547
rect 48055 -24836 48227 -24646
rect 48894 -24727 48928 -24310
rect 49090 -24727 49124 -24310
rect 49286 -24677 49320 -24310
rect 49503 -24677 49537 -24511
rect 49699 -24677 49733 -24511
rect 49895 -24677 49929 -24511
rect 50091 -24677 50125 -24511
rect 49286 -24727 50173 -24677
rect 48884 -24776 50173 -24727
rect 48884 -24790 49326 -24776
rect 48883 -24819 49326 -24790
rect 48883 -24836 49501 -24819
rect 47885 -24870 49996 -24836
rect 47084 -24936 49996 -24870
rect 50151 -24911 50230 -24880
rect 47885 -24947 49996 -24936
rect 50051 -24947 50230 -24911
rect 47885 -24989 50230 -24947
rect 48287 -24996 48513 -24989
rect 48324 -25003 48513 -24996
rect 49331 -24994 50230 -24989
rect 49331 -25013 50100 -24994
rect 47885 -25052 48327 -25037
rect 47885 -25101 49174 -25052
rect 47895 -25518 47929 -25101
rect 48091 -25518 48125 -25101
rect 48287 -25151 49174 -25101
rect 49337 -25139 49382 -25013
rect 48287 -25518 48321 -25151
rect 48504 -25317 48538 -25151
rect 48700 -25317 48734 -25151
rect 48896 -25317 48930 -25151
rect 49092 -25317 49126 -25151
rect 47810 -25567 47945 -25561
rect 47790 -25569 47945 -25567
rect 47376 -25605 47945 -25569
rect 43777 -26601 43960 -26587
rect 47376 -26601 47512 -25605
rect 47790 -25607 47945 -25605
rect 47810 -25615 47945 -25607
rect 49342 -25729 49376 -25139
rect 49532 -25136 49577 -25013
rect 49538 -25729 49572 -25136
rect 49954 -25137 49999 -25013
rect 50151 -25019 50230 -24994
rect 49961 -25729 49995 -25137
rect 50491 -24865 50613 -23869
rect 50401 -25004 50613 -24865
rect 50401 -25032 50540 -25004
rect 43777 -26737 47512 -26601
rect 43824 -28345 43960 -26737
rect 54880 -22211 54914 -21621
rect 55070 -21618 55115 -21495
rect 55076 -22211 55110 -21618
rect 55492 -21619 55537 -21495
rect 55711 -21502 55773 -21488
rect 55499 -22211 55533 -21619
rect 62213 -20963 62247 -20697
rect 62409 -20963 62443 -20697
rect 62605 -20963 62639 -20697
rect 62801 -20963 62835 -20697
rect 62165 -21000 62883 -20963
rect 58214 -21062 62883 -21000
rect 58214 -21194 62519 -21062
rect 63186 -21143 63220 -20726
rect 63382 -21143 63416 -20726
rect 63578 -21093 63612 -20726
rect 63795 -21093 63829 -20927
rect 63991 -21093 64025 -20927
rect 64187 -21093 64221 -20927
rect 64383 -21093 64417 -20927
rect 63578 -21143 64465 -21093
rect 56869 -21252 62519 -21194
rect 63176 -21192 64465 -21143
rect 63176 -21206 63618 -21192
rect 63175 -21235 63618 -21206
rect 63175 -21252 63793 -21235
rect 56869 -21264 64288 -21252
rect 56502 -21317 64288 -21264
rect 56502 -21381 56907 -21317
rect 55939 -21391 56037 -21388
rect 56502 -21391 56619 -21381
rect 55939 -21508 56619 -21391
rect 56869 -21476 56907 -21381
rect 55939 -21514 56037 -21508
rect 56872 -21969 56906 -21476
rect 57066 -21474 57104 -21317
rect 57068 -21969 57102 -21474
rect 57658 -21497 57708 -21317
rect 57784 -21494 57834 -21317
rect 57663 -21969 57697 -21497
rect 57793 -21969 57827 -21494
rect 58015 -21479 58058 -21317
rect 58212 -21363 64288 -21317
rect 58212 -21370 64392 -21363
rect 64465 -21370 64527 -21342
rect 58212 -21379 64527 -21370
rect 58021 -21769 58055 -21479
rect 58212 -21477 58255 -21379
rect 58217 -21769 58251 -21477
rect 55946 -23506 56348 -23440
rect 53451 -24482 53485 -24216
rect 53647 -24482 53681 -24216
rect 53843 -24482 53877 -24216
rect 54039 -24482 54073 -24216
rect 53403 -24581 54121 -24482
rect 53585 -24771 53757 -24581
rect 54424 -24662 54458 -24245
rect 54620 -24662 54654 -24245
rect 54816 -24612 54850 -24245
rect 55033 -24612 55067 -24446
rect 55229 -24612 55263 -24446
rect 55425 -24612 55459 -24446
rect 55621 -24612 55655 -24446
rect 54816 -24662 55703 -24612
rect 54414 -24711 55703 -24662
rect 54414 -24725 54856 -24711
rect 54413 -24754 54856 -24725
rect 54413 -24771 55031 -24754
rect 53415 -24882 55526 -24771
rect 53415 -24924 55630 -24882
rect 53817 -24931 54043 -24924
rect 53854 -24938 54043 -24931
rect 54861 -24948 55630 -24924
rect 53415 -24987 53857 -24972
rect 53415 -25036 54704 -24987
rect 53425 -25453 53459 -25036
rect 53621 -25453 53655 -25036
rect 53817 -25086 54704 -25036
rect 54867 -25074 54912 -24948
rect 53817 -25453 53851 -25086
rect 54034 -25252 54068 -25086
rect 54230 -25252 54264 -25086
rect 54426 -25252 54460 -25086
rect 54622 -25252 54656 -25086
rect 53340 -25502 53475 -25496
rect 53320 -25504 53475 -25502
rect 52792 -25540 53475 -25504
rect 52975 -26567 53111 -25540
rect 53320 -25542 53475 -25540
rect 53340 -25550 53475 -25542
rect 54872 -25664 54906 -25074
rect 55062 -25071 55107 -24948
rect 55068 -25664 55102 -25071
rect 55484 -25072 55529 -24948
rect 55491 -25664 55525 -25072
rect 55946 -24807 56012 -23506
rect 55929 -24920 56013 -24807
rect 56282 -24836 56348 -23506
rect 59179 -23713 59301 -21379
rect 62177 -21405 64527 -21379
rect 62579 -21412 62805 -21405
rect 62616 -21419 62805 -21412
rect 63623 -21422 64527 -21405
rect 63623 -21429 64392 -21422
rect 62177 -21468 62619 -21453
rect 62177 -21517 63466 -21468
rect 62187 -21934 62221 -21517
rect 62383 -21934 62417 -21517
rect 62579 -21567 63466 -21517
rect 63629 -21555 63674 -21429
rect 62579 -21934 62613 -21567
rect 62796 -21733 62830 -21567
rect 62992 -21733 63026 -21567
rect 63188 -21733 63222 -21567
rect 63384 -21733 63418 -21567
rect 59179 -23835 59811 -23713
rect 57119 -24513 57153 -24247
rect 57315 -24513 57349 -24247
rect 57511 -24513 57545 -24247
rect 57707 -24513 57741 -24247
rect 57071 -24612 57789 -24513
rect 57253 -24802 57425 -24612
rect 58092 -24693 58126 -24276
rect 58288 -24693 58322 -24276
rect 58484 -24643 58518 -24276
rect 58701 -24643 58735 -24477
rect 58897 -24643 58931 -24477
rect 59093 -24643 59127 -24477
rect 59289 -24643 59323 -24477
rect 58484 -24693 59371 -24643
rect 58082 -24742 59371 -24693
rect 58082 -24756 58524 -24742
rect 58081 -24785 58524 -24756
rect 58081 -24802 58699 -24785
rect 57083 -24836 59194 -24802
rect 56282 -24902 59194 -24836
rect 59349 -24877 59428 -24846
rect 57083 -24913 59194 -24902
rect 59249 -24913 59428 -24877
rect 57083 -24955 59428 -24913
rect 57485 -24962 57711 -24955
rect 57522 -24969 57711 -24962
rect 58529 -24960 59428 -24955
rect 58529 -24979 59298 -24960
rect 57083 -25018 57525 -25003
rect 57083 -25067 58372 -25018
rect 57093 -25484 57127 -25067
rect 57289 -25484 57323 -25067
rect 57485 -25117 58372 -25067
rect 58535 -25105 58580 -24979
rect 57485 -25484 57519 -25117
rect 57702 -25283 57736 -25117
rect 57898 -25283 57932 -25117
rect 58094 -25283 58128 -25117
rect 58290 -25283 58324 -25117
rect 57008 -25533 57143 -25527
rect 56988 -25535 57143 -25533
rect 56574 -25571 57143 -25535
rect 56574 -26567 56710 -25571
rect 56988 -25573 57143 -25571
rect 57008 -25581 57143 -25573
rect 58540 -25695 58574 -25105
rect 58730 -25102 58775 -24979
rect 58736 -25695 58770 -25102
rect 59152 -25103 59197 -24979
rect 59349 -24985 59428 -24960
rect 59159 -25695 59193 -25103
rect 59689 -24831 59811 -23835
rect 59599 -24970 59811 -24831
rect 59599 -24998 59738 -24970
rect 52975 -26703 56710 -26567
rect -32538 -28481 43960 -28345
rect 52975 -28600 53111 -26703
rect 63634 -22145 63668 -21555
rect 63824 -21552 63869 -21429
rect 63830 -22145 63864 -21552
rect 64246 -21553 64291 -21429
rect 64465 -21436 64527 -21422
rect 64253 -22145 64287 -21553
rect 71366 -20946 71400 -20680
rect 71562 -20946 71596 -20680
rect 71758 -20946 71792 -20680
rect 71954 -20946 71988 -20680
rect 71318 -21021 72036 -20946
rect 66961 -21045 72036 -21021
rect 66961 -21128 71672 -21045
rect 72339 -21126 72373 -20709
rect 72535 -21126 72569 -20709
rect 72731 -21076 72765 -20709
rect 72948 -21076 72982 -20910
rect 73144 -21076 73178 -20910
rect 73340 -21076 73374 -20910
rect 73536 -21076 73570 -20910
rect 72731 -21126 73618 -21076
rect 65623 -21198 71672 -21128
rect 72329 -21175 73618 -21126
rect 72329 -21189 72771 -21175
rect 65256 -21235 71672 -21198
rect 72328 -21218 72771 -21189
rect 72328 -21235 72946 -21218
rect 65256 -21251 73441 -21235
rect 65256 -21315 65661 -21251
rect 64693 -21325 64791 -21322
rect 65256 -21325 65373 -21315
rect 64693 -21442 65373 -21325
rect 65623 -21410 65661 -21315
rect 64693 -21448 64791 -21442
rect 65626 -21903 65660 -21410
rect 65820 -21408 65858 -21251
rect 65822 -21903 65856 -21408
rect 66412 -21431 66462 -21251
rect 66538 -21428 66588 -21251
rect 66417 -21903 66451 -21431
rect 66547 -21903 66581 -21428
rect 66769 -21413 66812 -21251
rect 66961 -21285 73441 -21251
rect 66775 -21703 66809 -21413
rect 66966 -21411 67009 -21285
rect 66971 -21703 67005 -21411
rect 64700 -23440 65102 -23374
rect 62205 -24416 62239 -24150
rect 62401 -24416 62435 -24150
rect 62597 -24416 62631 -24150
rect 62793 -24416 62827 -24150
rect 62157 -24515 62875 -24416
rect 62339 -24705 62511 -24515
rect 63178 -24596 63212 -24179
rect 63374 -24596 63408 -24179
rect 63570 -24546 63604 -24179
rect 63787 -24546 63821 -24380
rect 63983 -24546 64017 -24380
rect 64179 -24546 64213 -24380
rect 64375 -24546 64409 -24380
rect 63570 -24596 64457 -24546
rect 63168 -24645 64457 -24596
rect 63168 -24659 63610 -24645
rect 63167 -24688 63610 -24659
rect 63167 -24705 63785 -24688
rect 62169 -24816 64280 -24705
rect 62169 -24858 64384 -24816
rect 62571 -24865 62797 -24858
rect 62608 -24872 62797 -24865
rect 63615 -24882 64384 -24858
rect 62169 -24921 62611 -24906
rect 62169 -24970 63458 -24921
rect 62179 -25387 62213 -24970
rect 62375 -25387 62409 -24970
rect 62571 -25020 63458 -24970
rect 63621 -25008 63666 -24882
rect 62571 -25387 62605 -25020
rect 62788 -25186 62822 -25020
rect 62984 -25186 63018 -25020
rect 63180 -25186 63214 -25020
rect 63376 -25186 63410 -25020
rect 62094 -25436 62229 -25430
rect 62074 -25438 62229 -25436
rect 61546 -25474 62229 -25438
rect 61729 -26501 61865 -25474
rect 62074 -25476 62229 -25474
rect 62094 -25484 62229 -25476
rect 63626 -25598 63660 -25008
rect 63816 -25005 63861 -24882
rect 63822 -25598 63856 -25005
rect 64238 -25006 64283 -24882
rect 64245 -25598 64279 -25006
rect 64700 -24741 64766 -23440
rect 64683 -24854 64767 -24741
rect 65036 -24770 65102 -23440
rect 67933 -23647 68055 -21285
rect 71330 -21346 73441 -21285
rect 71330 -21353 73545 -21346
rect 73618 -21353 73680 -21325
rect 71330 -21388 73680 -21353
rect 71732 -21395 71958 -21388
rect 71769 -21402 71958 -21395
rect 72776 -21405 73680 -21388
rect 72776 -21412 73545 -21405
rect 71330 -21451 71772 -21436
rect 71330 -21500 72619 -21451
rect 71340 -21917 71374 -21500
rect 71536 -21917 71570 -21500
rect 71732 -21550 72619 -21500
rect 72782 -21538 72827 -21412
rect 71732 -21917 71766 -21550
rect 71949 -21716 71983 -21550
rect 72145 -21716 72179 -21550
rect 72341 -21716 72375 -21550
rect 72537 -21716 72571 -21550
rect 67933 -23769 68565 -23647
rect 65873 -24447 65907 -24181
rect 66069 -24447 66103 -24181
rect 66265 -24447 66299 -24181
rect 66461 -24447 66495 -24181
rect 65825 -24546 66543 -24447
rect 66007 -24736 66179 -24546
rect 66846 -24627 66880 -24210
rect 67042 -24627 67076 -24210
rect 67238 -24577 67272 -24210
rect 67455 -24577 67489 -24411
rect 67651 -24577 67685 -24411
rect 67847 -24577 67881 -24411
rect 68043 -24577 68077 -24411
rect 67238 -24627 68125 -24577
rect 66836 -24676 68125 -24627
rect 66836 -24690 67278 -24676
rect 66835 -24719 67278 -24690
rect 66835 -24736 67453 -24719
rect 65837 -24770 67948 -24736
rect 65036 -24836 67948 -24770
rect 68103 -24811 68182 -24780
rect 65837 -24847 67948 -24836
rect 68003 -24847 68182 -24811
rect 65837 -24889 68182 -24847
rect 66239 -24896 66465 -24889
rect 66276 -24903 66465 -24896
rect 67283 -24894 68182 -24889
rect 67283 -24913 68052 -24894
rect 65837 -24952 66279 -24937
rect 65837 -25001 67126 -24952
rect 65847 -25418 65881 -25001
rect 66043 -25418 66077 -25001
rect 66239 -25051 67126 -25001
rect 67289 -25039 67334 -24913
rect 66239 -25418 66273 -25051
rect 66456 -25217 66490 -25051
rect 66652 -25217 66686 -25051
rect 66848 -25217 66882 -25051
rect 67044 -25217 67078 -25051
rect 65762 -25467 65897 -25461
rect 65742 -25469 65897 -25467
rect 65328 -25505 65897 -25469
rect 65328 -26501 65464 -25505
rect 65742 -25507 65897 -25505
rect 65762 -25515 65897 -25507
rect 67294 -25629 67328 -25039
rect 67484 -25036 67529 -24913
rect 67490 -25629 67524 -25036
rect 67906 -25037 67951 -24913
rect 68103 -24919 68182 -24894
rect 67913 -25629 67947 -25037
rect 68443 -24765 68565 -23769
rect 68353 -24904 68565 -24765
rect 68353 -24932 68492 -24904
rect 61729 -26637 65464 -26501
rect -32592 -28736 53111 -28600
rect 8289 -28886 8425 -28884
rect 61729 -28886 61865 -26637
rect 72787 -22128 72821 -21538
rect 72977 -21535 73022 -21412
rect 72983 -22128 73017 -21535
rect 73399 -21536 73444 -21412
rect 73618 -21419 73680 -21405
rect 73406 -22128 73440 -21536
rect 80730 -20908 80764 -20642
rect 80926 -20908 80960 -20642
rect 81122 -20908 81156 -20642
rect 81318 -20908 81352 -20642
rect 80682 -20952 81400 -20908
rect 76123 -21007 81400 -20952
rect 76123 -21111 81036 -21007
rect 81703 -21088 81737 -20671
rect 81899 -21088 81933 -20671
rect 82095 -21038 82129 -20671
rect 82312 -21038 82346 -20872
rect 82508 -21038 82542 -20872
rect 82704 -21038 82738 -20872
rect 82900 -21038 82934 -20872
rect 82095 -21088 82982 -21038
rect 74776 -21181 81036 -21111
rect 81693 -21137 82982 -21088
rect 81693 -21151 82135 -21137
rect 74409 -21197 81036 -21181
rect 81692 -21180 82135 -21151
rect 81692 -21197 82310 -21180
rect 74409 -21234 82805 -21197
rect 74409 -21298 74814 -21234
rect 73846 -21308 73944 -21305
rect 74409 -21308 74526 -21298
rect 73846 -21425 74526 -21308
rect 74776 -21393 74814 -21298
rect 73846 -21431 73944 -21425
rect 74779 -21886 74813 -21393
rect 74973 -21391 75011 -21234
rect 74975 -21886 75009 -21391
rect 75565 -21414 75615 -21234
rect 75691 -21411 75741 -21234
rect 75570 -21886 75604 -21414
rect 75700 -21886 75734 -21411
rect 75922 -21396 75965 -21234
rect 76119 -21294 82805 -21234
rect 75928 -21686 75962 -21396
rect 76119 -21394 76162 -21294
rect 76124 -21686 76158 -21394
rect 73853 -23423 74255 -23357
rect 71358 -24399 71392 -24133
rect 71554 -24399 71588 -24133
rect 71750 -24399 71784 -24133
rect 71946 -24399 71980 -24133
rect 71310 -24498 72028 -24399
rect 71492 -24688 71664 -24498
rect 72331 -24579 72365 -24162
rect 72527 -24579 72561 -24162
rect 72723 -24529 72757 -24162
rect 72940 -24529 72974 -24363
rect 73136 -24529 73170 -24363
rect 73332 -24529 73366 -24363
rect 73528 -24529 73562 -24363
rect 72723 -24579 73610 -24529
rect 72321 -24628 73610 -24579
rect 72321 -24642 72763 -24628
rect 72320 -24671 72763 -24642
rect 72320 -24688 72938 -24671
rect 71322 -24799 73433 -24688
rect 71322 -24841 73537 -24799
rect 71724 -24848 71950 -24841
rect 71761 -24855 71950 -24848
rect 72768 -24865 73537 -24841
rect 71322 -24904 71764 -24889
rect 71322 -24953 72611 -24904
rect 71332 -25370 71366 -24953
rect 71528 -25370 71562 -24953
rect 71724 -25003 72611 -24953
rect 72774 -24991 72819 -24865
rect 71724 -25370 71758 -25003
rect 71941 -25169 71975 -25003
rect 72137 -25169 72171 -25003
rect 72333 -25169 72367 -25003
rect 72529 -25169 72563 -25003
rect 71247 -25419 71382 -25413
rect 71227 -25421 71382 -25419
rect 70699 -25457 71382 -25421
rect 70882 -26484 71018 -25457
rect 71227 -25459 71382 -25457
rect 71247 -25467 71382 -25459
rect 72779 -25581 72813 -24991
rect 72969 -24988 73014 -24865
rect 72975 -25581 73009 -24988
rect 73391 -24989 73436 -24865
rect 73398 -25581 73432 -24989
rect 73853 -24724 73919 -23423
rect 73836 -24837 73920 -24724
rect 74189 -24753 74255 -23423
rect 77086 -23630 77208 -21294
rect 80694 -21308 82805 -21294
rect 80694 -21315 82909 -21308
rect 82982 -21315 83044 -21287
rect 80694 -21350 83044 -21315
rect 81096 -21357 81322 -21350
rect 81133 -21364 81322 -21357
rect 82140 -21367 83044 -21350
rect 82140 -21374 82909 -21367
rect 80694 -21413 81136 -21398
rect 80694 -21462 81983 -21413
rect 80704 -21879 80738 -21462
rect 80900 -21879 80934 -21462
rect 81096 -21512 81983 -21462
rect 82146 -21500 82191 -21374
rect 81096 -21879 81130 -21512
rect 81313 -21678 81347 -21512
rect 81509 -21678 81543 -21512
rect 81705 -21678 81739 -21512
rect 81901 -21678 81935 -21512
rect 77086 -23752 77718 -23630
rect 75026 -24430 75060 -24164
rect 75222 -24430 75256 -24164
rect 75418 -24430 75452 -24164
rect 75614 -24430 75648 -24164
rect 74978 -24529 75696 -24430
rect 75160 -24719 75332 -24529
rect 75999 -24610 76033 -24193
rect 76195 -24610 76229 -24193
rect 76391 -24560 76425 -24193
rect 76608 -24560 76642 -24394
rect 76804 -24560 76838 -24394
rect 77000 -24560 77034 -24394
rect 77196 -24560 77230 -24394
rect 76391 -24610 77278 -24560
rect 75989 -24659 77278 -24610
rect 75989 -24673 76431 -24659
rect 75988 -24702 76431 -24673
rect 75988 -24719 76606 -24702
rect 74990 -24753 77101 -24719
rect 74189 -24819 77101 -24753
rect 77256 -24794 77335 -24763
rect 74990 -24830 77101 -24819
rect 77156 -24830 77335 -24794
rect 74990 -24872 77335 -24830
rect 75392 -24879 75618 -24872
rect 75429 -24886 75618 -24879
rect 76436 -24877 77335 -24872
rect 76436 -24896 77205 -24877
rect 74990 -24935 75432 -24920
rect 74990 -24984 76279 -24935
rect 75000 -25401 75034 -24984
rect 75196 -25401 75230 -24984
rect 75392 -25034 76279 -24984
rect 76442 -25022 76487 -24896
rect 75392 -25401 75426 -25034
rect 75609 -25200 75643 -25034
rect 75805 -25200 75839 -25034
rect 76001 -25200 76035 -25034
rect 76197 -25200 76231 -25034
rect 74915 -25450 75050 -25444
rect 74895 -25452 75050 -25450
rect 74481 -25488 75050 -25452
rect 74481 -26484 74617 -25488
rect 74895 -25490 75050 -25488
rect 74915 -25498 75050 -25490
rect 76447 -25612 76481 -25022
rect 76637 -25019 76682 -24896
rect 76643 -25612 76677 -25019
rect 77059 -25020 77104 -24896
rect 77256 -24902 77335 -24877
rect 77066 -25612 77100 -25020
rect 77596 -24748 77718 -23752
rect 77506 -24887 77718 -24748
rect 77506 -24915 77645 -24887
rect 70882 -26620 74617 -26484
rect -33001 -29022 61865 -28886
rect -33001 -29027 -22941 -29022
rect 70882 -29185 71018 -26620
rect 82151 -22090 82185 -21500
rect 82341 -21497 82386 -21374
rect 82347 -22090 82381 -21497
rect 82763 -21498 82808 -21374
rect 82982 -21381 83044 -21367
rect 82770 -22090 82804 -21498
rect 85898 -21073 86373 -17161
rect 90329 -18041 91702 -17504
rect 88428 -18579 91702 -18041
rect 90329 -18877 91702 -18579
rect 84140 -21143 86572 -21073
rect 83773 -21195 86572 -21143
rect 83773 -21196 85526 -21195
rect 83773 -21260 84178 -21196
rect 83210 -21270 83308 -21267
rect 83773 -21270 83890 -21260
rect 83210 -21387 83890 -21270
rect 84140 -21355 84178 -21260
rect 83210 -21393 83308 -21387
rect 84143 -21848 84177 -21355
rect 84337 -21353 84375 -21196
rect 84339 -21848 84373 -21353
rect 84929 -21376 84979 -21196
rect 85055 -21373 85105 -21196
rect 84934 -21848 84968 -21376
rect 85064 -21848 85098 -21373
rect 85286 -21358 85329 -21196
rect 85292 -21648 85326 -21358
rect 85483 -21356 85526 -21196
rect 85488 -21648 85522 -21356
rect 83217 -23385 83619 -23319
rect 80722 -24361 80756 -24095
rect 80918 -24361 80952 -24095
rect 81114 -24361 81148 -24095
rect 81310 -24361 81344 -24095
rect 80674 -24460 81392 -24361
rect 80856 -24650 81028 -24460
rect 81695 -24541 81729 -24124
rect 81891 -24541 81925 -24124
rect 82087 -24491 82121 -24124
rect 82304 -24491 82338 -24325
rect 82500 -24491 82534 -24325
rect 82696 -24491 82730 -24325
rect 82892 -24491 82926 -24325
rect 82087 -24541 82974 -24491
rect 81685 -24590 82974 -24541
rect 81685 -24604 82127 -24590
rect 81684 -24633 82127 -24604
rect 81684 -24650 82302 -24633
rect 80686 -24761 82797 -24650
rect 80686 -24803 82901 -24761
rect 81088 -24810 81314 -24803
rect 81125 -24817 81314 -24810
rect 82132 -24827 82901 -24803
rect 80686 -24866 81128 -24851
rect 80686 -24915 81975 -24866
rect 80696 -25332 80730 -24915
rect 80892 -25332 80926 -24915
rect 81088 -24965 81975 -24915
rect 82138 -24953 82183 -24827
rect 81088 -25332 81122 -24965
rect 81305 -25131 81339 -24965
rect 81501 -25131 81535 -24965
rect 81697 -25131 81731 -24965
rect 81893 -25131 81927 -24965
rect 80611 -25381 80746 -25375
rect 80591 -25383 80746 -25381
rect 80063 -25419 80746 -25383
rect 80246 -26446 80382 -25419
rect 80591 -25421 80746 -25419
rect 80611 -25429 80746 -25421
rect 82143 -25543 82177 -24953
rect 82333 -24950 82378 -24827
rect 82339 -25543 82373 -24950
rect 82755 -24951 82800 -24827
rect 82762 -25543 82796 -24951
rect 83217 -24686 83283 -23385
rect 83200 -24799 83284 -24686
rect 83553 -24715 83619 -23385
rect 86450 -23592 86572 -21195
rect 86450 -23714 87082 -23592
rect 84390 -24392 84424 -24126
rect 84586 -24392 84620 -24126
rect 84782 -24392 84816 -24126
rect 84978 -24392 85012 -24126
rect 84342 -24491 85060 -24392
rect 84524 -24681 84696 -24491
rect 85363 -24572 85397 -24155
rect 85559 -24572 85593 -24155
rect 85755 -24522 85789 -24155
rect 85972 -24522 86006 -24356
rect 86168 -24522 86202 -24356
rect 86364 -24522 86398 -24356
rect 86560 -24522 86594 -24356
rect 85755 -24572 86642 -24522
rect 85353 -24621 86642 -24572
rect 85353 -24635 85795 -24621
rect 85352 -24664 85795 -24635
rect 85352 -24681 85970 -24664
rect 84354 -24715 86465 -24681
rect 83553 -24781 86465 -24715
rect 86620 -24756 86699 -24725
rect 84354 -24792 86465 -24781
rect 86520 -24792 86699 -24756
rect 84354 -24834 86699 -24792
rect 84756 -24841 84982 -24834
rect 84793 -24848 84982 -24841
rect 85800 -24839 86699 -24834
rect 85800 -24858 86569 -24839
rect 84354 -24897 84796 -24882
rect 84354 -24946 85643 -24897
rect 84364 -25363 84398 -24946
rect 84560 -25363 84594 -24946
rect 84756 -24996 85643 -24946
rect 85806 -24984 85851 -24858
rect 84756 -25363 84790 -24996
rect 84973 -25162 85007 -24996
rect 85169 -25162 85203 -24996
rect 85365 -25162 85399 -24996
rect 85561 -25162 85595 -24996
rect 84279 -25412 84414 -25406
rect 84259 -25414 84414 -25412
rect 83845 -25450 84414 -25414
rect 83845 -26446 83981 -25450
rect 84259 -25452 84414 -25450
rect 84279 -25460 84414 -25452
rect 85811 -25574 85845 -24984
rect 86001 -24981 86046 -24858
rect 86007 -25574 86041 -24981
rect 86423 -24982 86468 -24858
rect 86620 -24864 86699 -24839
rect 86430 -25574 86464 -24982
rect 86960 -24710 87082 -23714
rect 86870 -24849 87082 -24710
rect 86870 -24877 87009 -24849
rect 80246 -26582 83981 -26446
rect -32755 -29321 71018 -29185
rect 80270 -29555 80406 -26582
rect 95829 -28339 98798 -15816
rect -32917 -29691 80406 -29555
rect 83333 -31308 98798 -28339
rect 83333 -32649 86302 -31308
rect 25923 -32870 87071 -32649
rect -32225 -33190 -26140 -32972
rect -26347 -33893 -26140 -33190
rect 6895 -33632 87071 -32870
rect -26196 -34019 -26162 -33893
rect -26196 -34053 -25608 -34019
rect -25569 -34137 -25521 -33971
rect -26016 -34171 -25521 -34137
rect -26016 -34289 -25608 -34255
rect -25569 -34373 -25521 -34171
rect -26016 -34407 -25521 -34373
rect -26016 -34525 -25608 -34491
rect -25569 -34609 -25521 -34407
rect -26016 -34643 -25521 -34609
rect -26016 -34761 -25608 -34727
rect -25569 -34845 -25521 -34643
rect -26016 -34879 -25521 -34845
rect -26016 -34997 -25608 -34963
rect -25569 -35069 -25521 -34879
rect -25449 -35069 -25383 -34081
rect 6895 -34786 7657 -33632
rect 25923 -33752 87071 -33632
rect -7334 -34797 8126 -34786
rect -9665 -34833 8126 -34797
rect -25569 -35081 -25383 -35069
rect -26016 -35115 -25383 -35081
rect -25569 -35128 -25383 -35115
rect -26016 -35233 -25608 -35199
rect -25569 -35317 -25521 -35128
rect -26016 -35351 -25521 -35317
rect -26016 -35469 -25608 -35435
rect -25569 -35546 -25521 -35351
rect -25449 -35460 -25383 -35128
rect -14690 -34886 8126 -34833
rect -14690 -34896 -9465 -34886
rect -14690 -34901 -13117 -34896
rect -12219 -34901 -10417 -34896
rect -14690 -35460 -14601 -34901
rect -14441 -35192 -14407 -34901
rect -14245 -35192 -14211 -34901
rect -14049 -35192 -14015 -34901
rect -13604 -35192 -13570 -34901
rect -25449 -35546 -14601 -35460
rect -25569 -35553 -14601 -35546
rect -26016 -35587 -14601 -35553
rect -25569 -35605 -14601 -35587
rect -26016 -35705 -25608 -35671
rect -25569 -35777 -25521 -35605
rect -25449 -35673 -14601 -35605
rect -25449 -35683 -21418 -35673
rect -25449 -35732 -23381 -35683
rect -25449 -35777 -25383 -35732
rect -25569 -35789 -25383 -35777
rect -26016 -35823 -25383 -35789
rect -25569 -35836 -25383 -35823
rect -26016 -35941 -25608 -35907
rect -25569 -36013 -25521 -35836
rect -25449 -36013 -25383 -35836
rect -25569 -36025 -25383 -36013
rect -26016 -36059 -25383 -36025
rect -25569 -36072 -25383 -36059
rect -26016 -36177 -25608 -36143
rect -25569 -36251 -25521 -36072
rect -25449 -36251 -25383 -36072
rect -25569 -36260 -25383 -36251
rect -23653 -36260 -23381 -35732
rect -23186 -36191 -23125 -35988
rect -22995 -36109 -22934 -35909
rect -22886 -36026 -22825 -35823
rect -22040 -35979 -22006 -35683
rect -21844 -35979 -21810 -35683
rect -21648 -35979 -21614 -35683
rect -21452 -35979 -21418 -35683
rect -20915 -35687 -20670 -35673
rect -20910 -35979 -20876 -35687
rect -22117 -36026 -21982 -36018
rect -22886 -36061 -21982 -36026
rect -22136 -36063 -21982 -36061
rect -22117 -36072 -21982 -36063
rect -21781 -36109 -21646 -36100
rect -22995 -36147 -21646 -36109
rect -21781 -36154 -21646 -36147
rect -21593 -36191 -21458 -36178
rect -23186 -36225 -21458 -36191
rect -23186 -36226 -23125 -36225
rect -21593 -36232 -21458 -36225
rect -25569 -36261 -23381 -36260
rect -26016 -36295 -23381 -36261
rect -25569 -36310 -23381 -36295
rect -26016 -36413 -25608 -36379
rect -25569 -36491 -25521 -36310
rect -25449 -36491 -23381 -36310
rect -25569 -36497 -23381 -36491
rect -26016 -36531 -23381 -36497
rect -25569 -36532 -23381 -36531
rect -25569 -36550 -25383 -36532
rect -26016 -36649 -25608 -36615
rect -25569 -36721 -25521 -36550
rect -25449 -36721 -25383 -36550
rect -25569 -36733 -25383 -36721
rect -26016 -36767 -25383 -36733
rect -25569 -36780 -25383 -36767
rect -26016 -36885 -25608 -36851
rect -25569 -36958 -25521 -36780
rect -25449 -36958 -25383 -36780
rect -25569 -36969 -25383 -36958
rect -26016 -37003 -25383 -36969
rect -25569 -37017 -25383 -37003
rect -26016 -37121 -25608 -37087
rect -25569 -37192 -25521 -37017
rect -25449 -37192 -25383 -37017
rect -25569 -37205 -25383 -37192
rect -26016 -37239 -25383 -37205
rect -25569 -37251 -25383 -37239
rect -26016 -37357 -25608 -37323
rect -25569 -37426 -25521 -37251
rect -25449 -37321 -25383 -37251
rect -23653 -37321 -23381 -36532
rect -20714 -35979 -20680 -35687
rect -20093 -35735 -18766 -35673
rect -20093 -35790 -18762 -35735
rect -20041 -36201 -20007 -35790
rect -19845 -36201 -19811 -35790
rect -19649 -35834 -18762 -35790
rect -19649 -36201 -19615 -35834
rect -19432 -36000 -19398 -35834
rect -19236 -36000 -19202 -35834
rect -19040 -36000 -19006 -35834
rect -18844 -36000 -18810 -35834
rect -20261 -36346 -20124 -36342
rect -20299 -36348 -20072 -36346
rect -19661 -36348 -19587 -36322
rect -20299 -36386 -19587 -36348
rect -20261 -36400 -20124 -36386
rect -20073 -36387 -19587 -36386
rect -20073 -36388 -20002 -36387
rect -19661 -36393 -19587 -36387
rect -18490 -36766 -18355 -36758
rect -18510 -36768 -18355 -36766
rect -18901 -36804 -18355 -36768
rect -22787 -37065 -22727 -36989
rect -22787 -37105 -22719 -37065
rect -25449 -37424 -23381 -37321
rect -23334 -37320 -23233 -37147
rect -22787 -37182 -22727 -37105
rect -20370 -37182 -20238 -37173
rect -22787 -37222 -20238 -37182
rect -22787 -37226 -22727 -37222
rect -20370 -37226 -20238 -37222
rect -18824 -37320 -18767 -36804
rect -18510 -36806 -18355 -36804
rect -18490 -36812 -18355 -36806
rect -18405 -37272 -18371 -36855
rect -18209 -37272 -18175 -36855
rect -18013 -37222 -17979 -36855
rect -17796 -37222 -17762 -37056
rect -17600 -37222 -17566 -37056
rect -17404 -37222 -17370 -37056
rect -17208 -37222 -17174 -37056
rect -18013 -37272 -17126 -37222
rect -16958 -37234 -16924 -36644
rect -23334 -37383 -18767 -37320
rect -18415 -37321 -17126 -37272
rect -18415 -37336 -17973 -37321
rect -16963 -37360 -16918 -37234
rect -16762 -37237 -16728 -36644
rect -16768 -37360 -16723 -37237
rect -16339 -37236 -16305 -36644
rect -16346 -37360 -16301 -37236
rect -17976 -37377 -17787 -37370
rect -23334 -37390 -23233 -37383
rect -18013 -37384 -17787 -37377
rect -16969 -37384 -16200 -37360
rect -18415 -37424 -16200 -37384
rect -25449 -37426 -16200 -37424
rect -25569 -37441 -16304 -37426
rect -26016 -37475 -16304 -37441
rect -25569 -37485 -16304 -37475
rect -26016 -37593 -25608 -37559
rect -25569 -37677 -25521 -37485
rect -26016 -37711 -25521 -37677
rect -26824 -37809 -26416 -37775
rect -26824 -38045 -26416 -38011
rect -26016 -37829 -25608 -37795
rect -25569 -37925 -25521 -37711
rect -26016 -37959 -25521 -37925
rect -25569 -38151 -25521 -37959
rect -25449 -37537 -16304 -37485
rect -25449 -37593 -18840 -37537
rect -25449 -38151 -25383 -37593
rect -23653 -37623 -18840 -37593
rect -23653 -37656 -18850 -37623
rect -21993 -37693 -20704 -37656
rect -25569 -38161 -25383 -38151
rect -26016 -38195 -25383 -38161
rect -25569 -38210 -25383 -38195
rect -21983 -38110 -21949 -37693
rect -21787 -38110 -21753 -37693
rect -21591 -37743 -20704 -37693
rect -21591 -38110 -21557 -37743
rect -21374 -37909 -21340 -37743
rect -21178 -37909 -21144 -37743
rect -20982 -37909 -20948 -37743
rect -20786 -37909 -20752 -37743
rect -20210 -37915 -20176 -37656
rect -20014 -37915 -19980 -37656
rect -19818 -37915 -19784 -37656
rect -19622 -37915 -19588 -37656
rect -19080 -37915 -19046 -37656
rect -26824 -38281 -26416 -38247
rect -25569 -38382 -25521 -38210
rect -25449 -38382 -25383 -38210
rect -25569 -38397 -25383 -38382
rect -26016 -38431 -25383 -38397
rect -25569 -38441 -25383 -38431
rect -26824 -38517 -26416 -38483
rect -25569 -38618 -25521 -38441
rect -25449 -38618 -25383 -38441
rect -25569 -38633 -25383 -38618
rect -26016 -38667 -25383 -38633
rect -25569 -38677 -25383 -38667
rect -26824 -38753 -26416 -38719
rect -25569 -38853 -25521 -38677
rect -25449 -38853 -25383 -38677
rect -18884 -37915 -18850 -37656
rect -18245 -37727 -18073 -37537
rect -17417 -37554 -16799 -37537
rect -17417 -37583 -16974 -37554
rect -17416 -37597 -16974 -37583
rect -17416 -37646 -16127 -37597
rect -18427 -37826 -17709 -37727
rect -18379 -38092 -18345 -37826
rect -18183 -38092 -18149 -37826
rect -17987 -38092 -17953 -37826
rect -17791 -38092 -17757 -37826
rect -17406 -38063 -17372 -37646
rect -17210 -38063 -17176 -37646
rect -17014 -37696 -16127 -37646
rect -17014 -38063 -16980 -37696
rect -16797 -37862 -16763 -37696
rect -16601 -37862 -16567 -37696
rect -16405 -37862 -16371 -37696
rect -16209 -37862 -16175 -37696
rect -25569 -38869 -25383 -38853
rect -26016 -38903 -25383 -38869
rect -25569 -38912 -25383 -38903
rect -26824 -38989 -26416 -38955
rect -25569 -39092 -25521 -38912
rect -25449 -39092 -25383 -38912
rect -25569 -39105 -25383 -39092
rect -26016 -39139 -25383 -39105
rect -25569 -39151 -25383 -39139
rect -26824 -39225 -26416 -39191
rect -25569 -39321 -25521 -39151
rect -25449 -39321 -25383 -39151
rect -25569 -39341 -25383 -39321
rect -26016 -39375 -25383 -39341
rect -25569 -39380 -25383 -39375
rect -26824 -39461 -26416 -39427
rect -25569 -39577 -25521 -39380
rect -26016 -39611 -25521 -39577
rect -25569 -39813 -25521 -39611
rect -26016 -39847 -25521 -39813
rect -25569 -39927 -25521 -39847
rect -25449 -39927 -25383 -39380
rect -25569 -39943 -25383 -39927
rect -26016 -39977 -25383 -39943
rect -25569 -39986 -25383 -39977
rect -25569 -40159 -25521 -39986
rect -25449 -40159 -25383 -39986
rect -25569 -40179 -25383 -40159
rect -26016 -40213 -25383 -40179
rect -25569 -40218 -25383 -40213
rect -25569 -40400 -25521 -40218
rect -25449 -40400 -25383 -40218
rect -25569 -40415 -25383 -40400
rect -26016 -40449 -25383 -40415
rect -25569 -40459 -25383 -40449
rect -25569 -40651 -25521 -40459
rect -26016 -40671 -25521 -40651
rect -25449 -40671 -25383 -40459
rect -26016 -40685 -25383 -40671
rect -25569 -40730 -25383 -40685
rect -25569 -40887 -25521 -40730
rect -26016 -40921 -25521 -40887
rect -25569 -41017 -25521 -40921
rect -26016 -41051 -25521 -41017
rect -25569 -41253 -25521 -41051
rect -26016 -41259 -25521 -41253
rect -25449 -41259 -25383 -40730
rect -26016 -41287 -25383 -41259
rect -25569 -41318 -25383 -41287
rect -25569 -41489 -25521 -41318
rect -26016 -41523 -25521 -41489
rect -25449 -41519 -25383 -41318
rect -14690 -36596 -14601 -35673
rect -13408 -35192 -13374 -34901
rect -13212 -35192 -13178 -34901
rect -11741 -35192 -11707 -34901
rect -11545 -35192 -11511 -34901
rect -11349 -35192 -11315 -34901
rect -10904 -35192 -10870 -34901
rect -10708 -35192 -10674 -34901
rect -10512 -35192 -10478 -34901
rect -8083 -35010 -8038 -34886
rect -8079 -35602 -8045 -35010
rect -7661 -35009 -7616 -34886
rect -7656 -35602 -7622 -35009
rect -7466 -35012 -7421 -34886
rect -7336 -34979 8126 -34886
rect -7460 -35602 -7426 -35012
rect -14343 -36593 -14309 -36302
rect -14147 -36593 -14113 -36302
rect -13951 -36593 -13917 -36302
rect -12600 -36593 -12566 -36302
rect -12404 -36593 -12370 -36302
rect -12208 -36593 -12174 -36302
rect -11643 -36593 -11609 -36302
rect -11447 -36593 -11413 -36302
rect -11251 -36593 -11217 -36302
rect -9900 -36593 -9866 -36302
rect -9704 -36593 -9670 -36302
rect -9508 -36593 -9474 -36302
rect -9018 -36593 -8984 -36302
rect -8822 -36593 -8788 -36302
rect -8626 -36593 -8592 -36302
rect -14403 -36596 -13908 -36593
rect -12661 -36594 -11208 -36593
rect -14690 -36598 -13586 -36596
rect -12661 -36598 -10895 -36594
rect -9961 -36598 -8583 -36593
rect -14690 -36661 -8583 -36598
rect -14690 -36664 -13586 -36661
rect -11368 -36662 -10895 -36661
rect -14228 -38360 -14075 -36664
rect -13448 -37645 -13377 -37644
rect -13036 -37645 -12962 -37639
rect -13448 -37646 -12962 -37645
rect -13674 -37684 -12962 -37646
rect -13674 -37686 -13447 -37684
rect -13036 -37710 -12962 -37684
rect -13416 -38248 -13382 -37831
rect -13220 -38248 -13186 -37831
rect -13024 -38198 -12990 -37831
rect -12807 -38198 -12773 -38032
rect -12611 -38198 -12577 -38032
rect -12415 -38198 -12381 -38032
rect -12219 -38198 -12185 -38032
rect -13024 -38248 -12137 -38198
rect -11969 -38210 -11935 -37620
rect -13426 -38297 -12137 -38248
rect -13426 -38312 -12984 -38297
rect -11974 -38336 -11929 -38210
rect -11773 -38213 -11739 -37620
rect -11779 -38336 -11734 -38213
rect -11350 -38212 -11316 -37620
rect -11357 -38336 -11312 -38212
rect -12987 -38353 -12798 -38346
rect -13024 -38360 -12798 -38353
rect -11980 -38360 -11211 -38336
rect -14228 -38402 -11211 -38360
rect -14228 -38513 -11315 -38402
rect -14228 -39760 -14075 -38513
rect -13256 -38703 -13084 -38513
rect -12428 -38530 -11810 -38513
rect -12428 -38559 -11985 -38530
rect -12427 -38573 -11985 -38559
rect -12427 -38622 -11138 -38573
rect -13438 -38802 -12720 -38703
rect -13390 -39068 -13356 -38802
rect -13194 -39068 -13160 -38802
rect -12998 -39068 -12964 -38802
rect -12802 -39068 -12768 -38802
rect -12417 -39039 -12383 -38622
rect -12221 -39039 -12187 -38622
rect -12025 -38672 -11138 -38622
rect -12025 -39039 -11991 -38672
rect -11808 -38838 -11774 -38672
rect -11612 -38838 -11578 -38672
rect -11416 -38838 -11382 -38672
rect -11220 -38838 -11186 -38672
rect -5971 -35086 -4919 -34979
rect -5971 -35215 -5931 -35086
rect -5971 -35398 -5937 -35215
rect -5782 -35215 -5736 -35086
rect -5775 -35398 -5741 -35215
rect -5584 -35211 -5538 -35086
rect -5579 -35398 -5545 -35211
rect -5471 -35215 -5425 -35086
rect -5465 -35398 -5431 -35215
rect -5275 -35210 -5229 -35086
rect -5269 -35398 -5235 -35210
rect -5162 -35220 -5116 -35086
rect -5156 -35398 -5122 -35220
rect -4965 -35208 -4919 -35086
rect -4960 -35398 -4926 -35208
rect -4644 -35816 -4529 -34979
rect -3157 -35017 -2564 -34979
rect -4649 -35952 -4526 -35816
rect -3471 -35086 -2419 -35017
rect -3471 -35215 -3431 -35086
rect -3471 -35398 -3437 -35215
rect -3282 -35215 -3236 -35086
rect -3275 -35398 -3241 -35215
rect -3084 -35211 -3038 -35086
rect -3079 -35398 -3045 -35211
rect -2971 -35215 -2925 -35086
rect -2965 -35398 -2931 -35215
rect -2775 -35210 -2729 -35086
rect -2769 -35398 -2735 -35210
rect -2662 -35220 -2616 -35086
rect -2656 -35398 -2622 -35220
rect -2465 -35208 -2419 -35086
rect -2460 -35398 -2426 -35208
rect -2076 -35851 -1962 -34979
rect -641 -35017 -48 -34979
rect -971 -35086 81 -35017
rect -971 -35215 -931 -35086
rect -971 -35398 -937 -35215
rect -782 -35215 -736 -35086
rect -775 -35398 -741 -35215
rect -584 -35211 -538 -35086
rect -579 -35398 -545 -35211
rect -471 -35215 -425 -35086
rect -465 -35398 -431 -35215
rect -275 -35210 -229 -35086
rect -2082 -35987 -1959 -35851
rect -269 -35398 -235 -35210
rect -162 -35220 -116 -35086
rect -156 -35398 -122 -35220
rect 35 -35208 81 -35086
rect 40 -35398 74 -35208
rect 406 -35851 521 -34979
rect 1893 -35017 2486 -34979
rect 4306 -35017 4899 -34979
rect 1529 -35086 2581 -35017
rect 1529 -35215 1569 -35086
rect 1529 -35398 1563 -35215
rect 1718 -35215 1764 -35086
rect 1725 -35398 1759 -35215
rect 1916 -35211 1962 -35086
rect 1921 -35398 1955 -35211
rect 2029 -35215 2075 -35086
rect 2035 -35398 2069 -35215
rect 2225 -35210 2271 -35086
rect 401 -35987 524 -35851
rect 2231 -35398 2265 -35210
rect 2338 -35220 2384 -35086
rect 2344 -35398 2378 -35220
rect 2535 -35208 2581 -35086
rect 2540 -35398 2574 -35208
rect 4029 -35086 5081 -35017
rect 4029 -35215 4069 -35086
rect 4029 -35398 4063 -35215
rect 4218 -35215 4264 -35086
rect 4225 -35398 4259 -35215
rect 4416 -35211 4462 -35086
rect 4421 -35398 4455 -35211
rect 4529 -35215 4575 -35086
rect 4535 -35398 4569 -35215
rect 4725 -35210 4771 -35086
rect 3634 -35706 3773 -35652
rect 4731 -35398 4765 -35210
rect 4838 -35220 4884 -35086
rect 4844 -35398 4878 -35220
rect 5035 -35208 5081 -35086
rect 5040 -35398 5074 -35208
rect 4712 -35712 4851 -35658
rect 7029 -35086 8081 -34979
rect 7029 -35215 7069 -35086
rect 7029 -35398 7063 -35215
rect 7218 -35215 7264 -35086
rect 7225 -35398 7259 -35215
rect 7416 -35211 7462 -35086
rect 7421 -35398 7455 -35211
rect 7529 -35215 7575 -35086
rect 7535 -35398 7569 -35215
rect 7725 -35210 7771 -35086
rect 6634 -35706 6773 -35652
rect 7731 -35398 7765 -35210
rect 7838 -35220 7884 -35086
rect 7844 -35398 7878 -35220
rect 8035 -35208 8081 -35086
rect 8040 -35398 8074 -35208
rect 7712 -35712 7851 -35658
rect -6442 -36455 -6254 -36381
rect 400 -36405 523 -36404
rect -6310 -36810 -6276 -36519
rect -6114 -36810 -6080 -36519
rect -5918 -36810 -5884 -36519
rect -4650 -36719 -4527 -36583
rect -2083 -36575 -1960 -36439
rect 400 -36467 706 -36405
rect -6319 -36878 -5824 -36810
rect -6303 -37268 -6215 -36878
rect -6120 -37268 -6032 -36878
rect -5938 -37268 -5850 -36878
rect -6816 -37271 -5712 -37268
rect -4645 -37271 -4530 -36719
rect -3494 -37271 -3021 -37270
rect -2079 -37271 -1964 -36575
rect -665 -37145 -528 -37094
rect -824 -37271 -701 -37249
rect -6816 -37334 -701 -37271
rect -6816 -37336 -5712 -37334
rect -13584 -39115 -13454 -39098
rect -13410 -39115 -13337 -39102
rect -13584 -39156 -13337 -39115
rect -6816 -39031 -6727 -37336
rect -6529 -37339 -6034 -37336
rect -4787 -37338 -3021 -37334
rect -4787 -37339 -3334 -37338
rect -2087 -37339 -701 -37334
rect -6469 -37630 -6435 -37339
rect -6273 -37630 -6239 -37339
rect -6077 -37630 -6043 -37339
rect -4726 -37630 -4692 -37339
rect -4530 -37630 -4496 -37339
rect -4334 -37630 -4300 -37339
rect -3769 -37630 -3735 -37339
rect -3573 -37630 -3539 -37339
rect -3377 -37630 -3343 -37339
rect -2026 -37630 -1992 -37339
rect -1830 -37630 -1796 -37339
rect -1634 -37630 -1600 -37339
rect -1144 -37630 -1110 -37339
rect -948 -37630 -914 -37339
rect -824 -37385 -701 -37339
rect -752 -37630 -718 -37385
rect -2259 -37953 -2185 -37794
rect -5950 -38076 -5818 -38063
rect -2259 -38076 -2184 -37953
rect -1656 -37705 -1488 -37694
rect -1656 -37763 -1453 -37705
rect -665 -37694 -626 -37145
rect -530 -37275 -407 -37248
rect 405 -37275 520 -36467
rect 2448 -37275 2571 -37261
rect -530 -37354 2571 -37275
rect -530 -37355 -175 -37354
rect -530 -37384 -376 -37355
rect -410 -37647 -376 -37384
rect -1656 -37768 -1488 -37763
rect -774 -37768 -606 -37694
rect -665 -38076 -626 -37768
rect -214 -37647 -180 -37355
rect 328 -37647 362 -37354
rect 524 -37647 558 -37354
rect 720 -37647 754 -37354
rect 916 -37647 950 -37354
rect 1275 -37394 2162 -37354
rect 1323 -37560 1357 -37394
rect 1519 -37560 1553 -37394
rect 1715 -37560 1749 -37394
rect 1911 -37560 1945 -37394
rect -6356 -38115 -626 -38076
rect -5950 -38123 -5818 -38115
rect -5914 -38602 -5854 -38458
rect -5914 -38664 -5674 -38602
rect -5877 -38665 -5674 -38664
rect -5842 -38676 -5674 -38665
rect -6567 -39031 -6533 -38740
rect -6371 -39031 -6337 -38740
rect -6175 -39031 -6141 -38740
rect -5730 -39031 -5696 -38740
rect -5534 -39031 -5500 -38740
rect -5338 -39031 -5304 -38740
rect -3867 -39031 -3833 -38740
rect -3671 -39031 -3637 -38740
rect -3475 -39031 -3441 -38740
rect -3030 -39031 -2996 -38740
rect -2834 -39031 -2800 -38740
rect -2638 -39031 -2604 -38740
rect 2128 -37761 2162 -37394
rect 2324 -37761 2358 -37354
rect 2448 -37397 2571 -37354
rect 2520 -37761 2554 -37397
rect 2837 -37297 2960 -37260
rect 4065 -37282 4188 -37237
rect 3727 -37297 4188 -37282
rect 2837 -37346 4188 -37297
rect 2837 -37396 3767 -37346
rect 2928 -37562 2962 -37396
rect 3124 -37562 3158 -37396
rect 3320 -37562 3354 -37396
rect 3516 -37562 3550 -37396
rect 3733 -37763 3767 -37396
rect 3929 -37763 3963 -37346
rect 4065 -37373 4188 -37346
rect 4125 -37763 4159 -37373
rect 4466 -37268 4589 -37235
rect 4466 -37273 5362 -37268
rect 5822 -37273 5945 -37240
rect 4466 -37341 5945 -37273
rect 4466 -37346 4787 -37341
rect 5290 -37342 5945 -37341
rect 4466 -37371 4589 -37346
rect 4552 -37638 4586 -37371
rect 4748 -37638 4782 -37346
rect 5290 -37638 5324 -37342
rect 5486 -37638 5520 -37342
rect 5682 -37638 5716 -37342
rect 5822 -37376 5945 -37342
rect 5878 -37638 5912 -37376
rect 7038 -37268 7161 -37241
rect 7038 -37337 8091 -37268
rect 7038 -37377 7161 -37337
rect 7039 -37466 7079 -37377
rect 7039 -37649 7073 -37466
rect 7228 -37466 7274 -37337
rect 7235 -37649 7269 -37466
rect 7426 -37462 7472 -37337
rect 7431 -37649 7465 -37462
rect 7539 -37466 7585 -37337
rect 7545 -37649 7579 -37466
rect 7735 -37461 7781 -37337
rect 6644 -37957 6783 -37903
rect 7741 -37649 7775 -37461
rect 7848 -37471 7894 -37337
rect 7854 -37649 7888 -37471
rect 8045 -37459 8091 -37337
rect 8050 -37649 8084 -37459
rect 7722 -37963 7861 -37909
rect 15965 -36705 16200 -36682
rect 10557 -36950 16200 -36705
rect 10557 -36952 16076 -36950
rect 25923 -35141 27026 -33752
rect 17736 -36885 17954 -36639
rect 17775 -37742 17917 -36885
rect 25977 -36745 26307 -36662
rect 25977 -36924 27156 -36745
rect 25977 -36956 26307 -36924
rect 28544 -37278 28679 -37270
rect 28524 -37280 28679 -37278
rect 28317 -37316 28679 -37280
rect 28524 -37318 28679 -37316
rect 28544 -37324 28679 -37318
rect 20271 -37603 25496 -37540
rect 21223 -37608 23025 -37603
rect 23923 -37608 25496 -37603
rect 27656 -37604 27690 -37338
rect 27852 -37604 27886 -37338
rect 28048 -37604 28082 -37338
rect 28244 -37604 28278 -37338
rect 17738 -37931 17917 -37742
rect -6816 -39036 -5243 -39031
rect -4345 -39036 -2543 -39031
rect -6816 -39099 -1591 -39036
rect -13584 -39248 -13454 -39156
rect -13410 -39162 -13337 -39156
rect -6816 -39738 -6727 -39099
rect -10612 -39760 -6727 -39738
rect -14690 -39823 -6727 -39760
rect -14690 -39828 -13117 -39823
rect -12219 -39828 -10417 -39823
rect -14690 -40453 -14601 -39828
rect -14441 -40119 -14407 -39828
rect -14245 -40119 -14211 -39828
rect -14049 -40119 -14015 -39828
rect -13604 -40119 -13570 -39828
rect -13408 -40119 -13374 -39828
rect -13212 -40119 -13178 -39828
rect -22237 -40620 -14600 -40453
rect -21867 -40759 -21085 -40620
rect -20709 -40746 -20191 -40620
rect -21927 -40892 -21059 -40759
rect -20724 -40815 -20170 -40746
rect -19820 -40747 -19267 -40620
rect -19820 -40788 -19265 -40747
rect -21927 -41004 -21874 -40892
rect -23186 -41711 -23126 -41530
rect -21918 -41604 -21884 -41004
rect -21731 -41020 -21678 -40892
rect -20719 -40942 -20671 -40815
rect -21722 -41604 -21688 -41020
rect -20712 -41333 -20678 -40942
rect -20522 -40948 -20474 -40815
rect -19819 -40816 -19265 -40788
rect -20892 -41449 -20834 -41354
rect -20516 -41333 -20482 -40948
rect -19814 -40943 -19766 -40816
rect -20485 -41449 -20342 -41442
rect -20892 -41485 -20342 -41449
rect -20892 -41491 -20834 -41485
rect -20485 -41502 -20342 -41485
rect -19807 -41334 -19773 -40943
rect -19617 -40949 -19569 -40816
rect -19611 -41334 -19577 -40949
rect -23186 -41752 -21297 -41711
rect -23186 -41767 -23126 -41752
rect -21357 -41757 -21297 -41752
rect -22995 -41800 -22935 -41787
rect -21677 -41800 -21532 -41789
rect -22995 -41841 -21532 -41800
rect -21357 -41813 -21212 -41757
rect -22995 -42024 -22935 -41841
rect -21677 -41845 -21532 -41841
rect -22885 -41892 -22825 -41890
rect -22006 -41892 -21861 -41884
rect -22885 -41933 -21861 -41892
rect -22885 -42127 -22825 -41933
rect -22006 -41940 -21861 -41933
rect -18405 -42272 -18371 -41855
rect -18209 -42272 -18175 -41855
rect -18013 -42222 -17979 -41855
rect -17796 -42222 -17762 -42056
rect -17600 -42222 -17566 -42056
rect -17404 -42222 -17370 -42056
rect -17208 -42222 -17174 -42056
rect -18013 -42272 -17126 -42222
rect -16958 -42234 -16924 -41644
rect -18415 -42321 -17126 -42272
rect -18415 -42336 -17973 -42321
rect -16963 -42360 -16918 -42234
rect -16762 -42237 -16728 -41644
rect -16768 -42360 -16723 -42237
rect -16339 -42236 -16305 -41644
rect -14690 -41523 -14601 -40620
rect -11741 -40119 -11707 -39828
rect -11545 -40119 -11511 -39828
rect -11349 -40119 -11315 -39828
rect -10904 -40119 -10870 -39828
rect -10708 -40119 -10674 -39828
rect -10512 -40119 -10478 -39828
rect -8056 -39944 -8011 -39823
rect -8052 -40536 -8018 -39944
rect -7634 -39943 -7589 -39823
rect -7629 -40536 -7595 -39943
rect -7439 -39946 -7394 -39823
rect -6816 -39938 -6727 -39823
rect -7433 -40536 -7399 -39946
rect -6816 -40027 -6726 -39938
rect -6528 -40027 -6259 -39099
rect -5982 -40027 -5713 -39099
rect -5105 -40027 -4836 -39099
rect -4243 -40027 -3974 -39099
rect -3340 -40027 -3071 -39099
rect -2309 -40027 -2040 -39099
rect 18077 -39089 18111 -38489
rect 18068 -39201 18121 -39089
rect 18273 -39073 18307 -38489
rect 18264 -39201 18317 -39073
rect 18068 -39334 18936 -39201
rect -6816 -40090 -1591 -40027
rect -6816 -40095 -5243 -40090
rect -4345 -40095 -2543 -40090
rect -14343 -41520 -14309 -41229
rect -14147 -41520 -14113 -41229
rect -13951 -41520 -13917 -41229
rect -12600 -41520 -12566 -41229
rect -12404 -41520 -12370 -41229
rect -12208 -41520 -12174 -41229
rect -11643 -41520 -11609 -41229
rect -11447 -41520 -11413 -41229
rect -11251 -41520 -11217 -41229
rect -9900 -41520 -9866 -41229
rect -9704 -41520 -9670 -41229
rect -9508 -41520 -9474 -41229
rect -9018 -41520 -8984 -41229
rect -8822 -41520 -8788 -41229
rect -8626 -41520 -8592 -41229
rect -14403 -41523 -13908 -41520
rect -12661 -41521 -11208 -41520
rect -14690 -41525 -13586 -41523
rect -12661 -41525 -10895 -41521
rect -9961 -41525 -8583 -41520
rect -14690 -41588 -8583 -41525
rect -16346 -42360 -16301 -42236
rect -17976 -42377 -17787 -42370
rect -22787 -42496 -22729 -42400
rect -18013 -42384 -17787 -42377
rect -16969 -42384 -16200 -42360
rect -20912 -42496 -20854 -42400
rect -19649 -42426 -16200 -42384
rect -22787 -42537 -20854 -42496
rect -19649 -42537 -16304 -42426
rect -19649 -42556 -18073 -42537
rect -22255 -44106 -22221 -43814
rect -19649 -43551 -19477 -42556
rect -18245 -42727 -18073 -42556
rect -17417 -42554 -16799 -42537
rect -17417 -42583 -16974 -42554
rect -17416 -42597 -16974 -42583
rect -17416 -42646 -16127 -42597
rect -18427 -42826 -17709 -42727
rect -18379 -43092 -18345 -42826
rect -18183 -43092 -18149 -42826
rect -17987 -43092 -17953 -42826
rect -17791 -43092 -17757 -42826
rect -17406 -43063 -17372 -42646
rect -17210 -43063 -17176 -42646
rect -17014 -42696 -16127 -42646
rect -17014 -43063 -16980 -42696
rect -16797 -42862 -16763 -42696
rect -16601 -42862 -16567 -42696
rect -16405 -42862 -16371 -42696
rect -16209 -42862 -16175 -42696
rect -14690 -41591 -13586 -41588
rect -11368 -41589 -10895 -41588
rect -6816 -41790 -6727 -40095
rect -6567 -40386 -6533 -40095
rect -6371 -40386 -6337 -40095
rect -6175 -40386 -6141 -40095
rect -5730 -40386 -5696 -40095
rect -5534 -40386 -5500 -40095
rect -5338 -40386 -5304 -40095
rect -3867 -40386 -3833 -40095
rect -3671 -40386 -3637 -40095
rect -3475 -40386 -3441 -40095
rect -3030 -40386 -2996 -40095
rect -2834 -40386 -2800 -40095
rect -2638 -40386 -2604 -40095
rect -3142 -40461 -2974 -40450
rect -3202 -40524 -2974 -40461
rect -3202 -40683 -3142 -40524
rect -4177 -40925 -4040 -40914
rect -3231 -40925 -3099 -40915
rect -6356 -40964 -626 -40925
rect -4177 -40974 -4040 -40964
rect -3231 -40975 -3099 -40964
rect -6469 -41787 -6435 -41496
rect -6273 -41787 -6239 -41496
rect -6077 -41787 -6043 -41496
rect -4356 -41363 -4188 -41358
rect -4128 -41363 -4068 -41290
rect -4356 -41421 -4068 -41363
rect -4356 -41432 -4188 -41421
rect -4128 -41422 -4068 -41421
rect -4726 -41787 -4692 -41496
rect -4530 -41787 -4496 -41496
rect -4334 -41787 -4300 -41496
rect -3769 -41787 -3735 -41496
rect -3573 -41787 -3539 -41496
rect -3377 -41787 -3343 -41496
rect -665 -41358 -626 -40964
rect -774 -41432 -606 -41358
rect -2026 -41787 -1992 -41496
rect -1830 -41787 -1796 -41496
rect -1634 -41787 -1600 -41496
rect -1144 -41787 -1110 -41496
rect -948 -41787 -914 -41496
rect -752 -41741 -718 -41496
rect -824 -41787 -701 -41741
rect -6529 -41790 -6034 -41787
rect -4787 -41788 -3334 -41787
rect -6816 -41792 -5712 -41790
rect -4787 -41792 -3021 -41788
rect -2087 -41792 -701 -41787
rect -6816 -41855 -701 -41792
rect -6816 -41858 -5712 -41855
rect -19651 -43638 -19475 -43551
rect -4645 -42407 -4530 -41855
rect -3494 -41856 -3021 -41855
rect -4650 -42543 -4527 -42407
rect -2079 -42551 -1964 -41855
rect -824 -41877 -701 -41855
rect -665 -41981 -626 -41432
rect -410 -41742 -376 -41479
rect -530 -41771 -376 -41742
rect -214 -41771 -180 -41479
rect -530 -41772 -175 -41771
rect 328 -41772 362 -41479
rect 524 -41772 558 -41479
rect 720 -41772 754 -41479
rect 916 -41772 950 -41479
rect 1323 -41732 1357 -41566
rect 1519 -41732 1553 -41566
rect 1715 -41732 1749 -41566
rect 1911 -41732 1945 -41566
rect 2128 -41732 2162 -41365
rect 1275 -41772 2162 -41732
rect 2324 -41772 2358 -41365
rect 2520 -41729 2554 -41365
rect 2448 -41772 2571 -41729
rect -530 -41851 2571 -41772
rect -530 -41878 -407 -41851
rect -665 -42032 -528 -41981
rect -2083 -42687 -1960 -42551
rect 405 -42659 520 -41851
rect 2448 -41865 2571 -41851
rect 2928 -41730 2962 -41564
rect 3124 -41730 3158 -41564
rect 3320 -41730 3354 -41564
rect 3516 -41730 3550 -41564
rect 3733 -41730 3767 -41363
rect 2837 -41780 3767 -41730
rect 3929 -41780 3963 -41363
rect 4125 -41753 4159 -41363
rect 4065 -41780 4188 -41753
rect 2837 -41829 4188 -41780
rect 2837 -41866 2960 -41829
rect 3727 -41844 4188 -41829
rect 4065 -41889 4188 -41844
rect 400 -42721 706 -42659
rect 400 -42722 523 -42721
rect 4552 -41755 4586 -41488
rect 19306 -38103 19438 -37968
rect 19306 -38438 19412 -38103
rect 21284 -37899 21318 -37608
rect 21480 -37899 21514 -37608
rect 21676 -37899 21710 -37608
rect 22121 -37899 22155 -37608
rect 22317 -37899 22351 -37608
rect 22513 -37899 22547 -37608
rect 21654 -37974 21822 -37963
rect 21654 -38037 21882 -37974
rect 21822 -38196 21882 -38037
rect 23984 -37899 24018 -37608
rect 24180 -37899 24214 -37608
rect 24376 -37899 24410 -37608
rect 24821 -37899 24855 -37608
rect 25017 -37899 25051 -37608
rect 25213 -37899 25247 -37608
rect 25407 -37668 25496 -37608
rect 27608 -37668 28326 -37604
rect 25407 -37703 28326 -37668
rect 25407 -37893 27962 -37703
rect 28629 -37784 28663 -37367
rect 28825 -37784 28859 -37367
rect 29021 -37734 29055 -37367
rect 29238 -37734 29272 -37568
rect 29434 -37734 29468 -37568
rect 29630 -37734 29664 -37568
rect 29826 -37734 29860 -37568
rect 29021 -37784 29908 -37734
rect 28619 -37833 29908 -37784
rect 28619 -37847 29061 -37833
rect 28618 -37876 29061 -37847
rect 28618 -37893 29236 -37876
rect 25407 -37962 29731 -37893
rect 21779 -38438 21911 -38428
rect 22720 -38438 22857 -38427
rect 19306 -38477 25036 -38438
rect 19306 -38871 19345 -38477
rect 21779 -38488 21911 -38477
rect 22720 -38487 22857 -38477
rect 19286 -38945 19454 -38871
rect 19398 -39300 19432 -39009
rect 19594 -39300 19628 -39009
rect 19790 -39300 19824 -39009
rect 20280 -39300 20314 -39009
rect 20476 -39300 20510 -39009
rect 20672 -39300 20706 -39009
rect 22748 -38876 22808 -38803
rect 22868 -38876 23036 -38871
rect 22748 -38934 23036 -38876
rect 22748 -38935 22808 -38934
rect 22023 -39300 22057 -39009
rect 22219 -39300 22253 -39009
rect 22415 -39300 22449 -39009
rect 22868 -38945 23036 -38934
rect 22980 -39300 23014 -39009
rect 23176 -39300 23210 -39009
rect 23372 -39300 23406 -39009
rect 24723 -39300 24757 -39009
rect 24919 -39300 24953 -39009
rect 25115 -39300 25149 -39009
rect 19389 -39305 20767 -39300
rect 22014 -39301 23467 -39300
rect 21701 -39305 23467 -39301
rect 24714 -39303 25209 -39300
rect 25407 -39303 25496 -37962
rect 27620 -38004 29731 -37962
rect 27620 -38011 29835 -38004
rect 29908 -38011 29970 -37983
rect 27620 -38046 29970 -38011
rect 28022 -38053 28248 -38046
rect 28059 -38060 28248 -38053
rect 29066 -38063 29970 -38046
rect 29066 -38070 29835 -38063
rect 27620 -38109 28062 -38094
rect 27620 -38158 28909 -38109
rect 26896 -38515 27155 -38472
rect 26030 -38626 27155 -38515
rect 27630 -38575 27664 -38158
rect 27826 -38575 27860 -38158
rect 28022 -38208 28909 -38158
rect 29072 -38196 29117 -38070
rect 28022 -38575 28056 -38208
rect 28239 -38374 28273 -38208
rect 28435 -38374 28469 -38208
rect 28631 -38374 28665 -38208
rect 28827 -38374 28861 -38208
rect 27545 -38624 27680 -38618
rect 27525 -38626 27680 -38624
rect 26030 -38662 27680 -38626
rect 26030 -38720 27155 -38662
rect 27525 -38664 27680 -38662
rect 27545 -38672 27680 -38664
rect 26896 -38735 27155 -38720
rect 24392 -39305 25496 -39303
rect 19389 -39368 25496 -39305
rect 21701 -39369 22174 -39368
rect 21891 -39588 22123 -39369
rect 24392 -39371 25496 -39368
rect 21833 -39652 22275 -39588
rect 21843 -40169 21877 -39652
rect 22039 -40169 22073 -39652
rect 22235 -40169 22269 -39652
rect 6644 -41223 6783 -41169
rect 4466 -41780 4589 -41755
rect 4748 -41780 4782 -41488
rect 4466 -41785 4787 -41780
rect 5290 -41784 5324 -41488
rect 5486 -41784 5520 -41488
rect 5682 -41784 5716 -41488
rect 5878 -41750 5912 -41488
rect 5822 -41784 5945 -41750
rect 5290 -41785 5945 -41784
rect 4466 -41853 5945 -41785
rect 4466 -41858 5362 -41853
rect 4466 -41891 4589 -41858
rect 5822 -41886 5945 -41853
rect 7039 -41660 7073 -41477
rect 7039 -41749 7079 -41660
rect 7235 -41660 7269 -41477
rect 7038 -41789 7161 -41749
rect 7228 -41789 7274 -41660
rect 7431 -41664 7465 -41477
rect 7545 -41660 7579 -41477
rect 7722 -41217 7861 -41163
rect 7426 -41789 7472 -41664
rect 7539 -41789 7585 -41660
rect 7741 -41665 7775 -41477
rect 7854 -41655 7888 -41477
rect 7735 -41789 7781 -41665
rect 7848 -41789 7894 -41655
rect 8050 -41667 8084 -41477
rect 8045 -41789 8091 -41667
rect 7038 -41858 8091 -41789
rect 7038 -41885 7161 -41858
rect 8833 -41228 8978 -41093
rect 8550 -42243 8673 -42242
rect -6366 -43474 -6227 -43420
rect -22059 -44090 -22025 -43814
rect -21517 -44090 -21483 -43814
rect -21321 -44090 -21287 -43814
rect -21125 -44090 -21091 -43814
rect -20929 -44090 -20895 -43814
rect -5971 -43911 -5937 -43728
rect -5971 -44040 -5931 -43911
rect -5775 -43911 -5741 -43728
rect -5782 -44040 -5736 -43911
rect -5579 -43915 -5545 -43728
rect -5465 -43911 -5431 -43728
rect -5288 -43468 -5149 -43414
rect -4649 -43310 -4526 -43174
rect -5584 -44040 -5538 -43915
rect -5471 -44040 -5425 -43911
rect -5269 -43916 -5235 -43728
rect -5156 -43906 -5122 -43728
rect -5275 -44040 -5229 -43916
rect -5162 -44040 -5116 -43906
rect -4960 -43918 -4926 -43728
rect -4965 -44040 -4919 -43918
rect -22077 -44106 -19475 -44090
rect -22265 -44173 -19475 -44106
rect -22077 -44182 -19475 -44173
rect -5971 -44147 -4919 -44040
rect -4644 -44147 -4529 -43310
rect -3471 -43911 -3437 -43728
rect -3471 -44040 -3431 -43911
rect -3275 -43911 -3241 -43728
rect -3282 -44040 -3236 -43911
rect -3079 -43915 -3045 -43728
rect -2965 -43911 -2931 -43728
rect -2082 -43275 -1959 -43139
rect -3084 -44040 -3038 -43915
rect -2971 -44040 -2925 -43911
rect -2769 -43916 -2735 -43728
rect -2656 -43906 -2622 -43728
rect -2775 -44040 -2729 -43916
rect -2662 -44040 -2616 -43906
rect -2460 -43918 -2426 -43728
rect -2465 -44040 -2419 -43918
rect -3471 -44109 -2419 -44040
rect -3157 -44147 -2564 -44109
rect -2076 -44147 -1962 -43275
rect -971 -43911 -937 -43728
rect -971 -44040 -931 -43911
rect -775 -43911 -741 -43728
rect -782 -44040 -736 -43911
rect -579 -43915 -545 -43728
rect -465 -43911 -431 -43728
rect 401 -43275 524 -43139
rect -584 -44040 -538 -43915
rect -471 -44040 -425 -43911
rect -269 -43916 -235 -43728
rect -156 -43906 -122 -43728
rect -275 -44040 -229 -43916
rect -162 -44040 -116 -43906
rect 40 -43918 74 -43728
rect 35 -44040 81 -43918
rect -971 -44109 81 -44040
rect -641 -44147 -48 -44109
rect 406 -44147 521 -43275
rect 1529 -43911 1563 -43728
rect 1529 -44040 1569 -43911
rect 1725 -43911 1759 -43728
rect 1718 -44040 1764 -43911
rect 1921 -43915 1955 -43728
rect 2035 -43911 2069 -43728
rect 1916 -44040 1962 -43915
rect 2029 -44040 2075 -43911
rect 2231 -43916 2265 -43728
rect 2344 -43906 2378 -43728
rect 3634 -43474 3773 -43420
rect 2225 -44040 2271 -43916
rect 2338 -44040 2384 -43906
rect 2540 -43918 2574 -43728
rect 2535 -44040 2581 -43918
rect 1529 -44109 2581 -44040
rect 4029 -43911 4063 -43728
rect 4029 -44040 4069 -43911
rect 4225 -43911 4259 -43728
rect 4218 -44040 4264 -43911
rect 4421 -43915 4455 -43728
rect 4535 -43911 4569 -43728
rect 4712 -43468 4851 -43414
rect 8549 -42286 8673 -42243
rect 4416 -44040 4462 -43915
rect 4529 -44040 4575 -43911
rect 4731 -43916 4765 -43728
rect 4844 -43906 4878 -43728
rect 8549 -43094 8607 -42286
rect 8693 -42844 8816 -42800
rect 6634 -43474 6773 -43420
rect 4725 -44040 4771 -43916
rect 4838 -44040 4884 -43906
rect 5040 -43918 5074 -43728
rect 5035 -44040 5081 -43918
rect 4029 -44109 5081 -44040
rect 7029 -43911 7063 -43728
rect 7029 -44040 7069 -43911
rect 7225 -43911 7259 -43728
rect 7218 -44040 7264 -43911
rect 7421 -43915 7455 -43728
rect 7535 -43911 7569 -43728
rect 7712 -43468 7851 -43414
rect 7416 -44040 7462 -43915
rect 7529 -44040 7575 -43911
rect 7731 -43916 7765 -43728
rect 7844 -43906 7878 -43728
rect 7725 -44040 7771 -43916
rect 7838 -44040 7884 -43906
rect 8040 -43918 8074 -43728
rect 8035 -44040 8081 -43918
rect 1893 -44147 2486 -44109
rect 4306 -44147 4899 -44109
rect 7029 -44147 8081 -44040
rect -6836 -44340 8126 -44147
rect 8550 -44504 8606 -43094
rect 8649 -43472 8714 -43335
rect 8652 -44232 8706 -43472
rect 8757 -44232 8811 -42844
rect 8856 -44449 8912 -41228
rect 18072 -41426 18106 -41035
rect 18065 -41553 18113 -41426
rect 18268 -41420 18302 -41035
rect 18262 -41553 18310 -41420
rect 19018 -41426 19052 -41035
rect 19011 -41553 19059 -41426
rect 19214 -41420 19248 -41035
rect 19208 -41553 19256 -41420
rect 19689 -41553 19775 -41545
rect 17242 -41565 19775 -41553
rect 19934 -41565 19968 -41269
rect 20130 -41565 20164 -41269
rect 20326 -41565 20360 -41269
rect 20522 -41565 20556 -41269
rect 20809 -41561 20872 -41547
rect 21064 -41561 21098 -41269
rect 21260 -41561 21294 -41269
rect 21490 -41553 21564 -41547
rect 21793 -41553 21827 -41262
rect 21989 -41553 22023 -41262
rect 22185 -41526 22219 -41262
rect 22673 -41526 22707 -40691
rect 22869 -41526 22903 -40691
rect 23073 -41526 23107 -40691
rect 23269 -41526 23303 -40691
rect 23673 -41526 23707 -40691
rect 23869 -41526 23903 -40691
rect 24073 -41526 24107 -40691
rect 24269 -41526 24303 -40691
rect 24673 -41526 24707 -40691
rect 24869 -41526 24903 -40691
rect 25073 -41526 25107 -40691
rect 25269 -41526 25303 -40691
rect 25407 -41526 25496 -39371
rect 29077 -38786 29111 -38196
rect 29267 -38193 29312 -38070
rect 29273 -38786 29307 -38193
rect 29689 -38194 29734 -38070
rect 29908 -38077 29970 -38063
rect 29696 -38786 29730 -38194
rect 36096 -37615 36130 -37349
rect 36292 -37615 36326 -37349
rect 36488 -37615 36522 -37349
rect 36684 -37615 36718 -37349
rect 36048 -37714 36766 -37615
rect 31066 -37839 33498 -37769
rect 30699 -37891 33498 -37839
rect 30699 -37892 32452 -37891
rect 30699 -37956 31104 -37892
rect 30136 -37966 30234 -37963
rect 30699 -37966 30816 -37956
rect 30136 -38083 30816 -37966
rect 31066 -38051 31104 -37956
rect 30136 -38089 30234 -38083
rect 31069 -38544 31103 -38051
rect 31263 -38049 31301 -37892
rect 31265 -38544 31299 -38049
rect 31855 -38072 31905 -37892
rect 31981 -38069 32031 -37892
rect 31860 -38544 31894 -38072
rect 31990 -38544 32024 -38069
rect 32212 -38054 32255 -37892
rect 32218 -38344 32252 -38054
rect 32409 -38052 32452 -37892
rect 33376 -37904 33498 -37891
rect 36230 -37904 36402 -37714
rect 37069 -37795 37103 -37378
rect 37265 -37795 37299 -37378
rect 37461 -37745 37495 -37378
rect 37678 -37745 37712 -37579
rect 37874 -37745 37908 -37579
rect 38070 -37745 38104 -37579
rect 38266 -37745 38300 -37579
rect 37461 -37795 38348 -37745
rect 37059 -37844 38348 -37795
rect 37059 -37858 37501 -37844
rect 37058 -37887 37501 -37858
rect 37058 -37904 37676 -37887
rect 33376 -38015 38171 -37904
rect 33376 -38022 38275 -38015
rect 38348 -38022 38410 -37994
rect 32414 -38344 32448 -38052
rect 33376 -38057 38410 -38022
rect 22185 -41553 25496 -41526
rect 21490 -41561 25496 -41553
rect 20809 -41565 25496 -41561
rect 17242 -41621 25496 -41565
rect 17242 -41622 21564 -41621
rect 9127 -42109 9318 -42103
rect 9127 -42192 9690 -42109
rect 9127 -42210 9318 -42192
rect 9607 -44057 9690 -42192
rect 17242 -42093 17368 -41622
rect 19689 -41628 21564 -41622
rect 19689 -41634 20872 -41628
rect 21490 -41634 21564 -41628
rect 22207 -41629 25496 -41621
rect 19689 -41638 19775 -41634
rect 20809 -41645 20872 -41634
rect 13573 -42096 14046 -42095
rect 16264 -42096 17368 -42093
rect 11261 -42159 17368 -42096
rect 11261 -42164 12639 -42159
rect 13573 -42163 15339 -42159
rect 16264 -42161 17368 -42159
rect 13886 -42164 15339 -42163
rect 16586 -42164 17081 -42161
rect 11270 -42455 11304 -42164
rect 11466 -42455 11500 -42164
rect 11662 -42455 11696 -42164
rect 12152 -42455 12186 -42164
rect 12348 -42455 12382 -42164
rect 12544 -42455 12578 -42164
rect 11158 -42593 11326 -42519
rect 10557 -42987 10852 -42889
rect 11178 -42987 11217 -42593
rect 13895 -42455 13929 -42164
rect 14091 -42455 14125 -42164
rect 14287 -42455 14321 -42164
rect 14852 -42455 14886 -42164
rect 15048 -42455 15082 -42164
rect 15244 -42455 15278 -42164
rect 14620 -42530 14680 -42529
rect 14740 -42530 14908 -42519
rect 14620 -42588 14908 -42530
rect 14620 -42661 14680 -42588
rect 14740 -42593 14908 -42588
rect 16595 -42455 16629 -42164
rect 16791 -42455 16825 -42164
rect 16987 -42455 17021 -42164
rect 13651 -42987 13783 -42976
rect 14592 -42987 14729 -42977
rect 10557 -43026 16908 -42987
rect 10557 -43092 10852 -43026
rect 13651 -43036 13783 -43026
rect 14592 -43037 14729 -43026
rect 13694 -43427 13754 -43268
rect 13526 -43490 13754 -43427
rect 13526 -43501 13694 -43490
rect 13156 -43856 13190 -43565
rect 13352 -43856 13386 -43565
rect 13548 -43856 13582 -43565
rect 13993 -43856 14027 -43565
rect 14189 -43856 14223 -43565
rect 14385 -43856 14419 -43565
rect 15856 -43856 15890 -43565
rect 16052 -43856 16086 -43565
rect 16248 -43856 16282 -43565
rect 16693 -43856 16727 -43565
rect 16889 -43856 16923 -43565
rect 17085 -43856 17119 -43565
rect 17279 -43856 17368 -42161
rect 30143 -40081 30545 -40015
rect 27648 -41057 27682 -40791
rect 27844 -41057 27878 -40791
rect 28040 -41057 28074 -40791
rect 28236 -41057 28270 -40791
rect 27600 -41156 28318 -41057
rect 27782 -41346 27954 -41156
rect 28621 -41237 28655 -40820
rect 28817 -41237 28851 -40820
rect 29013 -41187 29047 -40820
rect 29230 -41187 29264 -41021
rect 29426 -41187 29460 -41021
rect 29622 -41187 29656 -41021
rect 29818 -41187 29852 -41021
rect 29013 -41237 29900 -41187
rect 28611 -41286 29900 -41237
rect 28611 -41300 29053 -41286
rect 28610 -41329 29053 -41300
rect 28610 -41346 29228 -41329
rect 27612 -41457 29723 -41346
rect 27612 -41499 29827 -41457
rect 28014 -41506 28240 -41499
rect 28051 -41513 28240 -41506
rect 29058 -41523 29827 -41499
rect 27612 -41562 28054 -41547
rect 27612 -41611 28901 -41562
rect 27622 -42028 27656 -41611
rect 27818 -42028 27852 -41611
rect 28014 -41661 28901 -41611
rect 29064 -41649 29109 -41523
rect 28014 -42028 28048 -41661
rect 28231 -41827 28265 -41661
rect 28427 -41827 28461 -41661
rect 28623 -41827 28657 -41661
rect 28819 -41827 28853 -41661
rect 27537 -42077 27672 -42071
rect 27517 -42079 27672 -42077
rect 26989 -42115 27672 -42079
rect 13095 -43861 14897 -43856
rect 15795 -43861 17368 -43856
rect 12143 -43924 17368 -43861
rect 27172 -43142 27308 -42115
rect 27517 -42117 27672 -42115
rect 27537 -42125 27672 -42117
rect 29069 -42239 29103 -41649
rect 29259 -41646 29304 -41523
rect 29265 -42239 29299 -41646
rect 29681 -41647 29726 -41523
rect 29688 -42239 29722 -41647
rect 30143 -41382 30209 -40081
rect 30126 -41495 30210 -41382
rect 30479 -41411 30545 -40081
rect 33376 -40288 33498 -38057
rect 36462 -38064 36688 -38057
rect 36499 -38071 36688 -38064
rect 37506 -38074 38410 -38057
rect 37506 -38081 38275 -38074
rect 36060 -38120 36502 -38105
rect 36060 -38169 37349 -38120
rect 34897 -38637 35545 -38583
rect 36070 -38586 36104 -38169
rect 36266 -38586 36300 -38169
rect 36462 -38219 37349 -38169
rect 37512 -38207 37557 -38081
rect 36462 -38586 36496 -38219
rect 36679 -38385 36713 -38219
rect 36875 -38385 36909 -38219
rect 37071 -38385 37105 -38219
rect 37267 -38385 37301 -38219
rect 35985 -38635 36120 -38629
rect 35965 -38637 36120 -38635
rect 34897 -38673 36120 -38637
rect 34897 -38729 35545 -38673
rect 35965 -38675 36120 -38673
rect 35985 -38683 36120 -38675
rect 33376 -40410 34008 -40288
rect 31316 -41088 31350 -40822
rect 31512 -41088 31546 -40822
rect 31708 -41088 31742 -40822
rect 31904 -41088 31938 -40822
rect 31268 -41187 31986 -41088
rect 31450 -41377 31622 -41187
rect 32289 -41268 32323 -40851
rect 32485 -41268 32519 -40851
rect 32681 -41218 32715 -40851
rect 32898 -41218 32932 -41052
rect 33094 -41218 33128 -41052
rect 33290 -41218 33324 -41052
rect 33486 -41218 33520 -41052
rect 32681 -41268 33568 -41218
rect 32279 -41317 33568 -41268
rect 32279 -41331 32721 -41317
rect 32278 -41360 32721 -41331
rect 32278 -41377 32896 -41360
rect 31280 -41411 33391 -41377
rect 30479 -41477 33391 -41411
rect 33546 -41452 33625 -41421
rect 31280 -41488 33391 -41477
rect 33446 -41488 33625 -41452
rect 31280 -41530 33625 -41488
rect 31682 -41537 31908 -41530
rect 31719 -41544 31908 -41537
rect 32726 -41535 33625 -41530
rect 32726 -41554 33495 -41535
rect 31280 -41593 31722 -41578
rect 31280 -41642 32569 -41593
rect 31290 -42059 31324 -41642
rect 31486 -42059 31520 -41642
rect 31682 -41692 32569 -41642
rect 32732 -41680 32777 -41554
rect 31682 -42059 31716 -41692
rect 31899 -41858 31933 -41692
rect 32095 -41858 32129 -41692
rect 32291 -41858 32325 -41692
rect 32487 -41858 32521 -41692
rect 31205 -42108 31340 -42102
rect 31185 -42110 31340 -42108
rect 30771 -42146 31340 -42110
rect 30771 -43142 30907 -42146
rect 31185 -42148 31340 -42146
rect 31205 -42156 31340 -42148
rect 32737 -42270 32771 -41680
rect 32927 -41677 32972 -41554
rect 32933 -42270 32967 -41677
rect 33349 -41678 33394 -41554
rect 33546 -41560 33625 -41535
rect 33356 -42270 33390 -41678
rect 33886 -41406 34008 -40410
rect 33796 -41545 34008 -41406
rect 33796 -41573 33935 -41545
rect 27172 -43278 30907 -43142
rect 9583 -44236 9711 -44057
rect 26602 -44292 26823 -44097
rect 27172 -44504 27308 -43278
rect 34897 -44112 35043 -38729
rect 37517 -38797 37551 -38207
rect 37707 -38204 37752 -38081
rect 37713 -38797 37747 -38204
rect 38129 -38205 38174 -38081
rect 38348 -38088 38410 -38074
rect 38136 -38797 38170 -38205
rect 44959 -37654 44993 -37388
rect 45155 -37654 45189 -37388
rect 45351 -37654 45385 -37388
rect 45547 -37654 45581 -37388
rect 44911 -37738 45629 -37654
rect 40878 -37753 45629 -37738
rect 40878 -37780 45265 -37753
rect 39506 -37850 45265 -37780
rect 45932 -37834 45966 -37417
rect 46128 -37834 46162 -37417
rect 46324 -37784 46358 -37417
rect 46541 -37784 46575 -37618
rect 46737 -37784 46771 -37618
rect 46933 -37784 46967 -37618
rect 47129 -37784 47163 -37618
rect 46324 -37834 47211 -37784
rect 39139 -37903 45265 -37850
rect 45922 -37883 47211 -37834
rect 45922 -37897 46364 -37883
rect 39139 -37967 39544 -37903
rect 38576 -37977 38674 -37974
rect 39139 -37977 39256 -37967
rect 38576 -38094 39256 -37977
rect 39506 -38062 39544 -37967
rect 38576 -38100 38674 -38094
rect 39509 -38555 39543 -38062
rect 39703 -38060 39741 -37903
rect 39705 -38555 39739 -38060
rect 40295 -38083 40345 -37903
rect 40421 -38080 40471 -37903
rect 40300 -38555 40334 -38083
rect 40430 -38555 40464 -38080
rect 40652 -38065 40695 -37903
rect 40849 -37943 45265 -37903
rect 45921 -37926 46364 -37897
rect 45921 -37943 46539 -37926
rect 40849 -37992 47034 -37943
rect 40658 -38355 40692 -38065
rect 40849 -38063 40892 -37992
rect 40854 -38355 40888 -38063
rect 38583 -40092 38985 -40026
rect 36088 -41068 36122 -40802
rect 36284 -41068 36318 -40802
rect 36480 -41068 36514 -40802
rect 36676 -41068 36710 -40802
rect 36040 -41167 36758 -41068
rect 36222 -41357 36394 -41167
rect 37061 -41248 37095 -40831
rect 37257 -41248 37291 -40831
rect 37453 -41198 37487 -40831
rect 37670 -41198 37704 -41032
rect 37866 -41198 37900 -41032
rect 38062 -41198 38096 -41032
rect 38258 -41198 38292 -41032
rect 37453 -41248 38340 -41198
rect 37051 -41297 38340 -41248
rect 37051 -41311 37493 -41297
rect 37050 -41340 37493 -41311
rect 37050 -41357 37668 -41340
rect 36052 -41468 38163 -41357
rect 36052 -41510 38267 -41468
rect 36454 -41517 36680 -41510
rect 36491 -41524 36680 -41517
rect 37498 -41534 38267 -41510
rect 36052 -41573 36494 -41558
rect 36052 -41622 37341 -41573
rect 36062 -42039 36096 -41622
rect 36258 -42039 36292 -41622
rect 36454 -41672 37341 -41622
rect 37504 -41660 37549 -41534
rect 36454 -42039 36488 -41672
rect 36671 -41838 36705 -41672
rect 36867 -41838 36901 -41672
rect 37063 -41838 37097 -41672
rect 37259 -41838 37293 -41672
rect 35977 -42088 36112 -42082
rect 35957 -42090 36112 -42088
rect 35429 -42126 36112 -42090
rect 35612 -43153 35748 -42126
rect 35957 -42128 36112 -42126
rect 35977 -42136 36112 -42128
rect 37509 -42250 37543 -41660
rect 37699 -41657 37744 -41534
rect 37705 -42250 37739 -41657
rect 38121 -41658 38166 -41534
rect 38128 -42250 38162 -41658
rect 38583 -41393 38649 -40092
rect 38566 -41506 38650 -41393
rect 38919 -41422 38985 -40092
rect 41816 -40299 41938 -37992
rect 44923 -38054 47034 -37992
rect 44923 -38061 47138 -38054
rect 47211 -38061 47273 -38033
rect 44923 -38096 47273 -38061
rect 45325 -38103 45551 -38096
rect 45362 -38110 45551 -38103
rect 46369 -38113 47273 -38096
rect 46369 -38120 47138 -38113
rect 44923 -38159 45365 -38144
rect 44923 -38208 46212 -38159
rect 44933 -38625 44967 -38208
rect 45129 -38625 45163 -38208
rect 45325 -38258 46212 -38208
rect 46375 -38246 46420 -38120
rect 45325 -38625 45359 -38258
rect 45542 -38424 45576 -38258
rect 45738 -38424 45772 -38258
rect 45934 -38424 45968 -38258
rect 46130 -38424 46164 -38258
rect 43579 -38676 44346 -38669
rect 44848 -38674 44983 -38668
rect 44828 -38676 44983 -38674
rect 43579 -38712 44983 -38676
rect 43579 -38815 44346 -38712
rect 44828 -38714 44983 -38712
rect 44848 -38722 44983 -38714
rect 41816 -40421 42448 -40299
rect 39756 -41099 39790 -40833
rect 39952 -41099 39986 -40833
rect 40148 -41099 40182 -40833
rect 40344 -41099 40378 -40833
rect 39708 -41198 40426 -41099
rect 39890 -41388 40062 -41198
rect 40729 -41279 40763 -40862
rect 40925 -41279 40959 -40862
rect 41121 -41229 41155 -40862
rect 41338 -41229 41372 -41063
rect 41534 -41229 41568 -41063
rect 41730 -41229 41764 -41063
rect 41926 -41229 41960 -41063
rect 41121 -41279 42008 -41229
rect 40719 -41328 42008 -41279
rect 40719 -41342 41161 -41328
rect 40718 -41371 41161 -41342
rect 40718 -41388 41336 -41371
rect 39720 -41422 41831 -41388
rect 38919 -41488 41831 -41422
rect 41986 -41463 42065 -41432
rect 39720 -41499 41831 -41488
rect 41886 -41499 42065 -41463
rect 39720 -41541 42065 -41499
rect 40122 -41548 40348 -41541
rect 40159 -41555 40348 -41548
rect 41166 -41546 42065 -41541
rect 41166 -41565 41935 -41546
rect 39720 -41604 40162 -41589
rect 39720 -41653 41009 -41604
rect 39730 -42070 39764 -41653
rect 39926 -42070 39960 -41653
rect 40122 -41703 41009 -41653
rect 41172 -41691 41217 -41565
rect 40122 -42070 40156 -41703
rect 40339 -41869 40373 -41703
rect 40535 -41869 40569 -41703
rect 40731 -41869 40765 -41703
rect 40927 -41869 40961 -41703
rect 39645 -42119 39780 -42113
rect 39625 -42121 39780 -42119
rect 39211 -42157 39780 -42121
rect 39211 -43153 39347 -42157
rect 39625 -42159 39780 -42157
rect 39645 -42167 39780 -42159
rect 41177 -42281 41211 -41691
rect 41367 -41688 41412 -41565
rect 41373 -42281 41407 -41688
rect 41789 -41689 41834 -41565
rect 41986 -41571 42065 -41546
rect 41796 -42281 41830 -41689
rect 42326 -41417 42448 -40421
rect 42236 -41556 42448 -41417
rect 42236 -41584 42375 -41556
rect 35612 -43289 39347 -43153
rect 34828 -44315 35102 -44112
rect -32434 -44640 27308 -44504
rect 35612 -44703 35748 -43289
rect -32450 -44839 35748 -44703
rect 43579 -44130 43725 -38815
rect 46380 -38836 46414 -38246
rect 46570 -38243 46615 -38120
rect 46576 -38836 46610 -38243
rect 46992 -38244 47037 -38120
rect 47211 -38127 47273 -38113
rect 46999 -38836 47033 -38244
rect 54157 -37620 54191 -37354
rect 54353 -37620 54387 -37354
rect 54549 -37620 54583 -37354
rect 54745 -37620 54779 -37354
rect 54109 -37688 54827 -37620
rect 49729 -37719 54827 -37688
rect 49729 -37819 54463 -37719
rect 55130 -37800 55164 -37383
rect 55326 -37800 55360 -37383
rect 55522 -37750 55556 -37383
rect 55739 -37750 55773 -37584
rect 55935 -37750 55969 -37584
rect 56131 -37750 56165 -37584
rect 56327 -37750 56361 -37584
rect 55522 -37800 56409 -37750
rect 48369 -37889 54463 -37819
rect 55120 -37849 56409 -37800
rect 55120 -37863 55562 -37849
rect 48002 -37909 54463 -37889
rect 55119 -37892 55562 -37863
rect 55119 -37909 55737 -37892
rect 48002 -37942 56232 -37909
rect 48002 -38006 48407 -37942
rect 47439 -38016 47537 -38013
rect 48002 -38016 48119 -38006
rect 47439 -38133 48119 -38016
rect 48369 -38101 48407 -38006
rect 47439 -38139 47537 -38133
rect 48372 -38594 48406 -38101
rect 48566 -38099 48604 -37942
rect 48568 -38594 48602 -38099
rect 49158 -38122 49208 -37942
rect 49284 -38119 49334 -37942
rect 49163 -38594 49197 -38122
rect 49293 -38594 49327 -38119
rect 49515 -38104 49558 -37942
rect 49712 -38002 56232 -37942
rect 49521 -38394 49555 -38104
rect 49712 -38102 49755 -38002
rect 49717 -38394 49751 -38102
rect 47446 -40131 47848 -40065
rect 44951 -41107 44985 -40841
rect 45147 -41107 45181 -40841
rect 45343 -41107 45377 -40841
rect 45539 -41107 45573 -40841
rect 44903 -41206 45621 -41107
rect 45085 -41396 45257 -41206
rect 45924 -41287 45958 -40870
rect 46120 -41287 46154 -40870
rect 46316 -41237 46350 -40870
rect 46533 -41237 46567 -41071
rect 46729 -41237 46763 -41071
rect 46925 -41237 46959 -41071
rect 47121 -41237 47155 -41071
rect 46316 -41287 47203 -41237
rect 45914 -41336 47203 -41287
rect 45914 -41350 46356 -41336
rect 45913 -41379 46356 -41350
rect 45913 -41396 46531 -41379
rect 44915 -41507 47026 -41396
rect 44915 -41549 47130 -41507
rect 45317 -41556 45543 -41549
rect 45354 -41563 45543 -41556
rect 46361 -41573 47130 -41549
rect 44915 -41612 45357 -41597
rect 44915 -41661 46204 -41612
rect 44925 -42078 44959 -41661
rect 45121 -42078 45155 -41661
rect 45317 -41711 46204 -41661
rect 46367 -41699 46412 -41573
rect 45317 -42078 45351 -41711
rect 45534 -41877 45568 -41711
rect 45730 -41877 45764 -41711
rect 45926 -41877 45960 -41711
rect 46122 -41877 46156 -41711
rect 44840 -42127 44975 -42121
rect 44820 -42129 44975 -42127
rect 44292 -42165 44975 -42129
rect 44475 -43178 44611 -42165
rect 44820 -42167 44975 -42165
rect 44840 -42175 44975 -42167
rect 46372 -42289 46406 -41699
rect 46562 -41696 46607 -41573
rect 46568 -42289 46602 -41696
rect 46984 -41697 47029 -41573
rect 46991 -42289 47025 -41697
rect 47446 -41432 47512 -40131
rect 47429 -41545 47513 -41432
rect 47782 -41461 47848 -40131
rect 50679 -40338 50801 -38002
rect 54121 -38020 56232 -38002
rect 54121 -38027 56336 -38020
rect 56409 -38027 56471 -37999
rect 54121 -38062 56471 -38027
rect 54523 -38069 54749 -38062
rect 54560 -38076 54749 -38069
rect 55567 -38079 56471 -38062
rect 55567 -38086 56336 -38079
rect 54121 -38125 54563 -38110
rect 54121 -38174 55410 -38125
rect 52898 -38642 53627 -38577
rect 54131 -38591 54165 -38174
rect 54327 -38591 54361 -38174
rect 54523 -38224 55410 -38174
rect 55573 -38212 55618 -38086
rect 54523 -38591 54557 -38224
rect 54740 -38390 54774 -38224
rect 54936 -38390 54970 -38224
rect 55132 -38390 55166 -38224
rect 55328 -38390 55362 -38224
rect 54046 -38640 54181 -38634
rect 54026 -38642 54181 -38640
rect 52898 -38678 54181 -38642
rect 52898 -38723 53627 -38678
rect 54026 -38680 54181 -38678
rect 54046 -38688 54181 -38680
rect 50679 -40460 51311 -40338
rect 48619 -41138 48653 -40872
rect 48815 -41138 48849 -40872
rect 49011 -41138 49045 -40872
rect 49207 -41138 49241 -40872
rect 48571 -41237 49289 -41138
rect 48753 -41427 48925 -41237
rect 49592 -41318 49626 -40901
rect 49788 -41318 49822 -40901
rect 49984 -41268 50018 -40901
rect 50201 -41268 50235 -41102
rect 50397 -41268 50431 -41102
rect 50593 -41268 50627 -41102
rect 50789 -41268 50823 -41102
rect 49984 -41318 50871 -41268
rect 49582 -41367 50871 -41318
rect 49582 -41381 50024 -41367
rect 49581 -41410 50024 -41381
rect 49581 -41427 50199 -41410
rect 48583 -41461 50694 -41427
rect 47782 -41527 50694 -41461
rect 50849 -41502 50928 -41471
rect 48583 -41538 50694 -41527
rect 50749 -41538 50928 -41502
rect 48583 -41580 50928 -41538
rect 48985 -41587 49211 -41580
rect 49022 -41594 49211 -41587
rect 50029 -41585 50928 -41580
rect 50029 -41604 50798 -41585
rect 48583 -41643 49025 -41628
rect 48583 -41692 49872 -41643
rect 48593 -42109 48627 -41692
rect 48789 -42109 48823 -41692
rect 48985 -41742 49872 -41692
rect 50035 -41730 50080 -41604
rect 48985 -42109 49019 -41742
rect 49202 -41908 49236 -41742
rect 49398 -41908 49432 -41742
rect 49594 -41908 49628 -41742
rect 49790 -41908 49824 -41742
rect 48508 -42158 48643 -42152
rect 48488 -42160 48643 -42158
rect 48074 -42196 48643 -42160
rect 44475 -43192 44658 -43178
rect 48074 -43192 48210 -42196
rect 48488 -42198 48643 -42196
rect 48508 -42206 48643 -42198
rect 50040 -42320 50074 -41730
rect 50230 -41727 50275 -41604
rect 50236 -42320 50270 -41727
rect 50652 -41728 50697 -41604
rect 50849 -41610 50928 -41585
rect 50659 -42320 50693 -41728
rect 51189 -41456 51311 -40460
rect 51099 -41595 51311 -41456
rect 51099 -41623 51238 -41595
rect 44475 -43328 48210 -43192
rect 43525 -44269 43777 -44130
rect 44522 -44936 44658 -43328
rect 52898 -44091 53044 -38723
rect 55578 -38802 55612 -38212
rect 55768 -38209 55813 -38086
rect 55774 -38802 55808 -38209
rect 56190 -38210 56235 -38086
rect 56409 -38093 56471 -38079
rect 56197 -38802 56231 -38210
rect 62911 -37554 62945 -37288
rect 63107 -37554 63141 -37288
rect 63303 -37554 63337 -37288
rect 63499 -37554 63533 -37288
rect 62863 -37591 63581 -37554
rect 58912 -37653 63581 -37591
rect 58912 -37785 63217 -37653
rect 63884 -37734 63918 -37317
rect 64080 -37734 64114 -37317
rect 64276 -37684 64310 -37317
rect 64493 -37684 64527 -37518
rect 64689 -37684 64723 -37518
rect 64885 -37684 64919 -37518
rect 65081 -37684 65115 -37518
rect 64276 -37734 65163 -37684
rect 57567 -37843 63217 -37785
rect 63874 -37783 65163 -37734
rect 63874 -37797 64316 -37783
rect 63873 -37826 64316 -37797
rect 63873 -37843 64491 -37826
rect 57567 -37855 64986 -37843
rect 57200 -37908 64986 -37855
rect 57200 -37972 57605 -37908
rect 56637 -37982 56735 -37979
rect 57200 -37982 57317 -37972
rect 56637 -38099 57317 -37982
rect 57567 -38067 57605 -37972
rect 56637 -38105 56735 -38099
rect 57570 -38560 57604 -38067
rect 57764 -38065 57802 -37908
rect 57766 -38560 57800 -38065
rect 58356 -38088 58406 -37908
rect 58482 -38085 58532 -37908
rect 58361 -38560 58395 -38088
rect 58491 -38560 58525 -38085
rect 58713 -38070 58756 -37908
rect 58910 -37954 64986 -37908
rect 58910 -37961 65090 -37954
rect 65163 -37961 65225 -37933
rect 58910 -37970 65225 -37961
rect 58719 -38360 58753 -38070
rect 58910 -38068 58953 -37970
rect 58915 -38360 58949 -38068
rect 56644 -40097 57046 -40031
rect 54149 -41073 54183 -40807
rect 54345 -41073 54379 -40807
rect 54541 -41073 54575 -40807
rect 54737 -41073 54771 -40807
rect 54101 -41172 54819 -41073
rect 54283 -41362 54455 -41172
rect 55122 -41253 55156 -40836
rect 55318 -41253 55352 -40836
rect 55514 -41203 55548 -40836
rect 55731 -41203 55765 -41037
rect 55927 -41203 55961 -41037
rect 56123 -41203 56157 -41037
rect 56319 -41203 56353 -41037
rect 55514 -41253 56401 -41203
rect 55112 -41302 56401 -41253
rect 55112 -41316 55554 -41302
rect 55111 -41345 55554 -41316
rect 55111 -41362 55729 -41345
rect 54113 -41473 56224 -41362
rect 54113 -41515 56328 -41473
rect 54515 -41522 54741 -41515
rect 54552 -41529 54741 -41522
rect 55559 -41539 56328 -41515
rect 54113 -41578 54555 -41563
rect 54113 -41627 55402 -41578
rect 54123 -42044 54157 -41627
rect 54319 -42044 54353 -41627
rect 54515 -41677 55402 -41627
rect 55565 -41665 55610 -41539
rect 54515 -42044 54549 -41677
rect 54732 -41843 54766 -41677
rect 54928 -41843 54962 -41677
rect 55124 -41843 55158 -41677
rect 55320 -41843 55354 -41677
rect 54038 -42093 54173 -42087
rect 54018 -42095 54173 -42093
rect 53490 -42131 54173 -42095
rect 53673 -43158 53809 -42131
rect 54018 -42133 54173 -42131
rect 54038 -42141 54173 -42133
rect 55570 -42255 55604 -41665
rect 55760 -41662 55805 -41539
rect 55766 -42255 55800 -41662
rect 56182 -41663 56227 -41539
rect 56189 -42255 56223 -41663
rect 56644 -41398 56710 -40097
rect 56627 -41511 56711 -41398
rect 56980 -41427 57046 -40097
rect 59877 -40304 59999 -37970
rect 62875 -37996 65225 -37970
rect 63277 -38003 63503 -37996
rect 63314 -38010 63503 -38003
rect 64321 -38013 65225 -37996
rect 64321 -38020 65090 -38013
rect 62875 -38059 63317 -38044
rect 62875 -38108 64164 -38059
rect 61425 -38576 62351 -38452
rect 62885 -38525 62919 -38108
rect 63081 -38525 63115 -38108
rect 63277 -38158 64164 -38108
rect 64327 -38146 64372 -38020
rect 63277 -38525 63311 -38158
rect 63494 -38324 63528 -38158
rect 63690 -38324 63724 -38158
rect 63886 -38324 63920 -38158
rect 64082 -38324 64116 -38158
rect 62800 -38574 62935 -38568
rect 62780 -38576 62935 -38574
rect 61425 -38612 62935 -38576
rect 61425 -38691 62351 -38612
rect 62780 -38614 62935 -38612
rect 62800 -38622 62935 -38614
rect 59877 -40426 60509 -40304
rect 57817 -41104 57851 -40838
rect 58013 -41104 58047 -40838
rect 58209 -41104 58243 -40838
rect 58405 -41104 58439 -40838
rect 57769 -41203 58487 -41104
rect 57951 -41393 58123 -41203
rect 58790 -41284 58824 -40867
rect 58986 -41284 59020 -40867
rect 59182 -41234 59216 -40867
rect 59399 -41234 59433 -41068
rect 59595 -41234 59629 -41068
rect 59791 -41234 59825 -41068
rect 59987 -41234 60021 -41068
rect 59182 -41284 60069 -41234
rect 58780 -41333 60069 -41284
rect 58780 -41347 59222 -41333
rect 58779 -41376 59222 -41347
rect 58779 -41393 59397 -41376
rect 57781 -41427 59892 -41393
rect 56980 -41493 59892 -41427
rect 60047 -41468 60126 -41437
rect 57781 -41504 59892 -41493
rect 59947 -41504 60126 -41468
rect 57781 -41546 60126 -41504
rect 58183 -41553 58409 -41546
rect 58220 -41560 58409 -41553
rect 59227 -41551 60126 -41546
rect 59227 -41570 59996 -41551
rect 57781 -41609 58223 -41594
rect 57781 -41658 59070 -41609
rect 57791 -42075 57825 -41658
rect 57987 -42075 58021 -41658
rect 58183 -41708 59070 -41658
rect 59233 -41696 59278 -41570
rect 58183 -42075 58217 -41708
rect 58400 -41874 58434 -41708
rect 58596 -41874 58630 -41708
rect 58792 -41874 58826 -41708
rect 58988 -41874 59022 -41708
rect 57706 -42124 57841 -42118
rect 57686 -42126 57841 -42124
rect 57272 -42162 57841 -42126
rect 57272 -43158 57408 -42162
rect 57686 -42164 57841 -42162
rect 57706 -42172 57841 -42164
rect 59238 -42286 59272 -41696
rect 59428 -41693 59473 -41570
rect 59434 -42286 59468 -41693
rect 59850 -41694 59895 -41570
rect 60047 -41576 60126 -41551
rect 59857 -42286 59891 -41694
rect 60387 -41422 60509 -40426
rect 60297 -41561 60509 -41422
rect 60297 -41589 60436 -41561
rect 53673 -43294 57408 -43158
rect 52864 -44296 53096 -44091
rect -32458 -45072 44658 -44936
rect 53673 -45191 53809 -43294
rect 61425 -44076 61664 -38691
rect 64332 -38736 64366 -38146
rect 64522 -38143 64567 -38020
rect 64528 -38736 64562 -38143
rect 64944 -38144 64989 -38020
rect 65163 -38027 65225 -38013
rect 64951 -38736 64985 -38144
rect 72064 -37537 72098 -37271
rect 72260 -37537 72294 -37271
rect 72456 -37537 72490 -37271
rect 72652 -37537 72686 -37271
rect 72016 -37612 72734 -37537
rect 67659 -37636 72734 -37612
rect 67659 -37719 72370 -37636
rect 73037 -37717 73071 -37300
rect 73233 -37717 73267 -37300
rect 73429 -37667 73463 -37300
rect 73646 -37667 73680 -37501
rect 73842 -37667 73876 -37501
rect 74038 -37667 74072 -37501
rect 74234 -37667 74268 -37501
rect 73429 -37717 74316 -37667
rect 66321 -37789 72370 -37719
rect 73027 -37766 74316 -37717
rect 73027 -37780 73469 -37766
rect 65954 -37826 72370 -37789
rect 73026 -37809 73469 -37780
rect 73026 -37826 73644 -37809
rect 65954 -37842 74139 -37826
rect 65954 -37906 66359 -37842
rect 65391 -37916 65489 -37913
rect 65954 -37916 66071 -37906
rect 65391 -38033 66071 -37916
rect 66321 -38001 66359 -37906
rect 65391 -38039 65489 -38033
rect 66324 -38494 66358 -38001
rect 66518 -37999 66556 -37842
rect 66520 -38494 66554 -37999
rect 67110 -38022 67160 -37842
rect 67236 -38019 67286 -37842
rect 67115 -38494 67149 -38022
rect 67245 -38494 67279 -38019
rect 67467 -38004 67510 -37842
rect 67659 -37876 74139 -37842
rect 67473 -38294 67507 -38004
rect 67664 -38002 67707 -37876
rect 67669 -38294 67703 -38002
rect 61363 -44308 61711 -44076
rect 65398 -40031 65800 -39965
rect 62903 -41007 62937 -40741
rect 63099 -41007 63133 -40741
rect 63295 -41007 63329 -40741
rect 63491 -41007 63525 -40741
rect 62855 -41106 63573 -41007
rect 63037 -41296 63209 -41106
rect 63876 -41187 63910 -40770
rect 64072 -41187 64106 -40770
rect 64268 -41137 64302 -40770
rect 64485 -41137 64519 -40971
rect 64681 -41137 64715 -40971
rect 64877 -41137 64911 -40971
rect 65073 -41137 65107 -40971
rect 64268 -41187 65155 -41137
rect 63866 -41236 65155 -41187
rect 63866 -41250 64308 -41236
rect 63865 -41279 64308 -41250
rect 63865 -41296 64483 -41279
rect 62867 -41407 64978 -41296
rect 62867 -41449 65082 -41407
rect 63269 -41456 63495 -41449
rect 63306 -41463 63495 -41456
rect 64313 -41473 65082 -41449
rect 62867 -41512 63309 -41497
rect 62867 -41561 64156 -41512
rect 62877 -41978 62911 -41561
rect 63073 -41978 63107 -41561
rect 63269 -41611 64156 -41561
rect 64319 -41599 64364 -41473
rect 63269 -41978 63303 -41611
rect 63486 -41777 63520 -41611
rect 63682 -41777 63716 -41611
rect 63878 -41777 63912 -41611
rect 64074 -41777 64108 -41611
rect 64324 -42189 64358 -41599
rect 64514 -41596 64559 -41473
rect 64520 -42189 64554 -41596
rect 64936 -41597 64981 -41473
rect 64943 -42189 64977 -41597
rect 65398 -41332 65464 -40031
rect 65381 -41445 65465 -41332
rect 65734 -41361 65800 -40031
rect 68631 -40238 68753 -37876
rect 72028 -37937 74139 -37876
rect 72028 -37944 74243 -37937
rect 74316 -37944 74378 -37916
rect 72028 -37979 74378 -37944
rect 72430 -37986 72656 -37979
rect 72467 -37993 72656 -37986
rect 73474 -37996 74378 -37979
rect 73474 -38003 74243 -37996
rect 72028 -38042 72470 -38027
rect 72028 -38091 73317 -38042
rect 70753 -38559 71417 -38480
rect 72038 -38508 72072 -38091
rect 72234 -38508 72268 -38091
rect 72430 -38141 73317 -38091
rect 73480 -38129 73525 -38003
rect 72430 -38508 72464 -38141
rect 72647 -38307 72681 -38141
rect 72843 -38307 72877 -38141
rect 73039 -38307 73073 -38141
rect 73235 -38307 73269 -38141
rect 71953 -38557 72088 -38551
rect 71933 -38559 72088 -38557
rect 70753 -38595 72088 -38559
rect 70753 -38665 71417 -38595
rect 71933 -38597 72088 -38595
rect 71953 -38605 72088 -38597
rect 68631 -40360 69263 -40238
rect 66571 -41038 66605 -40772
rect 66767 -41038 66801 -40772
rect 66963 -41038 66997 -40772
rect 67159 -41038 67193 -40772
rect 66523 -41137 67241 -41038
rect 66705 -41327 66877 -41137
rect 67544 -41218 67578 -40801
rect 67740 -41218 67774 -40801
rect 67936 -41168 67970 -40801
rect 68153 -41168 68187 -41002
rect 68349 -41168 68383 -41002
rect 68545 -41168 68579 -41002
rect 68741 -41168 68775 -41002
rect 67936 -41218 68823 -41168
rect 67534 -41267 68823 -41218
rect 67534 -41281 67976 -41267
rect 67533 -41310 67976 -41281
rect 67533 -41327 68151 -41310
rect 66535 -41361 68646 -41327
rect 65734 -41427 68646 -41361
rect 68801 -41402 68880 -41371
rect 66535 -41438 68646 -41427
rect 68701 -41438 68880 -41402
rect 66535 -41480 68880 -41438
rect 66937 -41487 67163 -41480
rect 66974 -41494 67163 -41487
rect 67981 -41485 68880 -41480
rect 67981 -41504 68750 -41485
rect 66535 -41543 66977 -41528
rect 66535 -41592 67824 -41543
rect 66545 -42009 66579 -41592
rect 66741 -42009 66775 -41592
rect 66937 -41642 67824 -41592
rect 67987 -41630 68032 -41504
rect 66937 -42009 66971 -41642
rect 67154 -41808 67188 -41642
rect 67350 -41808 67384 -41642
rect 67546 -41808 67580 -41642
rect 67742 -41808 67776 -41642
rect 67992 -42220 68026 -41630
rect 68182 -41627 68227 -41504
rect 68188 -42220 68222 -41627
rect 68604 -41628 68649 -41504
rect 68801 -41510 68880 -41485
rect 68611 -42220 68645 -41628
rect 69141 -41356 69263 -40360
rect 69051 -41495 69263 -41356
rect 69051 -41523 69190 -41495
rect -32482 -45327 53809 -45191
rect -29580 -46390 -28157 -45411
rect 70753 -44073 70938 -38665
rect 73485 -38719 73519 -38129
rect 73675 -38126 73720 -38003
rect 73681 -38719 73715 -38126
rect 74097 -38127 74142 -38003
rect 74316 -38010 74378 -37996
rect 74104 -38719 74138 -38127
rect 81428 -37499 81462 -37233
rect 81624 -37499 81658 -37233
rect 81820 -37499 81854 -37233
rect 82016 -37499 82050 -37233
rect 81380 -37543 82098 -37499
rect 76821 -37598 82098 -37543
rect 76821 -37702 81734 -37598
rect 82401 -37679 82435 -37262
rect 82597 -37679 82631 -37262
rect 82793 -37629 82827 -37262
rect 83010 -37629 83044 -37463
rect 83206 -37629 83240 -37463
rect 83402 -37629 83436 -37463
rect 83598 -37629 83632 -37463
rect 82793 -37679 83680 -37629
rect 75474 -37772 81734 -37702
rect 82391 -37728 83680 -37679
rect 82391 -37742 82833 -37728
rect 75107 -37788 81734 -37772
rect 82390 -37771 82833 -37742
rect 82390 -37788 83008 -37771
rect 75107 -37825 83503 -37788
rect 75107 -37889 75512 -37825
rect 74544 -37899 74642 -37896
rect 75107 -37899 75224 -37889
rect 74544 -38016 75224 -37899
rect 75474 -37984 75512 -37889
rect 74544 -38022 74642 -38016
rect 75477 -38477 75511 -37984
rect 75671 -37982 75709 -37825
rect 75673 -38477 75707 -37982
rect 76263 -38005 76313 -37825
rect 76389 -38002 76439 -37825
rect 76268 -38477 76302 -38005
rect 76398 -38477 76432 -38002
rect 76620 -37987 76663 -37825
rect 76817 -37885 83503 -37825
rect 76626 -38277 76660 -37987
rect 76817 -37985 76860 -37885
rect 76822 -38277 76856 -37985
rect 74551 -40014 74953 -39948
rect 72056 -40990 72090 -40724
rect 72252 -40990 72286 -40724
rect 72448 -40990 72482 -40724
rect 72644 -40990 72678 -40724
rect 72008 -41089 72726 -40990
rect 72190 -41279 72362 -41089
rect 73029 -41170 73063 -40753
rect 73225 -41170 73259 -40753
rect 73421 -41120 73455 -40753
rect 73638 -41120 73672 -40954
rect 73834 -41120 73868 -40954
rect 74030 -41120 74064 -40954
rect 74226 -41120 74260 -40954
rect 73421 -41170 74308 -41120
rect 73019 -41219 74308 -41170
rect 73019 -41233 73461 -41219
rect 73018 -41262 73461 -41233
rect 73018 -41279 73636 -41262
rect 72020 -41390 74131 -41279
rect 72020 -41432 74235 -41390
rect 72422 -41439 72648 -41432
rect 72459 -41446 72648 -41439
rect 73466 -41456 74235 -41432
rect 72020 -41495 72462 -41480
rect 72020 -41544 73309 -41495
rect 72030 -41961 72064 -41544
rect 72226 -41961 72260 -41544
rect 72422 -41594 73309 -41544
rect 73472 -41582 73517 -41456
rect 72422 -41961 72456 -41594
rect 72639 -41760 72673 -41594
rect 72835 -41760 72869 -41594
rect 73031 -41760 73065 -41594
rect 73227 -41760 73261 -41594
rect 73477 -42172 73511 -41582
rect 73667 -41579 73712 -41456
rect 73673 -42172 73707 -41579
rect 74089 -41580 74134 -41456
rect 74096 -42172 74130 -41580
rect 74551 -41315 74617 -40014
rect 74534 -41428 74618 -41315
rect 74887 -41344 74953 -40014
rect 77784 -40221 77906 -37885
rect 81392 -37899 83503 -37885
rect 81392 -37906 83607 -37899
rect 83680 -37906 83742 -37878
rect 81392 -37941 83742 -37906
rect 81794 -37948 82020 -37941
rect 81831 -37955 82020 -37948
rect 82838 -37958 83742 -37941
rect 82838 -37965 83607 -37958
rect 81392 -38004 81834 -37989
rect 81392 -38053 82681 -38004
rect 79670 -38521 80878 -38338
rect 81402 -38470 81436 -38053
rect 81598 -38470 81632 -38053
rect 81794 -38103 82681 -38053
rect 82844 -38091 82889 -37965
rect 81794 -38470 81828 -38103
rect 82011 -38269 82045 -38103
rect 82207 -38269 82241 -38103
rect 82403 -38269 82437 -38103
rect 82599 -38269 82633 -38103
rect 81317 -38519 81452 -38513
rect 81297 -38521 81452 -38519
rect 79670 -38557 81452 -38521
rect 79670 -38632 80878 -38557
rect 81297 -38559 81452 -38557
rect 81317 -38567 81452 -38559
rect 77784 -40343 78416 -40221
rect 75724 -41021 75758 -40755
rect 75920 -41021 75954 -40755
rect 76116 -41021 76150 -40755
rect 76312 -41021 76346 -40755
rect 75676 -41120 76394 -41021
rect 75858 -41310 76030 -41120
rect 76697 -41201 76731 -40784
rect 76893 -41201 76927 -40784
rect 77089 -41151 77123 -40784
rect 77306 -41151 77340 -40985
rect 77502 -41151 77536 -40985
rect 77698 -41151 77732 -40985
rect 77894 -41151 77928 -40985
rect 77089 -41201 77976 -41151
rect 76687 -41250 77976 -41201
rect 76687 -41264 77129 -41250
rect 76686 -41293 77129 -41264
rect 76686 -41310 77304 -41293
rect 75688 -41344 77799 -41310
rect 74887 -41410 77799 -41344
rect 77954 -41385 78033 -41354
rect 75688 -41421 77799 -41410
rect 77854 -41421 78033 -41385
rect 75688 -41463 78033 -41421
rect 76090 -41470 76316 -41463
rect 76127 -41477 76316 -41470
rect 77134 -41468 78033 -41463
rect 77134 -41487 77903 -41468
rect 75688 -41526 76130 -41511
rect 75688 -41575 76977 -41526
rect 75698 -41992 75732 -41575
rect 75894 -41992 75928 -41575
rect 76090 -41625 76977 -41575
rect 77140 -41613 77185 -41487
rect 76090 -41992 76124 -41625
rect 76307 -41791 76341 -41625
rect 76503 -41791 76537 -41625
rect 76699 -41791 76733 -41625
rect 76895 -41791 76929 -41625
rect 77145 -42203 77179 -41613
rect 77335 -41610 77380 -41487
rect 77341 -42203 77375 -41610
rect 77757 -41611 77802 -41487
rect 77954 -41493 78033 -41468
rect 77764 -42203 77798 -41611
rect 78294 -41339 78416 -40343
rect 78204 -41478 78416 -41339
rect 78204 -41506 78343 -41478
rect 70668 -44318 71050 -44073
rect 79670 -44076 79964 -38632
rect 82849 -38681 82883 -38091
rect 83039 -38088 83084 -37965
rect 83045 -38681 83079 -38088
rect 83461 -38089 83506 -37965
rect 83680 -37972 83742 -37958
rect 83468 -38681 83502 -38089
rect 86596 -37664 87071 -33752
rect 90604 -34632 92221 -33888
rect 88763 -35170 92221 -34632
rect 90604 -35414 92221 -35170
rect 84838 -37734 87270 -37664
rect 84471 -37786 87270 -37734
rect 84471 -37787 86224 -37786
rect 84471 -37851 84876 -37787
rect 83908 -37861 84006 -37858
rect 84471 -37861 84588 -37851
rect 83908 -37978 84588 -37861
rect 84838 -37946 84876 -37851
rect 83908 -37984 84006 -37978
rect 84841 -38439 84875 -37946
rect 85035 -37944 85073 -37787
rect 85037 -38439 85071 -37944
rect 85627 -37967 85677 -37787
rect 85753 -37964 85803 -37787
rect 85632 -38439 85666 -37967
rect 85762 -38439 85796 -37964
rect 85984 -37949 86027 -37787
rect 85990 -38239 86024 -37949
rect 86181 -37947 86224 -37787
rect 86186 -38239 86220 -37947
rect 79621 -44314 80021 -44076
rect 83915 -39976 84317 -39910
rect 81420 -40952 81454 -40686
rect 81616 -40952 81650 -40686
rect 81812 -40952 81846 -40686
rect 82008 -40952 82042 -40686
rect 81372 -41051 82090 -40952
rect 81554 -41241 81726 -41051
rect 82393 -41132 82427 -40715
rect 82589 -41132 82623 -40715
rect 82785 -41082 82819 -40715
rect 83002 -41082 83036 -40916
rect 83198 -41082 83232 -40916
rect 83394 -41082 83428 -40916
rect 83590 -41082 83624 -40916
rect 82785 -41132 83672 -41082
rect 82383 -41181 83672 -41132
rect 82383 -41195 82825 -41181
rect 82382 -41224 82825 -41195
rect 82382 -41241 83000 -41224
rect 81384 -41352 83495 -41241
rect 81384 -41394 83599 -41352
rect 81786 -41401 82012 -41394
rect 81823 -41408 82012 -41401
rect 82830 -41418 83599 -41394
rect 81384 -41457 81826 -41442
rect 81384 -41506 82673 -41457
rect 81394 -41923 81428 -41506
rect 81590 -41923 81624 -41506
rect 81786 -41556 82673 -41506
rect 82836 -41544 82881 -41418
rect 81786 -41923 81820 -41556
rect 82003 -41722 82037 -41556
rect 82199 -41722 82233 -41556
rect 82395 -41722 82429 -41556
rect 82591 -41722 82625 -41556
rect 82841 -42134 82875 -41544
rect 83031 -41541 83076 -41418
rect 83037 -42134 83071 -41541
rect 83453 -41542 83498 -41418
rect 83460 -42134 83494 -41542
rect 83915 -41277 83981 -39976
rect 83898 -41390 83982 -41277
rect 84251 -41306 84317 -39976
rect 87148 -40183 87270 -37786
rect 87148 -40305 87780 -40183
rect 85088 -40983 85122 -40717
rect 85284 -40983 85318 -40717
rect 85480 -40983 85514 -40717
rect 85676 -40983 85710 -40717
rect 85040 -41082 85758 -40983
rect 85222 -41272 85394 -41082
rect 86061 -41163 86095 -40746
rect 86257 -41163 86291 -40746
rect 86453 -41113 86487 -40746
rect 86670 -41113 86704 -40947
rect 86866 -41113 86900 -40947
rect 87062 -41113 87096 -40947
rect 87258 -41113 87292 -40947
rect 86453 -41163 87340 -41113
rect 86051 -41212 87340 -41163
rect 86051 -41226 86493 -41212
rect 86050 -41255 86493 -41226
rect 86050 -41272 86668 -41255
rect 85052 -41306 87163 -41272
rect 84251 -41372 87163 -41306
rect 87318 -41347 87397 -41316
rect 85052 -41383 87163 -41372
rect 87218 -41383 87397 -41347
rect 85052 -41425 87397 -41383
rect 85454 -41432 85680 -41425
rect 85491 -41439 85680 -41432
rect 86498 -41430 87397 -41425
rect 86498 -41449 87267 -41430
rect 85052 -41488 85494 -41473
rect 85052 -41537 86341 -41488
rect 85062 -41954 85096 -41537
rect 85258 -41954 85292 -41537
rect 85454 -41587 86341 -41537
rect 86504 -41575 86549 -41449
rect 85454 -41954 85488 -41587
rect 85671 -41753 85705 -41587
rect 85867 -41753 85901 -41587
rect 86063 -41753 86097 -41587
rect 86259 -41753 86293 -41587
rect 86509 -42165 86543 -41575
rect 86699 -41572 86744 -41449
rect 86705 -42165 86739 -41572
rect 87121 -41573 87166 -41449
rect 87318 -41455 87397 -41430
rect 87128 -42165 87162 -41573
rect 87658 -41301 87780 -40305
rect 87568 -41440 87780 -41301
rect 87568 -41468 87707 -41440
rect 95829 -46113 98798 -31308
rect -23503 -46390 -23290 -46358
rect -29580 -46526 10852 -46390
rect -23503 -46536 -23290 -46526
rect 83333 -49082 98798 -46113
rect -32776 -50847 -27886 -50668
rect 83333 -50760 86302 -49082
rect -28065 -52016 -27886 -50847
rect 26626 -50981 87774 -50760
rect 7598 -51743 87774 -50981
rect -28016 -52164 -27982 -52016
rect -28016 -52198 -27428 -52164
rect -27389 -52282 -27341 -52116
rect -27836 -52316 -27341 -52282
rect -27836 -52434 -27428 -52400
rect -27389 -52518 -27341 -52316
rect -27836 -52552 -27341 -52518
rect -27836 -52670 -27428 -52636
rect -27389 -52754 -27341 -52552
rect -27836 -52788 -27341 -52754
rect -27836 -52906 -27428 -52872
rect -27389 -52990 -27341 -52788
rect -27836 -53024 -27341 -52990
rect -27836 -53142 -27428 -53108
rect -27389 -53214 -27341 -53024
rect -27269 -53214 -27203 -52226
rect 7598 -52897 8360 -51743
rect 26626 -51863 87774 -51743
rect -6631 -52908 8829 -52897
rect -8962 -52944 8829 -52908
rect -27389 -53226 -27203 -53214
rect -27836 -53260 -27203 -53226
rect -27389 -53273 -27203 -53260
rect -27836 -53378 -27428 -53344
rect -27389 -53462 -27341 -53273
rect -27836 -53496 -27341 -53462
rect -27836 -53614 -27428 -53580
rect -27389 -53691 -27341 -53496
rect -27269 -53691 -27203 -53273
rect -13987 -52997 8829 -52944
rect -13987 -53007 -8762 -52997
rect -13987 -53012 -12414 -53007
rect -11516 -53012 -9714 -53007
rect -13987 -53571 -13898 -53012
rect -13738 -53303 -13704 -53012
rect -13542 -53303 -13508 -53012
rect -13346 -53303 -13312 -53012
rect -12901 -53303 -12867 -53012
rect -27389 -53698 -27203 -53691
rect -27836 -53732 -27203 -53698
rect -27389 -53750 -27203 -53732
rect -27836 -53850 -27428 -53816
rect -27389 -53922 -27341 -53750
rect -27269 -53808 -27203 -53750
rect -22950 -53784 -13898 -53571
rect -22950 -53794 -20715 -53784
rect -22950 -53808 -22678 -53794
rect -27269 -53922 -22678 -53808
rect -27389 -53934 -22678 -53922
rect -27836 -53968 -22678 -53934
rect -27389 -53981 -22678 -53968
rect -27836 -54086 -27428 -54052
rect -27389 -54158 -27341 -53981
rect -27269 -54080 -22678 -53981
rect -27269 -54158 -27203 -54080
rect -27389 -54170 -27203 -54158
rect -27836 -54204 -27203 -54170
rect -27389 -54217 -27203 -54204
rect -27836 -54322 -27428 -54288
rect -27389 -54396 -27341 -54217
rect -27269 -54396 -27203 -54217
rect -27389 -54406 -27203 -54396
rect -27836 -54440 -27203 -54406
rect -27389 -54455 -27203 -54440
rect -27836 -54558 -27428 -54524
rect -27389 -54636 -27341 -54455
rect -27269 -54594 -27203 -54455
rect -22950 -54594 -22678 -54080
rect -22483 -54302 -22422 -54099
rect -22292 -54220 -22231 -54020
rect -22183 -54137 -22122 -53934
rect -21337 -54090 -21303 -53794
rect -21141 -54090 -21107 -53794
rect -20945 -54090 -20911 -53794
rect -20749 -54090 -20715 -53794
rect -20212 -53798 -19967 -53784
rect -20207 -54090 -20173 -53798
rect -21414 -54137 -21279 -54129
rect -22183 -54172 -21279 -54137
rect -21433 -54174 -21279 -54172
rect -21414 -54183 -21279 -54174
rect -21078 -54220 -20943 -54211
rect -22292 -54258 -20943 -54220
rect -21078 -54265 -20943 -54258
rect -20890 -54302 -20755 -54289
rect -22483 -54336 -20755 -54302
rect -22483 -54337 -22422 -54336
rect -20890 -54343 -20755 -54336
rect -27269 -54636 -22678 -54594
rect -27389 -54642 -22678 -54636
rect -27836 -54676 -22678 -54642
rect -27389 -54695 -22678 -54676
rect -27836 -54794 -27428 -54760
rect -27389 -54866 -27341 -54695
rect -27269 -54866 -22678 -54695
rect -27389 -54878 -27203 -54866
rect -27836 -54912 -27203 -54878
rect -27389 -54925 -27203 -54912
rect -27836 -55030 -27428 -54996
rect -27389 -55103 -27341 -54925
rect -27269 -55103 -27203 -54925
rect -27389 -55114 -27203 -55103
rect -27836 -55148 -27203 -55114
rect -27389 -55162 -27203 -55148
rect -27836 -55266 -27428 -55232
rect -27389 -55337 -27341 -55162
rect -27269 -55328 -27203 -55162
rect -22950 -55328 -22678 -54866
rect -20011 -54090 -19977 -53798
rect -19390 -53846 -18063 -53784
rect -19390 -53901 -18059 -53846
rect -19338 -54312 -19304 -53901
rect -19142 -54312 -19108 -53901
rect -18946 -53945 -18059 -53901
rect -18946 -54312 -18912 -53945
rect -18729 -54111 -18695 -53945
rect -18533 -54111 -18499 -53945
rect -18337 -54111 -18303 -53945
rect -18141 -54111 -18107 -53945
rect -19558 -54457 -19421 -54453
rect -19596 -54459 -19369 -54457
rect -18958 -54459 -18884 -54433
rect -19596 -54497 -18884 -54459
rect -19558 -54511 -19421 -54497
rect -19370 -54498 -18884 -54497
rect -19370 -54499 -19299 -54498
rect -18958 -54504 -18884 -54498
rect -17787 -54877 -17652 -54869
rect -17807 -54879 -17652 -54877
rect -18198 -54915 -17652 -54879
rect -22084 -55176 -22024 -55100
rect -22084 -55216 -22016 -55176
rect -27269 -55337 -22678 -55328
rect -27389 -55350 -22678 -55337
rect -27836 -55384 -22678 -55350
rect -27389 -55396 -22678 -55384
rect -27836 -55502 -27428 -55468
rect -27389 -55571 -27341 -55396
rect -27269 -55535 -22678 -55396
rect -22631 -55431 -22530 -55258
rect -22084 -55293 -22024 -55216
rect -19667 -55293 -19535 -55284
rect -22084 -55333 -19535 -55293
rect -22084 -55337 -22024 -55333
rect -19667 -55337 -19535 -55333
rect -18121 -55431 -18064 -54915
rect -17807 -54917 -17652 -54915
rect -17787 -54923 -17652 -54917
rect -17702 -55383 -17668 -54966
rect -17506 -55383 -17472 -54966
rect -17310 -55333 -17276 -54966
rect -17093 -55333 -17059 -55167
rect -16897 -55333 -16863 -55167
rect -16701 -55333 -16667 -55167
rect -16505 -55333 -16471 -55167
rect -17310 -55383 -16423 -55333
rect -16255 -55345 -16221 -54755
rect -22631 -55494 -18064 -55431
rect -17712 -55432 -16423 -55383
rect -17712 -55447 -17270 -55432
rect -16260 -55471 -16215 -55345
rect -16059 -55348 -16025 -54755
rect -16065 -55471 -16020 -55348
rect -15636 -55347 -15602 -54755
rect -15643 -55471 -15598 -55347
rect -17273 -55488 -17084 -55481
rect -22631 -55501 -22530 -55494
rect -17310 -55495 -17084 -55488
rect -16266 -55495 -15497 -55471
rect -17712 -55535 -15497 -55495
rect -27269 -55537 -15497 -55535
rect -27269 -55571 -15601 -55537
rect -27389 -55586 -15601 -55571
rect -27836 -55600 -15601 -55586
rect -27836 -55620 -27203 -55600
rect -27389 -55630 -27203 -55620
rect -27836 -55738 -27428 -55704
rect -27389 -55822 -27341 -55630
rect -27836 -55856 -27341 -55822
rect -28644 -55954 -28236 -55920
rect -28644 -56190 -28236 -56156
rect -27836 -55974 -27428 -55940
rect -27389 -56070 -27341 -55856
rect -27836 -56104 -27341 -56070
rect -27389 -56296 -27341 -56104
rect -27269 -56296 -27203 -55630
rect -22950 -55648 -15601 -55600
rect -22950 -55734 -18137 -55648
rect -22950 -55767 -18147 -55734
rect -21290 -55804 -20001 -55767
rect -27389 -56306 -27203 -56296
rect -27836 -56340 -27203 -56306
rect -21280 -56221 -21246 -55804
rect -21084 -56221 -21050 -55804
rect -20888 -55854 -20001 -55804
rect -20888 -56221 -20854 -55854
rect -20671 -56020 -20637 -55854
rect -20475 -56020 -20441 -55854
rect -20279 -56020 -20245 -55854
rect -20083 -56020 -20049 -55854
rect -19507 -56026 -19473 -55767
rect -19311 -56026 -19277 -55767
rect -19115 -56026 -19081 -55767
rect -18919 -56026 -18885 -55767
rect -18377 -56026 -18343 -55767
rect -27389 -56355 -27203 -56340
rect -28644 -56426 -28236 -56392
rect -27389 -56527 -27341 -56355
rect -27269 -56527 -27203 -56355
rect -27389 -56542 -27203 -56527
rect -27836 -56576 -27203 -56542
rect -27389 -56586 -27203 -56576
rect -28644 -56662 -28236 -56628
rect -27389 -56763 -27341 -56586
rect -27269 -56763 -27203 -56586
rect -27389 -56778 -27203 -56763
rect -27836 -56812 -27203 -56778
rect -18181 -56026 -18147 -55767
rect -17542 -55838 -17370 -55648
rect -16714 -55665 -16096 -55648
rect -16714 -55694 -16271 -55665
rect -16713 -55708 -16271 -55694
rect -16713 -55757 -15424 -55708
rect -17724 -55937 -17006 -55838
rect -17676 -56203 -17642 -55937
rect -17480 -56203 -17446 -55937
rect -17284 -56203 -17250 -55937
rect -17088 -56203 -17054 -55937
rect -16703 -56174 -16669 -55757
rect -16507 -56174 -16473 -55757
rect -16311 -55807 -15424 -55757
rect -16311 -56174 -16277 -55807
rect -16094 -55973 -16060 -55807
rect -15898 -55973 -15864 -55807
rect -15702 -55973 -15668 -55807
rect -15506 -55973 -15472 -55807
rect -27389 -56822 -27203 -56812
rect -28644 -56898 -28236 -56864
rect -27389 -56998 -27341 -56822
rect -27269 -56998 -27203 -56822
rect -27389 -57014 -27203 -56998
rect -27836 -57048 -27203 -57014
rect -27389 -57057 -27203 -57048
rect -13987 -54707 -13898 -53784
rect -12705 -53303 -12671 -53012
rect -12509 -53303 -12475 -53012
rect -11038 -53303 -11004 -53012
rect -10842 -53303 -10808 -53012
rect -10646 -53303 -10612 -53012
rect -10201 -53303 -10167 -53012
rect -10005 -53303 -9971 -53012
rect -9809 -53303 -9775 -53012
rect -7380 -53121 -7335 -52997
rect -7376 -53713 -7342 -53121
rect -6958 -53120 -6913 -52997
rect -6953 -53713 -6919 -53120
rect -6763 -53123 -6718 -52997
rect -6633 -53090 8829 -52997
rect -6757 -53713 -6723 -53123
rect -13640 -54704 -13606 -54413
rect -13444 -54704 -13410 -54413
rect -13248 -54704 -13214 -54413
rect -11897 -54704 -11863 -54413
rect -11701 -54704 -11667 -54413
rect -11505 -54704 -11471 -54413
rect -10940 -54704 -10906 -54413
rect -10744 -54704 -10710 -54413
rect -10548 -54704 -10514 -54413
rect -9197 -54704 -9163 -54413
rect -9001 -54704 -8967 -54413
rect -8805 -54704 -8771 -54413
rect -8315 -54704 -8281 -54413
rect -8119 -54704 -8085 -54413
rect -7923 -54704 -7889 -54413
rect -13700 -54707 -13205 -54704
rect -11958 -54705 -10505 -54704
rect -13987 -54709 -12883 -54707
rect -11958 -54709 -10192 -54705
rect -9258 -54709 -7880 -54704
rect -13987 -54772 -7880 -54709
rect -13987 -54775 -12883 -54772
rect -10665 -54773 -10192 -54772
rect -28644 -57134 -28236 -57100
rect -27389 -57237 -27341 -57057
rect -27269 -57237 -27203 -57057
rect -27389 -57250 -27203 -57237
rect -27836 -57284 -27203 -57250
rect -27389 -57296 -27203 -57284
rect -28644 -57370 -28236 -57336
rect -27389 -57466 -27341 -57296
rect -27269 -57466 -27203 -57296
rect -27389 -57486 -27203 -57466
rect -27836 -57520 -27203 -57486
rect -27389 -57525 -27203 -57520
rect -28644 -57606 -28236 -57572
rect -27389 -57722 -27341 -57525
rect -27836 -57756 -27341 -57722
rect -27389 -57958 -27341 -57756
rect -27836 -57992 -27341 -57958
rect -27389 -58072 -27341 -57992
rect -27269 -58072 -27203 -57525
rect -27389 -58088 -27203 -58072
rect -27836 -58122 -27203 -58088
rect -27389 -58131 -27203 -58122
rect -27389 -58304 -27341 -58131
rect -27269 -58304 -27203 -58131
rect -27389 -58324 -27203 -58304
rect -27836 -58358 -27203 -58324
rect -27389 -58363 -27203 -58358
rect -27389 -58545 -27341 -58363
rect -27269 -58545 -27203 -58363
rect -27389 -58560 -27203 -58545
rect -27836 -58594 -27203 -58560
rect -27389 -58604 -27203 -58594
rect -27389 -58796 -27341 -58604
rect -27836 -58816 -27341 -58796
rect -27269 -58816 -27203 -58604
rect -27836 -58830 -27203 -58816
rect -27389 -58875 -27203 -58830
rect -27389 -59032 -27341 -58875
rect -27836 -59066 -27341 -59032
rect -27389 -59162 -27341 -59066
rect -27836 -59196 -27341 -59162
rect -27389 -59398 -27341 -59196
rect -27836 -59404 -27341 -59398
rect -27269 -59404 -27203 -58875
rect -27836 -59432 -27203 -59404
rect -27389 -59463 -27203 -59432
rect -27389 -59634 -27341 -59463
rect -27836 -59668 -27341 -59634
rect -27269 -59664 -27203 -59463
rect -13525 -56471 -13372 -54775
rect -12745 -55756 -12674 -55755
rect -12333 -55756 -12259 -55750
rect -12745 -55757 -12259 -55756
rect -12971 -55795 -12259 -55757
rect -12971 -55797 -12744 -55795
rect -12333 -55821 -12259 -55795
rect -12713 -56359 -12679 -55942
rect -12517 -56359 -12483 -55942
rect -12321 -56309 -12287 -55942
rect -12104 -56309 -12070 -56143
rect -11908 -56309 -11874 -56143
rect -11712 -56309 -11678 -56143
rect -11516 -56309 -11482 -56143
rect -12321 -56359 -11434 -56309
rect -11266 -56321 -11232 -55731
rect -12723 -56408 -11434 -56359
rect -12723 -56423 -12281 -56408
rect -11271 -56447 -11226 -56321
rect -11070 -56324 -11036 -55731
rect -11076 -56447 -11031 -56324
rect -10647 -56323 -10613 -55731
rect -10654 -56447 -10609 -56323
rect -12284 -56464 -12095 -56457
rect -12321 -56471 -12095 -56464
rect -11277 -56471 -10508 -56447
rect -13525 -56513 -10508 -56471
rect -13525 -56624 -10612 -56513
rect -13525 -57871 -13372 -56624
rect -12553 -56814 -12381 -56624
rect -11725 -56641 -11107 -56624
rect -11725 -56670 -11282 -56641
rect -11724 -56684 -11282 -56670
rect -11724 -56733 -10435 -56684
rect -12735 -56913 -12017 -56814
rect -12687 -57179 -12653 -56913
rect -12491 -57179 -12457 -56913
rect -12295 -57179 -12261 -56913
rect -12099 -57179 -12065 -56913
rect -11714 -57150 -11680 -56733
rect -11518 -57150 -11484 -56733
rect -11322 -56783 -10435 -56733
rect -11322 -57150 -11288 -56783
rect -11105 -56949 -11071 -56783
rect -10909 -56949 -10875 -56783
rect -10713 -56949 -10679 -56783
rect -10517 -56949 -10483 -56783
rect -5268 -53197 -4216 -53090
rect -5268 -53326 -5228 -53197
rect -5268 -53509 -5234 -53326
rect -5079 -53326 -5033 -53197
rect -5072 -53509 -5038 -53326
rect -4881 -53322 -4835 -53197
rect -4876 -53509 -4842 -53322
rect -4768 -53326 -4722 -53197
rect -4762 -53509 -4728 -53326
rect -4572 -53321 -4526 -53197
rect -4566 -53509 -4532 -53321
rect -4459 -53331 -4413 -53197
rect -4453 -53509 -4419 -53331
rect -4262 -53319 -4216 -53197
rect -4257 -53509 -4223 -53319
rect -3941 -53927 -3826 -53090
rect -2454 -53128 -1861 -53090
rect -3946 -54063 -3823 -53927
rect -2768 -53197 -1716 -53128
rect -2768 -53326 -2728 -53197
rect -2768 -53509 -2734 -53326
rect -2579 -53326 -2533 -53197
rect -2572 -53509 -2538 -53326
rect -2381 -53322 -2335 -53197
rect -2376 -53509 -2342 -53322
rect -2268 -53326 -2222 -53197
rect -2262 -53509 -2228 -53326
rect -2072 -53321 -2026 -53197
rect -2066 -53509 -2032 -53321
rect -1959 -53331 -1913 -53197
rect -1953 -53509 -1919 -53331
rect -1762 -53319 -1716 -53197
rect -1757 -53509 -1723 -53319
rect -1373 -53962 -1259 -53090
rect 62 -53128 655 -53090
rect -268 -53197 784 -53128
rect -268 -53326 -228 -53197
rect -268 -53509 -234 -53326
rect -79 -53326 -33 -53197
rect -72 -53509 -38 -53326
rect 119 -53322 165 -53197
rect 124 -53509 158 -53322
rect 232 -53326 278 -53197
rect 238 -53509 272 -53326
rect 428 -53321 474 -53197
rect -1379 -54098 -1256 -53962
rect 434 -53509 468 -53321
rect 541 -53331 587 -53197
rect 547 -53509 581 -53331
rect 738 -53319 784 -53197
rect 743 -53509 777 -53319
rect 1109 -53962 1224 -53090
rect 2596 -53128 3189 -53090
rect 5009 -53128 5602 -53090
rect 2232 -53197 3284 -53128
rect 2232 -53326 2272 -53197
rect 2232 -53509 2266 -53326
rect 2421 -53326 2467 -53197
rect 2428 -53509 2462 -53326
rect 2619 -53322 2665 -53197
rect 2624 -53509 2658 -53322
rect 2732 -53326 2778 -53197
rect 2738 -53509 2772 -53326
rect 2928 -53321 2974 -53197
rect 1104 -54098 1227 -53962
rect 2934 -53509 2968 -53321
rect 3041 -53331 3087 -53197
rect 3047 -53509 3081 -53331
rect 3238 -53319 3284 -53197
rect 3243 -53509 3277 -53319
rect 4732 -53197 5784 -53128
rect 4732 -53326 4772 -53197
rect 4732 -53509 4766 -53326
rect 4921 -53326 4967 -53197
rect 4928 -53509 4962 -53326
rect 5119 -53322 5165 -53197
rect 5124 -53509 5158 -53322
rect 5232 -53326 5278 -53197
rect 5238 -53509 5272 -53326
rect 5428 -53321 5474 -53197
rect 4337 -53817 4476 -53763
rect 5434 -53509 5468 -53321
rect 5541 -53331 5587 -53197
rect 5547 -53509 5581 -53331
rect 5738 -53319 5784 -53197
rect 5743 -53509 5777 -53319
rect 5415 -53823 5554 -53769
rect 7732 -53197 8784 -53090
rect 7732 -53326 7772 -53197
rect 7732 -53509 7766 -53326
rect 7921 -53326 7967 -53197
rect 7928 -53509 7962 -53326
rect 8119 -53322 8165 -53197
rect 8124 -53509 8158 -53322
rect 8232 -53326 8278 -53197
rect 8238 -53509 8272 -53326
rect 8428 -53321 8474 -53197
rect 7337 -53817 7476 -53763
rect 8434 -53509 8468 -53321
rect 8541 -53331 8587 -53197
rect 8547 -53509 8581 -53331
rect 8738 -53319 8784 -53197
rect 8743 -53509 8777 -53319
rect 8415 -53823 8554 -53769
rect -5739 -54566 -5551 -54492
rect 1103 -54516 1226 -54515
rect -5607 -54921 -5573 -54630
rect -5411 -54921 -5377 -54630
rect -5215 -54921 -5181 -54630
rect -3947 -54830 -3824 -54694
rect -1380 -54686 -1257 -54550
rect 1103 -54578 1409 -54516
rect -5616 -54989 -5121 -54921
rect -5600 -55379 -5512 -54989
rect -5417 -55379 -5329 -54989
rect -5235 -55379 -5147 -54989
rect -6113 -55382 -5009 -55379
rect -3942 -55382 -3827 -54830
rect -2791 -55382 -2318 -55381
rect -1376 -55382 -1261 -54686
rect 38 -55256 175 -55205
rect -121 -55382 2 -55360
rect -6113 -55445 2 -55382
rect -6113 -55447 -5009 -55445
rect -12881 -57226 -12751 -57209
rect -12707 -57226 -12634 -57213
rect -12881 -57267 -12634 -57226
rect -6113 -57142 -6024 -55447
rect -5826 -55450 -5331 -55447
rect -4084 -55449 -2318 -55445
rect -4084 -55450 -2631 -55449
rect -1384 -55450 2 -55445
rect -5766 -55741 -5732 -55450
rect -5570 -55741 -5536 -55450
rect -5374 -55741 -5340 -55450
rect -4023 -55741 -3989 -55450
rect -3827 -55741 -3793 -55450
rect -3631 -55741 -3597 -55450
rect -3066 -55741 -3032 -55450
rect -2870 -55741 -2836 -55450
rect -2674 -55741 -2640 -55450
rect -1323 -55741 -1289 -55450
rect -1127 -55741 -1093 -55450
rect -931 -55741 -897 -55450
rect -441 -55741 -407 -55450
rect -245 -55741 -211 -55450
rect -121 -55496 2 -55450
rect -49 -55741 -15 -55496
rect -1556 -56064 -1482 -55905
rect -5247 -56187 -5115 -56174
rect -1556 -56187 -1481 -56064
rect -953 -55816 -785 -55805
rect -953 -55874 -750 -55816
rect 38 -55805 77 -55256
rect 173 -55386 296 -55359
rect 1108 -55386 1223 -54578
rect 3151 -55386 3274 -55372
rect 173 -55465 3274 -55386
rect 173 -55466 528 -55465
rect 173 -55495 327 -55466
rect 293 -55758 327 -55495
rect -953 -55879 -785 -55874
rect -71 -55879 97 -55805
rect 38 -56187 77 -55879
rect 489 -55758 523 -55466
rect 1031 -55758 1065 -55465
rect 1227 -55758 1261 -55465
rect 1423 -55758 1457 -55465
rect 1619 -55758 1653 -55465
rect 1978 -55505 2865 -55465
rect 2026 -55671 2060 -55505
rect 2222 -55671 2256 -55505
rect 2418 -55671 2452 -55505
rect 2614 -55671 2648 -55505
rect -5653 -56226 77 -56187
rect -5247 -56234 -5115 -56226
rect -5211 -56713 -5151 -56569
rect -5211 -56775 -4971 -56713
rect -5174 -56776 -4971 -56775
rect -5139 -56787 -4971 -56776
rect -5864 -57142 -5830 -56851
rect -5668 -57142 -5634 -56851
rect -5472 -57142 -5438 -56851
rect -5027 -57142 -4993 -56851
rect -4831 -57142 -4797 -56851
rect -4635 -57142 -4601 -56851
rect -3164 -57142 -3130 -56851
rect -2968 -57142 -2934 -56851
rect -2772 -57142 -2738 -56851
rect -2327 -57142 -2293 -56851
rect -2131 -57142 -2097 -56851
rect -1935 -57142 -1901 -56851
rect 2831 -55872 2865 -55505
rect 3027 -55872 3061 -55465
rect 3151 -55508 3274 -55465
rect 3223 -55872 3257 -55508
rect 3540 -55408 3663 -55371
rect 4768 -55393 4891 -55348
rect 4430 -55408 4891 -55393
rect 3540 -55457 4891 -55408
rect 3540 -55507 4470 -55457
rect 3631 -55673 3665 -55507
rect 3827 -55673 3861 -55507
rect 4023 -55673 4057 -55507
rect 4219 -55673 4253 -55507
rect 4436 -55874 4470 -55507
rect 4632 -55874 4666 -55457
rect 4768 -55484 4891 -55457
rect 4828 -55874 4862 -55484
rect 5169 -55379 5292 -55346
rect 5169 -55384 6065 -55379
rect 6525 -55384 6648 -55351
rect 5169 -55452 6648 -55384
rect 5169 -55457 5490 -55452
rect 5993 -55453 6648 -55452
rect 5169 -55482 5292 -55457
rect 5255 -55749 5289 -55482
rect 5451 -55749 5485 -55457
rect 5993 -55749 6027 -55453
rect 6189 -55749 6223 -55453
rect 6385 -55749 6419 -55453
rect 6525 -55487 6648 -55453
rect 6581 -55749 6615 -55487
rect 7741 -55379 7864 -55352
rect 7741 -55448 8794 -55379
rect 7741 -55488 7864 -55448
rect 7742 -55577 7782 -55488
rect 7742 -55760 7776 -55577
rect 7931 -55577 7977 -55448
rect 7938 -55760 7972 -55577
rect 8129 -55573 8175 -55448
rect 8134 -55760 8168 -55573
rect 8242 -55577 8288 -55448
rect 8248 -55760 8282 -55577
rect 8438 -55572 8484 -55448
rect 7347 -56068 7486 -56014
rect 8444 -55760 8478 -55572
rect 8551 -55582 8597 -55448
rect 8557 -55760 8591 -55582
rect 8748 -55570 8794 -55448
rect 8753 -55760 8787 -55570
rect 8425 -56074 8564 -56020
rect 16668 -54816 16903 -54793
rect 11260 -55061 16903 -54816
rect 11260 -55063 16779 -55061
rect 26626 -53252 27729 -51863
rect 18439 -54996 18657 -54750
rect 18478 -55853 18620 -54996
rect 26680 -54856 27010 -54773
rect 26680 -55035 27859 -54856
rect 26680 -55067 27010 -55035
rect 29247 -55389 29382 -55381
rect 29227 -55391 29382 -55389
rect 29020 -55427 29382 -55391
rect 29227 -55429 29382 -55427
rect 29247 -55435 29382 -55429
rect 20974 -55714 26199 -55651
rect 21926 -55719 23728 -55714
rect 24626 -55719 26199 -55714
rect 28359 -55715 28393 -55449
rect 28555 -55715 28589 -55449
rect 28751 -55715 28785 -55449
rect 28947 -55715 28981 -55449
rect 18441 -56042 18620 -55853
rect -6113 -57147 -4540 -57142
rect -3642 -57147 -1840 -57142
rect -6113 -57210 -888 -57147
rect -12881 -57359 -12751 -57267
rect -12707 -57273 -12634 -57267
rect -6113 -57849 -6024 -57210
rect -9909 -57871 -6024 -57849
rect -13987 -57934 -6024 -57871
rect -13987 -57939 -12414 -57934
rect -11516 -57939 -9714 -57934
rect -13987 -58564 -13898 -57939
rect -13738 -58230 -13704 -57939
rect -13542 -58230 -13508 -57939
rect -13346 -58230 -13312 -57939
rect -12901 -58230 -12867 -57939
rect -12705 -58230 -12671 -57939
rect -12509 -58230 -12475 -57939
rect -21534 -58731 -13897 -58564
rect -21164 -58870 -20382 -58731
rect -20006 -58857 -19488 -58731
rect -21224 -59003 -20356 -58870
rect -20021 -58926 -19467 -58857
rect -19117 -58858 -18564 -58731
rect -19117 -58899 -18562 -58858
rect -21224 -59115 -21171 -59003
rect -22483 -59822 -22423 -59641
rect -21215 -59715 -21181 -59115
rect -21028 -59131 -20975 -59003
rect -20016 -59053 -19968 -58926
rect -21019 -59715 -20985 -59131
rect -20009 -59444 -19975 -59053
rect -19819 -59059 -19771 -58926
rect -19116 -58927 -18562 -58899
rect -20189 -59560 -20131 -59465
rect -19813 -59444 -19779 -59059
rect -19111 -59054 -19063 -58927
rect -19782 -59560 -19639 -59553
rect -20189 -59596 -19639 -59560
rect -20189 -59602 -20131 -59596
rect -19782 -59613 -19639 -59596
rect -19104 -59445 -19070 -59054
rect -18914 -59060 -18866 -58927
rect -18908 -59445 -18874 -59060
rect -22483 -59863 -20594 -59822
rect -22483 -59878 -22423 -59863
rect -20654 -59868 -20594 -59863
rect -22292 -59911 -22232 -59898
rect -20974 -59911 -20829 -59900
rect -22292 -59952 -20829 -59911
rect -20654 -59924 -20509 -59868
rect -22292 -60135 -22232 -59952
rect -20974 -59956 -20829 -59952
rect -22182 -60003 -22122 -60001
rect -21303 -60003 -21158 -59995
rect -22182 -60044 -21158 -60003
rect -22182 -60238 -22122 -60044
rect -21303 -60051 -21158 -60044
rect -17702 -60383 -17668 -59966
rect -17506 -60383 -17472 -59966
rect -17310 -60333 -17276 -59966
rect -17093 -60333 -17059 -60167
rect -16897 -60333 -16863 -60167
rect -16701 -60333 -16667 -60167
rect -16505 -60333 -16471 -60167
rect -17310 -60383 -16423 -60333
rect -16255 -60345 -16221 -59755
rect -17712 -60432 -16423 -60383
rect -17712 -60447 -17270 -60432
rect -16260 -60471 -16215 -60345
rect -16059 -60348 -16025 -59755
rect -16065 -60471 -16020 -60348
rect -15636 -60347 -15602 -59755
rect -13987 -59634 -13898 -58731
rect -11038 -58230 -11004 -57939
rect -10842 -58230 -10808 -57939
rect -10646 -58230 -10612 -57939
rect -10201 -58230 -10167 -57939
rect -10005 -58230 -9971 -57939
rect -9809 -58230 -9775 -57939
rect -7353 -58055 -7308 -57934
rect -7349 -58647 -7315 -58055
rect -6931 -58054 -6886 -57934
rect -6926 -58647 -6892 -58054
rect -6736 -58057 -6691 -57934
rect -6113 -58049 -6024 -57934
rect -6730 -58647 -6696 -58057
rect -6113 -58138 -6023 -58049
rect -5825 -58138 -5556 -57210
rect -5279 -58138 -5010 -57210
rect -4402 -58138 -4133 -57210
rect -3540 -58138 -3271 -57210
rect -2637 -58138 -2368 -57210
rect -1606 -58138 -1337 -57210
rect 18780 -57200 18814 -56600
rect 18771 -57312 18824 -57200
rect 18976 -57184 19010 -56600
rect 18967 -57312 19020 -57184
rect 18771 -57445 19639 -57312
rect -6113 -58201 -888 -58138
rect -6113 -58206 -4540 -58201
rect -3642 -58206 -1840 -58201
rect -13640 -59631 -13606 -59340
rect -13444 -59631 -13410 -59340
rect -13248 -59631 -13214 -59340
rect -11897 -59631 -11863 -59340
rect -11701 -59631 -11667 -59340
rect -11505 -59631 -11471 -59340
rect -10940 -59631 -10906 -59340
rect -10744 -59631 -10710 -59340
rect -10548 -59631 -10514 -59340
rect -9197 -59631 -9163 -59340
rect -9001 -59631 -8967 -59340
rect -8805 -59631 -8771 -59340
rect -8315 -59631 -8281 -59340
rect -8119 -59631 -8085 -59340
rect -7923 -59631 -7889 -59340
rect -13700 -59634 -13205 -59631
rect -11958 -59632 -10505 -59631
rect -13987 -59636 -12883 -59634
rect -11958 -59636 -10192 -59632
rect -9258 -59636 -7880 -59631
rect -13987 -59699 -7880 -59636
rect -15643 -60471 -15598 -60347
rect -17273 -60488 -17084 -60481
rect -22084 -60607 -22026 -60511
rect -17310 -60495 -17084 -60488
rect -16266 -60495 -15497 -60471
rect -20209 -60607 -20151 -60511
rect -18946 -60537 -15497 -60495
rect -22084 -60648 -20151 -60607
rect -18946 -60648 -15601 -60537
rect -18946 -60667 -17370 -60648
rect -21552 -62217 -21518 -61925
rect -18946 -61662 -18774 -60667
rect -17542 -60838 -17370 -60667
rect -16714 -60665 -16096 -60648
rect -16714 -60694 -16271 -60665
rect -16713 -60708 -16271 -60694
rect -16713 -60757 -15424 -60708
rect -17724 -60937 -17006 -60838
rect -17676 -61203 -17642 -60937
rect -17480 -61203 -17446 -60937
rect -17284 -61203 -17250 -60937
rect -17088 -61203 -17054 -60937
rect -16703 -61174 -16669 -60757
rect -16507 -61174 -16473 -60757
rect -16311 -60807 -15424 -60757
rect -16311 -61174 -16277 -60807
rect -16094 -60973 -16060 -60807
rect -15898 -60973 -15864 -60807
rect -15702 -60973 -15668 -60807
rect -15506 -60973 -15472 -60807
rect -13987 -59702 -12883 -59699
rect -10665 -59700 -10192 -59699
rect -6113 -59901 -6024 -58206
rect -5864 -58497 -5830 -58206
rect -5668 -58497 -5634 -58206
rect -5472 -58497 -5438 -58206
rect -5027 -58497 -4993 -58206
rect -4831 -58497 -4797 -58206
rect -4635 -58497 -4601 -58206
rect -3164 -58497 -3130 -58206
rect -2968 -58497 -2934 -58206
rect -2772 -58497 -2738 -58206
rect -2327 -58497 -2293 -58206
rect -2131 -58497 -2097 -58206
rect -1935 -58497 -1901 -58206
rect -2439 -58572 -2271 -58561
rect -2499 -58635 -2271 -58572
rect -2499 -58794 -2439 -58635
rect -3474 -59036 -3337 -59025
rect -2528 -59036 -2396 -59026
rect -5653 -59075 77 -59036
rect -3474 -59085 -3337 -59075
rect -2528 -59086 -2396 -59075
rect -5766 -59898 -5732 -59607
rect -5570 -59898 -5536 -59607
rect -5374 -59898 -5340 -59607
rect -3653 -59474 -3485 -59469
rect -3425 -59474 -3365 -59401
rect -3653 -59532 -3365 -59474
rect -3653 -59543 -3485 -59532
rect -3425 -59533 -3365 -59532
rect -4023 -59898 -3989 -59607
rect -3827 -59898 -3793 -59607
rect -3631 -59898 -3597 -59607
rect -3066 -59898 -3032 -59607
rect -2870 -59898 -2836 -59607
rect -2674 -59898 -2640 -59607
rect 38 -59469 77 -59075
rect -71 -59543 97 -59469
rect -1323 -59898 -1289 -59607
rect -1127 -59898 -1093 -59607
rect -931 -59898 -897 -59607
rect -441 -59898 -407 -59607
rect -245 -59898 -211 -59607
rect -49 -59852 -15 -59607
rect -121 -59898 2 -59852
rect -5826 -59901 -5331 -59898
rect -4084 -59899 -2631 -59898
rect -6113 -59903 -5009 -59901
rect -4084 -59903 -2318 -59899
rect -1384 -59903 2 -59898
rect -6113 -59966 2 -59903
rect -6113 -59969 -5009 -59966
rect -18948 -61749 -18772 -61662
rect -3942 -60518 -3827 -59966
rect -2791 -59967 -2318 -59966
rect -3947 -60654 -3824 -60518
rect -1376 -60662 -1261 -59966
rect -121 -59988 2 -59966
rect 38 -60092 77 -59543
rect 293 -59853 327 -59590
rect 173 -59882 327 -59853
rect 489 -59882 523 -59590
rect 173 -59883 528 -59882
rect 1031 -59883 1065 -59590
rect 1227 -59883 1261 -59590
rect 1423 -59883 1457 -59590
rect 1619 -59883 1653 -59590
rect 2026 -59843 2060 -59677
rect 2222 -59843 2256 -59677
rect 2418 -59843 2452 -59677
rect 2614 -59843 2648 -59677
rect 2831 -59843 2865 -59476
rect 1978 -59883 2865 -59843
rect 3027 -59883 3061 -59476
rect 3223 -59840 3257 -59476
rect 3151 -59883 3274 -59840
rect 173 -59962 3274 -59883
rect 173 -59989 296 -59962
rect 38 -60143 175 -60092
rect -1380 -60798 -1257 -60662
rect 1108 -60770 1223 -59962
rect 3151 -59976 3274 -59962
rect 3631 -59841 3665 -59675
rect 3827 -59841 3861 -59675
rect 4023 -59841 4057 -59675
rect 4219 -59841 4253 -59675
rect 4436 -59841 4470 -59474
rect 3540 -59891 4470 -59841
rect 4632 -59891 4666 -59474
rect 4828 -59864 4862 -59474
rect 4768 -59891 4891 -59864
rect 3540 -59940 4891 -59891
rect 3540 -59977 3663 -59940
rect 4430 -59955 4891 -59940
rect 4768 -60000 4891 -59955
rect 1103 -60832 1409 -60770
rect 1103 -60833 1226 -60832
rect 5255 -59866 5289 -59599
rect 20009 -56214 20141 -56079
rect 20009 -56549 20115 -56214
rect 21987 -56010 22021 -55719
rect 22183 -56010 22217 -55719
rect 22379 -56010 22413 -55719
rect 22824 -56010 22858 -55719
rect 23020 -56010 23054 -55719
rect 23216 -56010 23250 -55719
rect 22357 -56085 22525 -56074
rect 22357 -56148 22585 -56085
rect 22525 -56307 22585 -56148
rect 24687 -56010 24721 -55719
rect 24883 -56010 24917 -55719
rect 25079 -56010 25113 -55719
rect 25524 -56010 25558 -55719
rect 25720 -56010 25754 -55719
rect 25916 -56010 25950 -55719
rect 26110 -55779 26199 -55719
rect 28311 -55779 29029 -55715
rect 26110 -55814 29029 -55779
rect 26110 -56004 28665 -55814
rect 29332 -55895 29366 -55478
rect 29528 -55895 29562 -55478
rect 29724 -55845 29758 -55478
rect 29941 -55845 29975 -55679
rect 30137 -55845 30171 -55679
rect 30333 -55845 30367 -55679
rect 30529 -55845 30563 -55679
rect 29724 -55895 30611 -55845
rect 29322 -55944 30611 -55895
rect 29322 -55958 29764 -55944
rect 29321 -55987 29764 -55958
rect 29321 -56004 29939 -55987
rect 26110 -56073 30434 -56004
rect 22482 -56549 22614 -56539
rect 23423 -56549 23560 -56538
rect 20009 -56588 25739 -56549
rect 20009 -56982 20048 -56588
rect 22482 -56599 22614 -56588
rect 23423 -56598 23560 -56588
rect 19989 -57056 20157 -56982
rect 20101 -57411 20135 -57120
rect 20297 -57411 20331 -57120
rect 20493 -57411 20527 -57120
rect 20983 -57411 21017 -57120
rect 21179 -57411 21213 -57120
rect 21375 -57411 21409 -57120
rect 23451 -56987 23511 -56914
rect 23571 -56987 23739 -56982
rect 23451 -57045 23739 -56987
rect 23451 -57046 23511 -57045
rect 22726 -57411 22760 -57120
rect 22922 -57411 22956 -57120
rect 23118 -57411 23152 -57120
rect 23571 -57056 23739 -57045
rect 23683 -57411 23717 -57120
rect 23879 -57411 23913 -57120
rect 24075 -57411 24109 -57120
rect 25426 -57411 25460 -57120
rect 25622 -57411 25656 -57120
rect 25818 -57411 25852 -57120
rect 20092 -57416 21470 -57411
rect 22717 -57412 24170 -57411
rect 22404 -57416 24170 -57412
rect 25417 -57414 25912 -57411
rect 26110 -57414 26199 -56073
rect 28323 -56115 30434 -56073
rect 28323 -56122 30538 -56115
rect 30611 -56122 30673 -56094
rect 28323 -56157 30673 -56122
rect 28725 -56164 28951 -56157
rect 28762 -56171 28951 -56164
rect 29769 -56174 30673 -56157
rect 29769 -56181 30538 -56174
rect 28323 -56220 28765 -56205
rect 28323 -56269 29612 -56220
rect 27599 -56626 27858 -56583
rect 26733 -56737 27858 -56626
rect 28333 -56686 28367 -56269
rect 28529 -56686 28563 -56269
rect 28725 -56319 29612 -56269
rect 29775 -56307 29820 -56181
rect 28725 -56686 28759 -56319
rect 28942 -56485 28976 -56319
rect 29138 -56485 29172 -56319
rect 29334 -56485 29368 -56319
rect 29530 -56485 29564 -56319
rect 28248 -56735 28383 -56729
rect 28228 -56737 28383 -56735
rect 26733 -56773 28383 -56737
rect 26733 -56831 27858 -56773
rect 28228 -56775 28383 -56773
rect 28248 -56783 28383 -56775
rect 27599 -56846 27858 -56831
rect 25095 -57416 26199 -57414
rect 20092 -57479 26199 -57416
rect 22404 -57480 22877 -57479
rect 22594 -57699 22826 -57480
rect 25095 -57482 26199 -57479
rect 22536 -57763 22978 -57699
rect 22546 -58280 22580 -57763
rect 22742 -58280 22776 -57763
rect 22938 -58280 22972 -57763
rect 7347 -59334 7486 -59280
rect 5169 -59891 5292 -59866
rect 5451 -59891 5485 -59599
rect 5169 -59896 5490 -59891
rect 5993 -59895 6027 -59599
rect 6189 -59895 6223 -59599
rect 6385 -59895 6419 -59599
rect 6581 -59861 6615 -59599
rect 6525 -59895 6648 -59861
rect 5993 -59896 6648 -59895
rect 5169 -59964 6648 -59896
rect 5169 -59969 6065 -59964
rect 5169 -60002 5292 -59969
rect 6525 -59997 6648 -59964
rect 7742 -59771 7776 -59588
rect 7742 -59860 7782 -59771
rect 7938 -59771 7972 -59588
rect 7741 -59900 7864 -59860
rect 7931 -59900 7977 -59771
rect 8134 -59775 8168 -59588
rect 8248 -59771 8282 -59588
rect 8425 -59328 8564 -59274
rect 8129 -59900 8175 -59775
rect 8242 -59900 8288 -59771
rect 8444 -59776 8478 -59588
rect 8557 -59766 8591 -59588
rect 8438 -59900 8484 -59776
rect 8551 -59900 8597 -59766
rect 8753 -59778 8787 -59588
rect 8748 -59900 8794 -59778
rect 7741 -59969 8794 -59900
rect 7741 -59996 7864 -59969
rect 9536 -59339 9681 -59204
rect 9253 -60354 9376 -60353
rect -5663 -61585 -5524 -61531
rect -21356 -62201 -21322 -61925
rect -20814 -62201 -20780 -61925
rect -20618 -62201 -20584 -61925
rect -20422 -62201 -20388 -61925
rect -20226 -62201 -20192 -61925
rect -5268 -62022 -5234 -61839
rect -5268 -62151 -5228 -62022
rect -5072 -62022 -5038 -61839
rect -5079 -62151 -5033 -62022
rect -4876 -62026 -4842 -61839
rect -4762 -62022 -4728 -61839
rect -4585 -61579 -4446 -61525
rect -3946 -61421 -3823 -61285
rect -4881 -62151 -4835 -62026
rect -4768 -62151 -4722 -62022
rect -4566 -62027 -4532 -61839
rect -4453 -62017 -4419 -61839
rect -4572 -62151 -4526 -62027
rect -4459 -62151 -4413 -62017
rect -4257 -62029 -4223 -61839
rect -4262 -62151 -4216 -62029
rect -21374 -62217 -18772 -62201
rect -21562 -62284 -18772 -62217
rect -21374 -62293 -18772 -62284
rect -5268 -62258 -4216 -62151
rect -3941 -62258 -3826 -61421
rect -2768 -62022 -2734 -61839
rect -2768 -62151 -2728 -62022
rect -2572 -62022 -2538 -61839
rect -2579 -62151 -2533 -62022
rect -2376 -62026 -2342 -61839
rect -2262 -62022 -2228 -61839
rect -1379 -61386 -1256 -61250
rect -2381 -62151 -2335 -62026
rect -2268 -62151 -2222 -62022
rect -2066 -62027 -2032 -61839
rect -1953 -62017 -1919 -61839
rect -2072 -62151 -2026 -62027
rect -1959 -62151 -1913 -62017
rect -1757 -62029 -1723 -61839
rect -1762 -62151 -1716 -62029
rect -2768 -62220 -1716 -62151
rect -2454 -62258 -1861 -62220
rect -1373 -62258 -1259 -61386
rect -268 -62022 -234 -61839
rect -268 -62151 -228 -62022
rect -72 -62022 -38 -61839
rect -79 -62151 -33 -62022
rect 124 -62026 158 -61839
rect 238 -62022 272 -61839
rect 1104 -61386 1227 -61250
rect 119 -62151 165 -62026
rect 232 -62151 278 -62022
rect 434 -62027 468 -61839
rect 547 -62017 581 -61839
rect 428 -62151 474 -62027
rect 541 -62151 587 -62017
rect 743 -62029 777 -61839
rect 738 -62151 784 -62029
rect -268 -62220 784 -62151
rect 62 -62258 655 -62220
rect 1109 -62258 1224 -61386
rect 2232 -62022 2266 -61839
rect 2232 -62151 2272 -62022
rect 2428 -62022 2462 -61839
rect 2421 -62151 2467 -62022
rect 2624 -62026 2658 -61839
rect 2738 -62022 2772 -61839
rect 2619 -62151 2665 -62026
rect 2732 -62151 2778 -62022
rect 2934 -62027 2968 -61839
rect 3047 -62017 3081 -61839
rect 4337 -61585 4476 -61531
rect 2928 -62151 2974 -62027
rect 3041 -62151 3087 -62017
rect 3243 -62029 3277 -61839
rect 3238 -62151 3284 -62029
rect 2232 -62220 3284 -62151
rect 4732 -62022 4766 -61839
rect 4732 -62151 4772 -62022
rect 4928 -62022 4962 -61839
rect 4921 -62151 4967 -62022
rect 5124 -62026 5158 -61839
rect 5238 -62022 5272 -61839
rect 5415 -61579 5554 -61525
rect 9252 -60397 9376 -60354
rect 5119 -62151 5165 -62026
rect 5232 -62151 5278 -62022
rect 5434 -62027 5468 -61839
rect 5547 -62017 5581 -61839
rect 9252 -61205 9310 -60397
rect 9396 -60955 9519 -60911
rect 7337 -61585 7476 -61531
rect 5428 -62151 5474 -62027
rect 5541 -62151 5587 -62017
rect 5743 -62029 5777 -61839
rect 5738 -62151 5784 -62029
rect 4732 -62220 5784 -62151
rect 7732 -62022 7766 -61839
rect 7732 -62151 7772 -62022
rect 7928 -62022 7962 -61839
rect 7921 -62151 7967 -62022
rect 8124 -62026 8158 -61839
rect 8238 -62022 8272 -61839
rect 8415 -61579 8554 -61525
rect 8119 -62151 8165 -62026
rect 8232 -62151 8278 -62022
rect 8434 -62027 8468 -61839
rect 8547 -62017 8581 -61839
rect 8428 -62151 8474 -62027
rect 8541 -62151 8587 -62017
rect 8743 -62029 8777 -61839
rect 8738 -62151 8784 -62029
rect 2596 -62258 3189 -62220
rect 5009 -62258 5602 -62220
rect 7732 -62258 8784 -62151
rect -6133 -62451 8829 -62258
rect 9253 -62615 9309 -61205
rect 9352 -61583 9417 -61446
rect 9355 -62343 9409 -61583
rect 9460 -62343 9514 -60955
rect 9559 -62560 9615 -59339
rect 18775 -59537 18809 -59146
rect 18768 -59664 18816 -59537
rect 18971 -59531 19005 -59146
rect 18965 -59664 19013 -59531
rect 19721 -59537 19755 -59146
rect 19714 -59664 19762 -59537
rect 19917 -59531 19951 -59146
rect 19911 -59664 19959 -59531
rect 20392 -59664 20478 -59656
rect 17945 -59676 20478 -59664
rect 20637 -59676 20671 -59380
rect 20833 -59676 20867 -59380
rect 21029 -59676 21063 -59380
rect 21225 -59676 21259 -59380
rect 21512 -59672 21575 -59658
rect 21767 -59672 21801 -59380
rect 21963 -59672 21997 -59380
rect 22193 -59664 22267 -59658
rect 22496 -59664 22530 -59373
rect 22692 -59664 22726 -59373
rect 22888 -59637 22922 -59373
rect 23376 -59637 23410 -58802
rect 23572 -59637 23606 -58802
rect 23776 -59637 23810 -58802
rect 23972 -59637 24006 -58802
rect 24376 -59637 24410 -58802
rect 24572 -59637 24606 -58802
rect 24776 -59637 24810 -58802
rect 24972 -59637 25006 -58802
rect 25376 -59637 25410 -58802
rect 25572 -59637 25606 -58802
rect 25776 -59637 25810 -58802
rect 25972 -59637 26006 -58802
rect 26110 -59637 26199 -57482
rect 29780 -56897 29814 -56307
rect 29970 -56304 30015 -56181
rect 29976 -56897 30010 -56304
rect 30392 -56305 30437 -56181
rect 30611 -56188 30673 -56174
rect 30399 -56897 30433 -56305
rect 36799 -55726 36833 -55460
rect 36995 -55726 37029 -55460
rect 37191 -55726 37225 -55460
rect 37387 -55726 37421 -55460
rect 36751 -55825 37469 -55726
rect 31769 -55950 34201 -55880
rect 31402 -56002 34201 -55950
rect 31402 -56003 33155 -56002
rect 31402 -56067 31807 -56003
rect 30839 -56077 30937 -56074
rect 31402 -56077 31519 -56067
rect 30839 -56194 31519 -56077
rect 31769 -56162 31807 -56067
rect 30839 -56200 30937 -56194
rect 31772 -56655 31806 -56162
rect 31966 -56160 32004 -56003
rect 31968 -56655 32002 -56160
rect 32558 -56183 32608 -56003
rect 32684 -56180 32734 -56003
rect 32563 -56655 32597 -56183
rect 32693 -56655 32727 -56180
rect 32915 -56165 32958 -56003
rect 32921 -56455 32955 -56165
rect 33112 -56163 33155 -56003
rect 34079 -56015 34201 -56002
rect 36933 -56015 37105 -55825
rect 37772 -55906 37806 -55489
rect 37968 -55906 38002 -55489
rect 38164 -55856 38198 -55489
rect 38381 -55856 38415 -55690
rect 38577 -55856 38611 -55690
rect 38773 -55856 38807 -55690
rect 38969 -55856 39003 -55690
rect 38164 -55906 39051 -55856
rect 37762 -55955 39051 -55906
rect 37762 -55969 38204 -55955
rect 37761 -55998 38204 -55969
rect 37761 -56015 38379 -55998
rect 34079 -56126 38874 -56015
rect 34079 -56133 38978 -56126
rect 39051 -56133 39113 -56105
rect 33117 -56455 33151 -56163
rect 34079 -56168 39113 -56133
rect 22888 -59664 26199 -59637
rect 22193 -59672 26199 -59664
rect 21512 -59676 26199 -59672
rect 17945 -59732 26199 -59676
rect 17945 -59733 22267 -59732
rect 9830 -60220 10021 -60214
rect 9830 -60303 10393 -60220
rect 9830 -60321 10021 -60303
rect 10310 -62168 10393 -60303
rect 17945 -60204 18071 -59733
rect 20392 -59739 22267 -59733
rect 20392 -59745 21575 -59739
rect 22193 -59745 22267 -59739
rect 22910 -59740 26199 -59732
rect 20392 -59749 20478 -59745
rect 21512 -59756 21575 -59745
rect 14276 -60207 14749 -60206
rect 16967 -60207 18071 -60204
rect 11964 -60270 18071 -60207
rect 11964 -60275 13342 -60270
rect 14276 -60274 16042 -60270
rect 16967 -60272 18071 -60270
rect 14589 -60275 16042 -60274
rect 17289 -60275 17784 -60272
rect 11973 -60566 12007 -60275
rect 12169 -60566 12203 -60275
rect 12365 -60566 12399 -60275
rect 12855 -60566 12889 -60275
rect 13051 -60566 13085 -60275
rect 13247 -60566 13281 -60275
rect 11861 -60704 12029 -60630
rect 11260 -61098 11555 -61000
rect 11881 -61098 11920 -60704
rect 14598 -60566 14632 -60275
rect 14794 -60566 14828 -60275
rect 14990 -60566 15024 -60275
rect 15555 -60566 15589 -60275
rect 15751 -60566 15785 -60275
rect 15947 -60566 15981 -60275
rect 15323 -60641 15383 -60640
rect 15443 -60641 15611 -60630
rect 15323 -60699 15611 -60641
rect 15323 -60772 15383 -60699
rect 15443 -60704 15611 -60699
rect 17298 -60566 17332 -60275
rect 17494 -60566 17528 -60275
rect 17690 -60566 17724 -60275
rect 14354 -61098 14486 -61087
rect 15295 -61098 15432 -61088
rect 11260 -61137 17611 -61098
rect 11260 -61203 11555 -61137
rect 14354 -61147 14486 -61137
rect 15295 -61148 15432 -61137
rect 14397 -61538 14457 -61379
rect 14229 -61601 14457 -61538
rect 14229 -61612 14397 -61601
rect 13859 -61967 13893 -61676
rect 14055 -61967 14089 -61676
rect 14251 -61967 14285 -61676
rect 14696 -61967 14730 -61676
rect 14892 -61967 14926 -61676
rect 15088 -61967 15122 -61676
rect 16559 -61967 16593 -61676
rect 16755 -61967 16789 -61676
rect 16951 -61967 16985 -61676
rect 17396 -61967 17430 -61676
rect 17592 -61967 17626 -61676
rect 17788 -61967 17822 -61676
rect 17982 -61967 18071 -60272
rect 30846 -58192 31248 -58126
rect 28351 -59168 28385 -58902
rect 28547 -59168 28581 -58902
rect 28743 -59168 28777 -58902
rect 28939 -59168 28973 -58902
rect 28303 -59267 29021 -59168
rect 28485 -59457 28657 -59267
rect 29324 -59348 29358 -58931
rect 29520 -59348 29554 -58931
rect 29716 -59298 29750 -58931
rect 29933 -59298 29967 -59132
rect 30129 -59298 30163 -59132
rect 30325 -59298 30359 -59132
rect 30521 -59298 30555 -59132
rect 29716 -59348 30603 -59298
rect 29314 -59397 30603 -59348
rect 29314 -59411 29756 -59397
rect 29313 -59440 29756 -59411
rect 29313 -59457 29931 -59440
rect 28315 -59568 30426 -59457
rect 28315 -59610 30530 -59568
rect 28717 -59617 28943 -59610
rect 28754 -59624 28943 -59617
rect 29761 -59634 30530 -59610
rect 28315 -59673 28757 -59658
rect 28315 -59722 29604 -59673
rect 28325 -60139 28359 -59722
rect 28521 -60139 28555 -59722
rect 28717 -59772 29604 -59722
rect 29767 -59760 29812 -59634
rect 28717 -60139 28751 -59772
rect 28934 -59938 28968 -59772
rect 29130 -59938 29164 -59772
rect 29326 -59938 29360 -59772
rect 29522 -59938 29556 -59772
rect 28240 -60188 28375 -60182
rect 28220 -60190 28375 -60188
rect 27692 -60226 28375 -60190
rect 13798 -61972 15600 -61967
rect 16498 -61972 18071 -61967
rect 12846 -62035 18071 -61972
rect 27875 -61253 28011 -60226
rect 28220 -60228 28375 -60226
rect 28240 -60236 28375 -60228
rect 29772 -60350 29806 -59760
rect 29962 -59757 30007 -59634
rect 29968 -60350 30002 -59757
rect 30384 -59758 30429 -59634
rect 30391 -60350 30425 -59758
rect 30846 -59493 30912 -58192
rect 30829 -59606 30913 -59493
rect 31182 -59522 31248 -58192
rect 34079 -58399 34201 -56168
rect 37165 -56175 37391 -56168
rect 37202 -56182 37391 -56175
rect 38209 -56185 39113 -56168
rect 38209 -56192 38978 -56185
rect 36763 -56231 37205 -56216
rect 36763 -56280 38052 -56231
rect 35600 -56748 36248 -56694
rect 36773 -56697 36807 -56280
rect 36969 -56697 37003 -56280
rect 37165 -56330 38052 -56280
rect 38215 -56318 38260 -56192
rect 37165 -56697 37199 -56330
rect 37382 -56496 37416 -56330
rect 37578 -56496 37612 -56330
rect 37774 -56496 37808 -56330
rect 37970 -56496 38004 -56330
rect 36688 -56746 36823 -56740
rect 36668 -56748 36823 -56746
rect 35600 -56784 36823 -56748
rect 35600 -56840 36248 -56784
rect 36668 -56786 36823 -56784
rect 36688 -56794 36823 -56786
rect 34079 -58521 34711 -58399
rect 32019 -59199 32053 -58933
rect 32215 -59199 32249 -58933
rect 32411 -59199 32445 -58933
rect 32607 -59199 32641 -58933
rect 31971 -59298 32689 -59199
rect 32153 -59488 32325 -59298
rect 32992 -59379 33026 -58962
rect 33188 -59379 33222 -58962
rect 33384 -59329 33418 -58962
rect 33601 -59329 33635 -59163
rect 33797 -59329 33831 -59163
rect 33993 -59329 34027 -59163
rect 34189 -59329 34223 -59163
rect 33384 -59379 34271 -59329
rect 32982 -59428 34271 -59379
rect 32982 -59442 33424 -59428
rect 32981 -59471 33424 -59442
rect 32981 -59488 33599 -59471
rect 31983 -59522 34094 -59488
rect 31182 -59588 34094 -59522
rect 34249 -59563 34328 -59532
rect 31983 -59599 34094 -59588
rect 34149 -59599 34328 -59563
rect 31983 -59641 34328 -59599
rect 32385 -59648 32611 -59641
rect 32422 -59655 32611 -59648
rect 33429 -59646 34328 -59641
rect 33429 -59665 34198 -59646
rect 31983 -59704 32425 -59689
rect 31983 -59753 33272 -59704
rect 31993 -60170 32027 -59753
rect 32189 -60170 32223 -59753
rect 32385 -59803 33272 -59753
rect 33435 -59791 33480 -59665
rect 32385 -60170 32419 -59803
rect 32602 -59969 32636 -59803
rect 32798 -59969 32832 -59803
rect 32994 -59969 33028 -59803
rect 33190 -59969 33224 -59803
rect 31908 -60219 32043 -60213
rect 31888 -60221 32043 -60219
rect 31474 -60257 32043 -60221
rect 31474 -61253 31610 -60257
rect 31888 -60259 32043 -60257
rect 31908 -60267 32043 -60259
rect 33440 -60381 33474 -59791
rect 33630 -59788 33675 -59665
rect 33636 -60381 33670 -59788
rect 34052 -59789 34097 -59665
rect 34249 -59671 34328 -59646
rect 34059 -60381 34093 -59789
rect 34589 -59517 34711 -58521
rect 34499 -59656 34711 -59517
rect 34499 -59684 34638 -59656
rect 27875 -61389 31610 -61253
rect 10286 -62347 10414 -62168
rect 27305 -62403 27526 -62208
rect 27875 -62615 28011 -61389
rect 35600 -62223 35746 -56840
rect 38220 -56908 38254 -56318
rect 38410 -56315 38455 -56192
rect 38416 -56908 38450 -56315
rect 38832 -56316 38877 -56192
rect 39051 -56199 39113 -56185
rect 38839 -56908 38873 -56316
rect 45662 -55765 45696 -55499
rect 45858 -55765 45892 -55499
rect 46054 -55765 46088 -55499
rect 46250 -55765 46284 -55499
rect 45614 -55849 46332 -55765
rect 41581 -55864 46332 -55849
rect 41581 -55891 45968 -55864
rect 40209 -55961 45968 -55891
rect 46635 -55945 46669 -55528
rect 46831 -55945 46865 -55528
rect 47027 -55895 47061 -55528
rect 47244 -55895 47278 -55729
rect 47440 -55895 47474 -55729
rect 47636 -55895 47670 -55729
rect 47832 -55895 47866 -55729
rect 47027 -55945 47914 -55895
rect 39842 -56014 45968 -55961
rect 46625 -55994 47914 -55945
rect 46625 -56008 47067 -55994
rect 39842 -56078 40247 -56014
rect 39279 -56088 39377 -56085
rect 39842 -56088 39959 -56078
rect 39279 -56205 39959 -56088
rect 40209 -56173 40247 -56078
rect 39279 -56211 39377 -56205
rect 40212 -56666 40246 -56173
rect 40406 -56171 40444 -56014
rect 40408 -56666 40442 -56171
rect 40998 -56194 41048 -56014
rect 41124 -56191 41174 -56014
rect 41003 -56666 41037 -56194
rect 41133 -56666 41167 -56191
rect 41355 -56176 41398 -56014
rect 41552 -56054 45968 -56014
rect 46624 -56037 47067 -56008
rect 46624 -56054 47242 -56037
rect 41552 -56103 47737 -56054
rect 41361 -56466 41395 -56176
rect 41552 -56174 41595 -56103
rect 41557 -56466 41591 -56174
rect 39286 -58203 39688 -58137
rect 36791 -59179 36825 -58913
rect 36987 -59179 37021 -58913
rect 37183 -59179 37217 -58913
rect 37379 -59179 37413 -58913
rect 36743 -59278 37461 -59179
rect 36925 -59468 37097 -59278
rect 37764 -59359 37798 -58942
rect 37960 -59359 37994 -58942
rect 38156 -59309 38190 -58942
rect 38373 -59309 38407 -59143
rect 38569 -59309 38603 -59143
rect 38765 -59309 38799 -59143
rect 38961 -59309 38995 -59143
rect 38156 -59359 39043 -59309
rect 37754 -59408 39043 -59359
rect 37754 -59422 38196 -59408
rect 37753 -59451 38196 -59422
rect 37753 -59468 38371 -59451
rect 36755 -59579 38866 -59468
rect 36755 -59621 38970 -59579
rect 37157 -59628 37383 -59621
rect 37194 -59635 37383 -59628
rect 38201 -59645 38970 -59621
rect 36755 -59684 37197 -59669
rect 36755 -59733 38044 -59684
rect 36765 -60150 36799 -59733
rect 36961 -60150 36995 -59733
rect 37157 -59783 38044 -59733
rect 38207 -59771 38252 -59645
rect 37157 -60150 37191 -59783
rect 37374 -59949 37408 -59783
rect 37570 -59949 37604 -59783
rect 37766 -59949 37800 -59783
rect 37962 -59949 37996 -59783
rect 36680 -60199 36815 -60193
rect 36660 -60201 36815 -60199
rect 36132 -60237 36815 -60201
rect 36315 -61264 36451 -60237
rect 36660 -60239 36815 -60237
rect 36680 -60247 36815 -60239
rect 38212 -60361 38246 -59771
rect 38402 -59768 38447 -59645
rect 38408 -60361 38442 -59768
rect 38824 -59769 38869 -59645
rect 38831 -60361 38865 -59769
rect 39286 -59504 39352 -58203
rect 39269 -59617 39353 -59504
rect 39622 -59533 39688 -58203
rect 42519 -58410 42641 -56103
rect 45626 -56165 47737 -56103
rect 45626 -56172 47841 -56165
rect 47914 -56172 47976 -56144
rect 45626 -56207 47976 -56172
rect 46028 -56214 46254 -56207
rect 46065 -56221 46254 -56214
rect 47072 -56224 47976 -56207
rect 47072 -56231 47841 -56224
rect 45626 -56270 46068 -56255
rect 45626 -56319 46915 -56270
rect 45636 -56736 45670 -56319
rect 45832 -56736 45866 -56319
rect 46028 -56369 46915 -56319
rect 47078 -56357 47123 -56231
rect 46028 -56736 46062 -56369
rect 46245 -56535 46279 -56369
rect 46441 -56535 46475 -56369
rect 46637 -56535 46671 -56369
rect 46833 -56535 46867 -56369
rect 44282 -56787 45049 -56780
rect 45551 -56785 45686 -56779
rect 45531 -56787 45686 -56785
rect 44282 -56823 45686 -56787
rect 44282 -56926 45049 -56823
rect 45531 -56825 45686 -56823
rect 45551 -56833 45686 -56825
rect 42519 -58532 43151 -58410
rect 40459 -59210 40493 -58944
rect 40655 -59210 40689 -58944
rect 40851 -59210 40885 -58944
rect 41047 -59210 41081 -58944
rect 40411 -59309 41129 -59210
rect 40593 -59499 40765 -59309
rect 41432 -59390 41466 -58973
rect 41628 -59390 41662 -58973
rect 41824 -59340 41858 -58973
rect 42041 -59340 42075 -59174
rect 42237 -59340 42271 -59174
rect 42433 -59340 42467 -59174
rect 42629 -59340 42663 -59174
rect 41824 -59390 42711 -59340
rect 41422 -59439 42711 -59390
rect 41422 -59453 41864 -59439
rect 41421 -59482 41864 -59453
rect 41421 -59499 42039 -59482
rect 40423 -59533 42534 -59499
rect 39622 -59599 42534 -59533
rect 42689 -59574 42768 -59543
rect 40423 -59610 42534 -59599
rect 42589 -59610 42768 -59574
rect 40423 -59652 42768 -59610
rect 40825 -59659 41051 -59652
rect 40862 -59666 41051 -59659
rect 41869 -59657 42768 -59652
rect 41869 -59676 42638 -59657
rect 40423 -59715 40865 -59700
rect 40423 -59764 41712 -59715
rect 40433 -60181 40467 -59764
rect 40629 -60181 40663 -59764
rect 40825 -59814 41712 -59764
rect 41875 -59802 41920 -59676
rect 40825 -60181 40859 -59814
rect 41042 -59980 41076 -59814
rect 41238 -59980 41272 -59814
rect 41434 -59980 41468 -59814
rect 41630 -59980 41664 -59814
rect 40348 -60230 40483 -60224
rect 40328 -60232 40483 -60230
rect 39914 -60268 40483 -60232
rect 39914 -61264 40050 -60268
rect 40328 -60270 40483 -60268
rect 40348 -60278 40483 -60270
rect 41880 -60392 41914 -59802
rect 42070 -59799 42115 -59676
rect 42076 -60392 42110 -59799
rect 42492 -59800 42537 -59676
rect 42689 -59682 42768 -59657
rect 42499 -60392 42533 -59800
rect 43029 -59528 43151 -58532
rect 42939 -59667 43151 -59528
rect 42939 -59695 43078 -59667
rect 36315 -61400 40050 -61264
rect 35531 -62426 35805 -62223
rect -33062 -62751 28011 -62615
rect 36315 -62814 36451 -61400
rect -33463 -62950 36451 -62814
rect 44282 -62241 44428 -56926
rect 47083 -56947 47117 -56357
rect 47273 -56354 47318 -56231
rect 47279 -56947 47313 -56354
rect 47695 -56355 47740 -56231
rect 47914 -56238 47976 -56224
rect 47702 -56947 47736 -56355
rect 54860 -55731 54894 -55465
rect 55056 -55731 55090 -55465
rect 55252 -55731 55286 -55465
rect 55448 -55731 55482 -55465
rect 54812 -55799 55530 -55731
rect 50432 -55830 55530 -55799
rect 50432 -55930 55166 -55830
rect 55833 -55911 55867 -55494
rect 56029 -55911 56063 -55494
rect 56225 -55861 56259 -55494
rect 56442 -55861 56476 -55695
rect 56638 -55861 56672 -55695
rect 56834 -55861 56868 -55695
rect 57030 -55861 57064 -55695
rect 56225 -55911 57112 -55861
rect 49072 -56000 55166 -55930
rect 55823 -55960 57112 -55911
rect 55823 -55974 56265 -55960
rect 48705 -56020 55166 -56000
rect 55822 -56003 56265 -55974
rect 55822 -56020 56440 -56003
rect 48705 -56053 56935 -56020
rect 48705 -56117 49110 -56053
rect 48142 -56127 48240 -56124
rect 48705 -56127 48822 -56117
rect 48142 -56244 48822 -56127
rect 49072 -56212 49110 -56117
rect 48142 -56250 48240 -56244
rect 49075 -56705 49109 -56212
rect 49269 -56210 49307 -56053
rect 49271 -56705 49305 -56210
rect 49861 -56233 49911 -56053
rect 49987 -56230 50037 -56053
rect 49866 -56705 49900 -56233
rect 49996 -56705 50030 -56230
rect 50218 -56215 50261 -56053
rect 50415 -56113 56935 -56053
rect 50224 -56505 50258 -56215
rect 50415 -56213 50458 -56113
rect 50420 -56505 50454 -56213
rect 48149 -58242 48551 -58176
rect 45654 -59218 45688 -58952
rect 45850 -59218 45884 -58952
rect 46046 -59218 46080 -58952
rect 46242 -59218 46276 -58952
rect 45606 -59317 46324 -59218
rect 45788 -59507 45960 -59317
rect 46627 -59398 46661 -58981
rect 46823 -59398 46857 -58981
rect 47019 -59348 47053 -58981
rect 47236 -59348 47270 -59182
rect 47432 -59348 47466 -59182
rect 47628 -59348 47662 -59182
rect 47824 -59348 47858 -59182
rect 47019 -59398 47906 -59348
rect 46617 -59447 47906 -59398
rect 46617 -59461 47059 -59447
rect 46616 -59490 47059 -59461
rect 46616 -59507 47234 -59490
rect 45618 -59618 47729 -59507
rect 45618 -59660 47833 -59618
rect 46020 -59667 46246 -59660
rect 46057 -59674 46246 -59667
rect 47064 -59684 47833 -59660
rect 45618 -59723 46060 -59708
rect 45618 -59772 46907 -59723
rect 45628 -60189 45662 -59772
rect 45824 -60189 45858 -59772
rect 46020 -59822 46907 -59772
rect 47070 -59810 47115 -59684
rect 46020 -60189 46054 -59822
rect 46237 -59988 46271 -59822
rect 46433 -59988 46467 -59822
rect 46629 -59988 46663 -59822
rect 46825 -59988 46859 -59822
rect 45543 -60238 45678 -60232
rect 45523 -60240 45678 -60238
rect 44995 -60276 45678 -60240
rect 45178 -61289 45314 -60276
rect 45523 -60278 45678 -60276
rect 45543 -60286 45678 -60278
rect 47075 -60400 47109 -59810
rect 47265 -59807 47310 -59684
rect 47271 -60400 47305 -59807
rect 47687 -59808 47732 -59684
rect 47694 -60400 47728 -59808
rect 48149 -59543 48215 -58242
rect 48132 -59656 48216 -59543
rect 48485 -59572 48551 -58242
rect 51382 -58449 51504 -56113
rect 54824 -56131 56935 -56113
rect 54824 -56138 57039 -56131
rect 57112 -56138 57174 -56110
rect 54824 -56173 57174 -56138
rect 55226 -56180 55452 -56173
rect 55263 -56187 55452 -56180
rect 56270 -56190 57174 -56173
rect 56270 -56197 57039 -56190
rect 54824 -56236 55266 -56221
rect 54824 -56285 56113 -56236
rect 53601 -56753 54330 -56688
rect 54834 -56702 54868 -56285
rect 55030 -56702 55064 -56285
rect 55226 -56335 56113 -56285
rect 56276 -56323 56321 -56197
rect 55226 -56702 55260 -56335
rect 55443 -56501 55477 -56335
rect 55639 -56501 55673 -56335
rect 55835 -56501 55869 -56335
rect 56031 -56501 56065 -56335
rect 54749 -56751 54884 -56745
rect 54729 -56753 54884 -56751
rect 53601 -56789 54884 -56753
rect 53601 -56834 54330 -56789
rect 54729 -56791 54884 -56789
rect 54749 -56799 54884 -56791
rect 51382 -58571 52014 -58449
rect 49322 -59249 49356 -58983
rect 49518 -59249 49552 -58983
rect 49714 -59249 49748 -58983
rect 49910 -59249 49944 -58983
rect 49274 -59348 49992 -59249
rect 49456 -59538 49628 -59348
rect 50295 -59429 50329 -59012
rect 50491 -59429 50525 -59012
rect 50687 -59379 50721 -59012
rect 50904 -59379 50938 -59213
rect 51100 -59379 51134 -59213
rect 51296 -59379 51330 -59213
rect 51492 -59379 51526 -59213
rect 50687 -59429 51574 -59379
rect 50285 -59478 51574 -59429
rect 50285 -59492 50727 -59478
rect 50284 -59521 50727 -59492
rect 50284 -59538 50902 -59521
rect 49286 -59572 51397 -59538
rect 48485 -59638 51397 -59572
rect 51552 -59613 51631 -59582
rect 49286 -59649 51397 -59638
rect 51452 -59649 51631 -59613
rect 49286 -59691 51631 -59649
rect 49688 -59698 49914 -59691
rect 49725 -59705 49914 -59698
rect 50732 -59696 51631 -59691
rect 50732 -59715 51501 -59696
rect 49286 -59754 49728 -59739
rect 49286 -59803 50575 -59754
rect 49296 -60220 49330 -59803
rect 49492 -60220 49526 -59803
rect 49688 -59853 50575 -59803
rect 50738 -59841 50783 -59715
rect 49688 -60220 49722 -59853
rect 49905 -60019 49939 -59853
rect 50101 -60019 50135 -59853
rect 50297 -60019 50331 -59853
rect 50493 -60019 50527 -59853
rect 49211 -60269 49346 -60263
rect 49191 -60271 49346 -60269
rect 48777 -60307 49346 -60271
rect 45178 -61303 45361 -61289
rect 48777 -61303 48913 -60307
rect 49191 -60309 49346 -60307
rect 49211 -60317 49346 -60309
rect 50743 -60431 50777 -59841
rect 50933 -59838 50978 -59715
rect 50939 -60431 50973 -59838
rect 51355 -59839 51400 -59715
rect 51552 -59721 51631 -59696
rect 51362 -60431 51396 -59839
rect 51892 -59567 52014 -58571
rect 51802 -59706 52014 -59567
rect 51802 -59734 51941 -59706
rect 45178 -61439 48913 -61303
rect 44228 -62380 44480 -62241
rect 45225 -63047 45361 -61439
rect 53601 -62202 53747 -56834
rect 56281 -56913 56315 -56323
rect 56471 -56320 56516 -56197
rect 56477 -56913 56511 -56320
rect 56893 -56321 56938 -56197
rect 57112 -56204 57174 -56190
rect 56900 -56913 56934 -56321
rect 63614 -55665 63648 -55399
rect 63810 -55665 63844 -55399
rect 64006 -55665 64040 -55399
rect 64202 -55665 64236 -55399
rect 63566 -55702 64284 -55665
rect 59615 -55764 64284 -55702
rect 59615 -55896 63920 -55764
rect 64587 -55845 64621 -55428
rect 64783 -55845 64817 -55428
rect 64979 -55795 65013 -55428
rect 65196 -55795 65230 -55629
rect 65392 -55795 65426 -55629
rect 65588 -55795 65622 -55629
rect 65784 -55795 65818 -55629
rect 64979 -55845 65866 -55795
rect 58270 -55954 63920 -55896
rect 64577 -55894 65866 -55845
rect 64577 -55908 65019 -55894
rect 64576 -55937 65019 -55908
rect 64576 -55954 65194 -55937
rect 58270 -55966 65689 -55954
rect 57903 -56019 65689 -55966
rect 57903 -56083 58308 -56019
rect 57340 -56093 57438 -56090
rect 57903 -56093 58020 -56083
rect 57340 -56210 58020 -56093
rect 58270 -56178 58308 -56083
rect 57340 -56216 57438 -56210
rect 58273 -56671 58307 -56178
rect 58467 -56176 58505 -56019
rect 58469 -56671 58503 -56176
rect 59059 -56199 59109 -56019
rect 59185 -56196 59235 -56019
rect 59064 -56671 59098 -56199
rect 59194 -56671 59228 -56196
rect 59416 -56181 59459 -56019
rect 59613 -56065 65689 -56019
rect 59613 -56072 65793 -56065
rect 65866 -56072 65928 -56044
rect 59613 -56081 65928 -56072
rect 59422 -56471 59456 -56181
rect 59613 -56179 59656 -56081
rect 59618 -56471 59652 -56179
rect 57347 -58208 57749 -58142
rect 54852 -59184 54886 -58918
rect 55048 -59184 55082 -58918
rect 55244 -59184 55278 -58918
rect 55440 -59184 55474 -58918
rect 54804 -59283 55522 -59184
rect 54986 -59473 55158 -59283
rect 55825 -59364 55859 -58947
rect 56021 -59364 56055 -58947
rect 56217 -59314 56251 -58947
rect 56434 -59314 56468 -59148
rect 56630 -59314 56664 -59148
rect 56826 -59314 56860 -59148
rect 57022 -59314 57056 -59148
rect 56217 -59364 57104 -59314
rect 55815 -59413 57104 -59364
rect 55815 -59427 56257 -59413
rect 55814 -59456 56257 -59427
rect 55814 -59473 56432 -59456
rect 54816 -59584 56927 -59473
rect 54816 -59626 57031 -59584
rect 55218 -59633 55444 -59626
rect 55255 -59640 55444 -59633
rect 56262 -59650 57031 -59626
rect 54816 -59689 55258 -59674
rect 54816 -59738 56105 -59689
rect 54826 -60155 54860 -59738
rect 55022 -60155 55056 -59738
rect 55218 -59788 56105 -59738
rect 56268 -59776 56313 -59650
rect 55218 -60155 55252 -59788
rect 55435 -59954 55469 -59788
rect 55631 -59954 55665 -59788
rect 55827 -59954 55861 -59788
rect 56023 -59954 56057 -59788
rect 54741 -60204 54876 -60198
rect 54721 -60206 54876 -60204
rect 54193 -60242 54876 -60206
rect 54376 -61269 54512 -60242
rect 54721 -60244 54876 -60242
rect 54741 -60252 54876 -60244
rect 56273 -60366 56307 -59776
rect 56463 -59773 56508 -59650
rect 56469 -60366 56503 -59773
rect 56885 -59774 56930 -59650
rect 56892 -60366 56926 -59774
rect 57347 -59509 57413 -58208
rect 57330 -59622 57414 -59509
rect 57683 -59538 57749 -58208
rect 60580 -58415 60702 -56081
rect 63578 -56107 65928 -56081
rect 63980 -56114 64206 -56107
rect 64017 -56121 64206 -56114
rect 65024 -56124 65928 -56107
rect 65024 -56131 65793 -56124
rect 63578 -56170 64020 -56155
rect 63578 -56219 64867 -56170
rect 62128 -56687 63054 -56563
rect 63588 -56636 63622 -56219
rect 63784 -56636 63818 -56219
rect 63980 -56269 64867 -56219
rect 65030 -56257 65075 -56131
rect 63980 -56636 64014 -56269
rect 64197 -56435 64231 -56269
rect 64393 -56435 64427 -56269
rect 64589 -56435 64623 -56269
rect 64785 -56435 64819 -56269
rect 63503 -56685 63638 -56679
rect 63483 -56687 63638 -56685
rect 62128 -56723 63638 -56687
rect 62128 -56802 63054 -56723
rect 63483 -56725 63638 -56723
rect 63503 -56733 63638 -56725
rect 60580 -58537 61212 -58415
rect 58520 -59215 58554 -58949
rect 58716 -59215 58750 -58949
rect 58912 -59215 58946 -58949
rect 59108 -59215 59142 -58949
rect 58472 -59314 59190 -59215
rect 58654 -59504 58826 -59314
rect 59493 -59395 59527 -58978
rect 59689 -59395 59723 -58978
rect 59885 -59345 59919 -58978
rect 60102 -59345 60136 -59179
rect 60298 -59345 60332 -59179
rect 60494 -59345 60528 -59179
rect 60690 -59345 60724 -59179
rect 59885 -59395 60772 -59345
rect 59483 -59444 60772 -59395
rect 59483 -59458 59925 -59444
rect 59482 -59487 59925 -59458
rect 59482 -59504 60100 -59487
rect 58484 -59538 60595 -59504
rect 57683 -59604 60595 -59538
rect 60750 -59579 60829 -59548
rect 58484 -59615 60595 -59604
rect 60650 -59615 60829 -59579
rect 58484 -59657 60829 -59615
rect 58886 -59664 59112 -59657
rect 58923 -59671 59112 -59664
rect 59930 -59662 60829 -59657
rect 59930 -59681 60699 -59662
rect 58484 -59720 58926 -59705
rect 58484 -59769 59773 -59720
rect 58494 -60186 58528 -59769
rect 58690 -60186 58724 -59769
rect 58886 -59819 59773 -59769
rect 59936 -59807 59981 -59681
rect 58886 -60186 58920 -59819
rect 59103 -59985 59137 -59819
rect 59299 -59985 59333 -59819
rect 59495 -59985 59529 -59819
rect 59691 -59985 59725 -59819
rect 58409 -60235 58544 -60229
rect 58389 -60237 58544 -60235
rect 57975 -60273 58544 -60237
rect 57975 -61269 58111 -60273
rect 58389 -60275 58544 -60273
rect 58409 -60283 58544 -60275
rect 59941 -60397 59975 -59807
rect 60131 -59804 60176 -59681
rect 60137 -60397 60171 -59804
rect 60553 -59805 60598 -59681
rect 60750 -59687 60829 -59662
rect 60560 -60397 60594 -59805
rect 61090 -59533 61212 -58537
rect 61000 -59672 61212 -59533
rect 61000 -59700 61139 -59672
rect 54376 -61405 58111 -61269
rect 53567 -62407 53799 -62202
rect -32991 -63183 45361 -63047
rect 54376 -63302 54512 -61405
rect 62128 -62187 62367 -56802
rect 65035 -56847 65069 -56257
rect 65225 -56254 65270 -56131
rect 65231 -56847 65265 -56254
rect 65647 -56255 65692 -56131
rect 65866 -56138 65928 -56124
rect 65654 -56847 65688 -56255
rect 72767 -55648 72801 -55382
rect 72963 -55648 72997 -55382
rect 73159 -55648 73193 -55382
rect 73355 -55648 73389 -55382
rect 72719 -55723 73437 -55648
rect 68362 -55747 73437 -55723
rect 68362 -55830 73073 -55747
rect 73740 -55828 73774 -55411
rect 73936 -55828 73970 -55411
rect 74132 -55778 74166 -55411
rect 74349 -55778 74383 -55612
rect 74545 -55778 74579 -55612
rect 74741 -55778 74775 -55612
rect 74937 -55778 74971 -55612
rect 74132 -55828 75019 -55778
rect 67024 -55900 73073 -55830
rect 73730 -55877 75019 -55828
rect 73730 -55891 74172 -55877
rect 66657 -55937 73073 -55900
rect 73729 -55920 74172 -55891
rect 73729 -55937 74347 -55920
rect 66657 -55953 74842 -55937
rect 66657 -56017 67062 -55953
rect 66094 -56027 66192 -56024
rect 66657 -56027 66774 -56017
rect 66094 -56144 66774 -56027
rect 67024 -56112 67062 -56017
rect 66094 -56150 66192 -56144
rect 67027 -56605 67061 -56112
rect 67221 -56110 67259 -55953
rect 67223 -56605 67257 -56110
rect 67813 -56133 67863 -55953
rect 67939 -56130 67989 -55953
rect 67818 -56605 67852 -56133
rect 67948 -56605 67982 -56130
rect 68170 -56115 68213 -55953
rect 68362 -55987 74842 -55953
rect 68176 -56405 68210 -56115
rect 68367 -56113 68410 -55987
rect 68372 -56405 68406 -56113
rect 62066 -62419 62414 -62187
rect 66101 -58142 66503 -58076
rect 63606 -59118 63640 -58852
rect 63802 -59118 63836 -58852
rect 63998 -59118 64032 -58852
rect 64194 -59118 64228 -58852
rect 63558 -59217 64276 -59118
rect 63740 -59407 63912 -59217
rect 64579 -59298 64613 -58881
rect 64775 -59298 64809 -58881
rect 64971 -59248 65005 -58881
rect 65188 -59248 65222 -59082
rect 65384 -59248 65418 -59082
rect 65580 -59248 65614 -59082
rect 65776 -59248 65810 -59082
rect 64971 -59298 65858 -59248
rect 64569 -59347 65858 -59298
rect 64569 -59361 65011 -59347
rect 64568 -59390 65011 -59361
rect 64568 -59407 65186 -59390
rect 63570 -59518 65681 -59407
rect 63570 -59560 65785 -59518
rect 63972 -59567 64198 -59560
rect 64009 -59574 64198 -59567
rect 65016 -59584 65785 -59560
rect 63570 -59623 64012 -59608
rect 63570 -59672 64859 -59623
rect 63580 -60089 63614 -59672
rect 63776 -60089 63810 -59672
rect 63972 -59722 64859 -59672
rect 65022 -59710 65067 -59584
rect 63972 -60089 64006 -59722
rect 64189 -59888 64223 -59722
rect 64385 -59888 64419 -59722
rect 64581 -59888 64615 -59722
rect 64777 -59888 64811 -59722
rect 65027 -60300 65061 -59710
rect 65217 -59707 65262 -59584
rect 65223 -60300 65257 -59707
rect 65639 -59708 65684 -59584
rect 65646 -60300 65680 -59708
rect 66101 -59443 66167 -58142
rect 66084 -59556 66168 -59443
rect 66437 -59472 66503 -58142
rect 69334 -58349 69456 -55987
rect 72731 -56048 74842 -55987
rect 72731 -56055 74946 -56048
rect 75019 -56055 75081 -56027
rect 72731 -56090 75081 -56055
rect 73133 -56097 73359 -56090
rect 73170 -56104 73359 -56097
rect 74177 -56107 75081 -56090
rect 74177 -56114 74946 -56107
rect 72731 -56153 73173 -56138
rect 72731 -56202 74020 -56153
rect 71456 -56670 72120 -56591
rect 72741 -56619 72775 -56202
rect 72937 -56619 72971 -56202
rect 73133 -56252 74020 -56202
rect 74183 -56240 74228 -56114
rect 73133 -56619 73167 -56252
rect 73350 -56418 73384 -56252
rect 73546 -56418 73580 -56252
rect 73742 -56418 73776 -56252
rect 73938 -56418 73972 -56252
rect 72656 -56668 72791 -56662
rect 72636 -56670 72791 -56668
rect 71456 -56706 72791 -56670
rect 71456 -56776 72120 -56706
rect 72636 -56708 72791 -56706
rect 72656 -56716 72791 -56708
rect 69334 -58471 69966 -58349
rect 67274 -59149 67308 -58883
rect 67470 -59149 67504 -58883
rect 67666 -59149 67700 -58883
rect 67862 -59149 67896 -58883
rect 67226 -59248 67944 -59149
rect 67408 -59438 67580 -59248
rect 68247 -59329 68281 -58912
rect 68443 -59329 68477 -58912
rect 68639 -59279 68673 -58912
rect 68856 -59279 68890 -59113
rect 69052 -59279 69086 -59113
rect 69248 -59279 69282 -59113
rect 69444 -59279 69478 -59113
rect 68639 -59329 69526 -59279
rect 68237 -59378 69526 -59329
rect 68237 -59392 68679 -59378
rect 68236 -59421 68679 -59392
rect 68236 -59438 68854 -59421
rect 67238 -59472 69349 -59438
rect 66437 -59538 69349 -59472
rect 69504 -59513 69583 -59482
rect 67238 -59549 69349 -59538
rect 69404 -59549 69583 -59513
rect 67238 -59591 69583 -59549
rect 67640 -59598 67866 -59591
rect 67677 -59605 67866 -59598
rect 68684 -59596 69583 -59591
rect 68684 -59615 69453 -59596
rect 67238 -59654 67680 -59639
rect 67238 -59703 68527 -59654
rect 67248 -60120 67282 -59703
rect 67444 -60120 67478 -59703
rect 67640 -59753 68527 -59703
rect 68690 -59741 68735 -59615
rect 67640 -60120 67674 -59753
rect 67857 -59919 67891 -59753
rect 68053 -59919 68087 -59753
rect 68249 -59919 68283 -59753
rect 68445 -59919 68479 -59753
rect 68695 -60331 68729 -59741
rect 68885 -59738 68930 -59615
rect 68891 -60331 68925 -59738
rect 69307 -59739 69352 -59615
rect 69504 -59621 69583 -59596
rect 69314 -60331 69348 -59739
rect 69844 -59467 69966 -58471
rect 69754 -59606 69966 -59467
rect 69754 -59634 69893 -59606
rect -32976 -63438 54512 -63302
rect 71456 -62184 71641 -56776
rect 74188 -56830 74222 -56240
rect 74378 -56237 74423 -56114
rect 74384 -56830 74418 -56237
rect 74800 -56238 74845 -56114
rect 75019 -56121 75081 -56107
rect 74807 -56830 74841 -56238
rect 82131 -55610 82165 -55344
rect 82327 -55610 82361 -55344
rect 82523 -55610 82557 -55344
rect 82719 -55610 82753 -55344
rect 82083 -55654 82801 -55610
rect 77524 -55709 82801 -55654
rect 77524 -55813 82437 -55709
rect 83104 -55790 83138 -55373
rect 83300 -55790 83334 -55373
rect 83496 -55740 83530 -55373
rect 83713 -55740 83747 -55574
rect 83909 -55740 83943 -55574
rect 84105 -55740 84139 -55574
rect 84301 -55740 84335 -55574
rect 83496 -55790 84383 -55740
rect 76177 -55883 82437 -55813
rect 83094 -55839 84383 -55790
rect 83094 -55853 83536 -55839
rect 75810 -55899 82437 -55883
rect 83093 -55882 83536 -55853
rect 83093 -55899 83711 -55882
rect 75810 -55936 84206 -55899
rect 75810 -56000 76215 -55936
rect 75247 -56010 75345 -56007
rect 75810 -56010 75927 -56000
rect 75247 -56127 75927 -56010
rect 76177 -56095 76215 -56000
rect 75247 -56133 75345 -56127
rect 76180 -56588 76214 -56095
rect 76374 -56093 76412 -55936
rect 76376 -56588 76410 -56093
rect 76966 -56116 77016 -55936
rect 77092 -56113 77142 -55936
rect 76971 -56588 77005 -56116
rect 77101 -56588 77135 -56113
rect 77323 -56098 77366 -55936
rect 77520 -55996 84206 -55936
rect 77329 -56388 77363 -56098
rect 77520 -56096 77563 -55996
rect 77525 -56388 77559 -56096
rect 75254 -58125 75656 -58059
rect 72759 -59101 72793 -58835
rect 72955 -59101 72989 -58835
rect 73151 -59101 73185 -58835
rect 73347 -59101 73381 -58835
rect 72711 -59200 73429 -59101
rect 72893 -59390 73065 -59200
rect 73732 -59281 73766 -58864
rect 73928 -59281 73962 -58864
rect 74124 -59231 74158 -58864
rect 74341 -59231 74375 -59065
rect 74537 -59231 74571 -59065
rect 74733 -59231 74767 -59065
rect 74929 -59231 74963 -59065
rect 74124 -59281 75011 -59231
rect 73722 -59330 75011 -59281
rect 73722 -59344 74164 -59330
rect 73721 -59373 74164 -59344
rect 73721 -59390 74339 -59373
rect 72723 -59501 74834 -59390
rect 72723 -59543 74938 -59501
rect 73125 -59550 73351 -59543
rect 73162 -59557 73351 -59550
rect 74169 -59567 74938 -59543
rect 72723 -59606 73165 -59591
rect 72723 -59655 74012 -59606
rect 72733 -60072 72767 -59655
rect 72929 -60072 72963 -59655
rect 73125 -59705 74012 -59655
rect 74175 -59693 74220 -59567
rect 73125 -60072 73159 -59705
rect 73342 -59871 73376 -59705
rect 73538 -59871 73572 -59705
rect 73734 -59871 73768 -59705
rect 73930 -59871 73964 -59705
rect 74180 -60283 74214 -59693
rect 74370 -59690 74415 -59567
rect 74376 -60283 74410 -59690
rect 74792 -59691 74837 -59567
rect 74799 -60283 74833 -59691
rect 75254 -59426 75320 -58125
rect 75237 -59539 75321 -59426
rect 75590 -59455 75656 -58125
rect 78487 -58332 78609 -55996
rect 82095 -56010 84206 -55996
rect 82095 -56017 84310 -56010
rect 84383 -56017 84445 -55989
rect 82095 -56052 84445 -56017
rect 82497 -56059 82723 -56052
rect 82534 -56066 82723 -56059
rect 83541 -56069 84445 -56052
rect 83541 -56076 84310 -56069
rect 82095 -56115 82537 -56100
rect 82095 -56164 83384 -56115
rect 80373 -56632 81581 -56449
rect 82105 -56581 82139 -56164
rect 82301 -56581 82335 -56164
rect 82497 -56214 83384 -56164
rect 83547 -56202 83592 -56076
rect 82497 -56581 82531 -56214
rect 82714 -56380 82748 -56214
rect 82910 -56380 82944 -56214
rect 83106 -56380 83140 -56214
rect 83302 -56380 83336 -56214
rect 82020 -56630 82155 -56624
rect 82000 -56632 82155 -56630
rect 80373 -56668 82155 -56632
rect 80373 -56743 81581 -56668
rect 82000 -56670 82155 -56668
rect 82020 -56678 82155 -56670
rect 78487 -58454 79119 -58332
rect 76427 -59132 76461 -58866
rect 76623 -59132 76657 -58866
rect 76819 -59132 76853 -58866
rect 77015 -59132 77049 -58866
rect 76379 -59231 77097 -59132
rect 76561 -59421 76733 -59231
rect 77400 -59312 77434 -58895
rect 77596 -59312 77630 -58895
rect 77792 -59262 77826 -58895
rect 78009 -59262 78043 -59096
rect 78205 -59262 78239 -59096
rect 78401 -59262 78435 -59096
rect 78597 -59262 78631 -59096
rect 77792 -59312 78679 -59262
rect 77390 -59361 78679 -59312
rect 77390 -59375 77832 -59361
rect 77389 -59404 77832 -59375
rect 77389 -59421 78007 -59404
rect 76391 -59455 78502 -59421
rect 75590 -59521 78502 -59455
rect 78657 -59496 78736 -59465
rect 76391 -59532 78502 -59521
rect 78557 -59532 78736 -59496
rect 76391 -59574 78736 -59532
rect 76793 -59581 77019 -59574
rect 76830 -59588 77019 -59581
rect 77837 -59579 78736 -59574
rect 77837 -59598 78606 -59579
rect 76391 -59637 76833 -59622
rect 76391 -59686 77680 -59637
rect 76401 -60103 76435 -59686
rect 76597 -60103 76631 -59686
rect 76793 -59736 77680 -59686
rect 77843 -59724 77888 -59598
rect 76793 -60103 76827 -59736
rect 77010 -59902 77044 -59736
rect 77206 -59902 77240 -59736
rect 77402 -59902 77436 -59736
rect 77598 -59902 77632 -59736
rect 77848 -60314 77882 -59724
rect 78038 -59721 78083 -59598
rect 78044 -60314 78078 -59721
rect 78460 -59722 78505 -59598
rect 78657 -59604 78736 -59579
rect 78467 -60314 78501 -59722
rect 78997 -59450 79119 -58454
rect 78907 -59589 79119 -59450
rect 78907 -59617 79046 -59589
rect 71371 -62429 71753 -62184
rect -31679 -63836 -30520 -63625
rect -31679 -64501 -30522 -63836
rect 80373 -62187 80667 -56743
rect 83552 -56792 83586 -56202
rect 83742 -56199 83787 -56076
rect 83748 -56792 83782 -56199
rect 84164 -56200 84209 -56076
rect 84383 -56083 84445 -56069
rect 84171 -56792 84205 -56200
rect 87299 -55775 87774 -51863
rect 91309 -52743 92592 -52202
rect 89400 -53281 92592 -52743
rect 91309 -53546 92592 -53281
rect 85541 -55845 87973 -55775
rect 85174 -55897 87973 -55845
rect 85174 -55898 86927 -55897
rect 85174 -55962 85579 -55898
rect 84611 -55972 84709 -55969
rect 85174 -55972 85291 -55962
rect 84611 -56089 85291 -55972
rect 85541 -56057 85579 -55962
rect 84611 -56095 84709 -56089
rect 85544 -56550 85578 -56057
rect 85738 -56055 85776 -55898
rect 85740 -56550 85774 -56055
rect 86330 -56078 86380 -55898
rect 86456 -56075 86506 -55898
rect 86335 -56550 86369 -56078
rect 86465 -56550 86499 -56075
rect 86687 -56060 86730 -55898
rect 86693 -56350 86727 -56060
rect 86884 -56058 86927 -55898
rect 86889 -56350 86923 -56058
rect 80324 -62425 80724 -62187
rect 84618 -58087 85020 -58021
rect 82123 -59063 82157 -58797
rect 82319 -59063 82353 -58797
rect 82515 -59063 82549 -58797
rect 82711 -59063 82745 -58797
rect 82075 -59162 82793 -59063
rect 82257 -59352 82429 -59162
rect 83096 -59243 83130 -58826
rect 83292 -59243 83326 -58826
rect 83488 -59193 83522 -58826
rect 83705 -59193 83739 -59027
rect 83901 -59193 83935 -59027
rect 84097 -59193 84131 -59027
rect 84293 -59193 84327 -59027
rect 83488 -59243 84375 -59193
rect 83086 -59292 84375 -59243
rect 83086 -59306 83528 -59292
rect 83085 -59335 83528 -59306
rect 83085 -59352 83703 -59335
rect 82087 -59463 84198 -59352
rect 82087 -59505 84302 -59463
rect 82489 -59512 82715 -59505
rect 82526 -59519 82715 -59512
rect 83533 -59529 84302 -59505
rect 82087 -59568 82529 -59553
rect 82087 -59617 83376 -59568
rect 82097 -60034 82131 -59617
rect 82293 -60034 82327 -59617
rect 82489 -59667 83376 -59617
rect 83539 -59655 83584 -59529
rect 82489 -60034 82523 -59667
rect 82706 -59833 82740 -59667
rect 82902 -59833 82936 -59667
rect 83098 -59833 83132 -59667
rect 83294 -59833 83328 -59667
rect 83544 -60245 83578 -59655
rect 83734 -59652 83779 -59529
rect 83740 -60245 83774 -59652
rect 84156 -59653 84201 -59529
rect 84163 -60245 84197 -59653
rect 84618 -59388 84684 -58087
rect 84601 -59501 84685 -59388
rect 84954 -59417 85020 -58087
rect 87851 -58294 87973 -55897
rect 87851 -58416 88483 -58294
rect 85791 -59094 85825 -58828
rect 85987 -59094 86021 -58828
rect 86183 -59094 86217 -58828
rect 86379 -59094 86413 -58828
rect 85743 -59193 86461 -59094
rect 85925 -59383 86097 -59193
rect 86764 -59274 86798 -58857
rect 86960 -59274 86994 -58857
rect 87156 -59224 87190 -58857
rect 87373 -59224 87407 -59058
rect 87569 -59224 87603 -59058
rect 87765 -59224 87799 -59058
rect 87961 -59224 87995 -59058
rect 87156 -59274 88043 -59224
rect 86754 -59323 88043 -59274
rect 86754 -59337 87196 -59323
rect 86753 -59366 87196 -59337
rect 86753 -59383 87371 -59366
rect 85755 -59417 87866 -59383
rect 84954 -59483 87866 -59417
rect 88021 -59458 88100 -59427
rect 85755 -59494 87866 -59483
rect 87921 -59494 88100 -59458
rect 85755 -59536 88100 -59494
rect 86157 -59543 86383 -59536
rect 86194 -59550 86383 -59543
rect 87201 -59541 88100 -59536
rect 87201 -59560 87970 -59541
rect 85755 -59599 86197 -59584
rect 85755 -59648 87044 -59599
rect 85765 -60065 85799 -59648
rect 85961 -60065 85995 -59648
rect 86157 -59698 87044 -59648
rect 87207 -59686 87252 -59560
rect 86157 -60065 86191 -59698
rect 86374 -59864 86408 -59698
rect 86570 -59864 86604 -59698
rect 86766 -59864 86800 -59698
rect 86962 -59864 86996 -59698
rect 87212 -60276 87246 -59686
rect 87402 -59683 87447 -59560
rect 87408 -60276 87442 -59683
rect 87824 -59684 87869 -59560
rect 88021 -59566 88100 -59541
rect 87831 -60276 87865 -59684
rect 88361 -59412 88483 -58416
rect 88271 -59551 88483 -59412
rect 88271 -59579 88410 -59551
rect -22800 -64501 -22587 -64469
rect -31679 -64637 11555 -64501
rect -31679 -64865 -30522 -64637
rect -22800 -64647 -22587 -64637
<< obsli1 >>
rect -12466 120695 -12123 121054
rect -12316 119883 -12273 120695
rect -12170 120147 -12098 120171
rect -12170 120077 -10691 120147
rect -12170 120066 -12098 120077
rect -12316 119875 -12029 119883
rect -12316 119841 -11435 119875
rect -12316 119840 -12029 119841
rect -12316 119798 -12273 119840
rect -12356 119792 -12273 119798
rect -12655 119758 -12273 119792
rect -12356 119754 -12273 119758
rect -12313 119706 -12273 119754
rect -12183 119668 -12128 119806
rect -12293 119625 -12077 119668
rect -11445 119663 -11367 119669
rect -12043 119629 -11367 119663
rect -11445 119627 -11367 119629
rect -12293 119359 -12253 119625
rect -12116 119569 -12077 119625
rect -12116 119565 -12023 119569
rect -12205 119383 -12150 119538
rect -12116 119531 -11435 119565
rect -12116 119527 -12023 119531
rect -12114 119467 -12025 119472
rect -11401 119471 -11367 119627
rect -11443 119467 -11367 119471
rect -12114 119433 -11367 119467
rect -12114 119430 -12025 119433
rect -12363 119354 -12253 119359
rect -12655 119320 -12253 119354
rect -12363 119314 -12253 119320
rect -12313 119113 -12258 119268
rect -12301 119076 -12267 119113
rect -12196 119048 -12160 119383
rect -12114 119260 -12078 119430
rect -11443 119429 -11367 119433
rect -10761 119809 -10691 120077
rect -10933 119775 -10691 119809
rect -10702 119677 -10594 119711
rect -10933 119579 -10825 119613
rect -10702 119481 -10594 119515
rect -10933 119383 -10825 119417
rect -12114 119256 -12019 119260
rect -12114 119222 -11435 119256
rect -12114 119218 -12019 119222
rect -10791 119265 -10731 119338
rect -10778 119204 -10737 119265
rect -10778 119193 -10558 119204
rect -10778 119165 -10550 119193
rect -10750 119143 -10550 119165
rect -11765 119048 -11695 119054
rect -12198 118978 -11695 119048
rect -11765 118810 -11695 118978
rect -11765 118776 -11523 118810
rect -11862 118678 -11754 118712
rect -11631 118580 -11523 118614
rect -11862 118482 -11754 118516
rect -11631 118384 -11523 118418
rect -11725 118266 -11665 118339
rect -10588 119004 -10550 119143
rect -10503 119056 -10432 119130
rect -10395 119068 -10087 119102
rect -10932 118970 -10550 119004
rect -10588 118808 -10550 118970
rect -10932 118774 -10550 118808
rect -10581 118591 -10527 118726
rect -10477 118715 -10438 119056
rect -10395 118970 -10087 119004
rect -10395 118872 -10087 118906
rect -10477 118645 -10437 118715
rect -10395 118676 -10087 118710
rect -10479 118644 -10437 118645
rect -10575 118571 -10535 118591
rect -11719 118205 -11678 118266
rect -11898 118194 -11678 118205
rect -11906 118166 -11678 118194
rect -11906 118144 -11706 118166
rect -12369 118069 -12061 118103
rect -12024 118057 -11953 118131
rect -12369 117971 -12061 118005
rect -12369 117873 -12061 117907
rect -12018 117716 -11979 118057
rect -11906 118005 -11868 118144
rect -11906 117971 -11524 118005
rect -11906 117809 -11868 117971
rect -11906 117775 -11524 117809
rect -12369 117677 -12061 117711
rect -12019 117646 -11979 117716
rect -12019 117645 -11977 117646
rect -12017 117419 -11977 117645
rect -10573 118364 -10537 118571
rect -10803 118193 -10595 118227
rect -10479 118129 -10439 118644
rect -9693 119055 -8722 119093
rect -10479 118096 -10265 118129
rect -10473 118095 -10265 118096
rect -10803 117997 -10595 118031
rect -10473 117899 -10265 117933
rect -10803 117801 -10595 117835
rect -12285 116919 -11993 116962
rect -12285 116215 -12242 116919
rect -12036 116720 -11993 116919
rect -10561 117683 -10501 117756
rect -10548 117639 -10507 117683
rect -10565 117612 -10415 117639
rect -10615 117536 -10415 117612
rect -10565 117509 -10415 117536
rect -10517 117080 -10441 117509
rect -10125 117344 -10071 117356
rect -9693 117344 -9655 119055
rect -8760 118839 -8722 119055
rect -8810 118835 -8192 118839
rect -9113 118801 -8192 118835
rect -8612 118686 -8553 118740
rect -8604 118634 -8570 118686
rect -8455 118634 -8401 118766
rect -8229 118739 -8192 118801
rect -8229 118737 -8099 118739
rect -8229 118703 -7809 118737
rect -8229 118702 -8099 118703
rect -8609 118607 -8323 118634
rect -9113 118600 -8323 118607
rect -9113 118573 -8575 118600
rect -8609 118572 -8575 118573
rect -9113 118475 -8605 118509
rect -8538 118508 -8400 118562
rect -8357 118509 -8323 118600
rect -8357 118475 -7809 118509
rect -8436 118298 -8382 118436
rect -9113 118149 -8574 118183
rect -8609 118058 -8574 118149
rect -8523 118123 -8469 118261
rect -8427 118183 -8393 118298
rect -8427 118149 -7809 118183
rect -9113 118024 -8574 118058
rect -8427 118057 -8393 118149
rect -8540 118023 -8393 118057
rect -7812 118053 -7739 118054
rect -8540 117960 -8506 118023
rect -8317 118019 -7739 118053
rect -9113 117926 -8506 117960
rect -8468 117955 -8310 117956
rect -8468 117921 -7809 117955
rect -8468 117918 -8310 117921
rect -8676 117821 -8538 117827
rect -8468 117821 -8430 117918
rect -7773 117857 -7739 118019
rect -8317 117823 -7739 117857
rect -7813 117822 -7739 117823
rect -8676 117783 -8430 117821
rect -8676 117773 -8538 117783
rect -8468 117588 -8430 117783
rect -7773 117773 -7739 117822
rect -9113 117554 -8430 117588
rect -8395 117733 -7739 117773
rect -8395 117588 -8355 117733
rect -8395 117554 -7809 117588
rect -8395 117553 -8309 117554
rect -10125 117306 -9655 117344
rect -10125 117283 -10071 117306
rect -10517 117004 -9661 117080
rect -8659 117373 -8605 117511
rect -8854 117235 -8775 117247
rect -8648 117235 -8614 117373
rect -8523 117317 -8469 117455
rect -8854 117168 -8614 117235
rect -8784 117163 -8614 117168
rect -10018 116720 -9933 116746
rect -12036 116677 -9933 116720
rect -10018 116654 -9933 116677
rect -12139 116479 -12067 116503
rect -12139 116409 -10660 116479
rect -12139 116398 -12067 116409
rect -12285 116207 -11998 116215
rect -12285 116173 -11404 116207
rect -12285 116172 -11998 116173
rect -12285 116130 -12242 116172
rect -12325 116124 -12242 116130
rect -12624 116090 -12242 116124
rect -12325 116086 -12242 116090
rect -12282 116038 -12242 116086
rect -12152 116000 -12097 116138
rect -12262 115957 -12046 116000
rect -11414 115995 -11336 116001
rect -12012 115961 -11336 115995
rect -11414 115959 -11336 115961
rect -12262 115691 -12222 115957
rect -12085 115901 -12046 115957
rect -12085 115897 -11992 115901
rect -12174 115715 -12119 115870
rect -12085 115863 -11404 115897
rect -12085 115859 -11992 115863
rect -12083 115799 -11994 115804
rect -11370 115803 -11336 115959
rect -11412 115799 -11336 115803
rect -12083 115765 -11336 115799
rect -12083 115762 -11994 115765
rect -12332 115686 -12222 115691
rect -12624 115652 -12222 115686
rect -12332 115646 -12222 115652
rect -12282 115445 -12227 115600
rect -12270 115408 -12236 115445
rect -12165 115380 -12129 115715
rect -12083 115592 -12047 115762
rect -11412 115761 -11336 115765
rect -10730 116141 -10660 116409
rect -10902 116107 -10660 116141
rect -10671 116009 -10563 116043
rect -10902 115911 -10794 115945
rect -10671 115813 -10563 115847
rect -10902 115715 -10794 115749
rect -12083 115588 -11988 115592
rect -12083 115554 -11404 115588
rect -12083 115550 -11988 115554
rect -10760 115597 -10700 115670
rect -10747 115536 -10706 115597
rect -10747 115525 -10527 115536
rect -10747 115497 -10519 115525
rect -10719 115475 -10519 115497
rect -11734 115380 -11664 115386
rect -12167 115310 -11664 115380
rect -11734 115142 -11664 115310
rect -11734 115108 -11492 115142
rect -11831 115010 -11723 115044
rect -11600 114912 -11492 114946
rect -11831 114814 -11723 114848
rect -11600 114716 -11492 114750
rect -11694 114598 -11634 114671
rect -10557 115336 -10519 115475
rect -10472 115388 -10401 115462
rect -10364 115400 -10056 115434
rect -10901 115302 -10519 115336
rect -10557 115140 -10519 115302
rect -10901 115106 -10519 115140
rect -10550 114923 -10496 115058
rect -10446 115047 -10407 115388
rect -10364 115302 -10056 115336
rect -10364 115204 -10056 115238
rect -10446 114977 -10406 115047
rect -10364 115008 -10056 115042
rect -10448 114976 -10406 114977
rect -10544 114903 -10504 114923
rect -11688 114537 -11647 114598
rect -11867 114526 -11647 114537
rect -11875 114498 -11647 114526
rect -11875 114476 -11675 114498
rect -12338 114401 -12030 114435
rect -11993 114389 -11922 114463
rect -12338 114303 -12030 114337
rect -12338 114205 -12030 114239
rect -11987 114048 -11948 114389
rect -11875 114337 -11837 114476
rect -11875 114303 -11493 114337
rect -11875 114141 -11837 114303
rect -11875 114107 -11493 114141
rect -12338 114009 -12030 114043
rect -11988 113978 -11948 114048
rect -11988 113977 -11946 113978
rect -11986 113751 -11946 113977
rect -10542 114696 -10506 114903
rect -10772 114525 -10564 114559
rect -10448 114461 -10408 114976
rect -10448 114428 -10234 114461
rect -10442 114427 -10234 114428
rect -10772 114329 -10564 114363
rect -10442 114231 -10234 114265
rect -10772 114133 -10564 114167
rect -10530 114015 -10470 114088
rect -10517 113971 -10476 114015
rect -10534 113912 -10384 113971
rect -10534 113846 -9919 113912
rect -9737 113888 -9661 117004
rect -8513 116970 -8479 117317
rect -8832 116927 -8479 116970
rect -8832 116223 -8789 116927
rect -8686 116487 -8614 116511
rect -8686 116417 -7207 116487
rect -8686 116406 -8614 116417
rect -8832 116215 -8545 116223
rect -8832 116181 -7951 116215
rect -8832 116180 -8545 116181
rect -8832 116138 -8789 116180
rect -8872 116132 -8789 116138
rect -9171 116098 -8789 116132
rect -8872 116094 -8789 116098
rect -8829 116046 -8789 116094
rect -8699 116008 -8644 116146
rect -8809 115965 -8593 116008
rect -7961 116003 -7883 116009
rect -8559 115969 -7883 116003
rect -7961 115967 -7883 115969
rect -8809 115699 -8769 115965
rect -8632 115909 -8593 115965
rect -8632 115905 -8539 115909
rect -8721 115723 -8666 115878
rect -8632 115871 -7951 115905
rect -8632 115867 -8539 115871
rect -8630 115807 -8541 115812
rect -7917 115811 -7883 115967
rect -7959 115807 -7883 115811
rect -8630 115773 -7883 115807
rect -8630 115770 -8541 115773
rect -8879 115694 -8769 115699
rect -9171 115660 -8769 115694
rect -8879 115654 -8769 115660
rect -8829 115453 -8774 115608
rect -8817 115416 -8783 115453
rect -8712 115388 -8676 115723
rect -8630 115600 -8594 115770
rect -7959 115769 -7883 115773
rect -7277 116149 -7207 116417
rect -7449 116115 -7207 116149
rect -7218 116017 -7110 116051
rect -7449 115919 -7341 115953
rect -7218 115821 -7110 115855
rect -7449 115723 -7341 115757
rect -8630 115596 -8535 115600
rect -8630 115562 -7951 115596
rect -8630 115558 -8535 115562
rect -7307 115605 -7247 115678
rect -7294 115544 -7253 115605
rect -7294 115533 -7074 115544
rect -7294 115505 -7066 115533
rect -7266 115483 -7066 115505
rect -8281 115388 -8211 115394
rect -8714 115318 -8211 115388
rect -8281 115150 -8211 115318
rect -8281 115116 -8039 115150
rect -8378 115018 -8270 115052
rect -8147 114920 -8039 114954
rect -8378 114822 -8270 114856
rect -8147 114724 -8039 114758
rect -8241 114606 -8181 114679
rect -7104 115344 -7066 115483
rect -7019 115396 -6948 115470
rect -6911 115408 -6603 115442
rect -7448 115310 -7066 115344
rect -7104 115148 -7066 115310
rect -7448 115114 -7066 115148
rect -7097 114931 -7043 115066
rect -6993 115055 -6954 115396
rect -6911 115310 -6603 115344
rect -6911 115212 -6603 115246
rect -6993 114985 -6953 115055
rect -6911 115016 -6603 115050
rect -6995 114984 -6953 114985
rect -7091 114911 -7051 114931
rect -8235 114545 -8194 114606
rect -8414 114534 -8194 114545
rect -8422 114506 -8194 114534
rect -8422 114484 -8222 114506
rect -8885 114409 -8577 114443
rect -8540 114397 -8469 114471
rect -8885 114311 -8577 114345
rect -8885 114213 -8577 114247
rect -8534 114056 -8495 114397
rect -8422 114345 -8384 114484
rect -8422 114311 -8040 114345
rect -8422 114149 -8384 114311
rect -8422 114115 -8040 114149
rect -8885 114017 -8577 114051
rect -8535 113986 -8495 114056
rect -8535 113985 -8493 113986
rect -9740 113846 -9514 113888
rect -8533 113846 -8493 113985
rect -7089 114704 -7053 114911
rect -7319 114533 -7111 114567
rect -6995 114469 -6955 114984
rect -6995 114436 -6781 114469
rect -6989 114435 -6781 114436
rect -7319 114337 -7111 114371
rect -6989 114239 -6781 114273
rect -7319 114141 -7111 114175
rect -7077 114023 -7017 114096
rect -10534 113841 -8493 113846
rect -10493 113836 -8493 113841
rect -9995 113770 -8493 113836
rect -16901 8556 -16766 43724
rect -16664 25306 -16528 50250
rect -14618 113233 -14342 113305
rect -9740 113233 -9514 113770
rect -8533 113759 -8493 113770
rect -14618 113007 -9514 113233
rect -14618 112918 -14342 113007
rect -12354 111406 -12311 111544
rect -12384 111304 -12273 111406
rect -12354 110519 -12311 111304
rect -12208 110783 -12136 110807
rect -12208 110713 -10729 110783
rect -12208 110702 -12136 110713
rect -12354 110511 -12067 110519
rect -12354 110477 -11473 110511
rect -12354 110476 -12067 110477
rect -12354 110434 -12311 110476
rect -12394 110428 -12311 110434
rect -12693 110394 -12311 110428
rect -12394 110390 -12311 110394
rect -12351 110342 -12311 110390
rect -12221 110304 -12166 110442
rect -12331 110261 -12115 110304
rect -11483 110299 -11405 110305
rect -12081 110265 -11405 110299
rect -11483 110263 -11405 110265
rect -12331 109995 -12291 110261
rect -12154 110205 -12115 110261
rect -12154 110201 -12061 110205
rect -12243 110019 -12188 110174
rect -12154 110167 -11473 110201
rect -12154 110163 -12061 110167
rect -12152 110103 -12063 110108
rect -11439 110107 -11405 110263
rect -11481 110103 -11405 110107
rect -12152 110069 -11405 110103
rect -12152 110066 -12063 110069
rect -12401 109990 -12291 109995
rect -12693 109956 -12291 109990
rect -12401 109950 -12291 109956
rect -12351 109749 -12296 109904
rect -12339 109712 -12305 109749
rect -12234 109684 -12198 110019
rect -12152 109896 -12116 110066
rect -11481 110065 -11405 110069
rect -10799 110445 -10729 110713
rect -10971 110411 -10729 110445
rect -10740 110313 -10632 110347
rect -7064 113979 -7023 114023
rect -7081 113849 -6931 113979
rect -6745 113223 -6472 113518
rect -6653 111480 -6514 113223
rect -6678 111210 -6393 111480
rect -10971 110215 -10863 110249
rect -10740 110117 -10632 110151
rect -10971 110019 -10863 110053
rect -12152 109892 -12057 109896
rect -12152 109858 -11473 109892
rect -12152 109854 -12057 109858
rect -10829 109901 -10769 109974
rect -10816 109840 -10775 109901
rect -10816 109829 -10596 109840
rect -10816 109801 -10588 109829
rect -10788 109779 -10588 109801
rect -11803 109684 -11733 109690
rect -12236 109614 -11733 109684
rect -11803 109446 -11733 109614
rect -11803 109412 -11561 109446
rect -11900 109314 -11792 109348
rect -11669 109216 -11561 109250
rect -11900 109118 -11792 109152
rect -11669 109020 -11561 109054
rect -11763 108902 -11703 108975
rect -10626 109640 -10588 109779
rect -10541 109692 -10470 109766
rect -10433 109704 -10125 109738
rect -10970 109606 -10588 109640
rect -10626 109444 -10588 109606
rect -10970 109410 -10588 109444
rect -10619 109227 -10565 109362
rect -10515 109351 -10476 109692
rect -10433 109606 -10125 109640
rect -10433 109508 -10125 109542
rect -10515 109281 -10475 109351
rect -10433 109312 -10125 109346
rect -10517 109280 -10475 109281
rect -10613 109207 -10573 109227
rect -11757 108841 -11716 108902
rect -11936 108830 -11716 108841
rect -11944 108802 -11716 108830
rect -11944 108780 -11744 108802
rect -12407 108705 -12099 108739
rect -12062 108693 -11991 108767
rect -12407 108607 -12099 108641
rect -12407 108509 -12099 108543
rect -12056 108352 -12017 108693
rect -11944 108641 -11906 108780
rect -11944 108607 -11562 108641
rect -11944 108445 -11906 108607
rect -11944 108411 -11562 108445
rect -12407 108313 -12099 108347
rect -12057 108282 -12017 108352
rect -12057 108281 -12015 108282
rect -12055 108055 -12015 108281
rect -10611 109000 -10575 109207
rect -10841 108829 -10633 108863
rect -10517 108765 -10477 109280
rect -9731 109691 -8760 109729
rect -10517 108732 -10303 108765
rect -10511 108731 -10303 108732
rect -10841 108633 -10633 108667
rect -10511 108535 -10303 108569
rect -10841 108437 -10633 108471
rect -12323 107555 -12031 107598
rect -12323 106851 -12280 107555
rect -12074 107356 -12031 107555
rect -10599 108319 -10539 108392
rect -10586 108275 -10545 108319
rect -10603 108248 -10453 108275
rect -10653 108172 -10453 108248
rect -10603 108145 -10453 108172
rect -10555 107716 -10479 108145
rect -10163 107980 -10109 107992
rect -9731 107980 -9693 109691
rect -8798 109475 -8760 109691
rect -8848 109471 -8230 109475
rect -9151 109437 -8230 109471
rect -8650 109322 -8591 109376
rect -8642 109270 -8608 109322
rect -8493 109270 -8439 109402
rect -8267 109375 -8230 109437
rect -8267 109373 -8137 109375
rect -8267 109339 -7847 109373
rect -8267 109338 -8137 109339
rect -8647 109243 -8361 109270
rect -9151 109236 -8361 109243
rect -9151 109209 -8613 109236
rect -8647 109208 -8613 109209
rect -9151 109111 -8643 109145
rect -8576 109144 -8438 109198
rect -8395 109145 -8361 109236
rect -8395 109111 -7847 109145
rect -8474 108934 -8420 109072
rect -9151 108785 -8612 108819
rect -8647 108694 -8612 108785
rect -8561 108759 -8507 108897
rect -8465 108819 -8431 108934
rect -8465 108785 -7847 108819
rect -9151 108660 -8612 108694
rect -8465 108693 -8431 108785
rect -8578 108659 -8431 108693
rect -7850 108689 -7777 108690
rect -8578 108596 -8544 108659
rect -8355 108655 -7777 108689
rect -9151 108562 -8544 108596
rect -8506 108591 -8348 108592
rect -8506 108557 -7847 108591
rect -8506 108554 -8348 108557
rect -8714 108457 -8576 108463
rect -8506 108457 -8468 108554
rect -7811 108493 -7777 108655
rect -8355 108459 -7777 108493
rect -7851 108458 -7777 108459
rect -8714 108419 -8468 108457
rect -8714 108409 -8576 108419
rect -8506 108224 -8468 108419
rect -7811 108409 -7777 108458
rect -9151 108190 -8468 108224
rect -8433 108369 -7777 108409
rect -8433 108224 -8393 108369
rect -8433 108190 -7847 108224
rect -8433 108189 -8347 108190
rect -10163 107942 -9693 107980
rect -10163 107919 -10109 107942
rect -10555 107640 -9699 107716
rect -8697 108009 -8643 108147
rect -8892 107871 -8813 107883
rect -8686 107871 -8652 108009
rect -8561 107953 -8507 108091
rect -8892 107804 -8652 107871
rect -8822 107799 -8652 107804
rect -10056 107356 -9971 107382
rect -12074 107313 -9971 107356
rect -10056 107290 -9971 107313
rect -12177 107115 -12105 107139
rect -12177 107045 -10698 107115
rect -12177 107034 -12105 107045
rect -12323 106843 -12036 106851
rect -12323 106809 -11442 106843
rect -12323 106808 -12036 106809
rect -12323 106766 -12280 106808
rect -12363 106760 -12280 106766
rect -12662 106726 -12280 106760
rect -12363 106722 -12280 106726
rect -12320 106674 -12280 106722
rect -12190 106636 -12135 106774
rect -12300 106593 -12084 106636
rect -11452 106631 -11374 106637
rect -12050 106597 -11374 106631
rect -11452 106595 -11374 106597
rect -12300 106327 -12260 106593
rect -12123 106537 -12084 106593
rect -12123 106533 -12030 106537
rect -12212 106351 -12157 106506
rect -12123 106499 -11442 106533
rect -12123 106495 -12030 106499
rect -12121 106435 -12032 106440
rect -11408 106439 -11374 106595
rect -11450 106435 -11374 106439
rect -12121 106401 -11374 106435
rect -12121 106398 -12032 106401
rect -12370 106322 -12260 106327
rect -12662 106288 -12260 106322
rect -12370 106282 -12260 106288
rect -12320 106081 -12265 106236
rect -12308 106044 -12274 106081
rect -12203 106016 -12167 106351
rect -12121 106228 -12085 106398
rect -11450 106397 -11374 106401
rect -10768 106777 -10698 107045
rect -10940 106743 -10698 106777
rect -10709 106645 -10601 106679
rect -10940 106547 -10832 106581
rect -10709 106449 -10601 106483
rect -10940 106351 -10832 106385
rect -12121 106224 -12026 106228
rect -12121 106190 -11442 106224
rect -12121 106186 -12026 106190
rect -10798 106233 -10738 106306
rect -10785 106172 -10744 106233
rect -10785 106161 -10565 106172
rect -10785 106133 -10557 106161
rect -10757 106111 -10557 106133
rect -11772 106016 -11702 106022
rect -12205 105946 -11702 106016
rect -11772 105778 -11702 105946
rect -11772 105744 -11530 105778
rect -11869 105646 -11761 105680
rect -11638 105548 -11530 105582
rect -11869 105450 -11761 105484
rect -11638 105352 -11530 105386
rect -11732 105234 -11672 105307
rect -10595 105972 -10557 106111
rect -10510 106024 -10439 106098
rect -10402 106036 -10094 106070
rect -10939 105938 -10557 105972
rect -10595 105776 -10557 105938
rect -10939 105742 -10557 105776
rect -10588 105559 -10534 105694
rect -10484 105683 -10445 106024
rect -10402 105938 -10094 105972
rect -10402 105840 -10094 105874
rect -10484 105613 -10444 105683
rect -10402 105644 -10094 105678
rect -10486 105612 -10444 105613
rect -10582 105539 -10542 105559
rect -11726 105173 -11685 105234
rect -11905 105162 -11685 105173
rect -11913 105134 -11685 105162
rect -11913 105112 -11713 105134
rect -12376 105037 -12068 105071
rect -12031 105025 -11960 105099
rect -12376 104939 -12068 104973
rect -12376 104841 -12068 104875
rect -12025 104684 -11986 105025
rect -11913 104973 -11875 105112
rect -11913 104939 -11531 104973
rect -11913 104777 -11875 104939
rect -11913 104743 -11531 104777
rect -12376 104645 -12068 104679
rect -12026 104614 -11986 104684
rect -12026 104613 -11984 104614
rect -12024 104387 -11984 104613
rect -10580 105332 -10544 105539
rect -10810 105161 -10602 105195
rect -10486 105097 -10446 105612
rect -10486 105064 -10272 105097
rect -10480 105063 -10272 105064
rect -10810 104965 -10602 104999
rect -10480 104867 -10272 104901
rect -10810 104769 -10602 104803
rect -10568 104651 -10508 104724
rect -10555 104607 -10514 104651
rect -10572 104548 -10422 104607
rect -10572 104482 -9957 104548
rect -9775 104482 -9699 107640
rect -8551 107606 -8517 107953
rect -8870 107563 -8517 107606
rect -8870 106859 -8827 107563
rect -8724 107123 -8652 107147
rect -8724 107053 -7245 107123
rect -8724 107042 -8652 107053
rect -8870 106851 -8583 106859
rect -8870 106817 -7989 106851
rect -8870 106816 -8583 106817
rect -8870 106774 -8827 106816
rect -8910 106768 -8827 106774
rect -9209 106734 -8827 106768
rect -8910 106730 -8827 106734
rect -8867 106682 -8827 106730
rect -8737 106644 -8682 106782
rect -8847 106601 -8631 106644
rect -7999 106639 -7921 106645
rect -8597 106605 -7921 106639
rect -7999 106603 -7921 106605
rect -8847 106335 -8807 106601
rect -8670 106545 -8631 106601
rect -8670 106541 -8577 106545
rect -8759 106359 -8704 106514
rect -8670 106507 -7989 106541
rect -8670 106503 -8577 106507
rect -8668 106443 -8579 106448
rect -7955 106447 -7921 106603
rect -7997 106443 -7921 106447
rect -8668 106409 -7921 106443
rect -8668 106406 -8579 106409
rect -8917 106330 -8807 106335
rect -9209 106296 -8807 106330
rect -8917 106290 -8807 106296
rect -8867 106089 -8812 106244
rect -8855 106052 -8821 106089
rect -8750 106024 -8714 106359
rect -8668 106236 -8632 106406
rect -7997 106405 -7921 106409
rect -7315 106785 -7245 107053
rect -7487 106751 -7245 106785
rect -7256 106653 -7148 106687
rect -7487 106555 -7379 106589
rect -7256 106457 -7148 106491
rect -7487 106359 -7379 106393
rect -8668 106232 -8573 106236
rect -8668 106198 -7989 106232
rect -8668 106194 -8573 106198
rect -7345 106241 -7285 106314
rect -7332 106180 -7291 106241
rect -7332 106169 -7112 106180
rect -7332 106141 -7104 106169
rect -7304 106119 -7104 106141
rect -8319 106024 -8249 106030
rect -8752 105954 -8249 106024
rect -8319 105786 -8249 105954
rect -8319 105752 -8077 105786
rect -8416 105654 -8308 105688
rect -8185 105556 -8077 105590
rect -8416 105458 -8308 105492
rect -8185 105360 -8077 105394
rect -8279 105242 -8219 105315
rect -7142 105980 -7104 106119
rect -7057 106032 -6986 106106
rect -6949 106044 -6641 106078
rect -7486 105946 -7104 105980
rect -7142 105784 -7104 105946
rect -7486 105750 -7104 105784
rect -7135 105567 -7081 105702
rect -7031 105691 -6992 106032
rect -6949 105946 -6641 105980
rect -6949 105848 -6641 105882
rect -7031 105621 -6991 105691
rect -6949 105652 -6641 105686
rect -7033 105620 -6991 105621
rect -7129 105547 -7089 105567
rect -8273 105181 -8232 105242
rect -8452 105170 -8232 105181
rect -8460 105142 -8232 105170
rect -8460 105120 -8260 105142
rect -8923 105045 -8615 105079
rect -8578 105033 -8507 105107
rect -8923 104947 -8615 104981
rect -8923 104849 -8615 104883
rect -8572 104692 -8533 105033
rect -8460 104981 -8422 105120
rect -8460 104947 -8078 104981
rect -8460 104785 -8422 104947
rect -8460 104751 -8078 104785
rect -8923 104653 -8615 104687
rect -8573 104622 -8533 104692
rect -8573 104621 -8531 104622
rect -8571 104482 -8531 104621
rect -7127 105340 -7091 105547
rect -7357 105169 -7149 105203
rect -7033 105105 -6993 105620
rect -7033 105072 -6819 105105
rect -7027 105071 -6819 105072
rect -7357 104973 -7149 105007
rect -7027 104875 -6819 104909
rect -7357 104777 -7149 104811
rect -7115 104659 -7055 104732
rect -10572 104477 -8531 104482
rect -10531 104472 -8531 104477
rect -10033 104406 -8531 104472
rect -13779 103901 -13599 103938
rect -9763 103901 -9593 104406
rect -8571 104395 -8531 104406
rect -13779 103731 -9593 103901
rect -13779 103692 -13599 103731
rect -12371 102279 -12328 102391
rect -12471 102018 -12167 102279
rect -12371 101366 -12328 102018
rect -12225 101630 -12153 101654
rect -12225 101560 -10746 101630
rect -12225 101549 -12153 101560
rect -12371 101358 -12084 101366
rect -12371 101324 -11490 101358
rect -12371 101323 -12084 101324
rect -12371 101281 -12328 101323
rect -12411 101275 -12328 101281
rect -12710 101241 -12328 101275
rect -12411 101237 -12328 101241
rect -12368 101189 -12328 101237
rect -12238 101151 -12183 101289
rect -12348 101108 -12132 101151
rect -11500 101146 -11422 101152
rect -12098 101112 -11422 101146
rect -11500 101110 -11422 101112
rect -12348 100842 -12308 101108
rect -12171 101052 -12132 101108
rect -12171 101048 -12078 101052
rect -12260 100866 -12205 101021
rect -12171 101014 -11490 101048
rect -12171 101010 -12078 101014
rect -12169 100950 -12080 100955
rect -11456 100954 -11422 101110
rect -11498 100950 -11422 100954
rect -12169 100916 -11422 100950
rect -12169 100913 -12080 100916
rect -12418 100837 -12308 100842
rect -12710 100803 -12308 100837
rect -12418 100797 -12308 100803
rect -12368 100596 -12313 100751
rect -12356 100559 -12322 100596
rect -12251 100531 -12215 100866
rect -12169 100743 -12133 100913
rect -11498 100912 -11422 100916
rect -10816 101292 -10746 101560
rect -10988 101258 -10746 101292
rect -10757 101160 -10649 101194
rect -7102 104615 -7061 104659
rect -7119 104485 -6969 104615
rect -6774 103968 -6534 104236
rect -6706 102318 -6575 103968
rect -6770 101980 -6479 102318
rect -10988 101062 -10880 101096
rect -10757 100964 -10649 100998
rect -10988 100866 -10880 100900
rect -12169 100739 -12074 100743
rect -12169 100705 -11490 100739
rect -12169 100701 -12074 100705
rect -10846 100748 -10786 100821
rect -10833 100687 -10792 100748
rect -10833 100676 -10613 100687
rect -10833 100648 -10605 100676
rect -10805 100626 -10605 100648
rect -11820 100531 -11750 100537
rect -12253 100461 -11750 100531
rect -11820 100293 -11750 100461
rect -11820 100259 -11578 100293
rect -11917 100161 -11809 100195
rect -11686 100063 -11578 100097
rect -11917 99965 -11809 99999
rect -11686 99867 -11578 99901
rect -11780 99749 -11720 99822
rect -10643 100487 -10605 100626
rect -10558 100539 -10487 100613
rect -10450 100551 -10142 100585
rect -10987 100453 -10605 100487
rect -10643 100291 -10605 100453
rect -10987 100257 -10605 100291
rect -10636 100074 -10582 100209
rect -10532 100198 -10493 100539
rect -10450 100453 -10142 100487
rect -10450 100355 -10142 100389
rect -10532 100128 -10492 100198
rect -10450 100159 -10142 100193
rect -10534 100127 -10492 100128
rect -10630 100054 -10590 100074
rect -11774 99688 -11733 99749
rect -11953 99677 -11733 99688
rect -11961 99649 -11733 99677
rect -11961 99627 -11761 99649
rect -12424 99552 -12116 99586
rect -12079 99540 -12008 99614
rect -12424 99454 -12116 99488
rect -12424 99356 -12116 99390
rect -12073 99199 -12034 99540
rect -11961 99488 -11923 99627
rect -11961 99454 -11579 99488
rect -11961 99292 -11923 99454
rect -11961 99258 -11579 99292
rect -12424 99160 -12116 99194
rect -12074 99129 -12034 99199
rect -12074 99128 -12032 99129
rect -12072 98902 -12032 99128
rect -10628 99847 -10592 100054
rect -10858 99676 -10650 99710
rect -10534 99612 -10494 100127
rect -9748 100538 -8777 100576
rect -10534 99579 -10320 99612
rect -10528 99578 -10320 99579
rect -10858 99480 -10650 99514
rect -10528 99382 -10320 99416
rect -10858 99284 -10650 99318
rect -12340 98402 -12048 98445
rect -12340 97698 -12297 98402
rect -12091 98203 -12048 98402
rect -10616 99166 -10556 99239
rect -10603 99122 -10562 99166
rect -10620 99095 -10470 99122
rect -10670 99019 -10470 99095
rect -10620 98992 -10470 99019
rect -10572 98563 -10496 98992
rect -10180 98827 -10126 98839
rect -9748 98827 -9710 100538
rect -8815 100322 -8777 100538
rect -8865 100318 -8247 100322
rect -9168 100284 -8247 100318
rect -8667 100169 -8608 100223
rect -8659 100117 -8625 100169
rect -8510 100117 -8456 100249
rect -8284 100222 -8247 100284
rect -8284 100220 -8154 100222
rect -8284 100186 -7864 100220
rect -8284 100185 -8154 100186
rect -8664 100090 -8378 100117
rect -9168 100083 -8378 100090
rect -9168 100056 -8630 100083
rect -8664 100055 -8630 100056
rect -9168 99958 -8660 99992
rect -8593 99991 -8455 100045
rect -8412 99992 -8378 100083
rect -8412 99958 -7864 99992
rect -8491 99781 -8437 99919
rect -9168 99632 -8629 99666
rect -8664 99541 -8629 99632
rect -8578 99606 -8524 99744
rect -8482 99666 -8448 99781
rect -8482 99632 -7864 99666
rect -9168 99507 -8629 99541
rect -8482 99540 -8448 99632
rect -8595 99506 -8448 99540
rect -7867 99536 -7794 99537
rect -8595 99443 -8561 99506
rect -8372 99502 -7794 99536
rect -9168 99409 -8561 99443
rect -8523 99438 -8365 99439
rect -8523 99404 -7864 99438
rect -8523 99401 -8365 99404
rect -8731 99304 -8593 99310
rect -8523 99304 -8485 99401
rect -7828 99340 -7794 99502
rect -8372 99306 -7794 99340
rect -7868 99305 -7794 99306
rect -8731 99266 -8485 99304
rect -8731 99256 -8593 99266
rect -8523 99071 -8485 99266
rect -7828 99256 -7794 99305
rect -9168 99037 -8485 99071
rect -8450 99216 -7794 99256
rect -8450 99071 -8410 99216
rect -8450 99037 -7864 99071
rect -8450 99036 -8364 99037
rect -10180 98789 -9710 98827
rect -10180 98766 -10126 98789
rect -10572 98487 -9716 98563
rect -8714 98856 -8660 98994
rect -8909 98718 -8830 98730
rect -8703 98718 -8669 98856
rect -8578 98800 -8524 98938
rect -8909 98651 -8669 98718
rect -8839 98646 -8669 98651
rect -10073 98203 -9988 98229
rect -12091 98160 -9988 98203
rect -10073 98137 -9988 98160
rect -12194 97962 -12122 97986
rect -12194 97892 -10715 97962
rect -12194 97881 -12122 97892
rect -12340 97690 -12053 97698
rect -12340 97656 -11459 97690
rect -12340 97655 -12053 97656
rect -12340 97613 -12297 97655
rect -12380 97607 -12297 97613
rect -12679 97573 -12297 97607
rect -12380 97569 -12297 97573
rect -12337 97521 -12297 97569
rect -12207 97483 -12152 97621
rect -12317 97440 -12101 97483
rect -11469 97478 -11391 97484
rect -12067 97444 -11391 97478
rect -11469 97442 -11391 97444
rect -12317 97174 -12277 97440
rect -12140 97384 -12101 97440
rect -12140 97380 -12047 97384
rect -12229 97198 -12174 97353
rect -12140 97346 -11459 97380
rect -12140 97342 -12047 97346
rect -12138 97282 -12049 97287
rect -11425 97286 -11391 97442
rect -11467 97282 -11391 97286
rect -12138 97248 -11391 97282
rect -12138 97245 -12049 97248
rect -12387 97169 -12277 97174
rect -12679 97135 -12277 97169
rect -12387 97129 -12277 97135
rect -12337 96928 -12282 97083
rect -12325 96891 -12291 96928
rect -12220 96863 -12184 97198
rect -12138 97075 -12102 97245
rect -11467 97244 -11391 97248
rect -10785 97624 -10715 97892
rect -10957 97590 -10715 97624
rect -10726 97492 -10618 97526
rect -10957 97394 -10849 97428
rect -10726 97296 -10618 97330
rect -10957 97198 -10849 97232
rect -12138 97071 -12043 97075
rect -12138 97037 -11459 97071
rect -12138 97033 -12043 97037
rect -10815 97080 -10755 97153
rect -10802 97019 -10761 97080
rect -10802 97008 -10582 97019
rect -10802 96980 -10574 97008
rect -10774 96958 -10574 96980
rect -11789 96863 -11719 96869
rect -12222 96793 -11719 96863
rect -11789 96625 -11719 96793
rect -11789 96591 -11547 96625
rect -11886 96493 -11778 96527
rect -11655 96395 -11547 96429
rect -11886 96297 -11778 96331
rect -11655 96199 -11547 96233
rect -11749 96081 -11689 96154
rect -10612 96819 -10574 96958
rect -10527 96871 -10456 96945
rect -10419 96883 -10111 96917
rect -10956 96785 -10574 96819
rect -10612 96623 -10574 96785
rect -10956 96589 -10574 96623
rect -10605 96406 -10551 96541
rect -10501 96530 -10462 96871
rect -10419 96785 -10111 96819
rect -10419 96687 -10111 96721
rect -10501 96460 -10461 96530
rect -10419 96491 -10111 96525
rect -10503 96459 -10461 96460
rect -10599 96386 -10559 96406
rect -11743 96020 -11702 96081
rect -11922 96009 -11702 96020
rect -11930 95981 -11702 96009
rect -11930 95959 -11730 95981
rect -12393 95884 -12085 95918
rect -12048 95872 -11977 95946
rect -12393 95786 -12085 95820
rect -12393 95688 -12085 95722
rect -12042 95531 -12003 95872
rect -11930 95820 -11892 95959
rect -11930 95786 -11548 95820
rect -11930 95624 -11892 95786
rect -11930 95590 -11548 95624
rect -12393 95492 -12085 95526
rect -12043 95461 -12003 95531
rect -12043 95460 -12001 95461
rect -12041 95234 -12001 95460
rect -10597 96179 -10561 96386
rect -10827 96008 -10619 96042
rect -10503 95944 -10463 96459
rect -10503 95911 -10289 95944
rect -10497 95910 -10289 95911
rect -10827 95812 -10619 95846
rect -10497 95714 -10289 95748
rect -10827 95616 -10619 95650
rect -10585 95498 -10525 95571
rect -10572 95454 -10531 95498
rect -10589 95395 -10439 95454
rect -10589 95329 -9974 95395
rect -9792 95329 -9716 98487
rect -8568 98453 -8534 98800
rect -8887 98410 -8534 98453
rect -8887 97706 -8844 98410
rect -8741 97970 -8669 97994
rect -8741 97900 -7262 97970
rect -8741 97889 -8669 97900
rect -8887 97698 -8600 97706
rect -8887 97664 -8006 97698
rect -8887 97663 -8600 97664
rect -8887 97621 -8844 97663
rect -8927 97615 -8844 97621
rect -9226 97581 -8844 97615
rect -8927 97577 -8844 97581
rect -8884 97529 -8844 97577
rect -8754 97491 -8699 97629
rect -8864 97448 -8648 97491
rect -8016 97486 -7938 97492
rect -8614 97452 -7938 97486
rect -8016 97450 -7938 97452
rect -8864 97182 -8824 97448
rect -8687 97392 -8648 97448
rect -8687 97388 -8594 97392
rect -8776 97206 -8721 97361
rect -8687 97354 -8006 97388
rect -8687 97350 -8594 97354
rect -8685 97290 -8596 97295
rect -7972 97294 -7938 97450
rect -8014 97290 -7938 97294
rect -8685 97256 -7938 97290
rect -8685 97253 -8596 97256
rect -8934 97177 -8824 97182
rect -9226 97143 -8824 97177
rect -8934 97137 -8824 97143
rect -8884 96936 -8829 97091
rect -8872 96899 -8838 96936
rect -8767 96871 -8731 97206
rect -8685 97083 -8649 97253
rect -8014 97252 -7938 97256
rect -7332 97632 -7262 97900
rect -7504 97598 -7262 97632
rect -7273 97500 -7165 97534
rect -7504 97402 -7396 97436
rect -7273 97304 -7165 97338
rect -7504 97206 -7396 97240
rect -8685 97079 -8590 97083
rect -8685 97045 -8006 97079
rect -8685 97041 -8590 97045
rect -7362 97088 -7302 97161
rect -7349 97027 -7308 97088
rect -7349 97016 -7129 97027
rect -7349 96988 -7121 97016
rect -7321 96966 -7121 96988
rect -8336 96871 -8266 96877
rect -8769 96801 -8266 96871
rect -8336 96633 -8266 96801
rect -8336 96599 -8094 96633
rect -8433 96501 -8325 96535
rect -8202 96403 -8094 96437
rect -8433 96305 -8325 96339
rect -8202 96207 -8094 96241
rect -8296 96089 -8236 96162
rect -7159 96827 -7121 96966
rect -7074 96879 -7003 96953
rect -6966 96891 -6658 96925
rect -7503 96793 -7121 96827
rect -7159 96631 -7121 96793
rect -7503 96597 -7121 96631
rect -7152 96414 -7098 96549
rect -7048 96538 -7009 96879
rect -6966 96793 -6658 96827
rect -6966 96695 -6658 96729
rect -7048 96468 -7008 96538
rect -6966 96499 -6658 96533
rect -7050 96467 -7008 96468
rect -7146 96394 -7106 96414
rect -8290 96028 -8249 96089
rect -8469 96017 -8249 96028
rect -8477 95989 -8249 96017
rect -8477 95967 -8277 95989
rect -8940 95892 -8632 95926
rect -8595 95880 -8524 95954
rect -8940 95794 -8632 95828
rect -8940 95696 -8632 95730
rect -8589 95539 -8550 95880
rect -8477 95828 -8439 95967
rect -8477 95794 -8095 95828
rect -8477 95632 -8439 95794
rect -8477 95598 -8095 95632
rect -8940 95500 -8632 95534
rect -8590 95469 -8550 95539
rect -8590 95468 -8548 95469
rect -8588 95329 -8548 95468
rect -7144 96187 -7108 96394
rect -7374 96016 -7166 96050
rect -7050 95952 -7010 96467
rect -7050 95919 -6836 95952
rect -7044 95918 -6836 95919
rect -7374 95820 -7166 95854
rect -7044 95722 -6836 95756
rect -7374 95624 -7166 95658
rect -7132 95506 -7072 95579
rect -10589 95324 -8548 95329
rect -10548 95319 -8548 95324
rect -10050 95253 -8548 95319
rect -14622 94757 -14339 94827
rect -9769 94757 -9552 95253
rect -8588 95242 -8548 95253
rect -14622 94540 -9552 94757
rect -14622 94483 -14339 94540
rect -12437 93545 -12394 93637
rect -12524 93253 -12225 93545
rect -12437 92612 -12394 93253
rect -12291 92876 -12219 92900
rect -12291 92806 -10812 92876
rect -12291 92795 -12219 92806
rect -12437 92604 -12150 92612
rect -12437 92570 -11556 92604
rect -12437 92569 -12150 92570
rect -12437 92527 -12394 92569
rect -12477 92521 -12394 92527
rect -12776 92487 -12394 92521
rect -12477 92483 -12394 92487
rect -12434 92435 -12394 92483
rect -12304 92397 -12249 92535
rect -12414 92354 -12198 92397
rect -11566 92392 -11488 92398
rect -12164 92358 -11488 92392
rect -11566 92356 -11488 92358
rect -12414 92088 -12374 92354
rect -12237 92298 -12198 92354
rect -12237 92294 -12144 92298
rect -12326 92112 -12271 92267
rect -12237 92260 -11556 92294
rect -12237 92256 -12144 92260
rect -12235 92196 -12146 92201
rect -11522 92200 -11488 92356
rect -11564 92196 -11488 92200
rect -12235 92162 -11488 92196
rect -12235 92159 -12146 92162
rect -12484 92083 -12374 92088
rect -12776 92049 -12374 92083
rect -12484 92043 -12374 92049
rect -12434 91842 -12379 91997
rect -12422 91805 -12388 91842
rect -12317 91777 -12281 92112
rect -12235 91989 -12199 92159
rect -11564 92158 -11488 92162
rect -10882 92538 -10812 92806
rect -11054 92504 -10812 92538
rect -10823 92406 -10715 92440
rect -7119 95462 -7078 95506
rect -7136 95332 -6986 95462
rect -6771 94805 -6542 95055
rect -6720 93580 -6569 94805
rect -6788 93204 -6474 93580
rect -11054 92308 -10946 92342
rect -10823 92210 -10715 92244
rect -11054 92112 -10946 92146
rect -12235 91985 -12140 91989
rect -12235 91951 -11556 91985
rect -12235 91947 -12140 91951
rect -10912 91994 -10852 92067
rect -10899 91933 -10858 91994
rect -10899 91922 -10679 91933
rect -10899 91894 -10671 91922
rect -10871 91872 -10671 91894
rect -11886 91777 -11816 91783
rect -12319 91707 -11816 91777
rect -11886 91539 -11816 91707
rect -11886 91505 -11644 91539
rect -11983 91407 -11875 91441
rect -11752 91309 -11644 91343
rect -11983 91211 -11875 91245
rect -11752 91113 -11644 91147
rect -11846 90995 -11786 91068
rect -10709 91733 -10671 91872
rect -10624 91785 -10553 91859
rect -10516 91797 -10208 91831
rect -11053 91699 -10671 91733
rect -10709 91537 -10671 91699
rect -11053 91503 -10671 91537
rect -10702 91320 -10648 91455
rect -10598 91444 -10559 91785
rect -10516 91699 -10208 91733
rect -10516 91601 -10208 91635
rect -10598 91374 -10558 91444
rect -10516 91405 -10208 91439
rect -10600 91373 -10558 91374
rect -10696 91300 -10656 91320
rect -11840 90934 -11799 90995
rect -12019 90923 -11799 90934
rect -12027 90895 -11799 90923
rect -12027 90873 -11827 90895
rect -12490 90798 -12182 90832
rect -12145 90786 -12074 90860
rect -12490 90700 -12182 90734
rect -12490 90602 -12182 90636
rect -12139 90445 -12100 90786
rect -12027 90734 -11989 90873
rect -12027 90700 -11645 90734
rect -12027 90538 -11989 90700
rect -12027 90504 -11645 90538
rect -12490 90406 -12182 90440
rect -12140 90375 -12100 90445
rect -12140 90374 -12098 90375
rect -12138 90148 -12098 90374
rect -10694 91093 -10658 91300
rect -10924 90922 -10716 90956
rect -10600 90858 -10560 91373
rect -9814 91784 -8843 91822
rect -10600 90825 -10386 90858
rect -10594 90824 -10386 90825
rect -10924 90726 -10716 90760
rect -10594 90628 -10386 90662
rect -10924 90530 -10716 90564
rect -12406 89648 -12114 89691
rect -12406 88944 -12363 89648
rect -12157 89449 -12114 89648
rect -10682 90412 -10622 90485
rect -10669 90368 -10628 90412
rect -10686 90341 -10536 90368
rect -10736 90265 -10536 90341
rect -10686 90238 -10536 90265
rect -10638 89809 -10562 90238
rect -10246 90073 -10192 90085
rect -9814 90073 -9776 91784
rect -8881 91568 -8843 91784
rect -8931 91564 -8313 91568
rect -9234 91530 -8313 91564
rect -8733 91415 -8674 91469
rect -8725 91363 -8691 91415
rect -8576 91363 -8522 91495
rect -8350 91468 -8313 91530
rect -8350 91466 -8220 91468
rect -8350 91432 -7930 91466
rect -8350 91431 -8220 91432
rect -8730 91336 -8444 91363
rect -9234 91329 -8444 91336
rect -9234 91302 -8696 91329
rect -8730 91301 -8696 91302
rect -9234 91204 -8726 91238
rect -8659 91237 -8521 91291
rect -8478 91238 -8444 91329
rect -8478 91204 -7930 91238
rect -8557 91027 -8503 91165
rect -9234 90878 -8695 90912
rect -8730 90787 -8695 90878
rect -8644 90852 -8590 90990
rect -8548 90912 -8514 91027
rect -8548 90878 -7930 90912
rect -9234 90753 -8695 90787
rect -8548 90786 -8514 90878
rect -8661 90752 -8514 90786
rect -7933 90782 -7860 90783
rect -8661 90689 -8627 90752
rect -8438 90748 -7860 90782
rect -9234 90655 -8627 90689
rect -8589 90684 -8431 90685
rect -8589 90650 -7930 90684
rect -8589 90647 -8431 90650
rect -8797 90550 -8659 90556
rect -8589 90550 -8551 90647
rect -7894 90586 -7860 90748
rect -8438 90552 -7860 90586
rect -7934 90551 -7860 90552
rect -8797 90512 -8551 90550
rect -8797 90502 -8659 90512
rect -8589 90317 -8551 90512
rect -7894 90502 -7860 90551
rect -9234 90283 -8551 90317
rect -8516 90462 -7860 90502
rect -8516 90317 -8476 90462
rect -8516 90283 -7930 90317
rect -8516 90282 -8430 90283
rect -10246 90035 -9776 90073
rect -10246 90012 -10192 90035
rect -10638 89733 -9782 89809
rect -8780 90102 -8726 90240
rect -8975 89964 -8896 89976
rect -8769 89964 -8735 90102
rect -8644 90046 -8590 90184
rect -8975 89897 -8735 89964
rect -8905 89892 -8735 89897
rect -10139 89449 -10054 89475
rect -12157 89406 -10054 89449
rect -10139 89383 -10054 89406
rect -12260 89208 -12188 89232
rect -12260 89138 -10781 89208
rect -12260 89127 -12188 89138
rect -12406 88936 -12119 88944
rect -12406 88902 -11525 88936
rect -12406 88901 -12119 88902
rect -12406 88859 -12363 88901
rect -12446 88853 -12363 88859
rect -12745 88819 -12363 88853
rect -12446 88815 -12363 88819
rect -12403 88767 -12363 88815
rect -12273 88729 -12218 88867
rect -12383 88686 -12167 88729
rect -11535 88724 -11457 88730
rect -12133 88690 -11457 88724
rect -11535 88688 -11457 88690
rect -12383 88420 -12343 88686
rect -12206 88630 -12167 88686
rect -12206 88626 -12113 88630
rect -12295 88444 -12240 88599
rect -12206 88592 -11525 88626
rect -12206 88588 -12113 88592
rect -12204 88528 -12115 88533
rect -11491 88532 -11457 88688
rect -11533 88528 -11457 88532
rect -12204 88494 -11457 88528
rect -12204 88491 -12115 88494
rect -12453 88415 -12343 88420
rect -12745 88381 -12343 88415
rect -12453 88375 -12343 88381
rect -12403 88174 -12348 88329
rect -12391 88137 -12357 88174
rect -12286 88109 -12250 88444
rect -12204 88321 -12168 88491
rect -11533 88490 -11457 88494
rect -10851 88870 -10781 89138
rect -11023 88836 -10781 88870
rect -10792 88738 -10684 88772
rect -11023 88640 -10915 88674
rect -10792 88542 -10684 88576
rect -11023 88444 -10915 88478
rect -12204 88317 -12109 88321
rect -12204 88283 -11525 88317
rect -12204 88279 -12109 88283
rect -10881 88326 -10821 88399
rect -10868 88265 -10827 88326
rect -10868 88254 -10648 88265
rect -10868 88226 -10640 88254
rect -10840 88204 -10640 88226
rect -11855 88109 -11785 88115
rect -12288 88039 -11785 88109
rect -11855 87871 -11785 88039
rect -11855 87837 -11613 87871
rect -11952 87739 -11844 87773
rect -11721 87641 -11613 87675
rect -11952 87543 -11844 87577
rect -11721 87445 -11613 87479
rect -11815 87327 -11755 87400
rect -10678 88065 -10640 88204
rect -10593 88117 -10522 88191
rect -10485 88129 -10177 88163
rect -11022 88031 -10640 88065
rect -10678 87869 -10640 88031
rect -11022 87835 -10640 87869
rect -10671 87652 -10617 87787
rect -10567 87776 -10528 88117
rect -10485 88031 -10177 88065
rect -10485 87933 -10177 87967
rect -10567 87706 -10527 87776
rect -10485 87737 -10177 87771
rect -10569 87705 -10527 87706
rect -10665 87632 -10625 87652
rect -11809 87266 -11768 87327
rect -11988 87255 -11768 87266
rect -11996 87227 -11768 87255
rect -11996 87205 -11796 87227
rect -12459 87130 -12151 87164
rect -12114 87118 -12043 87192
rect -12459 87032 -12151 87066
rect -12459 86934 -12151 86968
rect -12108 86777 -12069 87118
rect -11996 87066 -11958 87205
rect -11996 87032 -11614 87066
rect -11996 86870 -11958 87032
rect -11996 86836 -11614 86870
rect -12459 86738 -12151 86772
rect -12109 86707 -12069 86777
rect -12109 86706 -12067 86707
rect -12107 86480 -12067 86706
rect -10663 87425 -10627 87632
rect -10893 87254 -10685 87288
rect -10569 87190 -10529 87705
rect -10569 87157 -10355 87190
rect -10563 87156 -10355 87157
rect -10893 87058 -10685 87092
rect -10563 86960 -10355 86994
rect -10893 86862 -10685 86896
rect -10651 86744 -10591 86817
rect -10638 86700 -10597 86744
rect -10655 86641 -10505 86700
rect -10655 86575 -10040 86641
rect -9858 86575 -9782 89733
rect -8634 89699 -8600 90046
rect -8953 89656 -8600 89699
rect -8953 88952 -8910 89656
rect -8807 89216 -8735 89240
rect -8807 89146 -7328 89216
rect -8807 89135 -8735 89146
rect -8953 88944 -8666 88952
rect -8953 88910 -8072 88944
rect -8953 88909 -8666 88910
rect -8953 88867 -8910 88909
rect -8993 88861 -8910 88867
rect -9292 88827 -8910 88861
rect -8993 88823 -8910 88827
rect -8950 88775 -8910 88823
rect -8820 88737 -8765 88875
rect -8930 88694 -8714 88737
rect -8082 88732 -8004 88738
rect -8680 88698 -8004 88732
rect -8082 88696 -8004 88698
rect -8930 88428 -8890 88694
rect -8753 88638 -8714 88694
rect -8753 88634 -8660 88638
rect -8842 88452 -8787 88607
rect -8753 88600 -8072 88634
rect -8753 88596 -8660 88600
rect -8751 88536 -8662 88541
rect -8038 88540 -8004 88696
rect -8080 88536 -8004 88540
rect -8751 88502 -8004 88536
rect -8751 88499 -8662 88502
rect -9000 88423 -8890 88428
rect -9292 88389 -8890 88423
rect -9000 88383 -8890 88389
rect -8950 88182 -8895 88337
rect -8938 88145 -8904 88182
rect -8833 88117 -8797 88452
rect -8751 88329 -8715 88499
rect -8080 88498 -8004 88502
rect -7398 88878 -7328 89146
rect -7570 88844 -7328 88878
rect -7339 88746 -7231 88780
rect -7570 88648 -7462 88682
rect -7339 88550 -7231 88584
rect -7570 88452 -7462 88486
rect -8751 88325 -8656 88329
rect -8751 88291 -8072 88325
rect -8751 88287 -8656 88291
rect -7428 88334 -7368 88407
rect -7415 88273 -7374 88334
rect -7415 88262 -7195 88273
rect -7415 88234 -7187 88262
rect -7387 88212 -7187 88234
rect -8402 88117 -8332 88123
rect -8835 88047 -8332 88117
rect -8402 87879 -8332 88047
rect -8402 87845 -8160 87879
rect -8499 87747 -8391 87781
rect -8268 87649 -8160 87683
rect -8499 87551 -8391 87585
rect -8268 87453 -8160 87487
rect -8362 87335 -8302 87408
rect -7225 88073 -7187 88212
rect -7140 88125 -7069 88199
rect -7032 88137 -6724 88171
rect -7569 88039 -7187 88073
rect -7225 87877 -7187 88039
rect -7569 87843 -7187 87877
rect -7218 87660 -7164 87795
rect -7114 87784 -7075 88125
rect -7032 88039 -6724 88073
rect -7032 87941 -6724 87975
rect -7114 87714 -7074 87784
rect -7032 87745 -6724 87779
rect -7116 87713 -7074 87714
rect -7212 87640 -7172 87660
rect -8356 87274 -8315 87335
rect -8535 87263 -8315 87274
rect -8543 87235 -8315 87263
rect -8543 87213 -8343 87235
rect -9006 87138 -8698 87172
rect -8661 87126 -8590 87200
rect -9006 87040 -8698 87074
rect -9006 86942 -8698 86976
rect -8655 86785 -8616 87126
rect -8543 87074 -8505 87213
rect -8543 87040 -8161 87074
rect -8543 86878 -8505 87040
rect -8543 86844 -8161 86878
rect -9006 86746 -8698 86780
rect -8656 86715 -8616 86785
rect -8656 86714 -8614 86715
rect -8654 86575 -8614 86714
rect -7210 87433 -7174 87640
rect -7440 87262 -7232 87296
rect -7116 87198 -7076 87713
rect -7116 87165 -6902 87198
rect -7110 87164 -6902 87165
rect -7440 87066 -7232 87100
rect -7110 86968 -6902 87002
rect -7440 86870 -7232 86904
rect -7198 86752 -7138 86825
rect -10655 86570 -8614 86575
rect -10614 86565 -8614 86570
rect -10116 86499 -8614 86565
rect -13774 85949 -13607 85964
rect -9686 85949 -9525 86499
rect -8654 86488 -8614 86499
rect -13774 85788 -9525 85949
rect -13774 85770 -13607 85788
rect -12471 84341 -12428 84439
rect -12533 84127 -12313 84341
rect -12471 83414 -12428 84127
rect -12325 83678 -12253 83702
rect -12325 83608 -10846 83678
rect -12325 83597 -12253 83608
rect -12471 83406 -12184 83414
rect -12471 83372 -11590 83406
rect -12471 83371 -12184 83372
rect -12471 83329 -12428 83371
rect -12511 83323 -12428 83329
rect -12810 83289 -12428 83323
rect -12511 83285 -12428 83289
rect -12468 83237 -12428 83285
rect -12338 83199 -12283 83337
rect -12448 83156 -12232 83199
rect -11600 83194 -11522 83200
rect -12198 83160 -11522 83194
rect -11600 83158 -11522 83160
rect -12448 82890 -12408 83156
rect -12271 83100 -12232 83156
rect -12271 83096 -12178 83100
rect -12360 82914 -12305 83069
rect -12271 83062 -11590 83096
rect -12271 83058 -12178 83062
rect -12269 82998 -12180 83003
rect -11556 83002 -11522 83158
rect -11598 82998 -11522 83002
rect -12269 82964 -11522 82998
rect -12269 82961 -12180 82964
rect -12518 82885 -12408 82890
rect -12810 82851 -12408 82885
rect -12518 82845 -12408 82851
rect -12468 82644 -12413 82799
rect -12456 82607 -12422 82644
rect -12351 82579 -12315 82914
rect -12269 82791 -12233 82961
rect -11598 82960 -11522 82964
rect -10916 83340 -10846 83608
rect -11088 83306 -10846 83340
rect -10857 83208 -10749 83242
rect -7185 86708 -7144 86752
rect -7202 86578 -7052 86708
rect -6832 85766 -6612 86012
rect -6825 84339 -6692 85766
rect -6917 84113 -6683 84339
rect -11088 83110 -10980 83144
rect -10857 83012 -10749 83046
rect -11088 82914 -10980 82948
rect -12269 82787 -12174 82791
rect -12269 82753 -11590 82787
rect -12269 82749 -12174 82753
rect -10946 82796 -10886 82869
rect -10933 82735 -10892 82796
rect -10933 82724 -10713 82735
rect -10933 82696 -10705 82724
rect -10905 82674 -10705 82696
rect -11920 82579 -11850 82585
rect -12353 82509 -11850 82579
rect -11920 82341 -11850 82509
rect -11920 82307 -11678 82341
rect -12017 82209 -11909 82243
rect -11786 82111 -11678 82145
rect -12017 82013 -11909 82047
rect -11786 81915 -11678 81949
rect -11880 81797 -11820 81870
rect -10743 82535 -10705 82674
rect -10658 82587 -10587 82661
rect -10550 82599 -10242 82633
rect -11087 82501 -10705 82535
rect -10743 82339 -10705 82501
rect -11087 82305 -10705 82339
rect -10736 82122 -10682 82257
rect -10632 82246 -10593 82587
rect -10550 82501 -10242 82535
rect -10550 82403 -10242 82437
rect -10632 82176 -10592 82246
rect -10550 82207 -10242 82241
rect -10634 82175 -10592 82176
rect -10730 82102 -10690 82122
rect -11874 81736 -11833 81797
rect -12053 81725 -11833 81736
rect -12061 81697 -11833 81725
rect -12061 81675 -11861 81697
rect -12524 81600 -12216 81634
rect -12179 81588 -12108 81662
rect -12524 81502 -12216 81536
rect -12524 81404 -12216 81438
rect -12173 81247 -12134 81588
rect -12061 81536 -12023 81675
rect -12061 81502 -11679 81536
rect -12061 81340 -12023 81502
rect -12061 81306 -11679 81340
rect -12524 81208 -12216 81242
rect -12174 81177 -12134 81247
rect -12174 81176 -12132 81177
rect -12172 80950 -12132 81176
rect -10728 81895 -10692 82102
rect -10958 81724 -10750 81758
rect -10634 81660 -10594 82175
rect -9848 82586 -8877 82624
rect -10634 81627 -10420 81660
rect -10628 81626 -10420 81627
rect -10958 81528 -10750 81562
rect -10628 81430 -10420 81464
rect -10958 81332 -10750 81366
rect -12440 80450 -12148 80493
rect -12440 79746 -12397 80450
rect -12191 80251 -12148 80450
rect -10716 81214 -10656 81287
rect -10703 81170 -10662 81214
rect -10720 81143 -10570 81170
rect -10770 81067 -10570 81143
rect -10720 81040 -10570 81067
rect -10672 80611 -10596 81040
rect -10280 80875 -10226 80887
rect -9848 80875 -9810 82586
rect -8915 82370 -8877 82586
rect -8965 82366 -8347 82370
rect -9268 82332 -8347 82366
rect -8767 82217 -8708 82271
rect -8759 82165 -8725 82217
rect -8610 82165 -8556 82297
rect -8384 82270 -8347 82332
rect -8384 82268 -8254 82270
rect -8384 82234 -7964 82268
rect -8384 82233 -8254 82234
rect -8764 82138 -8478 82165
rect -9268 82131 -8478 82138
rect -9268 82104 -8730 82131
rect -8764 82103 -8730 82104
rect -9268 82006 -8760 82040
rect -8693 82039 -8555 82093
rect -8512 82040 -8478 82131
rect -8512 82006 -7964 82040
rect -8591 81829 -8537 81967
rect -9268 81680 -8729 81714
rect -8764 81589 -8729 81680
rect -8678 81654 -8624 81792
rect -8582 81714 -8548 81829
rect -8582 81680 -7964 81714
rect -9268 81555 -8729 81589
rect -8582 81588 -8548 81680
rect -8695 81554 -8548 81588
rect -7967 81584 -7894 81585
rect -8695 81491 -8661 81554
rect -8472 81550 -7894 81584
rect -9268 81457 -8661 81491
rect -8623 81486 -8465 81487
rect -8623 81452 -7964 81486
rect -8623 81449 -8465 81452
rect -8831 81352 -8693 81358
rect -8623 81352 -8585 81449
rect -7928 81388 -7894 81550
rect -8472 81354 -7894 81388
rect -7968 81353 -7894 81354
rect -8831 81314 -8585 81352
rect -8831 81304 -8693 81314
rect -8623 81119 -8585 81314
rect -7928 81304 -7894 81353
rect -9268 81085 -8585 81119
rect -8550 81264 -7894 81304
rect -8550 81119 -8510 81264
rect -8550 81085 -7964 81119
rect -8550 81084 -8464 81085
rect -10280 80837 -9810 80875
rect -10280 80814 -10226 80837
rect -10672 80535 -9816 80611
rect -8814 80904 -8760 81042
rect -9009 80766 -8930 80778
rect -8803 80766 -8769 80904
rect -8678 80848 -8624 80986
rect -9009 80699 -8769 80766
rect -8939 80694 -8769 80699
rect -10173 80251 -10088 80277
rect -12191 80208 -10088 80251
rect -10173 80185 -10088 80208
rect -12294 80010 -12222 80034
rect -12294 79940 -10815 80010
rect -12294 79929 -12222 79940
rect -12440 79738 -12153 79746
rect -12440 79704 -11559 79738
rect -12440 79703 -12153 79704
rect -12440 79661 -12397 79703
rect -12480 79655 -12397 79661
rect -12779 79621 -12397 79655
rect -12480 79617 -12397 79621
rect -12437 79569 -12397 79617
rect -12307 79531 -12252 79669
rect -12417 79488 -12201 79531
rect -11569 79526 -11491 79532
rect -12167 79492 -11491 79526
rect -11569 79490 -11491 79492
rect -12417 79222 -12377 79488
rect -12240 79432 -12201 79488
rect -12240 79428 -12147 79432
rect -12329 79246 -12274 79401
rect -12240 79394 -11559 79428
rect -12240 79390 -12147 79394
rect -12238 79330 -12149 79335
rect -11525 79334 -11491 79490
rect -11567 79330 -11491 79334
rect -12238 79296 -11491 79330
rect -12238 79293 -12149 79296
rect -12487 79217 -12377 79222
rect -12779 79183 -12377 79217
rect -12487 79177 -12377 79183
rect -12437 78976 -12382 79131
rect -12425 78939 -12391 78976
rect -12320 78911 -12284 79246
rect -12238 79123 -12202 79293
rect -11567 79292 -11491 79296
rect -10885 79672 -10815 79940
rect -11057 79638 -10815 79672
rect -10826 79540 -10718 79574
rect -11057 79442 -10949 79476
rect -10826 79344 -10718 79378
rect -11057 79246 -10949 79280
rect -12238 79119 -12143 79123
rect -12238 79085 -11559 79119
rect -12238 79081 -12143 79085
rect -10915 79128 -10855 79201
rect -10902 79067 -10861 79128
rect -10902 79056 -10682 79067
rect -10902 79028 -10674 79056
rect -10874 79006 -10674 79028
rect -11889 78911 -11819 78917
rect -12322 78841 -11819 78911
rect -11889 78673 -11819 78841
rect -11889 78639 -11647 78673
rect -11986 78541 -11878 78575
rect -11755 78443 -11647 78477
rect -11986 78345 -11878 78379
rect -11755 78247 -11647 78281
rect -11849 78129 -11789 78202
rect -10712 78867 -10674 79006
rect -10627 78919 -10556 78993
rect -10519 78931 -10211 78965
rect -11056 78833 -10674 78867
rect -10712 78671 -10674 78833
rect -11056 78637 -10674 78671
rect -10705 78454 -10651 78589
rect -10601 78578 -10562 78919
rect -10519 78833 -10211 78867
rect -10519 78735 -10211 78769
rect -10601 78508 -10561 78578
rect -10519 78539 -10211 78573
rect -10603 78507 -10561 78508
rect -10699 78434 -10659 78454
rect -11843 78068 -11802 78129
rect -12022 78057 -11802 78068
rect -12030 78029 -11802 78057
rect -12030 78007 -11830 78029
rect -12493 77932 -12185 77966
rect -12148 77920 -12077 77994
rect -12493 77834 -12185 77868
rect -12493 77736 -12185 77770
rect -12142 77579 -12103 77920
rect -12030 77868 -11992 78007
rect -12030 77834 -11648 77868
rect -12030 77672 -11992 77834
rect -12030 77638 -11648 77672
rect -12493 77540 -12185 77574
rect -12143 77509 -12103 77579
rect -12143 77508 -12101 77509
rect -12141 77282 -12101 77508
rect -10697 78227 -10661 78434
rect -10927 78056 -10719 78090
rect -10603 77992 -10563 78507
rect -10603 77959 -10389 77992
rect -10597 77958 -10389 77959
rect -10927 77860 -10719 77894
rect -10597 77762 -10389 77796
rect -10927 77664 -10719 77698
rect -10685 77546 -10625 77619
rect -10672 77502 -10631 77546
rect -10689 77443 -10539 77502
rect -10689 77377 -10074 77443
rect -9892 77377 -9816 80535
rect -8668 80501 -8634 80848
rect -8987 80458 -8634 80501
rect -8987 79754 -8944 80458
rect -8841 80018 -8769 80042
rect -8841 79948 -7362 80018
rect -8841 79937 -8769 79948
rect -8987 79746 -8700 79754
rect -8987 79712 -8106 79746
rect -8987 79711 -8700 79712
rect -8987 79669 -8944 79711
rect -9027 79663 -8944 79669
rect -9326 79629 -8944 79663
rect -9027 79625 -8944 79629
rect -8984 79577 -8944 79625
rect -8854 79539 -8799 79677
rect -8964 79496 -8748 79539
rect -8116 79534 -8038 79540
rect -8714 79500 -8038 79534
rect -8116 79498 -8038 79500
rect -8964 79230 -8924 79496
rect -8787 79440 -8748 79496
rect -8787 79436 -8694 79440
rect -8876 79254 -8821 79409
rect -8787 79402 -8106 79436
rect -8787 79398 -8694 79402
rect -8785 79338 -8696 79343
rect -8072 79342 -8038 79498
rect -8114 79338 -8038 79342
rect -8785 79304 -8038 79338
rect -8785 79301 -8696 79304
rect -9034 79225 -8924 79230
rect -9326 79191 -8924 79225
rect -9034 79185 -8924 79191
rect -8984 78984 -8929 79139
rect -8972 78947 -8938 78984
rect -8867 78919 -8831 79254
rect -8785 79131 -8749 79301
rect -8114 79300 -8038 79304
rect -7432 79680 -7362 79948
rect -7604 79646 -7362 79680
rect -7373 79548 -7265 79582
rect -7604 79450 -7496 79484
rect -7373 79352 -7265 79386
rect -7604 79254 -7496 79288
rect -8785 79127 -8690 79131
rect -8785 79093 -8106 79127
rect -8785 79089 -8690 79093
rect -7462 79136 -7402 79209
rect -7449 79075 -7408 79136
rect -7449 79064 -7229 79075
rect -7449 79036 -7221 79064
rect -7421 79014 -7221 79036
rect -8436 78919 -8366 78925
rect -8869 78849 -8366 78919
rect -8436 78681 -8366 78849
rect -8436 78647 -8194 78681
rect -8533 78549 -8425 78583
rect -8302 78451 -8194 78485
rect -8533 78353 -8425 78387
rect -8302 78255 -8194 78289
rect -8396 78137 -8336 78210
rect -7259 78875 -7221 79014
rect -7174 78927 -7103 79001
rect -7066 78939 -6758 78973
rect -7603 78841 -7221 78875
rect -7259 78679 -7221 78841
rect -7603 78645 -7221 78679
rect -7252 78462 -7198 78597
rect -7148 78586 -7109 78927
rect -7066 78841 -6758 78875
rect -7066 78743 -6758 78777
rect -7148 78516 -7108 78586
rect -7066 78547 -6758 78581
rect -7150 78515 -7108 78516
rect -7246 78442 -7206 78462
rect -8390 78076 -8349 78137
rect -8569 78065 -8349 78076
rect -8577 78037 -8349 78065
rect -8577 78015 -8377 78037
rect -9040 77940 -8732 77974
rect -8695 77928 -8624 78002
rect -9040 77842 -8732 77876
rect -9040 77744 -8732 77778
rect -8689 77587 -8650 77928
rect -8577 77876 -8539 78015
rect -8577 77842 -8195 77876
rect -8577 77680 -8539 77842
rect -8577 77646 -8195 77680
rect -9040 77548 -8732 77582
rect -8690 77517 -8650 77587
rect -8690 77516 -8648 77517
rect -8688 77377 -8648 77516
rect -7244 78235 -7208 78442
rect -7474 78064 -7266 78098
rect -7150 78000 -7110 78515
rect -7150 77967 -6936 78000
rect -7144 77966 -6936 77967
rect -7474 77868 -7266 77902
rect -7144 77770 -6936 77804
rect -7474 77672 -7266 77706
rect -7232 77554 -7172 77627
rect -10689 77372 -8648 77377
rect -10648 77367 -8648 77372
rect -10150 77301 -8648 77367
rect -9772 76797 -9626 77301
rect -8688 77290 -8648 77301
rect -13773 76651 -9626 76797
rect -12557 75249 -12226 75586
rect -13809 75173 -13518 75207
rect -14589 75164 -13518 75173
rect -14598 74924 -13518 75164
rect -14589 74907 -13518 74924
rect -13809 74890 -13518 74907
rect -12432 74551 -12389 75249
rect -12286 74815 -12214 74839
rect -12286 74745 -10807 74815
rect -12286 74734 -12214 74745
rect -12432 74543 -12145 74551
rect -12432 74509 -11551 74543
rect -12432 74508 -12145 74509
rect -12432 74466 -12389 74508
rect -12472 74460 -12389 74466
rect -12771 74426 -12389 74460
rect -12472 74422 -12389 74426
rect -12429 74374 -12389 74422
rect -12299 74336 -12244 74474
rect -12409 74293 -12193 74336
rect -11561 74331 -11483 74337
rect -12159 74297 -11483 74331
rect -11561 74295 -11483 74297
rect -12409 74027 -12369 74293
rect -12232 74237 -12193 74293
rect -12232 74233 -12139 74237
rect -12321 74051 -12266 74206
rect -12232 74199 -11551 74233
rect -12232 74195 -12139 74199
rect -12230 74135 -12141 74140
rect -11517 74139 -11483 74295
rect -11559 74135 -11483 74139
rect -12230 74101 -11483 74135
rect -12230 74098 -12141 74101
rect -12479 74022 -12369 74027
rect -12771 73988 -12369 74022
rect -12479 73982 -12369 73988
rect -12429 73781 -12374 73936
rect -12417 73744 -12383 73781
rect -12312 73716 -12276 74051
rect -12230 73928 -12194 74098
rect -11559 74097 -11483 74101
rect -10877 74477 -10807 74745
rect -11049 74443 -10807 74477
rect -10818 74345 -10710 74379
rect -7219 77510 -7178 77554
rect -7236 77380 -7086 77510
rect -6878 76775 -6656 77072
rect -6856 75514 -6689 76775
rect -6923 75249 -6658 75514
rect -11049 74247 -10941 74281
rect -10818 74149 -10710 74183
rect -11049 74051 -10941 74085
rect -12230 73924 -12135 73928
rect -12230 73890 -11551 73924
rect -12230 73886 -12135 73890
rect -10907 73933 -10847 74006
rect -10894 73872 -10853 73933
rect -10894 73861 -10674 73872
rect -10894 73833 -10666 73861
rect -10866 73811 -10666 73833
rect -11881 73716 -11811 73722
rect -12314 73646 -11811 73716
rect -11881 73478 -11811 73646
rect -11881 73444 -11639 73478
rect -11978 73346 -11870 73380
rect -11747 73248 -11639 73282
rect -11978 73150 -11870 73184
rect -11747 73052 -11639 73086
rect -11841 72934 -11781 73007
rect -10704 73672 -10666 73811
rect -10619 73724 -10548 73798
rect -10511 73736 -10203 73770
rect -11048 73638 -10666 73672
rect -10704 73476 -10666 73638
rect -11048 73442 -10666 73476
rect -10697 73259 -10643 73394
rect -10593 73383 -10554 73724
rect -10511 73638 -10203 73672
rect -10511 73540 -10203 73574
rect -10593 73313 -10553 73383
rect -10511 73344 -10203 73378
rect -10595 73312 -10553 73313
rect -10691 73239 -10651 73259
rect -11835 72873 -11794 72934
rect -12014 72862 -11794 72873
rect -12022 72834 -11794 72862
rect -12022 72812 -11822 72834
rect -12485 72737 -12177 72771
rect -12140 72725 -12069 72799
rect -12485 72639 -12177 72673
rect -12485 72541 -12177 72575
rect -12134 72384 -12095 72725
rect -12022 72673 -11984 72812
rect -12022 72639 -11640 72673
rect -12022 72477 -11984 72639
rect -12022 72443 -11640 72477
rect -12485 72345 -12177 72379
rect -12135 72314 -12095 72384
rect -12135 72313 -12093 72314
rect -12133 72087 -12093 72313
rect -10689 73032 -10653 73239
rect -10919 72861 -10711 72895
rect -10595 72797 -10555 73312
rect -9809 73723 -8838 73761
rect -10595 72764 -10381 72797
rect -10589 72763 -10381 72764
rect -10919 72665 -10711 72699
rect -10589 72567 -10381 72601
rect -10919 72469 -10711 72503
rect -12401 71587 -12109 71630
rect -12401 70883 -12358 71587
rect -12152 71388 -12109 71587
rect -10677 72351 -10617 72424
rect -10664 72307 -10623 72351
rect -10681 72280 -10531 72307
rect -10731 72204 -10531 72280
rect -10681 72177 -10531 72204
rect -10633 71748 -10557 72177
rect -10241 72012 -10187 72024
rect -9809 72012 -9771 73723
rect -8876 73507 -8838 73723
rect -8926 73503 -8308 73507
rect -9229 73469 -8308 73503
rect -8728 73354 -8669 73408
rect -8720 73302 -8686 73354
rect -8571 73302 -8517 73434
rect -8345 73407 -8308 73469
rect -8345 73405 -8215 73407
rect -8345 73371 -7925 73405
rect -8345 73370 -8215 73371
rect -8725 73275 -8439 73302
rect -9229 73268 -8439 73275
rect -9229 73241 -8691 73268
rect -8725 73240 -8691 73241
rect -9229 73143 -8721 73177
rect -8654 73176 -8516 73230
rect -8473 73177 -8439 73268
rect -8473 73143 -7925 73177
rect -8552 72966 -8498 73104
rect -9229 72817 -8690 72851
rect -8725 72726 -8690 72817
rect -8639 72791 -8585 72929
rect -8543 72851 -8509 72966
rect -8543 72817 -7925 72851
rect -9229 72692 -8690 72726
rect -8543 72725 -8509 72817
rect -8656 72691 -8509 72725
rect -7928 72721 -7855 72722
rect -8656 72628 -8622 72691
rect -8433 72687 -7855 72721
rect -9229 72594 -8622 72628
rect -8584 72623 -8426 72624
rect -8584 72589 -7925 72623
rect -8584 72586 -8426 72589
rect -8792 72489 -8654 72495
rect -8584 72489 -8546 72586
rect -7889 72525 -7855 72687
rect -8433 72491 -7855 72525
rect -7929 72490 -7855 72491
rect -8792 72451 -8546 72489
rect -8792 72441 -8654 72451
rect -8584 72256 -8546 72451
rect -7889 72441 -7855 72490
rect -9229 72222 -8546 72256
rect -8511 72401 -7855 72441
rect -8511 72256 -8471 72401
rect -8511 72222 -7925 72256
rect -8511 72221 -8425 72222
rect -10241 71974 -9771 72012
rect -10241 71951 -10187 71974
rect -10633 71672 -9777 71748
rect -8775 72041 -8721 72179
rect -8970 71903 -8891 71915
rect -8764 71903 -8730 72041
rect -8639 71985 -8585 72123
rect -8970 71836 -8730 71903
rect -8900 71831 -8730 71836
rect -10134 71388 -10049 71414
rect -12152 71345 -10049 71388
rect -10134 71322 -10049 71345
rect -12255 71147 -12183 71171
rect -12255 71077 -10776 71147
rect -12255 71066 -12183 71077
rect -12401 70875 -12114 70883
rect -12401 70841 -11520 70875
rect -12401 70840 -12114 70841
rect -12401 70798 -12358 70840
rect -12441 70792 -12358 70798
rect -12740 70758 -12358 70792
rect -12441 70754 -12358 70758
rect -12398 70706 -12358 70754
rect -12268 70668 -12213 70806
rect -12378 70625 -12162 70668
rect -11530 70663 -11452 70669
rect -12128 70629 -11452 70663
rect -11530 70627 -11452 70629
rect -12378 70359 -12338 70625
rect -12201 70569 -12162 70625
rect -12201 70565 -12108 70569
rect -12290 70383 -12235 70538
rect -12201 70531 -11520 70565
rect -12201 70527 -12108 70531
rect -12199 70467 -12110 70472
rect -11486 70471 -11452 70627
rect -11528 70467 -11452 70471
rect -12199 70433 -11452 70467
rect -12199 70430 -12110 70433
rect -12448 70354 -12338 70359
rect -12740 70320 -12338 70354
rect -12448 70314 -12338 70320
rect -12398 70113 -12343 70268
rect -12386 70076 -12352 70113
rect -12281 70048 -12245 70383
rect -12199 70260 -12163 70430
rect -11528 70429 -11452 70433
rect -10846 70809 -10776 71077
rect -11018 70775 -10776 70809
rect -10787 70677 -10679 70711
rect -11018 70579 -10910 70613
rect -10787 70481 -10679 70515
rect -11018 70383 -10910 70417
rect -12199 70256 -12104 70260
rect -12199 70222 -11520 70256
rect -12199 70218 -12104 70222
rect -10876 70265 -10816 70338
rect -10863 70204 -10822 70265
rect -10863 70193 -10643 70204
rect -10863 70165 -10635 70193
rect -10835 70143 -10635 70165
rect -11850 70048 -11780 70054
rect -12283 69978 -11780 70048
rect -11850 69810 -11780 69978
rect -11850 69776 -11608 69810
rect -11947 69678 -11839 69712
rect -11716 69580 -11608 69614
rect -11947 69482 -11839 69516
rect -11716 69384 -11608 69418
rect -11810 69266 -11750 69339
rect -10673 70004 -10635 70143
rect -10588 70056 -10517 70130
rect -10480 70068 -10172 70102
rect -11017 69970 -10635 70004
rect -10673 69808 -10635 69970
rect -11017 69774 -10635 69808
rect -10666 69591 -10612 69726
rect -10562 69715 -10523 70056
rect -10480 69970 -10172 70004
rect -10480 69872 -10172 69906
rect -10562 69645 -10522 69715
rect -10480 69676 -10172 69710
rect -10564 69644 -10522 69645
rect -10660 69571 -10620 69591
rect -11804 69205 -11763 69266
rect -11983 69194 -11763 69205
rect -11991 69166 -11763 69194
rect -11991 69144 -11791 69166
rect -12454 69069 -12146 69103
rect -12109 69057 -12038 69131
rect -12454 68971 -12146 69005
rect -12454 68873 -12146 68907
rect -12103 68716 -12064 69057
rect -11991 69005 -11953 69144
rect -11991 68971 -11609 69005
rect -11991 68809 -11953 68971
rect -11991 68775 -11609 68809
rect -12454 68677 -12146 68711
rect -12104 68646 -12064 68716
rect -12104 68645 -12062 68646
rect -12102 68419 -12062 68645
rect -10658 69364 -10622 69571
rect -10888 69193 -10680 69227
rect -10564 69129 -10524 69644
rect -10564 69096 -10350 69129
rect -10558 69095 -10350 69096
rect -10888 68997 -10680 69031
rect -10558 68899 -10350 68933
rect -10888 68801 -10680 68835
rect -10646 68683 -10586 68756
rect -10633 68639 -10592 68683
rect -10650 68580 -10500 68639
rect -10650 68514 -10035 68580
rect -9853 68514 -9777 71672
rect -8629 71638 -8595 71985
rect -8948 71595 -8595 71638
rect -8948 70891 -8905 71595
rect -8802 71155 -8730 71179
rect -8802 71085 -7323 71155
rect -8802 71074 -8730 71085
rect -8948 70883 -8661 70891
rect -8948 70849 -8067 70883
rect -8948 70848 -8661 70849
rect -8948 70806 -8905 70848
rect -8988 70800 -8905 70806
rect -9287 70766 -8905 70800
rect -8988 70762 -8905 70766
rect -8945 70714 -8905 70762
rect -8815 70676 -8760 70814
rect -8925 70633 -8709 70676
rect -8077 70671 -7999 70677
rect -8675 70637 -7999 70671
rect -8077 70635 -7999 70637
rect -8925 70367 -8885 70633
rect -8748 70577 -8709 70633
rect -8748 70573 -8655 70577
rect -8837 70391 -8782 70546
rect -8748 70539 -8067 70573
rect -8748 70535 -8655 70539
rect -8746 70475 -8657 70480
rect -8033 70479 -7999 70635
rect -8075 70475 -7999 70479
rect -8746 70441 -7999 70475
rect -8746 70438 -8657 70441
rect -8995 70362 -8885 70367
rect -9287 70328 -8885 70362
rect -8995 70322 -8885 70328
rect -8945 70121 -8890 70276
rect -8933 70084 -8899 70121
rect -8828 70056 -8792 70391
rect -8746 70268 -8710 70438
rect -8075 70437 -7999 70441
rect -7393 70817 -7323 71085
rect -7565 70783 -7323 70817
rect -7334 70685 -7226 70719
rect -7565 70587 -7457 70621
rect -7334 70489 -7226 70523
rect -7565 70391 -7457 70425
rect -8746 70264 -8651 70268
rect -8746 70230 -8067 70264
rect -8746 70226 -8651 70230
rect -7423 70273 -7363 70346
rect -7410 70212 -7369 70273
rect -7410 70201 -7190 70212
rect -7410 70173 -7182 70201
rect -7382 70151 -7182 70173
rect -8397 70056 -8327 70062
rect -8830 69986 -8327 70056
rect -8397 69818 -8327 69986
rect -8397 69784 -8155 69818
rect -8494 69686 -8386 69720
rect -8263 69588 -8155 69622
rect -8494 69490 -8386 69524
rect -8263 69392 -8155 69426
rect -8357 69274 -8297 69347
rect -7220 70012 -7182 70151
rect -7135 70064 -7064 70138
rect -7027 70076 -6719 70110
rect -7564 69978 -7182 70012
rect -7220 69816 -7182 69978
rect -7564 69782 -7182 69816
rect -7213 69599 -7159 69734
rect -7109 69723 -7070 70064
rect -7027 69978 -6719 70012
rect -7027 69880 -6719 69914
rect -7109 69653 -7069 69723
rect -7027 69684 -6719 69718
rect -7111 69652 -7069 69653
rect -7207 69579 -7167 69599
rect -8351 69213 -8310 69274
rect -8530 69202 -8310 69213
rect -8538 69174 -8310 69202
rect -8538 69152 -8338 69174
rect -9001 69077 -8693 69111
rect -8656 69065 -8585 69139
rect -9001 68979 -8693 69013
rect -9001 68881 -8693 68915
rect -8650 68724 -8611 69065
rect -8538 69013 -8500 69152
rect -8538 68979 -8156 69013
rect -8538 68817 -8500 68979
rect -8538 68783 -8156 68817
rect -9001 68685 -8693 68719
rect -8651 68654 -8611 68724
rect -8651 68653 -8609 68654
rect -8649 68514 -8609 68653
rect -7205 69372 -7169 69579
rect -7435 69201 -7227 69235
rect -7111 69137 -7071 69652
rect -7111 69104 -6897 69137
rect -7105 69103 -6897 69104
rect -7435 69005 -7227 69039
rect -7105 68907 -6897 68941
rect -10650 68509 -8609 68514
rect -10609 68504 -8609 68509
rect -10111 68438 -8609 68504
rect -13775 67928 -13628 67962
rect -9645 67928 -9499 68438
rect -8649 68427 -8609 68438
rect -13775 67782 -9499 67928
rect -13775 67759 -13628 67782
rect -12421 67023 -12378 67136
rect -12458 66800 -12288 67023
rect -12421 66111 -12378 66800
rect -12275 66375 -12203 66399
rect -12275 66305 -10796 66375
rect -12275 66294 -12203 66305
rect -12421 66103 -12134 66111
rect -12421 66069 -11540 66103
rect -12421 66068 -12134 66069
rect -12421 66026 -12378 66068
rect -12461 66020 -12378 66026
rect -12760 65986 -12378 66020
rect -12461 65982 -12378 65986
rect -12418 65934 -12378 65982
rect -12288 65896 -12233 66034
rect -12398 65853 -12182 65896
rect -11550 65891 -11472 65897
rect -12148 65857 -11472 65891
rect -11550 65855 -11472 65857
rect -12398 65587 -12358 65853
rect -12221 65797 -12182 65853
rect -12221 65793 -12128 65797
rect -12310 65611 -12255 65766
rect -12221 65759 -11540 65793
rect -12221 65755 -12128 65759
rect -12219 65695 -12130 65700
rect -11506 65699 -11472 65855
rect -11548 65695 -11472 65699
rect -12219 65661 -11472 65695
rect -12219 65658 -12130 65661
rect -12468 65582 -12358 65587
rect -12760 65548 -12358 65582
rect -12468 65542 -12358 65548
rect -12418 65341 -12363 65496
rect -12406 65304 -12372 65341
rect -12301 65276 -12265 65611
rect -12219 65488 -12183 65658
rect -11548 65657 -11472 65661
rect -10866 66037 -10796 66305
rect -11038 66003 -10796 66037
rect -10807 65905 -10699 65939
rect -7435 68809 -7227 68843
rect -7193 68691 -7133 68764
rect -7180 68647 -7139 68691
rect -7197 68517 -7047 68647
rect -6834 67871 -6567 68228
rect -6789 67050 -6600 67871
rect -6800 66693 -6533 67050
rect -11038 65807 -10930 65841
rect -10807 65709 -10699 65743
rect -11038 65611 -10930 65645
rect -12219 65484 -12124 65488
rect -12219 65450 -11540 65484
rect -12219 65446 -12124 65450
rect -10896 65493 -10836 65566
rect -10883 65432 -10842 65493
rect -10883 65421 -10663 65432
rect -10883 65393 -10655 65421
rect -10855 65371 -10655 65393
rect -11870 65276 -11800 65282
rect -12303 65206 -11800 65276
rect -11870 65038 -11800 65206
rect -11870 65004 -11628 65038
rect -11967 64906 -11859 64940
rect -11736 64808 -11628 64842
rect -11967 64710 -11859 64744
rect -11736 64612 -11628 64646
rect -11830 64494 -11770 64567
rect -10693 65232 -10655 65371
rect -10608 65284 -10537 65358
rect -10500 65296 -10192 65330
rect -11037 65198 -10655 65232
rect -10693 65036 -10655 65198
rect -11037 65002 -10655 65036
rect -10686 64819 -10632 64954
rect -10582 64943 -10543 65284
rect -10500 65198 -10192 65232
rect -10500 65100 -10192 65134
rect -10582 64873 -10542 64943
rect -10500 64904 -10192 64938
rect -10584 64872 -10542 64873
rect -10680 64799 -10640 64819
rect -11824 64433 -11783 64494
rect -12003 64422 -11783 64433
rect -12011 64394 -11783 64422
rect -12011 64372 -11811 64394
rect -12474 64297 -12166 64331
rect -12129 64285 -12058 64359
rect -12474 64199 -12166 64233
rect -12474 64101 -12166 64135
rect -12123 63944 -12084 64285
rect -12011 64233 -11973 64372
rect -12011 64199 -11629 64233
rect -12011 64037 -11973 64199
rect -12011 64003 -11629 64037
rect -12474 63905 -12166 63939
rect -12124 63874 -12084 63944
rect -12124 63873 -12082 63874
rect -12122 63647 -12082 63873
rect -10678 64592 -10642 64799
rect -10908 64421 -10700 64455
rect -10584 64357 -10544 64872
rect -9798 65283 -8827 65321
rect -10584 64324 -10370 64357
rect -10578 64323 -10370 64324
rect -10908 64225 -10700 64259
rect -10578 64127 -10370 64161
rect -10908 64029 -10700 64063
rect -12390 63147 -12098 63190
rect -12390 62443 -12347 63147
rect -12141 62948 -12098 63147
rect -10666 63911 -10606 63984
rect -10653 63867 -10612 63911
rect -10670 63840 -10520 63867
rect -10720 63764 -10520 63840
rect -10670 63737 -10520 63764
rect -10622 63308 -10546 63737
rect -10230 63572 -10176 63584
rect -9798 63572 -9760 65283
rect -8865 65067 -8827 65283
rect -8915 65063 -8297 65067
rect -9218 65029 -8297 65063
rect -8717 64914 -8658 64968
rect -8709 64862 -8675 64914
rect -8560 64862 -8506 64994
rect -8334 64967 -8297 65029
rect -8334 64965 -8204 64967
rect -8334 64931 -7914 64965
rect -8334 64930 -8204 64931
rect -8714 64835 -8428 64862
rect -9218 64828 -8428 64835
rect -9218 64801 -8680 64828
rect -8714 64800 -8680 64801
rect -9218 64703 -8710 64737
rect -8643 64736 -8505 64790
rect -8462 64737 -8428 64828
rect -8462 64703 -7914 64737
rect -8541 64526 -8487 64664
rect -9218 64377 -8679 64411
rect -8714 64286 -8679 64377
rect -8628 64351 -8574 64489
rect -8532 64411 -8498 64526
rect -8532 64377 -7914 64411
rect -9218 64252 -8679 64286
rect -8532 64285 -8498 64377
rect -8645 64251 -8498 64285
rect -7917 64281 -7844 64282
rect -8645 64188 -8611 64251
rect -8422 64247 -7844 64281
rect -9218 64154 -8611 64188
rect -8573 64183 -8415 64184
rect -8573 64149 -7914 64183
rect -8573 64146 -8415 64149
rect -8781 64049 -8643 64055
rect -8573 64049 -8535 64146
rect -7878 64085 -7844 64247
rect -8422 64051 -7844 64085
rect -7918 64050 -7844 64051
rect -8781 64011 -8535 64049
rect -8781 64001 -8643 64011
rect -8573 63816 -8535 64011
rect -7878 64001 -7844 64050
rect -9218 63782 -8535 63816
rect -8500 63961 -7844 64001
rect -8500 63816 -8460 63961
rect -8500 63782 -7914 63816
rect -8500 63781 -8414 63782
rect -10230 63534 -9760 63572
rect -10230 63511 -10176 63534
rect -10622 63232 -9766 63308
rect -8764 63601 -8710 63739
rect -8959 63463 -8880 63475
rect -8753 63463 -8719 63601
rect -8628 63545 -8574 63683
rect -8959 63396 -8719 63463
rect -8889 63391 -8719 63396
rect -10123 62948 -10038 62974
rect -12141 62905 -10038 62948
rect -10123 62882 -10038 62905
rect -12244 62707 -12172 62731
rect -12244 62637 -10765 62707
rect -12244 62626 -12172 62637
rect -12390 62435 -12103 62443
rect -12390 62401 -11509 62435
rect -12390 62400 -12103 62401
rect -12390 62358 -12347 62400
rect -12430 62352 -12347 62358
rect -12729 62318 -12347 62352
rect -12430 62314 -12347 62318
rect -12387 62266 -12347 62314
rect -12257 62228 -12202 62366
rect -12367 62185 -12151 62228
rect -11519 62223 -11441 62229
rect -12117 62189 -11441 62223
rect -11519 62187 -11441 62189
rect -12367 61919 -12327 62185
rect -12190 62129 -12151 62185
rect -12190 62125 -12097 62129
rect -12279 61943 -12224 62098
rect -12190 62091 -11509 62125
rect -12190 62087 -12097 62091
rect -12188 62027 -12099 62032
rect -11475 62031 -11441 62187
rect -11517 62027 -11441 62031
rect -12188 61993 -11441 62027
rect -12188 61990 -12099 61993
rect -12437 61914 -12327 61919
rect -12729 61880 -12327 61914
rect -12437 61874 -12327 61880
rect -12387 61673 -12332 61828
rect -12375 61636 -12341 61673
rect -12270 61608 -12234 61943
rect -12188 61820 -12152 61990
rect -11517 61989 -11441 61993
rect -10835 62369 -10765 62637
rect -11007 62335 -10765 62369
rect -10776 62237 -10668 62271
rect -11007 62139 -10899 62173
rect -10776 62041 -10668 62075
rect -11007 61943 -10899 61977
rect -12188 61816 -12093 61820
rect -12188 61782 -11509 61816
rect -12188 61778 -12093 61782
rect -10865 61825 -10805 61898
rect -10852 61764 -10811 61825
rect -10852 61753 -10632 61764
rect -10852 61725 -10624 61753
rect -10824 61703 -10624 61725
rect -11839 61608 -11769 61614
rect -12272 61538 -11769 61608
rect -11839 61370 -11769 61538
rect -11839 61336 -11597 61370
rect -11936 61238 -11828 61272
rect -11705 61140 -11597 61174
rect -11936 61042 -11828 61076
rect -11705 60944 -11597 60978
rect -11799 60826 -11739 60899
rect -10662 61564 -10624 61703
rect -10577 61616 -10506 61690
rect -10469 61628 -10161 61662
rect -11006 61530 -10624 61564
rect -10662 61368 -10624 61530
rect -11006 61334 -10624 61368
rect -10655 61151 -10601 61286
rect -10551 61275 -10512 61616
rect -10469 61530 -10161 61564
rect -10469 61432 -10161 61466
rect -10551 61205 -10511 61275
rect -10469 61236 -10161 61270
rect -10553 61204 -10511 61205
rect -10649 61131 -10609 61151
rect -11793 60765 -11752 60826
rect -11972 60754 -11752 60765
rect -11980 60726 -11752 60754
rect -11980 60704 -11780 60726
rect -12443 60629 -12135 60663
rect -12098 60617 -12027 60691
rect -12443 60531 -12135 60565
rect -12443 60433 -12135 60467
rect -12092 60276 -12053 60617
rect -11980 60565 -11942 60704
rect -11980 60531 -11598 60565
rect -11980 60369 -11942 60531
rect -11980 60335 -11598 60369
rect -12443 60237 -12135 60271
rect -12093 60206 -12053 60276
rect -12093 60205 -12051 60206
rect -12091 59979 -12051 60205
rect -10647 60924 -10611 61131
rect -10877 60753 -10669 60787
rect -10553 60689 -10513 61204
rect -10553 60656 -10339 60689
rect -10547 60655 -10339 60656
rect -10877 60557 -10669 60591
rect -10547 60459 -10339 60493
rect -10877 60361 -10669 60395
rect -10635 60243 -10575 60316
rect -10622 60199 -10581 60243
rect -10639 60140 -10489 60199
rect -10639 60074 -10024 60140
rect -9842 60074 -9766 63232
rect -8618 63198 -8584 63545
rect -8937 63155 -8584 63198
rect -8937 62451 -8894 63155
rect -8791 62715 -8719 62739
rect -8791 62645 -7312 62715
rect -8791 62634 -8719 62645
rect -8937 62443 -8650 62451
rect -8937 62409 -8056 62443
rect -8937 62408 -8650 62409
rect -8937 62366 -8894 62408
rect -8977 62360 -8894 62366
rect -9276 62326 -8894 62360
rect -8977 62322 -8894 62326
rect -8934 62274 -8894 62322
rect -8804 62236 -8749 62374
rect -8914 62193 -8698 62236
rect -8066 62231 -7988 62237
rect -8664 62197 -7988 62231
rect -8066 62195 -7988 62197
rect -8914 61927 -8874 62193
rect -8737 62137 -8698 62193
rect -8737 62133 -8644 62137
rect -8826 61951 -8771 62106
rect -8737 62099 -8056 62133
rect -8737 62095 -8644 62099
rect -8735 62035 -8646 62040
rect -8022 62039 -7988 62195
rect -8064 62035 -7988 62039
rect -8735 62001 -7988 62035
rect -8735 61998 -8646 62001
rect -8984 61922 -8874 61927
rect -9276 61888 -8874 61922
rect -8984 61882 -8874 61888
rect -8934 61681 -8879 61836
rect -8922 61644 -8888 61681
rect -8817 61616 -8781 61951
rect -8735 61828 -8699 61998
rect -8064 61997 -7988 62001
rect -7382 62377 -7312 62645
rect -7554 62343 -7312 62377
rect -7323 62245 -7215 62279
rect -7554 62147 -7446 62181
rect -7323 62049 -7215 62083
rect -7554 61951 -7446 61985
rect -8735 61824 -8640 61828
rect -8735 61790 -8056 61824
rect -8735 61786 -8640 61790
rect -7412 61833 -7352 61906
rect -7399 61772 -7358 61833
rect -7399 61761 -7179 61772
rect -7399 61733 -7171 61761
rect -7371 61711 -7171 61733
rect -8386 61616 -8316 61622
rect -8819 61546 -8316 61616
rect -8386 61378 -8316 61546
rect -8386 61344 -8144 61378
rect -8483 61246 -8375 61280
rect -8252 61148 -8144 61182
rect -8483 61050 -8375 61084
rect -8252 60952 -8144 60986
rect -8346 60834 -8286 60907
rect -7209 61572 -7171 61711
rect -7124 61624 -7053 61698
rect -7016 61636 -6708 61670
rect -7553 61538 -7171 61572
rect -7209 61376 -7171 61538
rect -7553 61342 -7171 61376
rect -7098 61283 -7059 61624
rect -7016 61538 -6708 61572
rect -7016 61440 -6708 61474
rect -7098 61213 -7058 61283
rect -7016 61244 -6708 61278
rect -7100 61212 -7058 61213
rect -8340 60773 -8299 60834
rect -8519 60762 -8299 60773
rect -8527 60734 -8299 60762
rect -8527 60712 -8327 60734
rect -8990 60637 -8682 60671
rect -8645 60625 -8574 60699
rect -8990 60539 -8682 60573
rect -8990 60441 -8682 60475
rect -8639 60284 -8600 60625
rect -8527 60573 -8489 60712
rect -8527 60539 -8145 60573
rect -8527 60377 -8489 60539
rect -8527 60343 -8145 60377
rect -8990 60245 -8682 60279
rect -8640 60214 -8600 60284
rect -8640 60213 -8598 60214
rect -8638 60074 -8598 60213
rect -7424 60761 -7216 60795
rect -7100 60697 -7060 61212
rect -7100 60664 -6886 60697
rect -7094 60663 -6886 60664
rect -7424 60565 -7216 60599
rect -7094 60467 -6886 60501
rect -7424 60369 -7216 60403
rect -7182 60251 -7122 60324
rect -10639 60069 -8598 60074
rect -10598 60064 -8598 60069
rect -10100 59998 -8598 60064
rect -13776 59348 -13608 59367
rect -9856 59348 -9710 59998
rect -8638 59987 -8598 59998
rect -13776 59291 -9710 59348
rect -13777 59202 -9710 59291
rect -13777 57336 -13606 59202
rect -7169 60207 -7128 60251
rect -7186 60077 -7036 60207
rect -10483 57985 -10449 57988
rect -10499 57867 -10441 57985
rect -10483 57820 -10449 57867
rect -11277 57786 -9684 57820
rect -10506 57611 -10452 57745
rect -10498 57420 -10459 57611
rect -11277 57386 -9684 57420
rect -10509 57226 -10455 57339
rect -10509 57156 -10268 57226
rect -10511 56971 -10453 57089
rect -10499 56820 -10465 56971
rect -11277 56786 -9684 56820
rect -10504 56618 -10450 56752
rect -8424 57981 -8287 57982
rect -8819 57980 -7871 57981
rect -8821 57974 -7871 57980
rect -8821 57933 -7841 57974
rect -8821 57898 -8782 57933
rect -8424 57922 -8287 57933
rect -8830 57868 -8760 57898
rect -8903 57862 -8699 57868
rect -9095 57828 -8607 57862
rect -8903 57822 -8699 57828
rect -8838 57672 -8792 57822
rect -8903 57666 -8699 57672
rect -9095 57632 -8607 57666
rect -8903 57626 -8699 57632
rect -8838 57476 -8792 57626
rect -7915 57806 -7841 57933
rect -7965 57764 -7573 57770
rect -8057 57730 -7569 57764
rect -7965 57724 -7573 57730
rect -9091 57470 -8699 57476
rect -9095 57436 -8607 57470
rect -9091 57430 -8699 57436
rect -8823 57226 -8749 57394
rect -8441 57245 -8402 57651
rect -8817 57029 -8764 57226
rect -8454 57113 -8394 57245
rect -8980 57028 -8694 57029
rect -8980 57024 -8651 57028
rect -10497 56420 -10458 56618
rect -11277 56386 -9684 56420
rect -10502 56235 -10448 56339
rect -10502 56165 -10267 56235
rect -10484 55894 -10426 56012
rect -10472 55820 -10438 55894
rect -11277 55786 -9684 55820
rect -10489 55618 -10435 55752
rect -10482 55420 -10448 55618
rect -11277 55386 -9684 55420
rect -10504 55191 -10450 55350
rect -11083 55121 -9716 55191
rect -11083 54938 -11013 55121
rect -9080 56990 -8557 57024
rect -8980 56987 -8651 56990
rect -9148 56926 -9063 56931
rect -9148 56892 -8972 56926
rect -9148 56889 -9063 56892
rect -9148 56735 -9114 56889
rect -8936 56854 -8701 56987
rect -8569 56926 -8477 56932
rect -8665 56892 -8477 56926
rect -8569 56888 -8477 56892
rect -8936 56829 -8902 56854
rect -8990 56828 -8902 56829
rect -9080 56794 -8902 56828
rect -8990 56793 -8902 56794
rect -9148 56730 -9058 56735
rect -9148 56696 -8972 56730
rect -9148 56693 -9058 56696
rect -9148 56541 -9114 56693
rect -8936 56635 -8902 56793
rect -8990 56632 -8902 56635
rect -9080 56599 -8902 56632
rect -9080 56598 -8972 56599
rect -9148 56534 -9059 56541
rect -9148 56500 -8972 56534
rect -9148 56499 -9059 56500
rect -9148 56339 -9114 56499
rect -8936 56437 -8902 56599
rect -8735 56831 -8701 56854
rect -8735 56828 -8652 56831
rect -8735 56794 -8557 56828
rect -8735 56790 -8652 56794
rect -8735 56637 -8701 56790
rect -8511 56735 -8477 56888
rect -8580 56730 -8477 56735
rect -8665 56696 -8477 56730
rect -8580 56691 -8477 56696
rect -8735 56632 -8652 56637
rect -8735 56598 -8557 56632
rect -8735 56596 -8652 56598
rect -8988 56436 -8902 56437
rect -9080 56402 -8902 56436
rect -8988 56401 -8902 56402
rect -8848 56345 -8774 56470
rect -8735 56439 -8701 56596
rect -8511 56539 -8477 56691
rect -8580 56534 -8477 56539
rect -8665 56500 -8477 56534
rect -8580 56495 -8477 56500
rect -8735 56436 -8660 56439
rect -8735 56402 -8557 56436
rect -8735 56398 -8660 56402
rect -9148 56338 -9069 56339
rect -8995 56338 -8639 56345
rect -8511 56343 -8477 56495
rect -8569 56338 -8477 56343
rect -9148 56304 -8477 56338
rect -9148 56303 -9069 56304
rect -8995 56298 -8639 56304
rect -8569 56299 -8477 56304
rect -9022 56253 -8854 56254
rect -9022 56180 -8760 56253
rect -8830 56125 -8760 56180
rect -8903 56119 -8699 56125
rect -9095 56085 -8607 56119
rect -8903 56079 -8699 56085
rect -8838 55929 -8792 56079
rect -8903 55923 -8699 55929
rect -9095 55889 -8607 55923
rect -8903 55883 -8699 55889
rect -8838 55733 -8792 55883
rect -9091 55727 -8699 55733
rect -9095 55693 -8607 55727
rect -9091 55687 -8699 55693
rect -9073 55472 -8909 55529
rect -8995 55313 -8950 55472
rect -8995 55308 -8771 55313
rect -8995 55268 -8656 55308
rect -8816 55248 -8656 55268
rect -8816 55198 -8771 55248
rect -8830 55168 -8760 55198
rect -8903 55162 -8699 55168
rect -9095 55128 -8607 55162
rect -8903 55122 -8699 55128
rect -11156 54932 -10952 54938
rect -11348 54898 -10860 54932
rect -11156 54892 -10952 54898
rect -11091 54742 -11045 54892
rect -10230 54896 -10096 54956
rect -10217 54800 -10156 54896
rect -11156 54736 -10952 54742
rect -11348 54702 -10860 54736
rect -11156 54696 -10952 54702
rect -11091 54546 -11045 54696
rect -10501 54786 -10084 54800
rect -10501 54766 -9639 54786
rect -10121 54752 -9639 54766
rect -11344 54540 -10952 54546
rect -11348 54506 -10860 54540
rect -11344 54500 -10952 54506
rect -10556 54668 -10293 54702
rect -10556 54590 -10521 54668
rect -10242 54591 -10188 54726
rect -10556 54556 -10293 54590
rect -10233 54497 -10194 54591
rect -10121 54590 -10083 54752
rect -8838 54972 -8792 55122
rect -8903 54966 -8699 54972
rect -9095 54932 -8607 54966
rect -8903 54926 -8699 54932
rect -8838 54776 -8792 54926
rect -9091 54770 -8699 54776
rect -9095 54736 -8607 54770
rect -9091 54730 -8699 54736
rect -10121 54556 -9639 54590
rect -11076 54296 -11002 54464
rect -10234 54443 -10194 54497
rect -10247 54442 -10189 54443
rect -10248 54283 -10188 54442
rect -10144 54373 -10090 54508
rect -8823 54526 -8749 54694
rect -10136 54353 -10096 54373
rect -10892 53923 -10832 54054
rect -10133 54062 -10097 54353
rect -8814 54329 -8757 54526
rect -8980 54328 -8694 54329
rect -8980 54327 -8651 54328
rect -8980 54324 -8529 54327
rect -9764 54178 -9632 54193
rect -9449 54178 -9317 54196
rect -10868 53811 -10832 53923
rect -11355 53777 -10439 53811
rect -10147 53930 -10087 54062
rect -9764 54043 -9317 54178
rect -9764 54033 -9632 54043
rect -9449 54036 -9317 54043
rect -10946 53607 -10892 53742
rect -10936 53202 -10899 53607
rect -10845 53364 -10439 53398
rect -10845 53202 -10811 53364
rect -10747 53266 -10307 53300
rect -11111 53168 -10439 53202
rect -11111 53165 -10811 53168
rect -11111 53073 -11074 53165
rect -11355 53039 -11074 53073
rect -11111 52877 -11074 53039
rect -10948 52996 -10894 53131
rect -10341 53090 -10307 53266
rect -10450 53089 -10307 53090
rect -10747 53055 -10307 53089
rect -11355 52843 -11074 52877
rect -11111 52681 -11074 52843
rect -11026 52808 -10972 52943
rect -11355 52647 -11074 52681
rect -11108 52472 -11054 52607
rect -11100 52453 -11063 52472
rect -11098 52400 -11063 52453
rect -11195 52340 -11063 52400
rect -11017 52285 -10979 52808
rect -10935 52494 -10901 52996
rect -10845 52991 -10747 52992
rect -10845 52957 -10439 52991
rect -10845 52779 -10810 52957
rect -10344 52894 -10307 53055
rect -10448 52893 -10307 52894
rect -10747 52859 -10307 52893
rect -10845 52745 -10440 52779
rect -10845 52583 -10811 52745
rect -10845 52549 -10440 52583
rect -9080 54290 -8529 54324
rect -8980 54287 -8529 54290
rect -9148 54226 -9063 54231
rect -9148 54192 -8972 54226
rect -9148 54189 -9063 54192
rect -9148 54035 -9114 54189
rect -8936 54154 -8701 54287
rect -8661 54281 -8529 54287
rect -8569 54226 -8477 54232
rect -8665 54192 -8477 54226
rect -8569 54188 -8477 54192
rect -8936 54129 -8902 54154
rect -8990 54128 -8902 54129
rect -9080 54094 -8902 54128
rect -8990 54093 -8902 54094
rect -9148 54030 -9058 54035
rect -9148 53996 -8972 54030
rect -9148 53993 -9058 53996
rect -9148 53841 -9114 53993
rect -8936 53935 -8902 54093
rect -8990 53932 -8902 53935
rect -9080 53899 -8902 53932
rect -9080 53898 -8972 53899
rect -9148 53834 -9059 53841
rect -9148 53800 -8972 53834
rect -9148 53799 -9059 53800
rect -9148 53639 -9114 53799
rect -8936 53737 -8902 53899
rect -8735 54131 -8701 54154
rect -8735 54128 -8652 54131
rect -8735 54094 -8557 54128
rect -8735 54090 -8652 54094
rect -8735 53937 -8701 54090
rect -8511 54035 -8477 54188
rect -8580 54030 -8477 54035
rect -8665 53996 -8477 54030
rect -8580 53991 -8477 53996
rect -8735 53932 -8652 53937
rect -8735 53898 -8557 53932
rect -8735 53896 -8652 53898
rect -8988 53736 -8902 53737
rect -9080 53702 -8902 53736
rect -8988 53701 -8902 53702
rect -8848 53645 -8774 53770
rect -8735 53739 -8701 53896
rect -8511 53839 -8477 53991
rect -8580 53834 -8477 53839
rect -8665 53800 -8477 53834
rect -8580 53795 -8477 53800
rect -8735 53736 -8660 53739
rect -8735 53702 -8557 53736
rect -8735 53698 -8660 53702
rect -9148 53638 -9069 53639
rect -8995 53638 -8639 53645
rect -8511 53643 -8477 53795
rect -8569 53638 -8477 53643
rect -9148 53604 -8477 53638
rect -9148 53603 -9069 53604
rect -8995 53598 -8639 53604
rect -8569 53599 -8477 53604
rect -9022 53553 -8854 53554
rect -9022 53480 -8760 53553
rect -8830 53425 -8760 53480
rect -8903 53419 -8699 53425
rect -9095 53385 -8607 53419
rect -8903 53379 -8699 53385
rect -8838 53229 -8792 53379
rect -8903 53223 -8699 53229
rect -9095 53189 -8607 53223
rect -8903 53183 -8699 53189
rect -8838 53033 -8792 53183
rect -9091 53027 -8699 53033
rect -9095 52993 -8607 53027
rect -9091 52987 -8699 52993
rect -10935 52460 -10669 52494
rect -10935 52455 -10901 52460
rect -11017 52225 -10813 52285
rect -10714 52185 -10669 52460
rect -11395 52172 -11293 52179
rect -10959 52172 -10669 52185
rect -11395 52138 -10669 52172
rect -11395 52133 -11293 52138
rect -10959 52135 -10669 52138
rect -11395 51981 -11357 52133
rect -10714 52079 -10669 52135
rect -10923 52074 -10843 52078
rect -11321 52040 -10843 52074
rect -10923 52033 -10843 52040
rect -11395 51976 -11293 51981
rect -11395 51942 -10913 51976
rect -11395 51935 -11293 51942
rect -10879 51766 -10843 52033
rect -10804 51860 -10744 52003
rect -10705 51869 -10669 52079
rect -9073 52772 -8909 52829
rect -8823 52783 -8749 52951
rect -8812 52748 -8754 52783
rect -8808 52691 -8766 52748
rect -8812 52631 -8680 52691
rect -8808 52573 -8766 52631
rect -8830 52543 -8760 52573
rect -8903 52537 -8699 52543
rect -9095 52503 -8607 52537
rect -8903 52497 -8699 52503
rect -8838 52347 -8792 52497
rect -8441 52722 -8402 57113
rect -7872 57574 -7826 57724
rect -7965 57568 -7761 57574
rect -8057 57534 -7569 57568
rect -7965 57528 -7761 57534
rect -7872 57378 -7826 57528
rect -7965 57372 -7761 57378
rect -8057 57338 -7569 57372
rect -7965 57332 -7761 57338
rect -7904 57291 -7834 57332
rect -7904 57245 -7655 57291
rect -8059 57172 -7853 57209
rect -8059 57149 -7852 57172
rect -7915 57137 -7852 57149
rect -7704 57148 -7655 57245
rect -7915 56969 -7841 57137
rect -7755 57091 -7591 57148
rect -7965 56927 -7573 56933
rect -8057 56893 -7569 56927
rect -7965 56887 -7573 56893
rect -7872 56737 -7826 56887
rect -7965 56731 -7761 56737
rect -8057 56697 -7569 56731
rect -7965 56691 -7761 56697
rect -7872 56541 -7826 56691
rect -7965 56535 -7761 56541
rect -8057 56501 -7569 56535
rect -7965 56495 -7761 56501
rect -7904 56440 -7834 56495
rect -7904 56367 -7642 56440
rect -7810 56366 -7642 56367
rect -8187 56316 -8095 56321
rect -8025 56316 -7669 56322
rect -7595 56316 -7516 56317
rect -8187 56282 -7516 56316
rect -8187 56277 -8095 56282
rect -8187 56125 -8153 56277
rect -8025 56275 -7669 56282
rect -7595 56281 -7516 56282
rect -8004 56218 -7929 56222
rect -8107 56184 -7929 56218
rect -8004 56181 -7929 56184
rect -8187 56120 -8084 56125
rect -8187 56086 -7999 56120
rect -8187 56081 -8084 56086
rect -8187 55929 -8153 56081
rect -7963 56024 -7929 56181
rect -7890 56150 -7816 56275
rect -7762 56218 -7676 56219
rect -7762 56184 -7584 56218
rect -7762 56183 -7676 56184
rect -8012 56022 -7929 56024
rect -8107 55988 -7929 56022
rect -8012 55983 -7929 55988
rect -8187 55924 -8084 55929
rect -8187 55890 -7999 55924
rect -8187 55885 -8084 55890
rect -8187 55732 -8153 55885
rect -7963 55830 -7929 55983
rect -8012 55826 -7929 55830
rect -8107 55792 -7929 55826
rect -8012 55789 -7929 55792
rect -7963 55766 -7929 55789
rect -7762 56021 -7728 56183
rect -7550 56121 -7516 56281
rect -7605 56120 -7516 56121
rect -7692 56086 -7516 56120
rect -7605 56079 -7516 56086
rect -7692 56021 -7584 56022
rect -7762 55988 -7584 56021
rect -7762 55985 -7674 55988
rect -7762 55827 -7728 55985
rect -7550 55927 -7516 56079
rect -7606 55924 -7516 55927
rect -7692 55890 -7516 55924
rect -7606 55885 -7516 55890
rect -7762 55826 -7674 55827
rect -7762 55792 -7584 55826
rect -7762 55791 -7674 55792
rect -7762 55766 -7728 55791
rect -8187 55728 -8095 55732
rect -8187 55694 -7999 55728
rect -8187 55688 -8095 55694
rect -7963 55633 -7728 55766
rect -7550 55731 -7516 55885
rect -7601 55728 -7516 55731
rect -7692 55694 -7516 55728
rect -7601 55689 -7516 55694
rect -8013 55630 -7684 55633
rect -8107 55596 -7584 55630
rect -8013 55592 -7684 55596
rect -7970 55591 -7684 55592
rect -7929 55500 -7869 55591
rect -7908 55274 -7848 55296
rect -7915 55106 -7841 55274
rect -7965 55064 -7573 55070
rect -8057 55030 -7569 55064
rect -7965 55024 -7573 55030
rect -8452 52590 -8392 52722
rect -8903 52341 -8699 52347
rect -9095 52307 -8607 52341
rect -8903 52301 -8699 52307
rect -8838 52151 -8792 52301
rect -9091 52145 -8699 52151
rect -9095 52111 -8607 52145
rect -9091 52105 -8699 52111
rect -10705 51863 -10620 51869
rect -10918 51765 -10843 51766
rect -11321 51731 -10843 51765
rect -10918 51730 -10843 51731
rect -10797 51577 -10761 51860
rect -10705 51829 -10421 51863
rect -7872 54874 -7826 55024
rect -7965 54868 -7761 54874
rect -8057 54834 -7569 54868
rect -7965 54828 -7761 54834
rect -7872 54678 -7826 54828
rect -7965 54672 -7761 54678
rect -8057 54638 -7569 54672
rect -7965 54632 -7761 54638
rect -7904 54596 -7834 54632
rect -7904 54534 -7643 54596
rect -7705 54448 -7643 54534
rect -7755 54391 -7591 54448
rect -7965 54227 -7573 54233
rect -8057 54193 -7569 54227
rect -7965 54187 -7573 54193
rect -7872 54037 -7826 54187
rect -7965 54031 -7761 54037
rect -8057 53997 -7569 54031
rect -7965 53991 -7761 53997
rect -7872 53841 -7826 53991
rect -7965 53835 -7761 53841
rect -8057 53801 -7569 53835
rect -7965 53795 -7761 53801
rect -7904 53740 -7834 53795
rect -7904 53667 -7642 53740
rect -7810 53666 -7642 53667
rect -8187 53616 -8095 53621
rect -8025 53616 -7669 53622
rect -7595 53616 -7516 53617
rect -8187 53582 -7516 53616
rect -8187 53577 -8095 53582
rect -8187 53425 -8153 53577
rect -8025 53575 -7669 53582
rect -7595 53581 -7516 53582
rect -8004 53518 -7929 53522
rect -8107 53484 -7929 53518
rect -8004 53481 -7929 53484
rect -8187 53420 -8084 53425
rect -8187 53386 -7999 53420
rect -8187 53381 -8084 53386
rect -8187 53229 -8153 53381
rect -7963 53324 -7929 53481
rect -7890 53450 -7816 53575
rect -7762 53518 -7676 53519
rect -7762 53484 -7584 53518
rect -7762 53483 -7676 53484
rect -8012 53322 -7929 53324
rect -8107 53288 -7929 53322
rect -8012 53283 -7929 53288
rect -8187 53224 -8084 53229
rect -8187 53190 -7999 53224
rect -8187 53185 -8084 53190
rect -8187 53032 -8153 53185
rect -7963 53130 -7929 53283
rect -8012 53126 -7929 53130
rect -8107 53092 -7929 53126
rect -8012 53089 -7929 53092
rect -7963 53066 -7929 53089
rect -7762 53321 -7728 53483
rect -7550 53421 -7516 53581
rect -7605 53420 -7516 53421
rect -7692 53386 -7516 53420
rect -7605 53379 -7516 53386
rect -7692 53321 -7584 53322
rect -7762 53288 -7584 53321
rect -7762 53285 -7674 53288
rect -7762 53127 -7728 53285
rect -7550 53227 -7516 53379
rect -7606 53224 -7516 53227
rect -7692 53190 -7516 53224
rect -7606 53185 -7516 53190
rect -7762 53126 -7674 53127
rect -7762 53092 -7584 53126
rect -7762 53091 -7674 53092
rect -7762 53066 -7728 53091
rect -8187 53028 -8095 53032
rect -8187 52994 -7999 53028
rect -8187 52988 -8095 52994
rect -7963 52933 -7728 53066
rect -7550 53031 -7516 53185
rect -7601 53028 -7516 53031
rect -7692 52994 -7516 53028
rect -7601 52989 -7516 52994
rect -8013 52930 -7684 52933
rect -8107 52896 -7584 52930
rect -8013 52892 -7684 52896
rect -7970 52891 -7684 52892
rect -7931 52816 -7871 52891
rect -10705 51824 -10620 51829
rect -10724 51637 -10664 51783
rect -10708 51578 -10672 51637
rect -10730 51272 -10670 51321
rect -10730 51239 -10669 51272
rect -11395 51226 -11293 51233
rect -10959 51226 -10669 51239
rect -11395 51192 -10669 51226
rect -11395 51187 -11293 51192
rect -10959 51189 -10669 51192
rect -11395 51035 -11357 51187
rect -10714 51133 -10669 51189
rect -10923 51128 -10843 51132
rect -11321 51094 -10843 51128
rect -10923 51087 -10843 51094
rect -11395 51030 -11293 51035
rect -11395 50996 -10913 51030
rect -11395 50989 -11293 50996
rect -10879 50820 -10843 51087
rect -10804 50914 -10744 51057
rect -10705 50923 -10669 51133
rect -8105 51573 -8045 51670
rect -10705 50917 -10620 50923
rect -10918 50819 -10843 50820
rect -11321 50785 -10843 50819
rect -10918 50784 -10843 50785
rect -10797 50492 -10761 50914
rect -10705 50883 -10421 50917
rect -10705 50878 -10620 50883
rect -10724 50691 -10664 50837
rect -11012 50456 -10761 50492
rect -12933 49853 -12796 49854
rect -13349 49852 -12401 49853
rect -13349 49846 -12399 49852
rect -13379 49805 -12399 49846
rect -13379 49678 -13305 49805
rect -12933 49794 -12796 49805
rect -12438 49770 -12399 49805
rect -12460 49740 -12390 49770
rect -13647 49636 -13255 49642
rect -13651 49602 -13163 49636
rect -13647 49596 -13255 49602
rect -13394 49446 -13348 49596
rect -12521 49734 -12317 49740
rect -12613 49700 -12125 49734
rect -12521 49694 -12317 49700
rect -13459 49440 -13255 49446
rect -13651 49406 -13163 49440
rect -13459 49400 -13255 49406
rect -13394 49250 -13348 49400
rect -13459 49244 -13255 49250
rect -13651 49210 -13163 49244
rect -13459 49204 -13255 49210
rect -13386 49163 -13316 49204
rect -13565 49117 -13316 49163
rect -13565 49020 -13516 49117
rect -13367 49044 -13161 49081
rect -13368 49021 -13161 49044
rect -13629 48963 -13465 49020
rect -13368 49009 -13305 49021
rect -13379 48841 -13305 49009
rect -13647 48799 -13255 48805
rect -13651 48765 -13163 48799
rect -13647 48759 -13255 48765
rect -13394 48609 -13348 48759
rect -13459 48603 -13255 48609
rect -13651 48569 -13163 48603
rect -13459 48563 -13255 48569
rect -13394 48413 -13348 48563
rect -13459 48407 -13255 48413
rect -13651 48373 -13163 48407
rect -13459 48367 -13255 48373
rect -13386 48312 -13316 48367
rect -13578 48239 -13316 48312
rect -13578 48238 -13410 48239
rect -13704 48188 -13625 48189
rect -13551 48188 -13195 48194
rect -13125 48188 -13033 48193
rect -13704 48154 -13033 48188
rect -13704 48153 -13625 48154
rect -13704 47993 -13670 48153
rect -13551 48147 -13195 48154
rect -13125 48149 -13033 48154
rect -13544 48090 -13458 48091
rect -13636 48056 -13458 48090
rect -13544 48055 -13458 48056
rect -13704 47992 -13615 47993
rect -13704 47958 -13528 47992
rect -13704 47951 -13615 47958
rect -13704 47799 -13670 47951
rect -13636 47893 -13528 47894
rect -13492 47893 -13458 48055
rect -13404 48022 -13330 48147
rect -13291 48090 -13216 48094
rect -13291 48056 -13113 48090
rect -13291 48053 -13216 48056
rect -13636 47860 -13458 47893
rect -13546 47857 -13458 47860
rect -13704 47796 -13614 47799
rect -13704 47762 -13528 47796
rect -13704 47757 -13614 47762
rect -13704 47603 -13670 47757
rect -13492 47699 -13458 47857
rect -13546 47698 -13458 47699
rect -13636 47664 -13458 47698
rect -13546 47663 -13458 47664
rect -13492 47638 -13458 47663
rect -13291 47896 -13257 48053
rect -13067 47997 -13033 48149
rect -13136 47992 -13033 47997
rect -13221 47958 -13033 47992
rect -13136 47953 -13033 47958
rect -13291 47894 -13208 47896
rect -13291 47860 -13113 47894
rect -13291 47855 -13208 47860
rect -13291 47702 -13257 47855
rect -13067 47801 -13033 47953
rect -13136 47796 -13033 47801
rect -13221 47762 -13033 47796
rect -13136 47757 -13033 47762
rect -13291 47698 -13208 47702
rect -13291 47664 -13113 47698
rect -13291 47661 -13208 47664
rect -13291 47638 -13257 47661
rect -13704 47600 -13619 47603
rect -13704 47566 -13528 47600
rect -13704 47561 -13619 47566
rect -13492 47505 -13257 47638
rect -13067 47604 -13033 47757
rect -13125 47600 -13033 47604
rect -13221 47566 -13033 47600
rect -13125 47560 -13033 47566
rect -13536 47502 -13207 47505
rect -13636 47468 -13113 47502
rect -13536 47464 -13207 47468
rect -13536 47463 -13250 47464
rect -13351 47372 -13291 47463
rect -13372 47146 -13312 47168
rect -13379 46978 -13305 47146
rect -13647 46936 -13255 46942
rect -13651 46902 -13163 46936
rect -13647 46896 -13255 46902
rect -13394 46746 -13348 46896
rect -12818 49117 -12779 49523
rect -12428 49544 -12382 49694
rect -12521 49538 -12317 49544
rect -12613 49504 -12125 49538
rect -12521 49498 -12317 49504
rect -12428 49348 -12382 49498
rect -12521 49342 -12129 49348
rect -12613 49308 -12125 49342
rect -12521 49302 -12129 49308
rect -12826 48985 -12766 49117
rect -12471 49098 -12397 49266
rect -13459 46740 -13255 46746
rect -13651 46706 -13163 46740
rect -13459 46700 -13255 46706
rect -13394 46550 -13348 46700
rect -13459 46544 -13255 46550
rect -13651 46510 -13163 46544
rect -13459 46504 -13255 46510
rect -13386 46468 -13316 46504
rect -13577 46406 -13316 46468
rect -13577 46320 -13515 46406
rect -13629 46263 -13465 46320
rect -13647 46099 -13255 46105
rect -13651 46065 -13163 46099
rect -13647 46059 -13255 46065
rect -13394 45909 -13348 46059
rect -13459 45903 -13255 45909
rect -13651 45869 -13163 45903
rect -13459 45863 -13255 45869
rect -13394 45713 -13348 45863
rect -13459 45707 -13255 45713
rect -13651 45673 -13163 45707
rect -13459 45667 -13255 45673
rect -13386 45612 -13316 45667
rect -13578 45539 -13316 45612
rect -13578 45538 -13410 45539
rect -13704 45488 -13625 45489
rect -13551 45488 -13195 45494
rect -13125 45488 -13033 45493
rect -13704 45454 -13033 45488
rect -13704 45453 -13625 45454
rect -13704 45293 -13670 45453
rect -13551 45447 -13195 45454
rect -13125 45449 -13033 45454
rect -13544 45390 -13458 45391
rect -13636 45356 -13458 45390
rect -13544 45355 -13458 45356
rect -13704 45292 -13615 45293
rect -13704 45258 -13528 45292
rect -13704 45251 -13615 45258
rect -13704 45099 -13670 45251
rect -13636 45193 -13528 45194
rect -13492 45193 -13458 45355
rect -13404 45322 -13330 45447
rect -13291 45390 -13216 45394
rect -13291 45356 -13113 45390
rect -13291 45353 -13216 45356
rect -13636 45160 -13458 45193
rect -13546 45157 -13458 45160
rect -13704 45096 -13614 45099
rect -13704 45062 -13528 45096
rect -13704 45057 -13614 45062
rect -13704 44903 -13670 45057
rect -13492 44999 -13458 45157
rect -13546 44998 -13458 44999
rect -13636 44964 -13458 44998
rect -13546 44963 -13458 44964
rect -13492 44938 -13458 44963
rect -13291 45196 -13257 45353
rect -13067 45297 -13033 45449
rect -13136 45292 -13033 45297
rect -13221 45258 -13033 45292
rect -13136 45253 -13033 45258
rect -13291 45194 -13208 45196
rect -13291 45160 -13113 45194
rect -13291 45155 -13208 45160
rect -13291 45002 -13257 45155
rect -13067 45101 -13033 45253
rect -13136 45096 -13033 45101
rect -13221 45062 -13033 45096
rect -13136 45057 -13033 45062
rect -13291 44998 -13208 45002
rect -13291 44964 -13113 44998
rect -13291 44961 -13208 44964
rect -13291 44938 -13257 44961
rect -13704 44900 -13619 44903
rect -13704 44866 -13528 44900
rect -13704 44861 -13619 44866
rect -13492 44805 -13257 44938
rect -13067 44904 -13033 45057
rect -13125 44900 -13033 44904
rect -13221 44866 -13033 44900
rect -13125 44860 -13033 44866
rect -13536 44802 -13207 44805
rect -13636 44768 -13113 44802
rect -13536 44764 -13207 44768
rect -13536 44763 -13250 44764
rect -13349 44688 -13289 44763
rect -12818 44594 -12779 48985
rect -12456 48901 -12403 49098
rect -12526 48900 -12240 48901
rect -12569 48896 -12240 48900
rect -12663 48862 -12140 48896
rect -12569 48859 -12240 48862
rect -12743 48798 -12651 48804
rect -12743 48764 -12555 48798
rect -12743 48760 -12651 48764
rect -12743 48607 -12709 48760
rect -12519 48726 -12284 48859
rect -12157 48798 -12072 48803
rect -12248 48764 -12072 48798
rect -12157 48761 -12072 48764
rect -12519 48703 -12485 48726
rect -12568 48700 -12485 48703
rect -12663 48666 -12485 48700
rect -12568 48662 -12485 48666
rect -12743 48602 -12640 48607
rect -12743 48568 -12555 48602
rect -12743 48563 -12640 48568
rect -12743 48411 -12709 48563
rect -12519 48509 -12485 48662
rect -12568 48504 -12485 48509
rect -12663 48470 -12485 48504
rect -12568 48468 -12485 48470
rect -12743 48406 -12640 48411
rect -12743 48372 -12555 48406
rect -12743 48367 -12640 48372
rect -12743 48215 -12709 48367
rect -12519 48311 -12485 48468
rect -12318 48701 -12284 48726
rect -12318 48700 -12230 48701
rect -12318 48666 -12140 48700
rect -12318 48665 -12230 48666
rect -12318 48507 -12284 48665
rect -12106 48607 -12072 48761
rect -12162 48602 -12072 48607
rect -12248 48568 -12072 48602
rect -12162 48565 -12072 48568
rect -12318 48504 -12230 48507
rect -12318 48471 -12140 48504
rect -12560 48308 -12485 48311
rect -12663 48274 -12485 48308
rect -12560 48270 -12485 48274
rect -12446 48217 -12372 48342
rect -12318 48309 -12284 48471
rect -12248 48470 -12140 48471
rect -12106 48413 -12072 48565
rect -12161 48406 -12072 48413
rect -12248 48372 -12072 48406
rect -12161 48371 -12072 48372
rect -12318 48308 -12232 48309
rect -12318 48274 -12140 48308
rect -12318 48273 -12232 48274
rect -12743 48210 -12651 48215
rect -12581 48210 -12225 48217
rect -12106 48211 -12072 48371
rect -12151 48210 -12072 48211
rect -12743 48176 -12072 48210
rect -12743 48171 -12651 48176
rect -12581 48170 -12225 48176
rect -12151 48175 -12072 48176
rect -12366 48125 -12198 48126
rect -12460 48052 -12198 48125
rect -12460 47997 -12390 48052
rect -12521 47991 -12317 47997
rect -12613 47957 -12125 47991
rect -12521 47951 -12317 47957
rect -12428 47801 -12382 47951
rect -12521 47795 -12317 47801
rect -12613 47761 -12125 47795
rect -12521 47755 -12317 47761
rect -12428 47605 -12382 47755
rect -12521 47599 -12129 47605
rect -12613 47565 -12125 47599
rect -12521 47559 -12129 47565
rect -11012 47557 -10850 50456
rect -10708 50353 -10672 50691
rect -9045 51541 -8969 51553
rect -9045 51507 -8367 51541
rect -8329 51531 -8045 51573
rect -9045 51497 -8969 51507
rect -9045 51355 -9011 51497
rect -8329 51447 -8287 51531
rect -8385 51443 -8287 51447
rect -8975 51409 -8287 51443
rect -8385 51405 -8287 51409
rect -9045 51345 -8969 51355
rect -9045 51311 -8367 51345
rect -8214 51313 -8158 51398
rect -9045 51299 -8969 51311
rect -9045 51143 -9011 51299
rect -8260 51253 -8158 51313
rect -8378 51232 -8296 51235
rect -8975 51198 -8296 51232
rect -8378 51193 -8296 51198
rect -9045 51134 -8969 51143
rect -9045 51100 -8367 51134
rect -9045 51090 -8969 51100
rect -8333 51039 -8296 51193
rect -8377 51036 -8296 51039
rect -8975 51002 -8296 51036
rect -8377 50997 -8296 51002
rect -8333 50827 -8296 50997
rect -8384 50824 -8296 50827
rect -8975 50790 -8296 50824
rect -8384 50786 -8296 50790
rect -12311 47344 -12147 47401
rect -12270 47185 -12225 47344
rect -12449 47180 -12225 47185
rect -12564 47140 -12225 47180
rect -12564 47120 -12404 47140
rect -12449 47070 -12404 47120
rect -12460 47040 -12390 47070
rect -12521 47034 -12317 47040
rect -12613 47000 -12125 47034
rect -12521 46994 -12317 47000
rect -12428 46844 -12382 46994
rect -12521 46838 -12317 46844
rect -12613 46804 -12125 46838
rect -12521 46798 -12317 46804
rect -12428 46648 -12382 46798
rect -11286 47446 -10850 47557
rect -12521 46642 -12129 46648
rect -12613 46608 -12125 46642
rect -12521 46602 -12129 46608
rect -12471 46398 -12397 46566
rect -12463 46201 -12406 46398
rect -12526 46200 -12240 46201
rect -12569 46199 -12240 46200
rect -12691 46196 -12240 46199
rect -12691 46162 -12140 46196
rect -12691 46159 -12240 46162
rect -12691 46153 -12559 46159
rect -12743 46098 -12651 46104
rect -12743 46064 -12555 46098
rect -12743 46060 -12651 46064
rect -12743 45907 -12709 46060
rect -12519 46026 -12284 46159
rect -12157 46098 -12072 46103
rect -12248 46064 -12072 46098
rect -12157 46061 -12072 46064
rect -12519 46003 -12485 46026
rect -12568 46000 -12485 46003
rect -12663 45966 -12485 46000
rect -12568 45962 -12485 45966
rect -12743 45902 -12640 45907
rect -12743 45868 -12555 45902
rect -12743 45863 -12640 45868
rect -12743 45711 -12709 45863
rect -12519 45809 -12485 45962
rect -12568 45804 -12485 45809
rect -12663 45770 -12485 45804
rect -12568 45768 -12485 45770
rect -12743 45706 -12640 45711
rect -12743 45672 -12555 45706
rect -12743 45667 -12640 45672
rect -12743 45515 -12709 45667
rect -12519 45611 -12485 45768
rect -12318 46001 -12284 46026
rect -12318 46000 -12230 46001
rect -12318 45966 -12140 46000
rect -12318 45965 -12230 45966
rect -12318 45807 -12284 45965
rect -12106 45907 -12072 46061
rect -12162 45902 -12072 45907
rect -12248 45868 -12072 45902
rect -12162 45865 -12072 45868
rect -12318 45804 -12230 45807
rect -12318 45771 -12140 45804
rect -12560 45608 -12485 45611
rect -12663 45574 -12485 45608
rect -12560 45570 -12485 45574
rect -12446 45517 -12372 45642
rect -12318 45609 -12284 45771
rect -12248 45770 -12140 45771
rect -12106 45713 -12072 45865
rect -12161 45706 -12072 45713
rect -12248 45672 -12072 45706
rect -12161 45671 -12072 45672
rect -12318 45608 -12232 45609
rect -12318 45574 -12140 45608
rect -12318 45573 -12232 45574
rect -12743 45510 -12651 45515
rect -12581 45510 -12225 45517
rect -12106 45511 -12072 45671
rect -12151 45510 -12072 45511
rect -12743 45476 -12072 45510
rect -12743 45471 -12651 45476
rect -12581 45470 -12225 45476
rect -12151 45475 -12072 45476
rect -12366 45425 -12198 45426
rect -12460 45352 -12198 45425
rect -12460 45297 -12390 45352
rect -12521 45291 -12317 45297
rect -12613 45257 -12125 45291
rect -12521 45251 -12317 45257
rect -12428 45101 -12382 45251
rect -12521 45095 -12317 45101
rect -12613 45061 -12125 45095
rect -12521 45055 -12317 45061
rect -12428 44905 -12382 45055
rect -12521 44899 -12129 44905
rect -12613 44865 -12125 44899
rect -12521 44859 -12129 44865
rect -12828 44462 -12768 44594
rect -12471 44655 -12397 44823
rect -12466 44620 -12408 44655
rect -12311 44644 -12147 44701
rect -12454 44563 -12412 44620
rect -12540 44503 -12408 44563
rect -12454 44445 -12412 44503
rect -12460 44415 -12390 44445
rect -12521 44409 -12317 44415
rect -12613 44375 -12125 44409
rect -12521 44369 -12317 44375
rect -12428 44219 -12382 44369
rect -12521 44213 -12317 44219
rect -12613 44179 -12125 44213
rect -12521 44173 -12317 44179
rect -12428 44023 -12382 44173
rect -12521 44017 -12129 44023
rect -12613 43983 -12125 44017
rect -12521 43977 -12129 43983
rect -11286 42302 -11175 47446
rect -11012 46375 -10850 47446
rect -10738 46056 -10644 50353
rect -8260 49120 -8219 51253
rect -8087 51122 -8045 51531
rect -8087 51118 -7994 51122
rect -8087 51084 -7803 51118
rect -8087 51080 -7994 51084
rect -8182 50933 -8126 51078
rect -8171 49377 -8130 50933
rect -8087 50926 -8045 51080
rect -8087 50922 -7994 50926
rect -8087 50888 -7803 50922
rect -8087 50884 -7994 50888
rect -8087 50604 -8031 50749
rect -8079 49576 -8038 50604
rect -7705 49576 -7554 49584
rect -4404 49576 -4223 49668
rect -8079 49487 -4223 49576
rect -4404 49471 -4223 49487
rect -4879 49377 -4670 49408
rect -8171 49245 -4670 49377
rect -5307 49120 -5036 49129
rect -4879 49127 -4670 49245
rect -8260 48992 -5036 49120
rect -9895 48623 -9715 48844
rect -7705 48757 -7554 48910
rect -9873 47849 -9743 48623
rect -7964 48075 -7800 48173
rect -10151 47766 -9743 47849
rect -10738 45973 -10372 46056
rect -10738 45678 -10644 45973
rect -10805 45393 -10586 45678
rect -11296 42233 -11157 42302
rect -10455 42139 -10372 45973
rect -10151 42465 -10068 47766
rect -9873 47377 -9743 47766
rect -10005 46863 -9580 47377
rect -7937 42613 -7814 48075
rect -7941 42563 -7808 42613
rect -7937 42554 -7814 42563
rect -10163 42401 -10045 42465
rect -10460 42080 -10365 42139
rect -7668 41799 -7593 48757
rect -7261 48494 -6963 48761
rect -7234 43149 -6999 48494
rect -6119 48527 -5979 48819
rect -5307 48767 -5036 48992
rect -7674 41581 -7585 41799
rect -6119 41553 -5980 48527
rect -5254 41541 -5082 48767
rect -5419 41341 -5048 41541
rect -13494 40640 -13440 40779
rect -13623 40591 -13189 40596
rect -13814 40557 -13000 40591
rect -13623 40553 -13189 40557
rect -13426 40453 -13380 40553
rect -13621 40282 -13191 40286
rect -13814 40248 -13000 40282
rect -13621 40243 -13191 40248
rect -13500 40025 -13446 40164
rect -13282 40147 -13236 40243
rect -13325 40036 -13000 40070
rect -11243 40650 -11189 40789
rect -11372 40601 -10938 40606
rect -11563 40567 -10749 40601
rect -11372 40563 -10938 40567
rect -11175 40463 -11129 40563
rect -11370 40292 -10940 40296
rect -11563 40258 -10749 40292
rect -11370 40253 -10940 40258
rect -13814 39938 -13463 39972
rect -13814 39742 -13537 39776
rect -13571 39596 -13537 39742
rect -13952 39562 -13537 39596
rect -13952 39098 -13918 39562
rect -13497 39526 -13463 39938
rect -13325 39776 -13291 40036
rect -13017 39972 -12927 39974
rect -13208 39938 -12927 39972
rect -13426 39616 -13372 39755
rect -13325 39742 -13000 39776
rect -13325 39543 -13291 39742
rect -13883 39492 -13463 39526
rect -13421 39509 -13291 39543
rect -13238 39644 -13000 39678
rect -13883 39414 -13849 39492
rect -13421 39431 -13387 39509
rect -13883 39380 -13606 39414
rect -13570 39397 -13387 39431
rect -13238 39414 -13199 39644
rect -13883 39218 -13849 39380
rect -13570 39316 -13536 39397
rect -13814 39282 -13536 39316
rect -13883 39184 -13606 39218
rect -13952 39064 -13606 39098
rect -13952 38902 -13918 39064
rect -13570 39000 -13536 39282
rect -13238 39380 -13000 39414
rect -13238 39378 -13199 39380
rect -13814 38966 -13536 39000
rect -13952 38868 -13606 38902
rect -13570 38584 -13536 38966
rect -13456 38867 -13402 39006
rect -12963 39000 -12927 39938
rect -13208 38966 -12927 39000
rect -11249 40035 -11195 40174
rect -11031 40157 -10985 40253
rect -11074 40046 -10749 40080
rect -11563 39948 -11212 39982
rect -11563 39752 -11286 39786
rect -11320 39606 -11286 39752
rect -11701 39572 -11286 39606
rect -11701 39108 -11667 39572
rect -11246 39536 -11212 39948
rect -11074 39786 -11040 40046
rect -10766 39982 -10676 39984
rect -10957 39948 -10676 39982
rect -11175 39626 -11121 39765
rect -11074 39752 -10749 39786
rect -11074 39553 -11040 39752
rect -11632 39502 -11212 39536
rect -11170 39519 -11040 39553
rect -10987 39654 -10749 39688
rect -11632 39424 -11598 39502
rect -11170 39441 -11136 39519
rect -11632 39390 -11355 39424
rect -11319 39407 -11136 39441
rect -10987 39424 -10948 39654
rect -11632 39228 -11598 39390
rect -11319 39326 -11285 39407
rect -11563 39292 -11285 39326
rect -11632 39194 -11355 39228
rect -11701 39074 -11355 39108
rect -11701 38912 -11667 39074
rect -11319 39010 -11285 39292
rect -10987 39390 -10749 39424
rect -10987 39388 -10948 39390
rect -11563 38976 -11285 39010
rect -11701 38878 -11355 38912
rect -13169 38584 -13033 38590
rect -13570 38550 -13033 38584
rect -13169 38544 -13033 38550
rect -13494 37640 -13440 37779
rect -11319 38827 -11285 38976
rect -11205 38877 -11151 39016
rect -10712 39010 -10676 39948
rect -10957 38976 -10676 39010
rect -7693 40650 -7639 40789
rect -7944 40601 -7510 40606
rect -8133 40567 -7319 40601
rect -7944 40563 -7510 40567
rect -7753 40463 -7707 40563
rect -7942 40292 -7512 40296
rect -8133 40258 -7319 40292
rect -7942 40253 -7512 40258
rect -7897 40157 -7851 40253
rect -8133 40046 -7808 40080
rect -12731 38730 -11120 38764
rect -12731 38628 -12697 38730
rect -12639 38660 -11198 38694
rect -12737 38492 -12691 38628
rect -12639 38388 -12605 38660
rect -11319 38604 -11282 38623
rect -11327 38469 -11273 38604
rect -11319 38468 -11273 38469
rect -12712 38354 -12605 38388
rect -13623 37591 -13189 37596
rect -13814 37557 -13000 37591
rect -13623 37553 -13189 37557
rect -13426 37453 -13380 37553
rect -13621 37282 -13191 37286
rect -13814 37248 -13000 37282
rect -13621 37243 -13191 37248
rect -13500 37025 -13446 37164
rect -13282 37147 -13236 37243
rect -13325 37036 -13000 37070
rect -13814 36938 -13463 36972
rect -13814 36742 -13537 36776
rect -13571 36596 -13537 36742
rect -13952 36562 -13537 36596
rect -13952 36098 -13918 36562
rect -13497 36526 -13463 36938
rect -13325 36776 -13291 37036
rect -13017 36972 -12927 36974
rect -13208 36938 -12927 36972
rect -13426 36616 -13372 36755
rect -13325 36742 -13000 36776
rect -13325 36543 -13291 36742
rect -13883 36492 -13463 36526
rect -13421 36509 -13291 36543
rect -13238 36644 -13000 36678
rect -13883 36414 -13849 36492
rect -13421 36431 -13387 36509
rect -13883 36380 -13606 36414
rect -13570 36397 -13387 36431
rect -13238 36414 -13199 36644
rect -13883 36218 -13849 36380
rect -13570 36316 -13536 36397
rect -13814 36282 -13536 36316
rect -13883 36184 -13606 36218
rect -13952 36064 -13606 36098
rect -13952 35902 -13918 36064
rect -13570 36000 -13536 36282
rect -13238 36380 -13000 36414
rect -13238 36378 -13199 36380
rect -13814 35966 -13536 36000
rect -13952 35868 -13606 35902
rect -13570 35678 -13536 35966
rect -13456 35867 -13402 36006
rect -12963 36000 -12927 36938
rect -13208 35966 -12927 36000
rect -13169 35679 -13033 35685
rect -13170 35678 -13033 35679
rect -13570 35644 -13033 35678
rect -13169 35639 -13033 35644
rect -13494 35140 -13440 35279
rect -12712 35723 -12678 38354
rect -11574 38395 -11293 38429
rect -11330 38233 -11293 38395
rect -11236 38268 -11198 38660
rect -11574 38199 -11293 38233
rect -11330 38037 -11293 38199
rect -11245 38133 -11191 38268
rect -11154 38080 -11120 38730
rect -11064 38493 -10659 38527
rect -11064 38331 -11030 38493
rect -11064 38297 -10659 38331
rect -11064 38119 -11029 38297
rect -10966 38183 -10526 38217
rect -10667 38182 -10526 38183
rect -11064 38085 -10658 38119
rect -11064 38084 -10966 38085
rect -11574 38003 -11293 38037
rect -11330 37911 -11293 38003
rect -11167 37945 -11113 38080
rect -10563 38021 -10526 38182
rect -10966 37987 -10526 38021
rect -10669 37986 -10526 37987
rect -11330 37908 -11030 37911
rect -11330 37874 -10658 37908
rect -11155 37469 -11118 37874
rect -11064 37712 -11030 37874
rect -10560 37810 -10526 37986
rect -10966 37776 -10526 37810
rect -11064 37678 -10658 37712
rect -11165 37334 -11111 37469
rect -8206 39982 -8116 39984
rect -8206 39948 -7925 39982
rect -8206 39010 -8170 39948
rect -7842 39786 -7808 40046
rect -7687 40035 -7633 40174
rect -5442 40640 -5388 40779
rect -5693 40591 -5259 40596
rect -5882 40557 -5068 40591
rect -5693 40553 -5259 40557
rect -5502 40453 -5456 40553
rect -5691 40282 -5261 40286
rect -5882 40248 -5068 40282
rect -5691 40243 -5261 40248
rect -5646 40147 -5600 40243
rect -8133 39752 -7808 39786
rect -7670 39948 -7319 39982
rect -8133 39654 -7895 39688
rect -7934 39424 -7895 39654
rect -7842 39553 -7808 39752
rect -7761 39626 -7707 39765
rect -7842 39519 -7712 39553
rect -8133 39390 -7895 39424
rect -7746 39441 -7712 39519
rect -7670 39536 -7636 39948
rect -7596 39752 -7319 39786
rect -7596 39606 -7562 39752
rect -7596 39572 -7181 39606
rect -7670 39502 -7250 39536
rect -7746 39407 -7563 39441
rect -7284 39424 -7250 39502
rect -7934 39388 -7895 39390
rect -7597 39326 -7563 39407
rect -7527 39390 -7250 39424
rect -7597 39292 -7319 39326
rect -8206 38976 -7925 39010
rect -7731 38877 -7677 39016
rect -7597 39010 -7563 39292
rect -7284 39228 -7250 39390
rect -7527 39194 -7250 39228
rect -7215 39108 -7181 39572
rect -7527 39074 -7181 39108
rect -7597 38976 -7319 39010
rect -7597 38827 -7563 38976
rect -7215 38912 -7181 39074
rect -7527 38878 -7181 38912
rect -5882 40036 -5557 40070
rect -5955 39972 -5865 39974
rect -5955 39938 -5674 39972
rect -5955 39000 -5919 39938
rect -5591 39776 -5557 40036
rect -5436 40025 -5382 40164
rect -5882 39742 -5557 39776
rect -5419 39938 -5068 39972
rect -5882 39644 -5644 39678
rect -5683 39414 -5644 39644
rect -5591 39543 -5557 39742
rect -5510 39616 -5456 39755
rect -5591 39509 -5461 39543
rect -5882 39380 -5644 39414
rect -5495 39431 -5461 39509
rect -5419 39526 -5385 39938
rect -5345 39742 -5068 39776
rect -5345 39596 -5311 39742
rect -5345 39562 -4930 39596
rect -5419 39492 -4999 39526
rect -5495 39397 -5312 39431
rect -5033 39414 -4999 39492
rect -5683 39378 -5644 39380
rect -5346 39316 -5312 39397
rect -5276 39380 -4999 39414
rect -5346 39282 -5068 39316
rect -5955 38966 -5674 39000
rect -5480 38867 -5426 39006
rect -5346 39000 -5312 39282
rect -5033 39218 -4999 39380
rect -5276 39184 -4999 39218
rect -4964 39098 -4930 39562
rect -5276 39064 -4930 39098
rect -5346 38966 -5068 39000
rect -7762 38730 -6151 38764
rect -8223 38493 -7818 38527
rect -7852 38331 -7818 38493
rect -8223 38297 -7818 38331
rect -8356 38183 -7916 38217
rect -8356 38182 -8215 38183
rect -8356 38021 -8319 38182
rect -7853 38119 -7818 38297
rect -8224 38085 -7818 38119
rect -7916 38084 -7818 38085
rect -7762 38080 -7728 38730
rect -7684 38660 -6243 38694
rect -7684 38268 -7646 38660
rect -7600 38604 -7563 38623
rect -7609 38469 -7555 38604
rect -7609 38468 -7563 38469
rect -7589 38395 -7308 38429
rect -7691 38133 -7637 38268
rect -7589 38233 -7552 38395
rect -6277 38388 -6243 38660
rect -6185 38628 -6151 38730
rect -6191 38492 -6145 38628
rect -6277 38354 -6170 38388
rect -7589 38199 -7308 38233
rect -8356 37987 -7916 38021
rect -8356 37986 -8213 37987
rect -8356 37810 -8322 37986
rect -7769 37945 -7715 38080
rect -7589 38037 -7552 38199
rect -7589 38003 -7308 38037
rect -7589 37911 -7552 38003
rect -7852 37908 -7552 37911
rect -8224 37874 -7552 37908
rect -8356 37776 -7916 37810
rect -7852 37712 -7818 37874
rect -8224 37678 -7818 37712
rect -7764 37469 -7727 37874
rect -11574 37265 -10658 37299
rect -10974 37114 -10916 37265
rect -10461 37114 -10415 37115
rect -10974 37049 -10415 37114
rect -12623 36970 -11056 37010
rect -10461 36979 -10415 37049
rect -12721 35587 -12675 35723
rect -12623 35542 -12589 36970
rect -12781 35508 -12589 35542
rect -12555 36911 -11154 36931
rect -12555 36895 -11152 36911
rect -13623 35091 -13189 35096
rect -13814 35057 -13000 35091
rect -13623 35053 -13189 35057
rect -13426 34953 -13380 35053
rect -13621 34782 -13191 34786
rect -13814 34748 -13000 34782
rect -13621 34743 -13191 34748
rect -13500 34525 -13446 34664
rect -13282 34647 -13236 34743
rect -13325 34536 -13000 34570
rect -13814 34438 -13463 34472
rect -13814 34242 -13537 34276
rect -13571 34096 -13537 34242
rect -13952 34062 -13537 34096
rect -13952 33598 -13918 34062
rect -13497 34026 -13463 34438
rect -13325 34276 -13291 34536
rect -13017 34472 -12927 34474
rect -13208 34438 -12927 34472
rect -13426 34116 -13372 34255
rect -13325 34242 -13000 34276
rect -13325 34043 -13291 34242
rect -13883 33992 -13463 34026
rect -13421 34009 -13291 34043
rect -13238 34144 -13000 34178
rect -13883 33914 -13849 33992
rect -13421 33931 -13387 34009
rect -13883 33880 -13606 33914
rect -13570 33897 -13387 33931
rect -13238 33914 -13199 34144
rect -13883 33718 -13849 33880
rect -13570 33816 -13536 33897
rect -13814 33782 -13536 33816
rect -13883 33684 -13606 33718
rect -13952 33564 -13606 33598
rect -13952 33402 -13918 33564
rect -13570 33500 -13536 33782
rect -13238 33880 -13000 33914
rect -13238 33878 -13199 33880
rect -13814 33466 -13536 33500
rect -13952 33368 -13606 33402
rect -13570 33262 -13536 33466
rect -13456 33367 -13402 33506
rect -12963 33500 -12927 34438
rect -13208 33466 -12927 33500
rect -12781 33540 -12747 35508
rect -12555 35446 -12519 36895
rect -11192 36859 -11152 36895
rect -11198 36724 -11144 36859
rect -11096 36806 -11056 36970
rect -11096 36805 -11054 36806
rect -11094 36735 -11054 36805
rect -11012 36740 -10704 36774
rect -11549 36642 -11167 36676
rect -11205 36480 -11167 36642
rect -11549 36446 -11167 36480
rect -11205 36307 -11167 36446
rect -11094 36394 -11055 36735
rect -11012 36544 -10704 36578
rect -11012 36446 -10704 36480
rect -7771 37334 -7717 37469
rect -8224 37265 -7308 37299
rect -8467 37114 -8421 37115
rect -7966 37114 -7908 37265
rect -8467 37049 -7908 37114
rect -8467 36979 -8421 37049
rect -7826 36970 -6259 37010
rect -7826 36806 -7786 36970
rect -7728 36911 -6327 36931
rect -7730 36895 -6327 36911
rect -7730 36859 -7690 36895
rect -7828 36805 -7786 36806
rect -8178 36740 -7870 36774
rect -7828 36735 -7788 36805
rect -8178 36544 -7870 36578
rect -11120 36320 -11049 36394
rect -11012 36348 -10704 36382
rect -8178 36446 -7870 36480
rect -7827 36394 -7788 36735
rect -7738 36724 -7684 36859
rect -7715 36642 -7333 36676
rect -7715 36480 -7677 36642
rect -7715 36446 -7333 36480
rect -8178 36348 -7870 36382
rect -11367 36285 -11167 36307
rect -11395 36257 -11167 36285
rect -11395 36246 -11175 36257
rect -11395 36185 -11354 36246
rect -11408 36112 -11348 36185
rect -11550 36033 -11442 36067
rect -11319 35935 -11211 35969
rect -11550 35837 -11442 35871
rect -11319 35739 -11211 35773
rect -11550 35641 -11308 35675
rect -11378 35547 -11308 35641
rect -11378 35477 -10527 35547
rect -12703 35410 -12519 35446
rect -10573 35411 -10527 35477
rect -12784 33404 -12738 33540
rect -12781 33371 -12747 33404
rect -13169 33262 -13033 33268
rect -13571 33228 -13033 33262
rect -13169 33222 -13033 33228
rect -13494 32640 -13440 32779
rect -13623 32591 -13189 32596
rect -13814 32557 -13000 32591
rect -13623 32553 -13189 32557
rect -13426 32453 -13380 32553
rect -13621 32282 -13191 32286
rect -13814 32248 -13000 32282
rect -13621 32243 -13191 32248
rect -13500 32025 -13446 32164
rect -13282 32147 -13236 32243
rect -13325 32036 -13000 32070
rect -13814 31938 -13463 31972
rect -13814 31742 -13537 31776
rect -13571 31596 -13537 31742
rect -13952 31562 -13537 31596
rect -13952 31098 -13918 31562
rect -13497 31526 -13463 31938
rect -13325 31776 -13291 32036
rect -13017 31972 -12927 31974
rect -13208 31938 -12927 31972
rect -13426 31616 -13372 31755
rect -13325 31742 -13000 31776
rect -13325 31543 -13291 31742
rect -13883 31492 -13463 31526
rect -13421 31509 -13291 31543
rect -13238 31644 -13000 31678
rect -13883 31414 -13849 31492
rect -13421 31431 -13387 31509
rect -13883 31380 -13606 31414
rect -13570 31397 -13387 31431
rect -13238 31414 -13199 31644
rect -13883 31218 -13849 31380
rect -13570 31316 -13536 31397
rect -13814 31282 -13536 31316
rect -13883 31184 -13606 31218
rect -13952 31064 -13606 31098
rect -13952 30902 -13918 31064
rect -13570 31000 -13536 31282
rect -13238 31380 -13000 31414
rect -13238 31378 -13199 31380
rect -13814 30966 -13536 31000
rect -13952 30868 -13606 30902
rect -13570 30782 -13536 30966
rect -13456 30867 -13402 31006
rect -12963 31000 -12927 31938
rect -13208 30966 -12927 31000
rect -12703 31043 -12667 35410
rect -12080 35342 -11058 35382
rect -12080 35246 -12034 35342
rect -11192 35297 -11156 35306
rect -11996 35284 -11156 35297
rect -11996 35261 -11152 35284
rect -11996 35142 -11950 35261
rect -11200 35254 -11152 35261
rect -11200 35119 -11146 35254
rect -11098 35201 -11058 35342
rect -11098 35200 -11056 35201
rect -11096 35130 -11056 35200
rect -11014 35135 -10706 35169
rect -11551 35037 -11169 35071
rect -11207 34875 -11169 35037
rect -11551 34841 -11169 34875
rect -11207 34702 -11169 34841
rect -11096 34789 -11057 35130
rect -7833 36320 -7762 36394
rect -7715 36307 -7677 36446
rect -7715 36285 -7515 36307
rect -7715 36257 -7487 36285
rect -7707 36246 -7487 36257
rect -7528 36185 -7487 36246
rect -7534 36112 -7474 36185
rect -7440 36033 -7332 36067
rect -7671 35935 -7563 35969
rect -7440 35837 -7332 35871
rect -7671 35739 -7563 35773
rect -7574 35641 -7332 35675
rect -7574 35547 -7504 35641
rect -8355 35477 -7504 35547
rect -8355 35411 -8309 35477
rect -6363 35446 -6327 36895
rect -6293 35542 -6259 36970
rect -6204 35723 -6170 38354
rect -5849 38584 -5713 38590
rect -5346 38584 -5312 38966
rect -4964 38902 -4930 39064
rect -5276 38868 -4930 38902
rect -5849 38550 -5312 38584
rect -5849 38544 -5713 38550
rect -5442 37640 -5388 37779
rect -5693 37591 -5259 37596
rect -5882 37557 -5068 37591
rect -5693 37553 -5259 37557
rect -5502 37453 -5456 37553
rect -5691 37282 -5261 37286
rect -5882 37248 -5068 37282
rect -5691 37243 -5261 37248
rect -5646 37147 -5600 37243
rect -5882 37036 -5557 37070
rect -5955 36972 -5865 36974
rect -5955 36938 -5674 36972
rect -5955 36000 -5919 36938
rect -5591 36776 -5557 37036
rect -5436 37025 -5382 37164
rect -5882 36742 -5557 36776
rect -5419 36938 -5068 36972
rect -5882 36644 -5644 36678
rect -5683 36414 -5644 36644
rect -5591 36543 -5557 36742
rect -5510 36616 -5456 36755
rect -5591 36509 -5461 36543
rect -5882 36380 -5644 36414
rect -5495 36431 -5461 36509
rect -5419 36526 -5385 36938
rect -5345 36742 -5068 36776
rect -5345 36596 -5311 36742
rect -5345 36562 -4930 36596
rect -5419 36492 -4999 36526
rect -5495 36397 -5312 36431
rect -5033 36414 -4999 36492
rect -5683 36378 -5644 36380
rect -5346 36316 -5312 36397
rect -5276 36380 -4999 36414
rect -5346 36282 -5068 36316
rect -5955 35966 -5674 36000
rect -5480 35867 -5426 36006
rect -5346 36000 -5312 36282
rect -5033 36218 -4999 36380
rect -5276 36184 -4999 36218
rect -4964 36098 -4930 36562
rect -5276 36064 -4930 36098
rect -5346 35966 -5068 36000
rect -6207 35587 -6161 35723
rect -6293 35508 -6101 35542
rect -6363 35410 -6179 35446
rect -7824 35342 -6802 35382
rect -7824 35201 -7784 35342
rect -7726 35297 -7690 35306
rect -7726 35284 -6886 35297
rect -7730 35261 -6886 35284
rect -7730 35254 -7682 35261
rect -7826 35200 -7784 35201
rect -8176 35135 -7868 35169
rect -7826 35130 -7786 35200
rect -11014 34939 -10706 34973
rect -11014 34841 -10706 34875
rect -8176 34939 -7868 34973
rect -8176 34841 -7868 34875
rect -11122 34715 -11051 34789
rect -11014 34743 -10706 34777
rect -7825 34789 -7786 35130
rect -7736 35119 -7682 35254
rect -6932 35142 -6886 35261
rect -6848 35246 -6802 35342
rect -7713 35037 -7331 35071
rect -7713 34875 -7675 35037
rect -7713 34841 -7331 34875
rect -11369 34680 -11169 34702
rect -11397 34652 -11169 34680
rect -11397 34641 -11177 34652
rect -11397 34580 -11356 34641
rect -11410 34507 -11350 34580
rect -11552 34428 -11444 34462
rect -11321 34330 -11213 34364
rect -11552 34232 -11444 34266
rect -11321 34134 -11213 34168
rect -11552 34036 -11310 34070
rect -11380 33939 -11310 34036
rect -8176 34743 -7868 34777
rect -7831 34715 -7760 34789
rect -7713 34702 -7675 34841
rect -7713 34680 -7513 34702
rect -7713 34652 -7485 34680
rect -7705 34641 -7485 34652
rect -7526 34580 -7485 34641
rect -7532 34507 -7472 34580
rect -7438 34428 -7330 34462
rect -7669 34330 -7561 34364
rect -7438 34232 -7330 34266
rect -7669 34134 -7561 34168
rect -7572 34036 -7330 34070
rect -11380 33905 -11111 33939
rect -11380 33899 -11310 33905
rect -11228 33734 -11182 33870
rect -11402 33653 -11264 33699
rect -11318 33507 -11264 33653
rect -11565 33433 -11284 33467
rect -11321 33271 -11284 33433
rect -11227 33306 -11189 33734
rect -11565 33237 -11284 33271
rect -11321 33075 -11284 33237
rect -11236 33171 -11182 33306
rect -11145 33118 -11111 33905
rect -7572 33939 -7502 34036
rect -11055 33531 -10650 33565
rect -11055 33369 -11021 33531
rect -11055 33335 -10650 33369
rect -11055 33157 -11020 33335
rect -10957 33221 -10517 33255
rect -10658 33220 -10517 33221
rect -11055 33123 -10649 33157
rect -11055 33122 -10957 33123
rect -11565 33041 -11284 33075
rect -11321 32949 -11284 33041
rect -11158 32983 -11104 33118
rect -10554 33059 -10517 33220
rect -10957 33025 -10517 33059
rect -10660 33024 -10517 33025
rect -11321 32946 -11021 32949
rect -11321 32912 -10649 32946
rect -11146 32507 -11109 32912
rect -11055 32750 -11021 32912
rect -10551 32848 -10517 33024
rect -10957 32814 -10517 32848
rect -7771 33905 -7502 33939
rect -8232 33531 -7827 33565
rect -7861 33369 -7827 33531
rect -8232 33335 -7827 33369
rect -11055 32716 -10649 32750
rect -11156 32372 -11102 32507
rect -11565 32303 -10649 32337
rect -11155 32152 -11102 32303
rect -11578 31799 -11186 31805
rect -12797 30994 -12667 31043
rect -11582 31765 -11094 31799
rect -11578 31759 -11186 31765
rect -11325 31609 -11279 31759
rect -11390 31603 -11186 31609
rect -11582 31569 -11094 31603
rect -11390 31563 -11186 31569
rect -11325 31413 -11279 31563
rect -11390 31407 -11186 31413
rect -11582 31373 -11094 31407
rect -11390 31367 -11186 31373
rect -11317 31337 -11247 31367
rect -11295 31279 -11253 31337
rect -11299 31219 -11167 31279
rect -11295 31162 -11253 31219
rect -11560 31081 -11396 31138
rect -11299 31127 -11241 31162
rect -12797 30907 -12751 30994
rect -13169 30782 -13033 30788
rect -13570 30748 -13033 30782
rect -13169 30742 -13033 30748
rect -13494 30140 -13440 30279
rect -11310 30959 -11236 31127
rect -10939 31188 -10879 31320
rect -11578 30917 -11186 30923
rect -11582 30883 -11094 30917
rect -11578 30877 -11186 30883
rect -11325 30727 -11279 30877
rect -11390 30721 -11186 30727
rect -11582 30687 -11094 30721
rect -11390 30681 -11186 30687
rect -11325 30531 -11279 30681
rect -13623 30091 -13189 30096
rect -13814 30057 -13000 30091
rect -13623 30053 -13189 30057
rect -13426 29953 -13380 30053
rect -13621 29782 -13191 29786
rect -13814 29748 -13000 29782
rect -13621 29743 -13191 29748
rect -13500 29525 -13446 29664
rect -13282 29647 -13236 29743
rect -13325 29536 -13000 29570
rect -11390 30525 -11186 30531
rect -11582 30491 -11094 30525
rect -11390 30485 -11186 30491
rect -11317 30430 -11247 30485
rect -11509 30357 -11247 30430
rect -11509 30356 -11341 30357
rect -11635 30306 -11556 30307
rect -11482 30306 -11126 30312
rect -11056 30306 -10964 30311
rect -11635 30272 -10964 30306
rect -11635 30271 -11556 30272
rect -11635 30111 -11601 30271
rect -11482 30265 -11126 30272
rect -11056 30267 -10964 30272
rect -11475 30208 -11389 30209
rect -11567 30174 -11389 30208
rect -11475 30173 -11389 30174
rect -11635 30110 -11546 30111
rect -11635 30076 -11459 30110
rect -11635 30069 -11546 30076
rect -11635 29917 -11601 30069
rect -11567 30011 -11459 30012
rect -11423 30011 -11389 30173
rect -11335 30140 -11261 30265
rect -11222 30208 -11147 30212
rect -11222 30174 -11044 30208
rect -11222 30171 -11147 30174
rect -11567 29978 -11389 30011
rect -11477 29975 -11389 29978
rect -11635 29914 -11545 29917
rect -11635 29880 -11459 29914
rect -11635 29875 -11545 29880
rect -11635 29721 -11601 29875
rect -11423 29817 -11389 29975
rect -11477 29816 -11389 29817
rect -11567 29782 -11389 29816
rect -11477 29781 -11389 29782
rect -11423 29756 -11389 29781
rect -11222 30014 -11188 30171
rect -10998 30115 -10964 30267
rect -11067 30110 -10964 30115
rect -11152 30076 -10964 30110
rect -11067 30071 -10964 30076
rect -11222 30012 -11139 30014
rect -11222 29978 -11044 30012
rect -11222 29973 -11139 29978
rect -11222 29820 -11188 29973
rect -10998 29919 -10964 30071
rect -11067 29914 -10964 29919
rect -11152 29880 -10964 29914
rect -11067 29875 -10964 29880
rect -11222 29816 -11139 29820
rect -11222 29782 -11044 29816
rect -11222 29779 -11139 29782
rect -11222 29756 -11188 29779
rect -11635 29718 -11550 29721
rect -11635 29684 -11459 29718
rect -11635 29679 -11550 29684
rect -11423 29623 -11188 29756
rect -10998 29722 -10964 29875
rect -11056 29718 -10964 29722
rect -11152 29684 -10964 29718
rect -11056 29678 -10964 29684
rect -11148 29623 -11016 29629
rect -11467 29620 -11016 29623
rect -13814 29438 -13463 29472
rect -13814 29242 -13537 29276
rect -13571 29096 -13537 29242
rect -13952 29062 -13537 29096
rect -13952 28598 -13918 29062
rect -13497 29026 -13463 29438
rect -13325 29276 -13291 29536
rect -13017 29472 -12927 29474
rect -13208 29438 -12927 29472
rect -13426 29116 -13372 29255
rect -13325 29242 -13000 29276
rect -13325 29043 -13291 29242
rect -13883 28992 -13463 29026
rect -13421 29009 -13291 29043
rect -13238 29144 -13000 29178
rect -13883 28914 -13849 28992
rect -13421 28931 -13387 29009
rect -13883 28880 -13606 28914
rect -13570 28897 -13387 28931
rect -13238 28914 -13199 29144
rect -13883 28718 -13849 28880
rect -13570 28816 -13536 28897
rect -13814 28782 -13536 28816
rect -13883 28684 -13606 28718
rect -13952 28564 -13606 28598
rect -13952 28402 -13918 28564
rect -13570 28500 -13536 28782
rect -13238 28880 -13000 28914
rect -13238 28878 -13199 28880
rect -13814 28466 -13536 28500
rect -13952 28368 -13606 28402
rect -13570 28234 -13536 28466
rect -13456 28367 -13402 28506
rect -12963 28500 -12927 29438
rect -13208 28466 -12927 28500
rect -11567 29586 -11016 29620
rect -11467 29583 -11016 29586
rect -11467 29582 -11138 29583
rect -11467 29581 -11181 29582
rect -11301 29384 -11244 29581
rect -11310 29216 -11236 29384
rect -11578 29174 -11186 29180
rect -11582 29140 -11094 29174
rect -11578 29134 -11186 29140
rect -11325 28984 -11279 29134
rect -11390 28978 -11186 28984
rect -11582 28944 -11094 28978
rect -11390 28938 -11186 28944
rect -13173 28234 -13037 28240
rect -13570 28200 -13037 28234
rect -13173 28194 -13037 28200
rect -13494 27640 -13440 27779
rect -12467 28237 -12331 28240
rect -12078 28237 -12032 28333
rect -12467 28197 -12032 28237
rect -11325 28788 -11279 28938
rect -11390 28782 -11186 28788
rect -11582 28748 -11094 28782
rect -11390 28742 -11186 28748
rect -11317 28712 -11247 28742
rect -11303 28662 -11258 28712
rect -11303 28642 -11143 28662
rect -11482 28602 -11143 28642
rect -11482 28597 -11258 28602
rect -11482 28438 -11437 28597
rect -11560 28381 -11396 28438
rect -12467 28194 -12331 28197
rect -11578 28217 -11186 28223
rect -11582 28183 -11094 28217
rect -11578 28177 -11186 28183
rect -11325 28027 -11279 28177
rect -11390 28021 -11186 28027
rect -11582 27987 -11094 28021
rect -11390 27981 -11186 27987
rect -11325 27831 -11279 27981
rect -13623 27591 -13189 27596
rect -13814 27557 -13000 27591
rect -13623 27553 -13189 27557
rect -13426 27453 -13380 27553
rect -13621 27282 -13191 27286
rect -13814 27248 -13000 27282
rect -13621 27243 -13191 27248
rect -13500 27025 -13446 27164
rect -13282 27147 -13236 27243
rect -13325 27036 -13000 27070
rect -13814 26938 -13463 26972
rect -13814 26742 -13537 26776
rect -13571 26596 -13537 26742
rect -13952 26562 -13537 26596
rect -13952 26098 -13918 26562
rect -13497 26526 -13463 26938
rect -13325 26776 -13291 27036
rect -13017 26972 -12927 26974
rect -13208 26938 -12927 26972
rect -13426 26616 -13372 26755
rect -13325 26742 -13000 26776
rect -13325 26543 -13291 26742
rect -13883 26492 -13463 26526
rect -13421 26509 -13291 26543
rect -13238 26644 -13000 26678
rect -13883 26414 -13849 26492
rect -13421 26431 -13387 26509
rect -13883 26380 -13606 26414
rect -13570 26397 -13387 26431
rect -13238 26414 -13199 26644
rect -13883 26218 -13849 26380
rect -13570 26316 -13536 26397
rect -13814 26282 -13536 26316
rect -13883 26184 -13606 26218
rect -13952 26064 -13606 26098
rect -13952 25902 -13918 26064
rect -13570 26000 -13536 26282
rect -13238 26380 -13000 26414
rect -13238 26378 -13199 26380
rect -13814 25966 -13536 26000
rect -13952 25868 -13606 25902
rect -13570 25791 -13536 25966
rect -13456 25867 -13402 26006
rect -12963 26000 -12927 26938
rect -13208 25966 -12927 26000
rect -11390 27825 -11186 27831
rect -11582 27791 -11094 27825
rect -11390 27785 -11186 27791
rect -11317 27730 -11247 27785
rect -11509 27657 -11247 27730
rect -11509 27656 -11341 27657
rect -11635 27606 -11556 27607
rect -11482 27606 -11126 27612
rect -11056 27606 -10964 27611
rect -11635 27572 -10964 27606
rect -11635 27571 -11556 27572
rect -11635 27411 -11601 27571
rect -11482 27565 -11126 27572
rect -11056 27567 -10964 27572
rect -11475 27508 -11389 27509
rect -11567 27474 -11389 27508
rect -11475 27473 -11389 27474
rect -11635 27410 -11546 27411
rect -11635 27376 -11459 27410
rect -11635 27369 -11546 27376
rect -11635 27217 -11601 27369
rect -11567 27311 -11459 27312
rect -11423 27311 -11389 27473
rect -11335 27440 -11261 27565
rect -11222 27508 -11147 27512
rect -11222 27474 -11044 27508
rect -11222 27471 -11147 27474
rect -11567 27278 -11389 27311
rect -11477 27275 -11389 27278
rect -11635 27214 -11545 27217
rect -11635 27180 -11459 27214
rect -11635 27175 -11545 27180
rect -11635 27021 -11601 27175
rect -11423 27117 -11389 27275
rect -11477 27116 -11389 27117
rect -11567 27082 -11389 27116
rect -11477 27081 -11389 27082
rect -11423 27056 -11389 27081
rect -11222 27314 -11188 27471
rect -10998 27415 -10964 27567
rect -11067 27410 -10964 27415
rect -11152 27376 -10964 27410
rect -11067 27371 -10964 27376
rect -11222 27312 -11139 27314
rect -11222 27278 -11044 27312
rect -11222 27273 -11139 27278
rect -11222 27120 -11188 27273
rect -10998 27219 -10964 27371
rect -11067 27214 -10964 27219
rect -11152 27180 -10964 27214
rect -11067 27175 -10964 27180
rect -11222 27116 -11139 27120
rect -11222 27082 -11044 27116
rect -11222 27079 -11139 27082
rect -11222 27056 -11188 27079
rect -11635 27018 -11550 27021
rect -11635 26984 -11459 27018
rect -11635 26979 -11550 26984
rect -11423 26923 -11188 27056
rect -10998 27022 -10964 27175
rect -11056 27018 -10964 27022
rect -11152 26984 -10964 27018
rect -11056 26978 -10964 26984
rect -11467 26920 -11138 26923
rect -11567 26886 -11044 26920
rect -11467 26882 -11138 26886
rect -11467 26881 -11181 26882
rect -11304 26684 -11251 26881
rect -10928 26797 -10889 31188
rect -8365 33221 -7925 33255
rect -8365 33220 -8224 33221
rect -8365 33059 -8328 33220
rect -7862 33157 -7827 33335
rect -8233 33123 -7827 33157
rect -7925 33122 -7827 33123
rect -7771 33118 -7737 33905
rect -7572 33899 -7502 33905
rect -7700 33734 -7654 33870
rect -7693 33306 -7655 33734
rect -7618 33653 -7480 33699
rect -7618 33507 -7564 33653
rect -7598 33433 -7317 33467
rect -7700 33171 -7646 33306
rect -7598 33271 -7561 33433
rect -7598 33237 -7317 33271
rect -8365 33025 -7925 33059
rect -8365 33024 -8222 33025
rect -8365 32848 -8331 33024
rect -7778 32983 -7724 33118
rect -7598 33075 -7561 33237
rect -7598 33041 -7317 33075
rect -7598 32949 -7561 33041
rect -7861 32946 -7561 32949
rect -8233 32912 -7561 32946
rect -8365 32814 -7925 32848
rect -7861 32750 -7827 32912
rect -8233 32716 -7827 32750
rect -7773 32507 -7736 32912
rect -7780 32372 -7726 32507
rect -8233 32303 -7317 32337
rect -7780 32152 -7727 32303
rect -8090 31398 -8030 31530
rect -10418 31019 -10358 31094
rect -10457 31018 -10171 31019
rect -10500 31014 -10171 31018
rect -10594 30980 -10071 31014
rect -10500 30977 -10171 30980
rect -10674 30916 -10582 30922
rect -10674 30882 -10486 30916
rect -10674 30878 -10582 30882
rect -10674 30725 -10640 30878
rect -10450 30844 -10215 30977
rect -10088 30916 -10003 30921
rect -10179 30882 -10003 30916
rect -10088 30879 -10003 30882
rect -10450 30821 -10416 30844
rect -10499 30818 -10416 30821
rect -10594 30784 -10416 30818
rect -10499 30780 -10416 30784
rect -10674 30720 -10571 30725
rect -10674 30686 -10486 30720
rect -10674 30681 -10571 30686
rect -10674 30529 -10640 30681
rect -10450 30627 -10416 30780
rect -10499 30622 -10416 30627
rect -10594 30588 -10416 30622
rect -10499 30586 -10416 30588
rect -10674 30524 -10571 30529
rect -10674 30490 -10486 30524
rect -10674 30485 -10571 30490
rect -10674 30333 -10640 30485
rect -10450 30429 -10416 30586
rect -10249 30819 -10215 30844
rect -10249 30818 -10161 30819
rect -10249 30784 -10071 30818
rect -10249 30783 -10161 30784
rect -10249 30625 -10215 30783
rect -10037 30725 -10003 30879
rect -10093 30720 -10003 30725
rect -10179 30686 -10003 30720
rect -10093 30683 -10003 30686
rect -10249 30622 -10161 30625
rect -10249 30589 -10071 30622
rect -10491 30426 -10416 30429
rect -10594 30392 -10416 30426
rect -10491 30388 -10416 30392
rect -10377 30335 -10303 30460
rect -10249 30427 -10215 30589
rect -10179 30588 -10071 30589
rect -10037 30531 -10003 30683
rect -10092 30524 -10003 30531
rect -10179 30490 -10003 30524
rect -10092 30489 -10003 30490
rect -10249 30426 -10163 30427
rect -10249 30392 -10071 30426
rect -10249 30391 -10163 30392
rect -10674 30328 -10582 30333
rect -10512 30328 -10156 30335
rect -10037 30329 -10003 30489
rect -10082 30328 -10003 30329
rect -10674 30294 -10003 30328
rect -10674 30289 -10582 30294
rect -10512 30288 -10156 30294
rect -10082 30293 -10003 30294
rect -8524 31019 -8464 31094
rect -8711 31018 -8425 31019
rect -8711 31014 -8382 31018
rect -8811 30980 -8288 31014
rect -8711 30977 -8382 30980
rect -10297 30243 -10129 30244
rect -10391 30170 -10129 30243
rect -10391 30115 -10321 30170
rect -10452 30109 -10248 30115
rect -10544 30075 -10056 30109
rect -10452 30069 -10248 30075
rect -10359 29919 -10313 30069
rect -10452 29913 -10248 29919
rect -10544 29879 -10056 29913
rect -10452 29873 -10248 29879
rect -10359 29723 -10313 29873
rect -10452 29717 -10060 29723
rect -10544 29683 -10056 29717
rect -10452 29677 -10060 29683
rect -8879 30916 -8794 30921
rect -8879 30882 -8703 30916
rect -8879 30879 -8794 30882
rect -8879 30725 -8845 30879
rect -8667 30844 -8432 30977
rect -8300 30916 -8208 30922
rect -8396 30882 -8208 30916
rect -8300 30878 -8208 30882
rect -8667 30819 -8633 30844
rect -8721 30818 -8633 30819
rect -8811 30784 -8633 30818
rect -8721 30783 -8633 30784
rect -8879 30720 -8789 30725
rect -8879 30686 -8703 30720
rect -8879 30683 -8789 30686
rect -8879 30531 -8845 30683
rect -8667 30625 -8633 30783
rect -8721 30622 -8633 30625
rect -8811 30589 -8633 30622
rect -8811 30588 -8703 30589
rect -8879 30524 -8790 30531
rect -8879 30490 -8703 30524
rect -8879 30489 -8790 30490
rect -8879 30329 -8845 30489
rect -8667 30427 -8633 30589
rect -8466 30821 -8432 30844
rect -8466 30818 -8383 30821
rect -8466 30784 -8288 30818
rect -8466 30780 -8383 30784
rect -8466 30627 -8432 30780
rect -8242 30725 -8208 30878
rect -8311 30720 -8208 30725
rect -8396 30686 -8208 30720
rect -8311 30681 -8208 30686
rect -8466 30622 -8383 30627
rect -8466 30588 -8288 30622
rect -8466 30586 -8383 30588
rect -8719 30426 -8633 30427
rect -8811 30392 -8633 30426
rect -8719 30391 -8633 30392
rect -8579 30335 -8505 30460
rect -8466 30429 -8432 30586
rect -8242 30529 -8208 30681
rect -8311 30524 -8208 30529
rect -8396 30490 -8208 30524
rect -8311 30485 -8208 30490
rect -8466 30426 -8391 30429
rect -8466 30392 -8288 30426
rect -8466 30388 -8391 30392
rect -8879 30328 -8800 30329
rect -8726 30328 -8370 30335
rect -8242 30333 -8208 30485
rect -8300 30328 -8208 30333
rect -8879 30294 -8208 30328
rect -8879 30293 -8800 30294
rect -8726 30288 -8370 30294
rect -8300 30289 -8208 30294
rect -8753 30243 -8585 30244
rect -8753 30170 -8491 30243
rect -8561 30115 -8491 30170
rect -8634 30109 -8430 30115
rect -8826 30075 -8338 30109
rect -8634 30069 -8430 30075
rect -8569 29919 -8523 30069
rect -8634 29913 -8430 29919
rect -8826 29879 -8338 29913
rect -8634 29873 -8430 29879
rect -8569 29723 -8523 29873
rect -8822 29717 -8430 29723
rect -8826 29683 -8338 29717
rect -8822 29677 -8430 29683
rect -10242 29462 -10078 29519
rect -10192 29376 -10130 29462
rect -10391 29314 -10130 29376
rect -10391 29278 -10321 29314
rect -10452 29272 -10248 29278
rect -8804 29462 -8640 29519
rect -8554 29473 -8480 29641
rect -8752 29376 -8690 29462
rect -8543 29413 -8321 29473
rect -8752 29314 -8491 29376
rect -8561 29278 -8491 29314
rect -10544 29238 -10056 29272
rect -10452 29232 -10248 29238
rect -10359 29082 -10313 29232
rect -10452 29076 -10248 29082
rect -10544 29042 -10056 29076
rect -10452 29036 -10248 29042
rect -11310 26516 -11236 26684
rect -10941 26665 -10881 26797
rect -11578 26474 -11186 26480
rect -11582 26440 -11094 26474
rect -11578 26434 -11186 26440
rect -11325 26284 -11279 26434
rect -11390 26278 -11186 26284
rect -11582 26244 -11094 26278
rect -11390 26238 -11186 26244
rect -11325 26088 -11279 26238
rect -10928 26259 -10889 26665
rect -10359 28886 -10313 29036
rect -10452 28880 -10060 28886
rect -10544 28846 -10056 28880
rect -10452 28840 -10060 28846
rect -10402 28636 -10328 28804
rect -8634 29272 -8430 29278
rect -8826 29238 -8338 29272
rect -8634 29232 -8430 29238
rect -8569 29082 -8523 29232
rect -8634 29076 -8430 29082
rect -8826 29042 -8338 29076
rect -8634 29036 -8430 29042
rect -8569 28886 -8523 29036
rect -8079 29516 -8040 31398
rect -7696 31799 -7304 31805
rect -7788 31765 -7300 31799
rect -7696 31759 -7304 31765
rect -7603 31609 -7557 31759
rect -7696 31603 -7492 31609
rect -7788 31569 -7300 31603
rect -7696 31563 -7492 31569
rect -7603 31413 -7557 31563
rect -7696 31407 -7492 31413
rect -7788 31373 -7300 31407
rect -7696 31367 -7492 31373
rect -7635 31337 -7565 31367
rect -7629 31279 -7587 31337
rect -7715 31219 -7583 31279
rect -7486 31081 -7322 31138
rect -6215 31043 -6179 35410
rect -6135 33540 -6101 35508
rect -5849 35679 -5713 35685
rect -5849 35678 -5712 35679
rect -5346 35678 -5312 35966
rect -4964 35902 -4930 36064
rect -5276 35868 -4930 35902
rect -5849 35644 -5312 35678
rect -5849 35639 -5713 35644
rect -5442 35140 -5388 35279
rect -5693 35091 -5259 35096
rect -5882 35057 -5068 35091
rect -5693 35053 -5259 35057
rect -5502 34953 -5456 35053
rect -5691 34782 -5261 34786
rect -5882 34748 -5068 34782
rect -5691 34743 -5261 34748
rect -5646 34647 -5600 34743
rect -6144 33404 -6098 33540
rect -6135 33371 -6101 33404
rect -5882 34536 -5557 34570
rect -5955 34472 -5865 34474
rect -5955 34438 -5674 34472
rect -5955 33500 -5919 34438
rect -5591 34276 -5557 34536
rect -5436 34525 -5382 34664
rect -5882 34242 -5557 34276
rect -5419 34438 -5068 34472
rect -5882 34144 -5644 34178
rect -5683 33914 -5644 34144
rect -5591 34043 -5557 34242
rect -5510 34116 -5456 34255
rect -5591 34009 -5461 34043
rect -5882 33880 -5644 33914
rect -5495 33931 -5461 34009
rect -5419 34026 -5385 34438
rect -5345 34242 -5068 34276
rect -5345 34096 -5311 34242
rect -5345 34062 -4930 34096
rect -5419 33992 -4999 34026
rect -5495 33897 -5312 33931
rect -5033 33914 -4999 33992
rect -5683 33878 -5644 33880
rect -5346 33816 -5312 33897
rect -5276 33880 -4999 33914
rect -5346 33782 -5068 33816
rect -5955 33466 -5674 33500
rect -5480 33367 -5426 33506
rect -5346 33500 -5312 33782
rect -5033 33718 -4999 33880
rect -5276 33684 -4999 33718
rect -4964 33598 -4930 34062
rect -5276 33564 -4930 33598
rect -5346 33466 -5068 33500
rect -5849 33262 -5713 33268
rect -5346 33262 -5312 33466
rect -4964 33402 -4930 33564
rect -5276 33368 -4930 33402
rect -5849 33228 -5311 33262
rect -5849 33222 -5713 33228
rect -5442 32640 -5388 32779
rect -5693 32591 -5259 32596
rect -5882 32557 -5068 32591
rect -5693 32553 -5259 32557
rect -5502 32453 -5456 32553
rect -5691 32282 -5261 32286
rect -5882 32248 -5068 32282
rect -5691 32243 -5261 32248
rect -5646 32147 -5600 32243
rect -6215 30994 -6085 31043
rect -7696 30917 -7304 30923
rect -7788 30883 -7300 30917
rect -7696 30877 -7304 30883
rect -7603 30727 -7557 30877
rect -6131 30907 -6085 30994
rect -7696 30721 -7492 30727
rect -7788 30687 -7300 30721
rect -7696 30681 -7492 30687
rect -7603 30531 -7557 30681
rect -5882 32036 -5557 32070
rect -5955 31972 -5865 31974
rect -5955 31938 -5674 31972
rect -5955 31000 -5919 31938
rect -5591 31776 -5557 32036
rect -5436 32025 -5382 32164
rect -5882 31742 -5557 31776
rect -5419 31938 -5068 31972
rect -5882 31644 -5644 31678
rect -5683 31414 -5644 31644
rect -5591 31543 -5557 31742
rect -5510 31616 -5456 31755
rect -5591 31509 -5461 31543
rect -5882 31380 -5644 31414
rect -5495 31431 -5461 31509
rect -5419 31526 -5385 31938
rect -5345 31742 -5068 31776
rect -5345 31596 -5311 31742
rect -5345 31562 -4930 31596
rect -5419 31492 -4999 31526
rect -5495 31397 -5312 31431
rect -5033 31414 -4999 31492
rect -5683 31378 -5644 31380
rect -5346 31316 -5312 31397
rect -5276 31380 -4999 31414
rect -5346 31282 -5068 31316
rect -5955 30966 -5674 31000
rect -5480 30867 -5426 31006
rect -5346 31000 -5312 31282
rect -5033 31218 -4999 31380
rect -5276 31184 -4999 31218
rect -4964 31098 -4930 31562
rect -5276 31064 -4930 31098
rect -5346 30966 -5068 31000
rect -7696 30525 -7492 30531
rect -7788 30491 -7300 30525
rect -7696 30485 -7492 30491
rect -7635 30430 -7565 30485
rect -7635 30357 -7373 30430
rect -7541 30356 -7373 30357
rect -8089 29384 -8029 29516
rect -8822 28880 -8430 28886
rect -8826 28846 -8338 28880
rect -8822 28840 -8430 28846
rect -10395 28614 -10335 28636
rect -10416 28319 -10356 28410
rect -8554 28636 -8480 28804
rect -8547 28614 -8487 28636
rect -10457 28318 -10171 28319
rect -10500 28314 -10171 28318
rect -10594 28280 -10071 28314
rect -10500 28277 -10171 28280
rect -10674 28216 -10582 28222
rect -10674 28182 -10486 28216
rect -10674 28178 -10582 28182
rect -10674 28025 -10640 28178
rect -10450 28144 -10215 28277
rect -10088 28216 -10003 28221
rect -10179 28182 -10003 28216
rect -10088 28179 -10003 28182
rect -10450 28121 -10416 28144
rect -10499 28118 -10416 28121
rect -10594 28084 -10416 28118
rect -10499 28080 -10416 28084
rect -10674 28020 -10571 28025
rect -10674 27986 -10486 28020
rect -10674 27981 -10571 27986
rect -10674 27829 -10640 27981
rect -10450 27927 -10416 28080
rect -10499 27922 -10416 27927
rect -10594 27888 -10416 27922
rect -10499 27886 -10416 27888
rect -10674 27824 -10571 27829
rect -10674 27790 -10486 27824
rect -10674 27785 -10571 27790
rect -10674 27633 -10640 27785
rect -10450 27729 -10416 27886
rect -10249 28119 -10215 28144
rect -10249 28118 -10161 28119
rect -10249 28084 -10071 28118
rect -10249 28083 -10161 28084
rect -10249 27925 -10215 28083
rect -10037 28025 -10003 28179
rect -10093 28020 -10003 28025
rect -10179 27986 -10003 28020
rect -10093 27983 -10003 27986
rect -10249 27922 -10161 27925
rect -10249 27889 -10071 27922
rect -10491 27726 -10416 27729
rect -10594 27692 -10416 27726
rect -10491 27688 -10416 27692
rect -10377 27635 -10303 27760
rect -10249 27727 -10215 27889
rect -10179 27888 -10071 27889
rect -10037 27831 -10003 27983
rect -10092 27824 -10003 27831
rect -10179 27790 -10003 27824
rect -10092 27789 -10003 27790
rect -10249 27726 -10163 27727
rect -10249 27692 -10071 27726
rect -10249 27691 -10163 27692
rect -10674 27628 -10582 27633
rect -10512 27628 -10156 27635
rect -10037 27629 -10003 27789
rect -10082 27628 -10003 27629
rect -10674 27594 -10003 27628
rect -10674 27589 -10582 27594
rect -10512 27588 -10156 27594
rect -10082 27593 -10003 27594
rect -8526 28319 -8466 28410
rect -8711 28318 -8425 28319
rect -8711 28314 -8382 28318
rect -8811 28280 -8288 28314
rect -8711 28277 -8382 28280
rect -10297 27543 -10129 27544
rect -10391 27470 -10129 27543
rect -8879 28216 -8794 28221
rect -8879 28182 -8703 28216
rect -8879 28179 -8794 28182
rect -8879 28025 -8845 28179
rect -8667 28144 -8432 28277
rect -8300 28216 -8208 28222
rect -8396 28182 -8208 28216
rect -8300 28178 -8208 28182
rect -8667 28119 -8633 28144
rect -8721 28118 -8633 28119
rect -8811 28084 -8633 28118
rect -8721 28083 -8633 28084
rect -8879 28020 -8789 28025
rect -8879 27986 -8703 28020
rect -8879 27983 -8789 27986
rect -8879 27831 -8845 27983
rect -8667 27925 -8633 28083
rect -8721 27922 -8633 27925
rect -8811 27889 -8633 27922
rect -8811 27888 -8703 27889
rect -8879 27824 -8790 27831
rect -8879 27790 -8703 27824
rect -8879 27789 -8790 27790
rect -8879 27629 -8845 27789
rect -8667 27727 -8633 27889
rect -8466 28121 -8432 28144
rect -8466 28118 -8383 28121
rect -8466 28084 -8288 28118
rect -8466 28080 -8383 28084
rect -8466 27927 -8432 28080
rect -8242 28025 -8208 28178
rect -8311 28020 -8208 28025
rect -8396 27986 -8208 28020
rect -8311 27981 -8208 27986
rect -8466 27922 -8383 27927
rect -8466 27888 -8288 27922
rect -8466 27886 -8383 27888
rect -8719 27726 -8633 27727
rect -8811 27692 -8633 27726
rect -8719 27691 -8633 27692
rect -8579 27635 -8505 27760
rect -8466 27729 -8432 27886
rect -8242 27829 -8208 27981
rect -8311 27824 -8208 27829
rect -8396 27790 -8208 27824
rect -8311 27785 -8208 27790
rect -8466 27726 -8391 27729
rect -8466 27692 -8288 27726
rect -8466 27688 -8391 27692
rect -8879 27628 -8800 27629
rect -8726 27628 -8370 27635
rect -8242 27633 -8208 27785
rect -8300 27628 -8208 27633
rect -8879 27594 -8208 27628
rect -8879 27593 -8800 27594
rect -8726 27588 -8370 27594
rect -8300 27589 -8208 27594
rect -10391 27415 -10321 27470
rect -10452 27409 -10248 27415
rect -10544 27375 -10056 27409
rect -10452 27369 -10248 27375
rect -10359 27219 -10313 27369
rect -10452 27213 -10248 27219
rect -10544 27179 -10056 27213
rect -10452 27173 -10248 27179
rect -10359 27023 -10313 27173
rect -10452 27017 -10060 27023
rect -10544 26983 -10056 27017
rect -10452 26977 -10060 26983
rect -10402 26773 -10328 26941
rect -8753 27543 -8585 27544
rect -8753 27470 -8491 27543
rect -8561 27415 -8491 27470
rect -8634 27409 -8430 27415
rect -8826 27375 -8338 27409
rect -8634 27369 -8430 27375
rect -8569 27219 -8523 27369
rect -8634 27213 -8430 27219
rect -8826 27179 -8338 27213
rect -8079 28575 -8040 29384
rect -8090 28438 -8030 28575
rect -8634 27173 -8430 27179
rect -8569 27023 -8523 27173
rect -8822 27017 -8430 27023
rect -8826 26983 -8338 27017
rect -8822 26977 -8430 26983
rect -10402 26761 -10339 26773
rect -10242 26762 -10078 26819
rect -10546 26738 -10339 26761
rect -10546 26701 -10340 26738
rect -10191 26665 -10142 26762
rect -10391 26619 -10142 26665
rect -8804 26762 -8640 26819
rect -10391 26578 -10321 26619
rect -10452 26572 -10248 26578
rect -10544 26538 -10056 26572
rect -10452 26532 -10248 26538
rect -10359 26382 -10313 26532
rect -10452 26376 -10248 26382
rect -10544 26342 -10056 26376
rect -8740 26665 -8691 26762
rect -8740 26619 -8491 26665
rect -8561 26578 -8491 26619
rect -8634 26572 -8430 26578
rect -8826 26538 -8338 26572
rect -8634 26532 -8430 26538
rect -8569 26382 -8523 26532
rect -8634 26376 -8430 26382
rect -10452 26336 -10248 26342
rect -11390 26082 -11186 26088
rect -11582 26048 -11094 26082
rect -11390 26042 -11186 26048
rect -10359 26186 -10313 26336
rect -8826 26342 -8338 26376
rect -8634 26336 -8430 26342
rect -10452 26180 -10060 26186
rect -10544 26146 -10056 26180
rect -10452 26140 -10060 26146
rect -11317 26012 -11247 26042
rect -11308 25977 -11269 26012
rect -10911 25977 -10774 25988
rect -10402 25977 -10328 26104
rect -8569 26186 -8523 26336
rect -8079 26259 -8040 28438
rect -7918 30306 -7826 30311
rect -7756 30306 -7400 30312
rect -7326 30306 -7247 30307
rect -7918 30272 -7247 30306
rect -7918 30267 -7826 30272
rect -7918 30115 -7884 30267
rect -7756 30265 -7400 30272
rect -7326 30271 -7247 30272
rect -7735 30208 -7660 30212
rect -7838 30174 -7660 30208
rect -7735 30171 -7660 30174
rect -7918 30110 -7815 30115
rect -7918 30076 -7730 30110
rect -7918 30071 -7815 30076
rect -7918 29919 -7884 30071
rect -7694 30014 -7660 30171
rect -7621 30140 -7547 30265
rect -7493 30208 -7407 30209
rect -7493 30174 -7315 30208
rect -7493 30173 -7407 30174
rect -7743 30012 -7660 30014
rect -7838 29978 -7660 30012
rect -7743 29973 -7660 29978
rect -7918 29914 -7815 29919
rect -7918 29880 -7730 29914
rect -7918 29875 -7815 29880
rect -7918 29722 -7884 29875
rect -7694 29820 -7660 29973
rect -7743 29816 -7660 29820
rect -7838 29782 -7660 29816
rect -7743 29779 -7660 29782
rect -7694 29756 -7660 29779
rect -7493 30011 -7459 30173
rect -7281 30111 -7247 30271
rect -7336 30110 -7247 30111
rect -7423 30076 -7247 30110
rect -7336 30069 -7247 30076
rect -7423 30011 -7315 30012
rect -7493 29978 -7315 30011
rect -7493 29975 -7405 29978
rect -7493 29817 -7459 29975
rect -7281 29917 -7247 30069
rect -7337 29914 -7247 29917
rect -7423 29880 -7247 29914
rect -7337 29875 -7247 29880
rect -7493 29816 -7405 29817
rect -7493 29782 -7315 29816
rect -7493 29781 -7405 29782
rect -7493 29756 -7459 29781
rect -7918 29718 -7826 29722
rect -7918 29684 -7730 29718
rect -7918 29678 -7826 29684
rect -7866 29623 -7734 29629
rect -7694 29623 -7459 29756
rect -7281 29721 -7247 29875
rect -7332 29718 -7247 29721
rect -7423 29684 -7247 29718
rect -7332 29679 -7247 29684
rect -7866 29620 -7415 29623
rect -7866 29586 -7315 29620
rect -5849 30782 -5713 30788
rect -5346 30782 -5312 30966
rect -4964 30902 -4930 31064
rect -5276 30868 -4930 30902
rect -5849 30748 -5312 30782
rect -5849 30742 -5713 30748
rect -5442 30140 -5388 30279
rect -5693 30091 -5259 30096
rect -5882 30057 -5068 30091
rect -5693 30053 -5259 30057
rect -7866 29583 -7415 29586
rect -7744 29582 -7415 29583
rect -7701 29581 -7415 29582
rect -7638 29384 -7581 29581
rect -7646 29216 -7572 29384
rect -5502 29953 -5456 30053
rect -5691 29782 -5261 29786
rect -5882 29748 -5068 29782
rect -5691 29743 -5261 29748
rect -5646 29647 -5600 29743
rect -7696 29174 -7304 29180
rect -7788 29140 -7300 29174
rect -7696 29134 -7304 29140
rect -7603 28984 -7557 29134
rect -7696 28978 -7492 28984
rect -7788 28944 -7300 28978
rect -7696 28938 -7492 28944
rect -7603 28788 -7557 28938
rect -7696 28782 -7492 28788
rect -7788 28748 -7300 28782
rect -7696 28742 -7492 28748
rect -7635 28712 -7565 28742
rect -7624 28662 -7579 28712
rect -7739 28642 -7579 28662
rect -7739 28602 -7400 28642
rect -7624 28597 -7400 28602
rect -7714 28487 -7582 28547
rect -7641 28427 -7583 28487
rect -7445 28438 -7400 28597
rect -7646 28259 -7572 28427
rect -7486 28381 -7322 28438
rect -5882 29536 -5557 29570
rect -5955 29472 -5865 29474
rect -5955 29438 -5674 29472
rect -5955 28500 -5919 29438
rect -5591 29276 -5557 29536
rect -5436 29525 -5382 29664
rect -5882 29242 -5557 29276
rect -5419 29438 -5068 29472
rect -5882 29144 -5644 29178
rect -5683 28914 -5644 29144
rect -5591 29043 -5557 29242
rect -5510 29116 -5456 29255
rect -5591 29009 -5461 29043
rect -5882 28880 -5644 28914
rect -5495 28931 -5461 29009
rect -5419 29026 -5385 29438
rect -5345 29242 -5068 29276
rect -5345 29096 -5311 29242
rect -5345 29062 -4930 29096
rect -5419 28992 -4999 29026
rect -5495 28897 -5312 28931
rect -5033 28914 -4999 28992
rect -5683 28878 -5644 28880
rect -5346 28816 -5312 28897
rect -5276 28880 -4999 28914
rect -5346 28782 -5068 28816
rect -5955 28466 -5674 28500
rect -5480 28367 -5426 28506
rect -5346 28500 -5312 28782
rect -5033 28718 -4999 28880
rect -5276 28684 -4999 28718
rect -4964 28598 -4930 29062
rect -5276 28564 -4930 28598
rect -5346 28466 -5068 28500
rect -7696 28217 -7304 28223
rect -7788 28183 -7300 28217
rect -7696 28177 -7304 28183
rect -7603 28027 -7557 28177
rect -6850 28237 -6804 28333
rect -6551 28237 -6415 28240
rect -6850 28197 -6415 28237
rect -6551 28194 -6415 28197
rect -7696 28021 -7492 28027
rect -7788 27987 -7300 28021
rect -7696 27981 -7492 27987
rect -7603 27831 -7557 27981
rect -7696 27825 -7492 27831
rect -7788 27791 -7300 27825
rect -7696 27785 -7492 27791
rect -7635 27730 -7565 27785
rect -7635 27657 -7373 27730
rect -7541 27656 -7373 27657
rect -7918 27606 -7826 27611
rect -7756 27606 -7400 27612
rect -7326 27606 -7247 27607
rect -7918 27572 -7247 27606
rect -7918 27567 -7826 27572
rect -7918 27415 -7884 27567
rect -7756 27565 -7400 27572
rect -7326 27571 -7247 27572
rect -7735 27508 -7660 27512
rect -7838 27474 -7660 27508
rect -7735 27471 -7660 27474
rect -7918 27410 -7815 27415
rect -7918 27376 -7730 27410
rect -7918 27371 -7815 27376
rect -7918 27219 -7884 27371
rect -7694 27314 -7660 27471
rect -7621 27440 -7547 27565
rect -7493 27508 -7407 27509
rect -7493 27474 -7315 27508
rect -7493 27473 -7407 27474
rect -7743 27312 -7660 27314
rect -7838 27278 -7660 27312
rect -7743 27273 -7660 27278
rect -7918 27214 -7815 27219
rect -7918 27180 -7730 27214
rect -7918 27175 -7815 27180
rect -7918 27022 -7884 27175
rect -7694 27120 -7660 27273
rect -7743 27116 -7660 27120
rect -7838 27082 -7660 27116
rect -7743 27079 -7660 27082
rect -7694 27056 -7660 27079
rect -7493 27311 -7459 27473
rect -7281 27411 -7247 27571
rect -7336 27410 -7247 27411
rect -7423 27376 -7247 27410
rect -7336 27369 -7247 27376
rect -7423 27311 -7315 27312
rect -7493 27278 -7315 27311
rect -7493 27275 -7405 27278
rect -7493 27117 -7459 27275
rect -7281 27217 -7247 27369
rect -7337 27214 -7247 27217
rect -7423 27180 -7247 27214
rect -7337 27175 -7247 27180
rect -7493 27116 -7405 27117
rect -7493 27082 -7315 27116
rect -7493 27081 -7405 27082
rect -7493 27056 -7459 27081
rect -7918 27018 -7826 27022
rect -7918 26984 -7730 27018
rect -7918 26978 -7826 26984
rect -7694 26923 -7459 27056
rect -7281 27021 -7247 27175
rect -7332 27018 -7247 27021
rect -7423 26984 -7247 27018
rect -7332 26979 -7247 26984
rect -7744 26920 -7415 26923
rect -7838 26886 -7315 26920
rect -6340 27812 -6204 27858
rect -7744 26882 -7415 26886
rect -7701 26881 -7415 26882
rect -7631 26684 -7578 26881
rect -6340 26835 -6270 27812
rect -5845 28234 -5709 28240
rect -5346 28234 -5312 28466
rect -4964 28402 -4930 28564
rect -5276 28368 -4930 28402
rect -5845 28200 -5312 28234
rect -5845 28194 -5709 28200
rect -5442 27640 -5388 27779
rect -5693 27591 -5259 27596
rect -5882 27557 -5068 27591
rect -5693 27553 -5259 27557
rect -5590 27327 -5536 27466
rect -5502 27453 -5456 27553
rect -5691 27282 -5261 27286
rect -5882 27248 -5068 27282
rect -5691 27243 -5261 27248
rect -5646 27147 -5600 27243
rect -6413 26829 -6209 26835
rect -5882 27036 -5557 27070
rect -6605 26795 -6117 26829
rect -6413 26789 -6209 26795
rect -7646 26516 -7572 26684
rect -6348 26639 -6302 26789
rect -6413 26633 -6209 26639
rect -6605 26599 -6117 26633
rect -6413 26593 -6209 26599
rect -7696 26474 -7304 26480
rect -7788 26440 -7300 26474
rect -7696 26434 -7304 26440
rect -8822 26180 -8430 26186
rect -8826 26146 -8338 26180
rect -8822 26140 -8430 26146
rect -11308 25936 -10328 25977
rect -11308 25930 -10358 25936
rect -11306 25929 -10358 25930
rect -10911 25928 -10774 25929
rect -8554 25977 -8480 26104
rect -7603 26284 -7557 26434
rect -6348 26443 -6302 26593
rect -6601 26437 -6209 26443
rect -6605 26403 -6117 26437
rect -6601 26397 -6209 26403
rect -7696 26278 -7492 26284
rect -7788 26244 -7300 26278
rect -7696 26238 -7492 26244
rect -7603 26088 -7557 26238
rect -7696 26082 -7492 26088
rect -7788 26048 -7300 26082
rect -7696 26042 -7492 26048
rect -7635 26012 -7565 26042
rect -8108 25977 -7971 25988
rect -7613 25977 -7574 26012
rect -8554 25936 -7574 25977
rect -8524 25930 -7574 25936
rect -8524 25929 -7576 25930
rect -8108 25928 -7971 25929
rect -12005 25791 -11959 25853
rect -5955 26972 -5865 26974
rect -5955 26938 -5674 26972
rect -5955 26000 -5919 26938
rect -5591 26776 -5557 27036
rect -5436 27025 -5382 27164
rect -5882 26742 -5557 26776
rect -5419 26938 -5068 26972
rect -5882 26644 -5644 26678
rect -5683 26414 -5644 26644
rect -5591 26543 -5557 26742
rect -5510 26616 -5456 26755
rect -5591 26509 -5461 26543
rect -5882 26380 -5644 26414
rect -5495 26431 -5461 26509
rect -5419 26526 -5385 26938
rect -5345 26742 -5068 26776
rect -5345 26596 -5311 26742
rect -5345 26562 -4930 26596
rect -5419 26492 -4999 26526
rect -5495 26397 -5312 26431
rect -5033 26414 -4999 26492
rect -5683 26378 -5644 26380
rect -5584 26249 -5530 26388
rect -5346 26316 -5312 26397
rect -5276 26380 -4999 26414
rect -5346 26282 -5068 26316
rect -5955 25966 -5674 26000
rect -5480 25867 -5426 26006
rect -5346 26000 -5312 26282
rect -5033 26218 -4999 26380
rect -5276 26184 -4999 26218
rect -4964 26098 -4930 26562
rect -5276 26064 -4930 26098
rect -5346 25966 -5068 26000
rect -13570 25757 -11959 25791
rect -12005 25717 -11959 25757
rect -10685 25590 -10621 25732
rect -14173 25304 -13998 25467
rect -14154 13747 -14018 25304
rect -10672 25227 -10638 25590
rect -10567 25315 -10479 25447
rect -10684 25072 -10629 25227
rect -10734 25020 -10624 25026
rect -11026 24986 -10624 25020
rect -10734 24981 -10624 24986
rect -10664 24715 -10624 24981
rect -10567 24957 -10531 25315
rect -6932 25791 -6886 25853
rect -5346 25791 -5312 25966
rect -4964 25902 -4930 26064
rect -5276 25868 -4930 25902
rect -6932 25757 -5312 25791
rect -8061 25607 -7997 25757
rect -6932 25717 -6886 25757
rect -8061 25594 -5704 25607
rect -8060 25573 -5704 25594
rect -5738 25200 -5704 25573
rect -5633 25315 -5526 25447
rect -10485 25118 -10390 25122
rect -10485 25084 -9806 25118
rect -10485 25080 -10390 25084
rect -10576 24802 -10521 24957
rect -10485 24910 -10449 25080
rect -10485 24907 -10396 24910
rect -9814 24907 -9738 24911
rect -10485 24873 -9738 24907
rect -10485 24868 -10396 24873
rect -9814 24869 -9738 24873
rect -10487 24809 -10394 24813
rect -10487 24775 -9806 24809
rect -10487 24771 -10394 24775
rect -10487 24715 -10448 24771
rect -10664 24672 -10448 24715
rect -9772 24713 -9738 24869
rect -9816 24711 -9738 24713
rect -10414 24677 -9738 24711
rect -10684 24586 -10644 24634
rect -10727 24582 -10644 24586
rect -11026 24548 -10644 24582
rect -10727 24542 -10644 24548
rect -10687 24500 -10644 24542
rect -10554 24534 -10499 24672
rect -9816 24671 -9738 24677
rect -10687 24499 -10400 24500
rect -10687 24465 -9806 24499
rect -10687 24457 -10400 24465
rect -13911 24167 -13740 24367
rect -13900 13786 -13764 24167
rect -11043 24115 -10969 24135
rect -10687 24115 -10644 24457
rect -11043 24076 -10536 24115
rect -11043 23967 -10969 24076
rect -11311 23925 -10919 23931
rect -11315 23891 -10827 23925
rect -11311 23885 -10919 23891
rect -11058 23735 -11012 23885
rect -11123 23729 -10919 23735
rect -11315 23695 -10827 23729
rect -11123 23689 -10919 23695
rect -11058 23539 -11012 23689
rect -11123 23533 -10919 23539
rect -11315 23499 -10827 23533
rect -11123 23493 -10919 23499
rect -11050 23463 -10980 23493
rect -11028 23405 -10986 23463
rect -11032 23345 -10900 23405
rect -11028 23288 -10986 23345
rect -11293 23207 -11129 23264
rect -11032 23253 -10974 23288
rect -11043 23085 -10969 23253
rect -10672 23314 -10612 23446
rect -11311 23043 -10919 23049
rect -11315 23009 -10827 23043
rect -11311 23003 -10919 23009
rect -11058 22853 -11012 23003
rect -11123 22847 -10919 22853
rect -11315 22813 -10827 22847
rect -11123 22807 -10919 22813
rect -11058 22657 -11012 22807
rect -11123 22651 -10919 22657
rect -11315 22617 -10827 22651
rect -11123 22611 -10919 22617
rect -11050 22556 -10980 22611
rect -11242 22483 -10980 22556
rect -11242 22482 -11074 22483
rect -11368 22432 -11289 22433
rect -11215 22432 -10859 22438
rect -10789 22432 -10697 22437
rect -11368 22398 -10697 22432
rect -11368 22397 -11289 22398
rect -11368 22237 -11334 22397
rect -11215 22391 -10859 22398
rect -10789 22393 -10697 22398
rect -11208 22334 -11122 22335
rect -11300 22300 -11122 22334
rect -11208 22299 -11122 22300
rect -11368 22236 -11279 22237
rect -11368 22202 -11192 22236
rect -11368 22195 -11279 22202
rect -11368 22043 -11334 22195
rect -11300 22137 -11192 22138
rect -11156 22137 -11122 22299
rect -11068 22266 -10994 22391
rect -10955 22334 -10880 22338
rect -10955 22300 -10777 22334
rect -10955 22297 -10880 22300
rect -11300 22104 -11122 22137
rect -11210 22101 -11122 22104
rect -11368 22040 -11278 22043
rect -11368 22006 -11192 22040
rect -11368 22001 -11278 22006
rect -11368 21847 -11334 22001
rect -11156 21943 -11122 22101
rect -11210 21942 -11122 21943
rect -11300 21908 -11122 21942
rect -11210 21907 -11122 21908
rect -11156 21882 -11122 21907
rect -10955 22140 -10921 22297
rect -10731 22241 -10697 22393
rect -10800 22236 -10697 22241
rect -10885 22202 -10697 22236
rect -10800 22197 -10697 22202
rect -10955 22138 -10872 22140
rect -10955 22104 -10777 22138
rect -10955 22099 -10872 22104
rect -10955 21946 -10921 22099
rect -10731 22045 -10697 22197
rect -10800 22040 -10697 22045
rect -10885 22006 -10697 22040
rect -10800 22001 -10697 22006
rect -10955 21942 -10872 21946
rect -10955 21908 -10777 21942
rect -10955 21905 -10872 21908
rect -10955 21882 -10921 21905
rect -11368 21844 -11283 21847
rect -11368 21810 -11192 21844
rect -11368 21805 -11283 21810
rect -11156 21749 -10921 21882
rect -10731 21848 -10697 22001
rect -10789 21844 -10697 21848
rect -10885 21810 -10697 21844
rect -10789 21804 -10697 21810
rect -10881 21749 -10749 21755
rect -11200 21746 -10749 21749
rect -11300 21712 -10749 21746
rect -11200 21709 -10749 21712
rect -11200 21708 -10871 21709
rect -11200 21707 -10914 21708
rect -11034 21510 -10977 21707
rect -11043 21342 -10969 21510
rect -11311 21300 -10919 21306
rect -11315 21266 -10827 21300
rect -11311 21260 -10919 21266
rect -11058 21110 -11012 21260
rect -11123 21104 -10919 21110
rect -11315 21070 -10827 21104
rect -11123 21064 -10919 21070
rect -11058 20914 -11012 21064
rect -11123 20908 -10919 20914
rect -11315 20874 -10827 20908
rect -11123 20868 -10919 20874
rect -11050 20838 -10980 20868
rect -11036 20788 -10991 20838
rect -11036 20768 -10876 20788
rect -11215 20728 -10876 20768
rect -11215 20723 -10991 20728
rect -11215 20564 -11170 20723
rect -11033 20613 -10901 20673
rect -11293 20507 -11129 20564
rect -11032 20553 -10974 20613
rect -11043 20385 -10969 20553
rect -11311 20343 -10919 20349
rect -11315 20309 -10827 20343
rect -11311 20303 -10919 20309
rect -11058 20153 -11012 20303
rect -11123 20147 -10919 20153
rect -11315 20113 -10827 20147
rect -11123 20107 -10919 20113
rect -11058 19957 -11012 20107
rect -11123 19951 -10919 19957
rect -11315 19917 -10827 19951
rect -11123 19911 -10919 19917
rect -11050 19856 -10980 19911
rect -11242 19783 -10980 19856
rect -11242 19782 -11074 19783
rect -11368 19732 -11289 19733
rect -11215 19732 -10859 19738
rect -10789 19732 -10697 19737
rect -11368 19698 -10697 19732
rect -11368 19697 -11289 19698
rect -11368 19537 -11334 19697
rect -11215 19691 -10859 19698
rect -10789 19693 -10697 19698
rect -11208 19634 -11122 19635
rect -11300 19600 -11122 19634
rect -11208 19599 -11122 19600
rect -11368 19536 -11279 19537
rect -11368 19502 -11192 19536
rect -11368 19495 -11279 19502
rect -11368 19343 -11334 19495
rect -11300 19437 -11192 19438
rect -11156 19437 -11122 19599
rect -11068 19566 -10994 19691
rect -10955 19634 -10880 19638
rect -10955 19600 -10777 19634
rect -10955 19597 -10880 19600
rect -11300 19404 -11122 19437
rect -11210 19401 -11122 19404
rect -11368 19340 -11278 19343
rect -11368 19306 -11192 19340
rect -11368 19301 -11278 19306
rect -11368 19147 -11334 19301
rect -11156 19243 -11122 19401
rect -11210 19242 -11122 19243
rect -11300 19208 -11122 19242
rect -11210 19207 -11122 19208
rect -11156 19182 -11122 19207
rect -10955 19440 -10921 19597
rect -10731 19541 -10697 19693
rect -10800 19536 -10697 19541
rect -10885 19502 -10697 19536
rect -10800 19497 -10697 19502
rect -10955 19438 -10872 19440
rect -10955 19404 -10777 19438
rect -10955 19399 -10872 19404
rect -10955 19246 -10921 19399
rect -10731 19345 -10697 19497
rect -10800 19340 -10697 19345
rect -10885 19306 -10697 19340
rect -10800 19301 -10697 19306
rect -10955 19242 -10872 19246
rect -10955 19208 -10777 19242
rect -10955 19205 -10872 19208
rect -10955 19182 -10921 19205
rect -11368 19144 -11283 19147
rect -11368 19110 -11192 19144
rect -11368 19105 -11283 19110
rect -11156 19049 -10921 19182
rect -10731 19148 -10697 19301
rect -10789 19144 -10697 19148
rect -10885 19110 -10697 19144
rect -10789 19104 -10697 19110
rect -11200 19046 -10871 19049
rect -11300 19012 -10777 19046
rect -11200 19008 -10871 19012
rect -11200 19007 -10914 19008
rect -11037 18810 -10984 19007
rect -10661 18923 -10622 23314
rect -10575 21642 -10536 24076
rect -10151 23145 -10091 23220
rect -10190 23144 -9904 23145
rect -10233 23140 -9904 23144
rect -10327 23106 -9804 23140
rect -10233 23103 -9904 23106
rect -10407 23042 -10315 23048
rect -10407 23008 -10219 23042
rect -10407 23004 -10315 23008
rect -10407 22851 -10373 23004
rect -10183 22970 -9948 23103
rect -9821 23042 -9736 23047
rect -9912 23008 -9736 23042
rect -9821 23005 -9736 23008
rect -10183 22947 -10149 22970
rect -10232 22944 -10149 22947
rect -10327 22910 -10149 22944
rect -10232 22906 -10149 22910
rect -10407 22846 -10304 22851
rect -10407 22812 -10219 22846
rect -10407 22807 -10304 22812
rect -10407 22655 -10373 22807
rect -10183 22753 -10149 22906
rect -10232 22748 -10149 22753
rect -10327 22714 -10149 22748
rect -10232 22712 -10149 22714
rect -10407 22650 -10304 22655
rect -10407 22616 -10219 22650
rect -10407 22611 -10304 22616
rect -10407 22459 -10373 22611
rect -10183 22555 -10149 22712
rect -9982 22945 -9948 22970
rect -9982 22944 -9894 22945
rect -9982 22910 -9804 22944
rect -9982 22909 -9894 22910
rect -9982 22751 -9948 22909
rect -9770 22851 -9736 23005
rect -9826 22846 -9736 22851
rect -9912 22812 -9736 22846
rect -9826 22809 -9736 22812
rect -9982 22748 -9894 22751
rect -9982 22715 -9804 22748
rect -10224 22552 -10149 22555
rect -10327 22518 -10149 22552
rect -10224 22514 -10149 22518
rect -10110 22461 -10036 22586
rect -9982 22553 -9948 22715
rect -9912 22714 -9804 22715
rect -9770 22657 -9736 22809
rect -9825 22650 -9736 22657
rect -9912 22616 -9736 22650
rect -9825 22615 -9736 22616
rect -9982 22552 -9896 22553
rect -9982 22518 -9804 22552
rect -9982 22517 -9896 22518
rect -10407 22454 -10315 22459
rect -10245 22454 -9889 22461
rect -9770 22455 -9736 22615
rect -9815 22454 -9736 22455
rect -10407 22420 -9736 22454
rect -10407 22415 -10315 22420
rect -10245 22414 -9889 22420
rect -9815 22419 -9736 22420
rect -10030 22369 -9862 22370
rect -10124 22296 -9862 22369
rect -10124 22241 -10054 22296
rect -10185 22235 -9981 22241
rect -10277 22201 -9789 22235
rect -10185 22195 -9981 22201
rect -5750 25045 -5695 25200
rect -5800 24993 -5690 24999
rect -6092 24959 -5690 24993
rect -5800 24954 -5690 24959
rect -5730 24688 -5690 24954
rect -5633 24930 -5597 25315
rect -5551 25091 -5456 25095
rect -5551 25057 -4872 25091
rect -5551 25053 -5456 25057
rect -5642 24775 -5587 24930
rect -5551 24883 -5515 25053
rect -5551 24880 -5462 24883
rect -4880 24880 -4804 24884
rect -5551 24846 -4804 24880
rect -5551 24841 -5462 24846
rect -4880 24842 -4804 24846
rect -5553 24782 -5460 24786
rect -5553 24748 -4872 24782
rect -5553 24744 -5460 24748
rect -5553 24688 -5514 24744
rect -5730 24645 -5514 24688
rect -4838 24686 -4804 24842
rect -4882 24684 -4804 24686
rect -5480 24650 -4804 24684
rect -5750 24559 -5710 24607
rect -5793 24555 -5710 24559
rect -6092 24521 -5710 24555
rect -5793 24515 -5710 24521
rect -5753 24473 -5710 24515
rect -5620 24507 -5565 24645
rect -4882 24644 -4804 24650
rect -5753 24472 -5466 24473
rect -7347 24180 -7225 24356
rect -5753 24438 -4872 24472
rect -5753 24430 -5466 24438
rect -10092 22045 -10046 22195
rect -10185 22039 -9981 22045
rect -10277 22005 -9789 22039
rect -10185 21999 -9981 22005
rect -10586 21510 -10526 21642
rect -10575 20701 -10536 21510
rect -10092 21849 -10046 21999
rect -10185 21843 -9793 21849
rect -10277 21809 -9789 21843
rect -10185 21803 -9793 21809
rect -10135 21599 -10061 21767
rect -10294 21539 -10072 21599
rect -9975 21588 -9811 21645
rect -9925 21502 -9863 21588
rect -10124 21440 -9863 21502
rect -10124 21404 -10054 21440
rect -10185 21398 -9981 21404
rect -10277 21364 -9789 21398
rect -10185 21358 -9981 21364
rect -10092 21208 -10046 21358
rect -7443 21669 -7371 21693
rect -8850 21599 -7371 21669
rect -10185 21202 -9981 21208
rect -10277 21168 -9789 21202
rect -10185 21162 -9981 21168
rect -10585 20564 -10525 20701
rect -11043 18642 -10969 18810
rect -10674 18791 -10614 18923
rect -11311 18600 -10919 18606
rect -11315 18566 -10827 18600
rect -11311 18560 -10919 18566
rect -11058 18410 -11012 18560
rect -11123 18404 -10919 18410
rect -11315 18370 -10827 18404
rect -11123 18364 -10919 18370
rect -11058 18214 -11012 18364
rect -10661 18385 -10622 18791
rect -10575 18385 -10536 20564
rect -10092 21012 -10046 21162
rect -8850 21331 -8780 21599
rect -7443 21588 -7371 21599
rect -7268 21405 -7225 24180
rect -6116 24115 -6042 24135
rect -5753 24115 -5710 24430
rect -6116 24076 -5609 24115
rect -6116 23967 -6042 24076
rect -5753 24072 -5710 24076
rect -6384 23925 -5992 23931
rect -6388 23891 -5900 23925
rect -6384 23885 -5992 23891
rect -6131 23735 -6085 23885
rect -6196 23729 -5992 23735
rect -6388 23695 -5900 23729
rect -6196 23689 -5992 23695
rect -6131 23539 -6085 23689
rect -6196 23533 -5992 23539
rect -6388 23499 -5900 23533
rect -6196 23493 -5992 23499
rect -6123 23463 -6053 23493
rect -6101 23405 -6059 23463
rect -6105 23345 -5973 23405
rect -6101 23288 -6059 23345
rect -6366 23207 -6202 23264
rect -6105 23253 -6047 23288
rect -6116 23085 -6042 23253
rect -5745 23314 -5685 23446
rect -6384 23043 -5992 23049
rect -6388 23009 -5900 23043
rect -6384 23003 -5992 23009
rect -6131 22853 -6085 23003
rect -6196 22847 -5992 22853
rect -6388 22813 -5900 22847
rect -6196 22807 -5992 22813
rect -6131 22657 -6085 22807
rect -6196 22651 -5992 22657
rect -6388 22617 -5900 22651
rect -6196 22611 -5992 22617
rect -6123 22556 -6053 22611
rect -6315 22483 -6053 22556
rect -6315 22482 -6147 22483
rect -6441 22432 -6362 22433
rect -6288 22432 -5932 22438
rect -5862 22432 -5770 22437
rect -6441 22398 -5770 22432
rect -6441 22397 -6362 22398
rect -6441 22237 -6407 22397
rect -6288 22391 -5932 22398
rect -5862 22393 -5770 22398
rect -6281 22334 -6195 22335
rect -6373 22300 -6195 22334
rect -6281 22299 -6195 22300
rect -6441 22236 -6352 22237
rect -6441 22202 -6265 22236
rect -6441 22195 -6352 22202
rect -6441 22043 -6407 22195
rect -6373 22137 -6265 22138
rect -6229 22137 -6195 22299
rect -6141 22266 -6067 22391
rect -6028 22334 -5953 22338
rect -6028 22300 -5850 22334
rect -6028 22297 -5953 22300
rect -6373 22104 -6195 22137
rect -6283 22101 -6195 22104
rect -6441 22040 -6351 22043
rect -6441 22006 -6265 22040
rect -6441 22001 -6351 22006
rect -6441 21847 -6407 22001
rect -6229 21943 -6195 22101
rect -6283 21942 -6195 21943
rect -6373 21908 -6195 21942
rect -6283 21907 -6195 21908
rect -6229 21882 -6195 21907
rect -6028 22140 -5994 22297
rect -5804 22241 -5770 22393
rect -5873 22236 -5770 22241
rect -5958 22202 -5770 22236
rect -5873 22197 -5770 22202
rect -6028 22138 -5945 22140
rect -6028 22104 -5850 22138
rect -6028 22099 -5945 22104
rect -6028 21946 -5994 22099
rect -5804 22045 -5770 22197
rect -5873 22040 -5770 22045
rect -5958 22006 -5770 22040
rect -5873 22001 -5770 22006
rect -6028 21942 -5945 21946
rect -6028 21908 -5850 21942
rect -6028 21905 -5945 21908
rect -6028 21882 -5994 21905
rect -6441 21844 -6356 21847
rect -6441 21810 -6265 21844
rect -6441 21805 -6356 21810
rect -6229 21749 -5994 21882
rect -5804 21848 -5770 22001
rect -5862 21844 -5770 21848
rect -5958 21810 -5770 21844
rect -5862 21804 -5770 21810
rect -5954 21749 -5822 21755
rect -6273 21746 -5822 21749
rect -8850 21297 -8608 21331
rect -7512 21397 -7225 21405
rect -8106 21363 -7225 21397
rect -7512 21362 -7225 21363
rect -8947 21199 -8839 21233
rect -8716 21101 -8608 21135
rect -10185 21006 -9793 21012
rect -10277 20972 -9789 21006
rect -10185 20966 -9793 20972
rect -10135 20762 -10061 20930
rect -10128 20740 -10068 20762
rect -10149 20445 -10089 20536
rect -10190 20444 -9904 20445
rect -10233 20440 -9904 20444
rect -10327 20406 -9804 20440
rect -10233 20403 -9904 20406
rect -10407 20342 -10315 20348
rect -10407 20308 -10219 20342
rect -10407 20304 -10315 20308
rect -10407 20151 -10373 20304
rect -10183 20270 -9948 20403
rect -8947 21003 -8839 21037
rect -8716 20905 -8608 20939
rect -8810 20787 -8750 20860
rect -8804 20726 -8763 20787
rect -8983 20715 -8763 20726
rect -9821 20342 -9736 20347
rect -9912 20308 -9736 20342
rect -9821 20305 -9736 20308
rect -10183 20247 -10149 20270
rect -10232 20244 -10149 20247
rect -10327 20210 -10149 20244
rect -10232 20206 -10149 20210
rect -10407 20146 -10304 20151
rect -10407 20112 -10219 20146
rect -10407 20107 -10304 20112
rect -10407 19955 -10373 20107
rect -10183 20053 -10149 20206
rect -10232 20048 -10149 20053
rect -10327 20014 -10149 20048
rect -10232 20012 -10149 20014
rect -10407 19950 -10304 19955
rect -10407 19916 -10219 19950
rect -10407 19911 -10304 19916
rect -10407 19759 -10373 19911
rect -10183 19855 -10149 20012
rect -9982 20245 -9948 20270
rect -9982 20244 -9894 20245
rect -9982 20210 -9804 20244
rect -9982 20209 -9894 20210
rect -9982 20051 -9948 20209
rect -9770 20151 -9736 20305
rect -9826 20146 -9736 20151
rect -9912 20112 -9736 20146
rect -9826 20109 -9736 20112
rect -9982 20048 -9894 20051
rect -9982 20015 -9804 20048
rect -10224 19852 -10149 19855
rect -10327 19818 -10149 19852
rect -10224 19814 -10149 19818
rect -10110 19761 -10036 19886
rect -9982 19853 -9948 20015
rect -9912 20014 -9804 20015
rect -9770 19957 -9736 20109
rect -9825 19950 -9736 19957
rect -9912 19916 -9736 19950
rect -9825 19915 -9736 19916
rect -9982 19852 -9896 19853
rect -9982 19818 -9804 19852
rect -9982 19817 -9896 19818
rect -10407 19754 -10315 19759
rect -10245 19754 -9889 19761
rect -9770 19755 -9736 19915
rect -9815 19754 -9736 19755
rect -10407 19720 -9736 19754
rect -10407 19715 -10315 19720
rect -10245 19714 -9889 19720
rect -9815 19719 -9736 19720
rect -10030 19669 -9862 19670
rect -10124 19596 -9862 19669
rect -10124 19541 -10054 19596
rect -10185 19535 -9981 19541
rect -10277 19501 -9789 19535
rect -10185 19495 -9981 19501
rect -8991 20687 -8763 20715
rect -8991 20665 -8791 20687
rect -9454 20590 -9146 20624
rect -9109 20578 -9038 20652
rect -9454 20492 -9146 20526
rect -9454 20394 -9146 20428
rect -9103 20237 -9064 20578
rect -8991 20526 -8953 20665
rect -8174 21185 -8096 21191
rect -7413 21190 -7358 21328
rect -7268 21320 -7225 21362
rect -7268 21314 -7185 21320
rect -7268 21280 -6886 21314
rect -7268 21276 -7185 21280
rect -7268 21228 -7228 21276
rect -6373 21712 -5822 21746
rect -6273 21709 -5822 21712
rect -6273 21708 -5944 21709
rect -6273 21707 -5987 21708
rect -6107 21510 -6050 21707
rect -6116 21342 -6042 21510
rect -6384 21300 -5992 21306
rect -6388 21266 -5900 21300
rect -6384 21260 -5992 21266
rect -8174 21151 -7498 21185
rect -8174 21149 -8096 21151
rect -8174 20993 -8140 21149
rect -7464 21147 -7248 21190
rect -7464 21091 -7425 21147
rect -7518 21087 -7425 21091
rect -8106 21053 -7425 21087
rect -7518 21049 -7425 21053
rect -8174 20989 -8098 20993
rect -7516 20989 -7427 20994
rect -8174 20955 -7427 20989
rect -8174 20951 -8098 20955
rect -7516 20952 -7427 20955
rect -7463 20782 -7427 20952
rect -7391 20905 -7336 21060
rect -7522 20778 -7427 20782
rect -8106 20744 -7427 20778
rect -7522 20740 -7427 20744
rect -8991 20492 -8609 20526
rect -8991 20330 -8953 20492
rect -7846 20570 -7776 20576
rect -7381 20570 -7345 20905
rect -7288 20881 -7248 21147
rect -7288 20876 -7178 20881
rect -7288 20842 -6886 20876
rect -7288 20836 -7178 20842
rect -7283 20635 -7228 20790
rect -7274 20598 -7240 20635
rect -7846 20500 -7343 20570
rect -8991 20296 -8609 20330
rect -9454 20198 -9146 20232
rect -9104 20167 -9064 20237
rect -9104 20166 -9062 20167
rect -10092 19345 -10046 19495
rect -10185 19339 -9981 19345
rect -10277 19305 -9789 19339
rect -10185 19299 -9981 19305
rect -10092 19149 -10046 19299
rect -10185 19143 -9793 19149
rect -10277 19109 -9789 19143
rect -10185 19103 -9793 19109
rect -10135 18899 -10061 19067
rect -9102 19651 -9062 20166
rect -9014 20113 -8960 20248
rect -9006 20093 -8966 20113
rect -9004 19886 -8968 20093
rect -8946 19715 -8738 19749
rect -9276 19618 -9062 19651
rect -9276 19617 -9068 19618
rect -8946 19519 -8738 19553
rect -7846 20332 -7776 20500
rect -8018 20298 -7776 20332
rect -7787 20200 -7679 20234
rect -8018 20102 -7910 20136
rect -7787 20004 -7679 20038
rect -6131 21110 -6085 21260
rect -6196 21104 -5992 21110
rect -6388 21070 -5900 21104
rect -6196 21064 -5992 21070
rect -6131 20914 -6085 21064
rect -6196 20908 -5992 20914
rect -6388 20874 -5900 20908
rect -6196 20868 -5992 20874
rect -6123 20838 -6053 20868
rect -6109 20788 -6064 20838
rect -6109 20768 -5949 20788
rect -6288 20728 -5949 20768
rect -6288 20723 -6064 20728
rect -6288 20564 -6243 20723
rect -6106 20613 -5974 20673
rect -6366 20507 -6202 20564
rect -6105 20553 -6047 20613
rect -6116 20385 -6042 20553
rect -6384 20343 -5992 20349
rect -6388 20309 -5900 20343
rect -6384 20303 -5992 20309
rect -6131 20153 -6085 20303
rect -6196 20147 -5992 20153
rect -6388 20113 -5900 20147
rect -6196 20107 -5992 20113
rect -8018 19906 -7910 19940
rect -7876 19788 -7816 19861
rect -7863 19727 -7822 19788
rect -7863 19716 -7643 19727
rect -7863 19688 -7635 19716
rect -7835 19666 -7635 19688
rect -9276 19421 -9068 19455
rect -8946 19323 -8738 19357
rect -10135 18887 -10072 18899
rect -9975 18888 -9811 18945
rect -10279 18864 -10072 18887
rect -10279 18827 -10073 18864
rect -9924 18791 -9875 18888
rect -10124 18745 -9875 18791
rect -10124 18704 -10054 18745
rect -10185 18698 -9981 18704
rect -10277 18664 -9789 18698
rect -10185 18658 -9981 18664
rect -10092 18508 -10046 18658
rect -7673 19527 -7635 19666
rect -6131 19957 -6085 20107
rect -7480 19591 -7172 19625
rect -8017 19493 -7635 19527
rect -7673 19331 -7635 19493
rect -8017 19297 -7635 19331
rect -7666 19114 -7612 19249
rect -7480 19493 -7172 19527
rect -7480 19395 -7172 19429
rect -7480 19199 -7172 19233
rect -7660 19094 -7620 19114
rect -7658 18840 -7622 19094
rect -6196 19951 -5992 19957
rect -6388 19917 -5900 19951
rect -6196 19911 -5992 19917
rect -6123 19856 -6053 19911
rect -6315 19783 -6053 19856
rect -6315 19782 -6147 19783
rect -6441 19732 -6362 19733
rect -6288 19732 -5932 19738
rect -5862 19732 -5770 19737
rect -6441 19698 -5770 19732
rect -6441 19697 -6362 19698
rect -6441 19537 -6407 19697
rect -6288 19691 -5932 19698
rect -5862 19693 -5770 19698
rect -6281 19634 -6195 19635
rect -6373 19600 -6195 19634
rect -6281 19599 -6195 19600
rect -6441 19536 -6352 19537
rect -6441 19502 -6265 19536
rect -6441 19495 -6352 19502
rect -6441 19343 -6407 19495
rect -6373 19437 -6265 19438
rect -6229 19437 -6195 19599
rect -6141 19566 -6067 19691
rect -6028 19634 -5953 19638
rect -6028 19600 -5850 19634
rect -6028 19597 -5953 19600
rect -6373 19404 -6195 19437
rect -6283 19401 -6195 19404
rect -6441 19340 -6351 19343
rect -6441 19306 -6265 19340
rect -6441 19301 -6351 19306
rect -6441 19147 -6407 19301
rect -6229 19243 -6195 19401
rect -6283 19242 -6195 19243
rect -6373 19208 -6195 19242
rect -6283 19207 -6195 19208
rect -6229 19182 -6195 19207
rect -6028 19440 -5994 19597
rect -5804 19541 -5770 19693
rect -5873 19536 -5770 19541
rect -5958 19502 -5770 19536
rect -5873 19497 -5770 19502
rect -6028 19438 -5945 19440
rect -6028 19404 -5850 19438
rect -6028 19399 -5945 19404
rect -6028 19246 -5994 19399
rect -5804 19345 -5770 19497
rect -5873 19340 -5770 19345
rect -5958 19306 -5770 19340
rect -5873 19301 -5770 19306
rect -6028 19242 -5945 19246
rect -6028 19208 -5850 19242
rect -6028 19205 -5945 19208
rect -6028 19182 -5994 19205
rect -6441 19144 -6356 19147
rect -6441 19110 -6265 19144
rect -6441 19105 -6356 19110
rect -6229 19049 -5994 19182
rect -5804 19148 -5770 19301
rect -5862 19144 -5770 19148
rect -5958 19110 -5770 19144
rect -5862 19104 -5770 19110
rect -6273 19046 -5944 19049
rect -7719 18654 -7565 18840
rect -6373 19012 -5850 19046
rect -6273 19008 -5944 19012
rect -6273 19007 -5987 19008
rect -6110 18810 -6057 19007
rect -5734 18923 -5695 23314
rect -5648 21642 -5609 24076
rect -5224 23145 -5164 23220
rect -5263 23144 -4977 23145
rect -5306 23140 -4977 23144
rect -5400 23106 -4877 23140
rect -5306 23103 -4977 23106
rect -5480 23042 -5388 23048
rect -5480 23008 -5292 23042
rect -5480 23004 -5388 23008
rect -5480 22851 -5446 23004
rect -5256 22970 -5021 23103
rect -4894 23042 -4809 23047
rect -4985 23008 -4809 23042
rect -4894 23005 -4809 23008
rect -5256 22947 -5222 22970
rect -5305 22944 -5222 22947
rect -5400 22910 -5222 22944
rect -5305 22906 -5222 22910
rect -5480 22846 -5377 22851
rect -5480 22812 -5292 22846
rect -5480 22807 -5377 22812
rect -5480 22655 -5446 22807
rect -5256 22753 -5222 22906
rect -5305 22748 -5222 22753
rect -5400 22714 -5222 22748
rect -5305 22712 -5222 22714
rect -5480 22650 -5377 22655
rect -5480 22616 -5292 22650
rect -5480 22611 -5377 22616
rect -5480 22459 -5446 22611
rect -5256 22555 -5222 22712
rect -5055 22945 -5021 22970
rect -5055 22944 -4967 22945
rect -5055 22910 -4877 22944
rect -5055 22909 -4967 22910
rect -5055 22751 -5021 22909
rect -4843 22851 -4809 23005
rect -4899 22846 -4809 22851
rect -4985 22812 -4809 22846
rect -4899 22809 -4809 22812
rect -5055 22748 -4967 22751
rect -5055 22715 -4877 22748
rect -5297 22552 -5222 22555
rect -5400 22518 -5222 22552
rect -5297 22514 -5222 22518
rect -5183 22461 -5109 22586
rect -5055 22553 -5021 22715
rect -4985 22714 -4877 22715
rect -4843 22657 -4809 22809
rect -4898 22650 -4809 22657
rect -4985 22616 -4809 22650
rect -4898 22615 -4809 22616
rect -5055 22552 -4969 22553
rect -5055 22518 -4877 22552
rect -5055 22517 -4969 22518
rect -5480 22454 -5388 22459
rect -5318 22454 -4962 22461
rect -4843 22455 -4809 22615
rect -4888 22454 -4809 22455
rect -5480 22420 -4809 22454
rect -5480 22415 -5388 22420
rect -5318 22414 -4962 22420
rect -4888 22419 -4809 22420
rect -5103 22369 -4935 22370
rect -5197 22296 -4935 22369
rect -5197 22241 -5127 22296
rect -5258 22235 -5054 22241
rect -5350 22201 -4862 22235
rect -5258 22195 -5054 22201
rect -5165 22045 -5119 22195
rect -5258 22039 -5054 22045
rect -5350 22005 -4862 22039
rect -5258 21999 -5054 22005
rect -5659 21510 -5599 21642
rect -5648 20701 -5609 21510
rect -5165 21849 -5119 21999
rect -5258 21843 -4866 21849
rect -5350 21809 -4862 21843
rect -5258 21803 -4866 21809
rect -5208 21599 -5134 21767
rect -5367 21539 -5145 21599
rect -5048 21588 -4884 21645
rect -4998 21502 -4936 21588
rect -5197 21440 -4936 21502
rect -5197 21404 -5127 21440
rect -5258 21398 -5054 21404
rect -5350 21364 -4862 21398
rect -5258 21358 -5054 21364
rect -5165 21208 -5119 21358
rect -5258 21202 -5054 21208
rect -5350 21168 -4862 21202
rect -5258 21162 -5054 21168
rect -5658 20564 -5598 20701
rect -6116 18642 -6042 18810
rect -5747 18791 -5687 18923
rect -6384 18600 -5992 18606
rect -6388 18566 -5900 18600
rect -6384 18560 -5992 18566
rect -10185 18502 -9981 18508
rect -10277 18468 -9789 18502
rect -10185 18462 -9981 18468
rect -11123 18208 -10919 18214
rect -11315 18174 -10827 18208
rect -11123 18168 -10919 18174
rect -10092 18312 -10046 18462
rect -6131 18410 -6085 18560
rect -6196 18404 -5992 18410
rect -10185 18306 -9793 18312
rect -10277 18272 -9789 18306
rect -10185 18266 -9793 18272
rect -11050 18138 -10980 18168
rect -11041 18103 -11002 18138
rect -10644 18103 -10507 18114
rect -10135 18103 -10061 18230
rect -11041 18062 -10061 18103
rect -11041 18056 -10091 18062
rect -11039 18055 -10091 18056
rect -10644 18054 -10507 18055
rect -6388 18370 -5900 18404
rect -6196 18364 -5992 18370
rect -6131 18214 -6085 18364
rect -5734 18385 -5695 18791
rect -5648 18385 -5609 20564
rect -5165 21012 -5119 21162
rect -5258 21006 -4866 21012
rect -5350 20972 -4862 21006
rect -5258 20966 -4866 20972
rect -5208 20762 -5134 20930
rect -5201 20740 -5141 20762
rect -5222 20445 -5162 20536
rect -5263 20444 -4977 20445
rect -5306 20440 -4977 20444
rect -5400 20406 -4877 20440
rect -5306 20403 -4977 20406
rect -5480 20342 -5388 20348
rect -5480 20308 -5292 20342
rect -5480 20304 -5388 20308
rect -5480 20151 -5446 20304
rect -5256 20270 -5021 20403
rect -4894 20342 -4809 20347
rect -4985 20308 -4809 20342
rect -4894 20305 -4809 20308
rect -5256 20247 -5222 20270
rect -5305 20244 -5222 20247
rect -5400 20210 -5222 20244
rect -5305 20206 -5222 20210
rect -5480 20146 -5377 20151
rect -5480 20112 -5292 20146
rect -5480 20107 -5377 20112
rect -5480 19955 -5446 20107
rect -5256 20053 -5222 20206
rect -5305 20048 -5222 20053
rect -5400 20014 -5222 20048
rect -5305 20012 -5222 20014
rect -5480 19950 -5377 19955
rect -5480 19916 -5292 19950
rect -5480 19911 -5377 19916
rect -5480 19759 -5446 19911
rect -5256 19855 -5222 20012
rect -5055 20245 -5021 20270
rect -5055 20244 -4967 20245
rect -5055 20210 -4877 20244
rect -5055 20209 -4967 20210
rect -5055 20051 -5021 20209
rect -4843 20151 -4809 20305
rect -4899 20146 -4809 20151
rect -4985 20112 -4809 20146
rect -4899 20109 -4809 20112
rect -5055 20048 -4967 20051
rect -5055 20015 -4877 20048
rect -5297 19852 -5222 19855
rect -5400 19818 -5222 19852
rect -5297 19814 -5222 19818
rect -5183 19761 -5109 19886
rect -5055 19853 -5021 20015
rect -4985 20014 -4877 20015
rect -4843 19957 -4809 20109
rect -4898 19950 -4809 19957
rect -4985 19916 -4809 19950
rect -4898 19915 -4809 19916
rect -5055 19852 -4969 19853
rect -5055 19818 -4877 19852
rect -5055 19817 -4969 19818
rect -5480 19754 -5388 19759
rect -5318 19754 -4962 19761
rect -4843 19755 -4809 19915
rect -4888 19754 -4809 19755
rect -5480 19720 -4809 19754
rect -5480 19715 -5388 19720
rect -5318 19714 -4962 19720
rect -4888 19719 -4809 19720
rect -5103 19669 -4935 19670
rect -5197 19596 -4935 19669
rect -5197 19541 -5127 19596
rect -5258 19535 -5054 19541
rect -5350 19501 -4862 19535
rect -5258 19495 -5054 19501
rect -5165 19345 -5119 19495
rect -5258 19339 -5054 19345
rect -5350 19305 -4862 19339
rect -5258 19299 -5054 19305
rect -5165 19149 -5119 19299
rect -5258 19143 -4866 19149
rect -5350 19109 -4862 19143
rect -5258 19103 -4866 19109
rect -5208 18899 -5134 19067
rect -5208 18887 -5145 18899
rect -5048 18888 -4884 18945
rect -5352 18864 -5145 18887
rect -5352 18827 -5146 18864
rect -4997 18791 -4948 18888
rect -5197 18745 -4948 18791
rect -5197 18704 -5127 18745
rect -5258 18698 -5054 18704
rect -5350 18664 -4862 18698
rect -5258 18658 -5054 18664
rect -5165 18508 -5119 18658
rect -5258 18502 -5054 18508
rect -5350 18468 -4862 18502
rect -5258 18462 -5054 18468
rect -6196 18208 -5992 18214
rect -6388 18174 -5900 18208
rect -6196 18168 -5992 18174
rect -5165 18312 -5119 18462
rect -5258 18306 -4866 18312
rect -5350 18272 -4862 18306
rect -5258 18266 -4866 18272
rect -6123 18138 -6053 18168
rect -6114 18103 -6075 18138
rect -5717 18103 -5580 18114
rect -5208 18103 -5134 18230
rect -6114 18062 -5134 18103
rect -6114 18056 -5164 18062
rect -6112 18055 -5164 18056
rect -5717 18054 -5580 18055
rect -11345 17179 -11179 17316
rect -11467 16680 -11395 16704
rect -12874 16610 -11395 16680
rect -12874 16342 -12804 16610
rect -11467 16599 -11395 16610
rect -11292 16416 -11249 17179
rect -12874 16308 -12632 16342
rect -11536 16408 -11249 16416
rect -12130 16374 -11249 16408
rect -11536 16373 -11249 16374
rect -12971 16210 -12863 16244
rect -12740 16112 -12632 16146
rect -12971 16014 -12863 16048
rect -12740 15916 -12632 15950
rect -12834 15798 -12774 15871
rect -12828 15737 -12787 15798
rect -13007 15726 -12787 15737
rect -13015 15698 -12787 15726
rect -13015 15676 -12815 15698
rect -13478 15601 -13170 15635
rect -13133 15589 -13062 15663
rect -13478 15503 -13170 15537
rect -13478 15405 -13170 15439
rect -13127 15248 -13088 15589
rect -13015 15537 -12977 15676
rect -12198 16196 -12120 16202
rect -11437 16201 -11382 16339
rect -11292 16331 -11249 16373
rect -11292 16325 -11209 16331
rect -11292 16291 -10910 16325
rect -11292 16287 -11209 16291
rect -11292 16239 -11252 16287
rect -12198 16162 -11522 16196
rect -12198 16160 -12120 16162
rect -12198 16004 -12164 16160
rect -11488 16158 -11272 16201
rect -11488 16102 -11449 16158
rect -11542 16098 -11449 16102
rect -12130 16064 -11449 16098
rect -11542 16060 -11449 16064
rect -12198 16000 -12122 16004
rect -11540 16000 -11451 16005
rect -12198 15966 -11451 16000
rect -12198 15962 -12122 15966
rect -11540 15963 -11451 15966
rect -11487 15793 -11451 15963
rect -11415 15916 -11360 16071
rect -11546 15789 -11451 15793
rect -12130 15755 -11451 15789
rect -11546 15751 -11451 15755
rect -13015 15503 -12633 15537
rect -13015 15341 -12977 15503
rect -11870 15581 -11800 15587
rect -11405 15581 -11369 15916
rect -11312 15892 -11272 16158
rect -11312 15887 -11202 15892
rect -11312 15853 -10910 15887
rect -11312 15847 -11202 15853
rect -11307 15646 -11252 15801
rect -11298 15609 -11264 15646
rect -11870 15511 -11367 15581
rect -13015 15307 -12633 15341
rect -13478 15209 -13170 15243
rect -13128 15178 -13088 15248
rect -13128 15177 -13086 15178
rect -13126 14662 -13086 15177
rect -13038 15124 -12984 15259
rect -13030 15104 -12990 15124
rect -13028 14897 -12992 15104
rect -12970 14726 -12762 14760
rect -13300 14629 -13086 14662
rect -13300 14628 -13092 14629
rect -12970 14530 -12762 14564
rect -11870 15343 -11800 15511
rect -12042 15309 -11800 15343
rect -11811 15211 -11703 15245
rect -12042 15113 -11934 15147
rect -11811 15015 -11703 15049
rect -12042 14917 -11934 14951
rect -11900 14799 -11840 14872
rect -11887 14738 -11846 14799
rect -11887 14727 -11667 14738
rect -11887 14699 -11659 14727
rect -11859 14677 -11659 14699
rect -13300 14432 -13092 14466
rect -12970 14334 -12762 14368
rect -13064 14216 -13004 14289
rect -13058 14172 -13017 14216
rect -13150 14042 -13000 14172
rect -14155 13609 -14018 13747
rect -14253 13471 -14195 13608
rect -13091 13565 -13023 14042
rect -13159 13507 -13022 13565
rect -14252 10561 -14200 13471
rect -13648 13422 -13511 13480
rect -13643 11816 -13608 13422
rect -11697 14538 -11659 14677
rect -11612 14590 -11541 14664
rect -11504 14602 -11196 14636
rect -12041 14504 -11659 14538
rect -11697 14342 -11659 14504
rect -12041 14308 -11659 14342
rect -11690 14125 -11636 14260
rect -11586 14249 -11547 14590
rect -11504 14504 -11196 14538
rect -11504 14406 -11196 14440
rect -11586 14179 -11546 14249
rect -11504 14210 -11196 14244
rect -11588 14178 -11546 14179
rect -11684 14105 -11644 14125
rect -11682 13723 -11646 14105
rect -11588 13952 -11548 14178
rect -11754 13606 -11631 13723
rect -11456 13360 -11398 13482
rect -11456 13347 -11166 13360
rect -10832 13347 -10730 13354
rect -11456 13313 -10730 13347
rect -11456 13310 -11166 13313
rect -11456 13254 -11411 13310
rect -10832 13308 -10730 13313
rect -11456 13044 -11420 13254
rect -11282 13249 -11202 13253
rect -11282 13215 -10804 13249
rect -11282 13208 -11202 13215
rect -11505 13038 -11420 13044
rect -11704 13004 -11420 13038
rect -11505 12999 -11420 13004
rect -13645 11797 -13608 11816
rect -13562 12497 -13425 12555
rect -13653 11662 -13599 11797
rect -13900 11588 -13619 11622
rect -13656 11426 -13619 11588
rect -13562 11461 -13524 12497
rect -13480 11767 -13343 11825
rect -13900 11392 -13619 11426
rect -13656 11230 -13619 11392
rect -13571 11326 -13517 11461
rect -13480 11273 -13446 11767
rect -13390 11686 -12985 11720
rect -13390 11524 -13356 11686
rect -13390 11490 -12985 11524
rect -13390 11312 -13355 11490
rect -13292 11376 -12852 11410
rect -12993 11375 -12852 11376
rect -13390 11278 -12984 11312
rect -13390 11277 -13292 11278
rect -13900 11196 -13619 11230
rect -13656 11104 -13619 11196
rect -13493 11138 -13439 11273
rect -12889 11214 -12852 11375
rect -13292 11180 -12852 11214
rect -12995 11179 -12852 11180
rect -13656 11101 -13356 11104
rect -13656 11067 -12984 11101
rect -13481 10662 -13444 11067
rect -13390 10905 -13356 11067
rect -12886 11003 -12852 11179
rect -13292 10969 -12852 11003
rect -13390 10871 -12984 10905
rect -14283 10403 -14167 10561
rect -13491 10527 -13437 10662
rect -13900 10458 -12984 10492
rect -11282 12941 -11246 13208
rect -10768 13156 -10730 13308
rect -10832 13151 -10730 13156
rect -11212 13117 -10730 13151
rect -10832 13110 -10730 13117
rect -9210 17158 -9002 17366
rect -9686 16219 -9421 16487
rect -11282 12940 -11207 12941
rect -11282 12906 -10804 12940
rect -11282 12905 -11207 12906
rect -11455 12455 -11397 12551
rect -11455 12442 -11165 12455
rect -10831 12442 -10729 12449
rect -11455 12408 -10729 12442
rect -11455 12405 -11165 12408
rect -11455 12349 -11410 12405
rect -10831 12403 -10729 12408
rect -11455 12139 -11419 12349
rect -11281 12344 -11201 12348
rect -11281 12310 -10803 12344
rect -11281 12303 -11201 12310
rect -11504 12133 -11419 12139
rect -11703 12099 -11419 12133
rect -11504 12094 -11419 12099
rect -11281 12036 -11245 12303
rect -10767 12251 -10729 12403
rect -10831 12246 -10729 12251
rect -11211 12212 -10729 12246
rect -10831 12205 -10729 12212
rect -11281 12035 -11206 12036
rect -11281 12001 -10803 12035
rect -11281 12000 -11206 12001
rect -11804 11578 -11746 11664
rect -11804 11536 -11520 11578
rect -10880 11546 -10804 11558
rect -11804 11527 -11746 11536
rect -11804 11127 -11762 11527
rect -11562 11452 -11520 11536
rect -11482 11512 -10804 11546
rect -10880 11502 -10804 11512
rect -11562 11448 -11464 11452
rect -11562 11414 -10874 11448
rect -11562 11410 -11464 11414
rect -10838 11360 -10804 11502
rect -10880 11350 -10804 11360
rect -11482 11316 -10804 11350
rect -10880 11304 -10804 11316
rect -11855 11123 -11762 11127
rect -12046 11089 -11762 11123
rect -11855 11085 -11762 11089
rect -11804 10931 -11762 11085
rect -11855 10927 -11762 10931
rect -12046 10893 -11762 10927
rect -11855 10889 -11762 10893
rect -11553 11237 -11471 11240
rect -11553 11203 -10874 11237
rect -11553 11198 -11471 11203
rect -11553 11044 -11516 11198
rect -10838 11148 -10804 11304
rect -10880 11139 -10804 11148
rect -11482 11105 -10804 11139
rect -10880 11095 -10804 11105
rect -11553 11041 -11472 11044
rect -11553 11007 -10874 11041
rect -11553 11002 -11472 11007
rect -11553 10832 -11516 11002
rect -11553 10829 -11465 10832
rect -11553 10795 -10874 10829
rect -11553 10791 -11465 10795
rect -9654 7738 -9468 16219
rect -9208 13828 -9002 17158
rect -8834 17244 -6249 17427
rect -8834 16482 -8651 17244
rect -6467 16680 -6395 16704
rect -7874 16610 -6395 16680
rect -8866 16214 -8601 16482
rect -7874 16342 -7804 16610
rect -6467 16599 -6395 16610
rect -6292 16416 -6249 17244
rect -7874 16308 -7632 16342
rect -6536 16408 -6249 16416
rect -7130 16374 -6249 16408
rect -6536 16373 -6249 16374
rect -7971 16210 -7863 16244
rect -7740 16112 -7632 16146
rect -7971 16014 -7863 16048
rect -7740 15916 -7632 15950
rect -7834 15798 -7774 15871
rect -7828 15737 -7787 15798
rect -8007 15726 -7787 15737
rect -8015 15698 -7787 15726
rect -8015 15676 -7815 15698
rect -8478 15601 -8170 15635
rect -8133 15589 -8062 15663
rect -8478 15503 -8170 15537
rect -8478 15405 -8170 15439
rect -8127 15248 -8088 15589
rect -8015 15537 -7977 15676
rect -7198 16196 -7120 16202
rect -6437 16201 -6382 16339
rect -6292 16331 -6249 16373
rect -6292 16325 -6209 16331
rect -6292 16291 -5910 16325
rect -6292 16287 -6209 16291
rect -6292 16239 -6252 16287
rect -7198 16162 -6522 16196
rect -7198 16160 -7120 16162
rect -7198 16004 -7164 16160
rect -6488 16158 -6272 16201
rect -6488 16102 -6449 16158
rect -6542 16098 -6449 16102
rect -7130 16064 -6449 16098
rect -6542 16060 -6449 16064
rect -7198 16000 -7122 16004
rect -6540 16000 -6451 16005
rect -7198 15966 -6451 16000
rect -7198 15962 -7122 15966
rect -6540 15963 -6451 15966
rect -6487 15793 -6451 15963
rect -6415 15916 -6360 16071
rect -6546 15789 -6451 15793
rect -7130 15755 -6451 15789
rect -6546 15751 -6451 15755
rect -8015 15503 -7633 15537
rect -8015 15341 -7977 15503
rect -6870 15581 -6800 15587
rect -6405 15581 -6369 15916
rect -6312 15892 -6272 16158
rect -6312 15887 -6202 15892
rect -6312 15853 -5910 15887
rect -6312 15847 -6202 15853
rect -6307 15646 -6252 15801
rect -6298 15609 -6264 15646
rect -6870 15511 -6367 15581
rect -8015 15307 -7633 15341
rect -8478 15209 -8170 15243
rect -8128 15178 -8088 15248
rect -8128 15177 -8086 15178
rect -8126 14662 -8086 15177
rect -8038 15124 -7984 15259
rect -8030 15104 -7990 15124
rect -8028 14897 -7992 15104
rect -7970 14726 -7762 14760
rect -8300 14629 -8086 14662
rect -8300 14628 -8092 14629
rect -7970 14530 -7762 14564
rect -6870 15343 -6800 15511
rect -7042 15309 -6800 15343
rect -6811 15211 -6703 15245
rect -7042 15113 -6934 15147
rect -6811 15015 -6703 15049
rect -7042 14917 -6934 14951
rect -6900 14799 -6840 14872
rect -6887 14738 -6846 14799
rect -6887 14727 -6667 14738
rect -6887 14699 -6659 14727
rect -6859 14677 -6659 14699
rect -8300 14432 -8092 14466
rect -7970 14334 -7762 14368
rect -8064 14216 -8004 14289
rect -8058 14172 -8017 14216
rect -6697 14538 -6659 14677
rect -6612 14590 -6541 14664
rect -6504 14602 -6196 14636
rect -7041 14504 -6659 14538
rect -6697 14342 -6659 14504
rect -7041 14308 -6659 14342
rect -8150 14042 -8000 14172
rect -8100 13667 -8066 14042
rect -6586 14249 -6547 14590
rect -6504 14504 -6196 14538
rect -6504 14406 -6196 14440
rect -6586 14179 -6546 14249
rect -6504 14210 -6196 14244
rect -6588 14178 -6546 14179
rect -6588 13952 -6548 14178
rect -8501 13633 -7585 13667
rect -8048 13463 -7994 13598
rect -8501 13220 -8095 13254
rect -8633 13122 -8193 13156
rect -8633 12946 -8599 13122
rect -8129 13058 -8095 13220
rect -8041 13058 -8004 13463
rect -8501 13024 -7829 13058
rect -8129 13021 -7829 13024
rect -8633 12945 -8490 12946
rect -8633 12911 -8193 12945
rect -8633 12750 -8596 12911
rect -8046 12852 -7992 12987
rect -7866 12929 -7829 13021
rect -7866 12895 -7585 12929
rect -8193 12847 -8095 12848
rect -8501 12813 -8095 12847
rect -8633 12749 -8492 12750
rect -8633 12715 -8193 12749
rect -8130 12635 -8095 12813
rect -8500 12601 -8095 12635
rect -8129 12439 -8095 12601
rect -8500 12405 -8095 12439
rect -8039 12345 -8005 12852
rect -7968 12664 -7914 12799
rect -7866 12733 -7829 12895
rect -7866 12699 -7585 12733
rect -8180 12311 -8005 12345
rect -8180 12174 -8146 12311
rect -7961 12271 -7923 12664
rect -7866 12537 -7829 12699
rect -7866 12503 -7585 12537
rect -7886 12328 -7832 12463
rect -7877 12309 -7840 12328
rect -8052 12213 -7915 12271
rect -7961 12187 -7923 12213
rect -8183 12116 -8046 12174
rect -7875 12009 -7840 12309
rect -7921 11968 -7840 12009
rect -8280 11902 -8143 11960
rect -7921 11765 -7851 11968
rect -7921 11731 -7679 11765
rect -8018 11633 -7910 11667
rect -7787 11535 -7679 11569
rect -8018 11437 -7910 11471
rect -7787 11339 -7679 11373
rect -7881 11221 -7821 11294
rect -7875 11160 -7834 11221
rect -8054 11149 -7834 11160
rect -8062 11121 -7834 11149
rect -8062 11099 -7862 11121
rect -8525 11024 -8217 11058
rect -8525 10926 -8217 10960
rect -8525 10828 -8217 10862
rect -8062 10960 -8024 11099
rect -8062 10926 -7680 10960
rect -8062 10764 -8024 10926
rect -8062 10730 -7680 10764
rect -8525 10632 -8217 10666
rect -6001 14077 -5943 14141
rect -6012 13707 -5942 14077
rect -6012 13673 -5770 13707
rect -6109 13575 -6001 13609
rect -5878 13477 -5770 13511
rect -6109 13379 -6001 13413
rect -5878 13281 -5770 13315
rect -5972 13163 -5912 13236
rect -5966 13102 -5925 13163
rect -6145 13091 -5925 13102
rect -6153 13063 -5925 13091
rect -6153 13041 -5953 13063
rect -6616 12966 -6308 13000
rect -6616 12868 -6308 12902
rect -6616 12770 -6308 12804
rect -6153 12902 -6115 13041
rect -6153 12868 -5771 12902
rect -6153 12706 -6115 12868
rect -6153 12672 -5771 12706
rect -6616 12574 -6308 12608
rect -6565 11803 -5649 11837
rect -6112 11633 -6058 11768
rect -6565 11390 -6159 11424
rect -6697 11292 -6257 11326
rect -6697 11116 -6663 11292
rect -6193 11228 -6159 11390
rect -6105 11228 -6068 11633
rect -6565 11194 -5893 11228
rect -6193 11191 -5893 11194
rect -6697 11115 -6554 11116
rect -6697 11081 -6257 11115
rect -6697 10920 -6660 11081
rect -5930 11099 -5893 11191
rect -5930 11065 -5649 11099
rect -6257 11017 -6159 11018
rect -6565 10983 -6159 11017
rect -6697 10919 -6556 10920
rect -6697 10885 -6257 10919
rect -6194 10805 -6159 10983
rect -6564 10771 -6159 10805
rect -6193 10609 -6159 10771
rect -6564 10575 -6159 10609
rect -5930 10903 -5893 11065
rect -5930 10869 -5649 10903
rect -5930 10707 -5893 10869
rect -5930 10673 -5649 10707
rect -117 10807 73 12397
rect 93931 12460 95152 38495
rect 14781 10133 15093 10167
rect 15184 10133 15392 10167
rect 16414 10138 16622 10172
rect 15059 10088 15093 10133
rect 15044 10007 15119 10088
rect 15184 9875 15792 9909
rect 15040 9651 15115 9674
rect 14781 9617 15115 9651
rect 15184 9617 15392 9651
rect 15040 9593 15115 9617
rect 15437 9393 15542 9875
rect 16282 9998 16360 10071
rect 15184 9359 15792 9393
rect -13709 7552 -9468 7738
rect -13709 2685 -13523 7552
rect 15018 9147 15088 9218
rect 15494 9206 15561 9273
rect 15018 9135 15071 9147
rect 14781 9101 15071 9135
rect 15184 9101 15392 9135
rect 14988 9100 15071 9101
rect 14586 8817 14773 8899
rect 15018 8817 15071 9100
rect 15504 8888 15538 9206
rect 15916 9880 16222 9914
rect 15916 9398 15950 9880
rect 16307 9790 16341 9998
rect 16414 9880 17022 9914
rect 16283 9717 16361 9790
rect 16307 9509 16341 9717
rect 16414 9622 16622 9656
rect 16288 9436 16366 9509
rect 16307 9398 16341 9436
rect 16669 9398 16703 9880
rect 69374 9778 69806 9916
rect 91774 9778 92206 9916
rect 15916 9364 16341 9398
rect 16414 9364 17022 9398
rect 15504 8854 15890 8888
rect 15927 8833 15995 8897
rect 16029 8854 16121 8888
rect 14586 8764 15071 8817
rect 6966 8691 7312 8756
rect 14586 8746 14773 8764
rect 15018 8739 15071 8764
rect 15942 8691 15978 8833
rect 16304 8743 16338 9364
rect 16716 9208 16784 9274
rect 16414 9106 16622 9140
rect 6966 8530 16005 8691
rect 16226 8605 16396 8743
rect 6966 8466 7312 8530
rect 7289 8261 7635 8307
rect 16722 8261 16775 9208
rect 7289 8079 16799 8261
rect 7289 8017 7635 8079
rect 9002 6558 9036 7500
rect 9234 6558 9350 6614
rect 9534 6558 9650 6614
rect 9834 6558 9950 6614
rect 10134 6558 10250 6614
rect 10434 6558 10550 6614
rect 10718 6558 10752 7500
rect 12164 6562 12198 7500
rect 14997 6931 15211 6970
rect 19201 6931 19643 7085
rect 22939 6931 23303 7116
rect 14997 6807 23303 6931
rect 14997 6756 15211 6807
rect 16227 6562 16406 6623
rect 19201 6620 19643 6807
rect 22939 6666 23303 6807
rect 9002 6524 10788 6558
rect 9038 5639 9072 6524
rect 10754 5639 10788 6524
rect 12164 6480 16406 6562
rect 16227 6444 16406 6480
rect 13866 5898 14130 5964
rect 12465 5641 14130 5898
rect 12470 4639 12504 5641
rect 18791 5216 19168 5573
rect -5845 2685 -5539 2764
rect -13709 2548 -5539 2685
rect -5845 2483 -5539 2548
rect 262 2542 1111 2595
rect -9731 1371 -9659 1425
rect -9385 1371 -9351 1979
rect -9149 1571 -9115 1979
rect -8913 1571 -8879 1979
rect -8677 1571 -8643 1979
rect -8441 1571 -8407 1979
rect -8205 1571 -8171 1979
rect -7969 1571 -7935 1979
rect -7733 1571 -7699 1979
rect -9731 1337 -9351 1371
rect -7843 1385 -7771 1459
rect -7367 1385 -7333 1979
rect -7131 1571 -7097 1979
rect -6895 1571 -6861 1979
rect -6659 1571 -6625 1979
rect -6293 1505 -6259 1979
rect -6057 1571 -6023 1979
rect -3486 2037 -3452 2041
rect -3492 1784 -3446 2037
rect -3290 1849 -3256 2041
rect -3296 1784 -3250 1849
rect -3094 1849 -3060 2041
rect -3100 1784 -3054 1849
rect -2636 2037 -2602 2041
rect -3492 1776 -3054 1784
rect -2642 1784 -2596 2037
rect -2440 1849 -2406 2041
rect -2446 1784 -2400 1849
rect -2042 2110 -1874 2150
rect -2168 2076 -1874 2110
rect -2244 1849 -2210 2041
rect -2250 1784 -2204 1849
rect -2642 1776 -2204 1784
rect -2168 1776 -2134 2076
rect -3492 1761 -2888 1776
rect -2846 1761 -2678 1769
rect -3492 1738 -2678 1761
rect -5642 1514 -5574 1521
rect -6467 1471 -6259 1505
rect -7843 1351 -7333 1385
rect -6912 1382 -6810 1430
rect -6467 1382 -6433 1471
rect -9731 1269 -9659 1337
rect -7843 1303 -7771 1351
rect -6912 1348 -6433 1382
rect -6310 1352 -6234 1412
rect -5779 1352 -5574 1514
rect -4212 1461 -4099 1535
rect -6912 1290 -6810 1348
rect -6310 1299 -5642 1352
rect -6310 1291 -5701 1299
rect -13337 1235 -9855 1263
rect -6310 1235 -6234 1291
rect -13337 1171 -9707 1235
rect -13311 763 -13277 1171
rect -13193 763 -13159 1171
rect -13075 763 -13041 1171
rect -12957 763 -12923 1171
rect -12839 763 -12805 1171
rect -12721 763 -12687 1171
rect -12603 763 -12569 1171
rect -12485 763 -12451 1171
rect -12367 763 -12333 1171
rect -12249 763 -12215 1171
rect -12131 763 -12097 1171
rect -12013 763 -11979 1171
rect -11895 763 -11861 1171
rect -11777 763 -11743 1171
rect -11659 763 -11625 1171
rect -11541 763 -11507 1171
rect -11423 763 -11389 1171
rect -11305 763 -11271 1171
rect -11187 763 -11153 1171
rect -11069 763 -11035 1171
rect -10951 763 -10917 1171
rect -10833 763 -10799 1171
rect -10715 763 -10681 1171
rect -10597 763 -10563 1171
rect -10479 763 -10445 1171
rect -10361 763 -10327 1171
rect -10243 763 -10209 1171
rect -10125 763 -10091 1171
rect -10007 763 -9973 1171
rect -9889 763 -9855 1171
rect -9771 692 -9737 1171
rect -9535 692 -9501 1171
rect -9299 692 -9265 1171
rect -9063 692 -9029 1171
rect -8827 692 -8793 1171
rect -8591 692 -8557 1171
rect -8355 692 -8321 1171
rect -8119 692 -8085 1171
rect -7883 692 -7849 1171
rect -7765 763 -7731 1171
rect -7647 692 -7613 1171
rect -7529 763 -7495 1171
rect -7411 692 -7377 1171
rect -7293 763 -7259 1171
rect -7175 692 -7141 1171
rect -7057 763 -7023 1171
rect -6939 692 -6905 1171
rect -6821 763 -6787 1171
rect -6703 692 -6669 1171
rect -6585 763 -6551 1171
rect -6467 692 -6433 1171
rect -6349 763 -6315 1171
rect -6231 692 -6197 1171
rect -13321 680 -6175 692
rect -4187 680 -4102 1461
rect -3584 1502 -3550 1661
rect -3492 1645 -3446 1738
rect -3486 1553 -3452 1645
rect -3388 1502 -3354 1661
rect -3296 1645 -3250 1738
rect -3100 1709 -2678 1738
rect -3100 1706 -2888 1709
rect -3290 1553 -3256 1645
rect -3192 1502 -3158 1661
rect -3100 1645 -3054 1706
rect -2846 1695 -2678 1709
rect -2642 1738 -2134 1776
rect -3094 1553 -3060 1645
rect -2734 1502 -2700 1661
rect -2642 1645 -2596 1738
rect -2636 1553 -2602 1645
rect -2538 1502 -2504 1661
rect -2446 1645 -2400 1738
rect -2250 1706 -2134 1738
rect -2088 1784 -2054 2041
rect -1990 1833 -1956 2041
rect -1892 1784 -1858 2041
rect -1794 1833 -1760 2041
rect -1696 1784 -1662 2041
rect -1598 1833 -1564 2041
rect -1500 1784 -1466 2041
rect -1402 1833 -1368 2041
rect -1304 1784 -1270 2041
rect -2088 1750 -1270 1784
rect -2440 1553 -2406 1645
rect -2342 1502 -2308 1661
rect -2250 1645 -2204 1706
rect -2244 1553 -2210 1645
rect -3593 1434 -2209 1502
rect -2088 1487 -2054 1750
rect -1990 1487 -1956 1695
rect -1892 1487 -1858 1750
rect -1794 1487 -1760 1695
rect -1696 1487 -1662 1750
rect -1598 1487 -1564 1695
rect -1500 1487 -1466 1750
rect -1402 1487 -1368 1695
rect -1304 1487 -1270 1750
rect -2743 1297 -2209 1434
rect -2734 1138 -2700 1297
rect -2636 1154 -2602 1246
rect -13321 678 -4102 680
rect -13342 595 -4102 678
rect -13342 558 -6155 595
rect -2642 1061 -2596 1154
rect -2538 1138 -2504 1297
rect -2440 1154 -2406 1246
rect -2446 1061 -2400 1154
rect -2342 1138 -2308 1297
rect -2244 1154 -2210 1246
rect -2250 1093 -2204 1154
rect -2250 1061 -2134 1093
rect -2642 1023 -2134 1061
rect -2642 1015 -2204 1023
rect -2642 762 -2596 1015
rect -2636 758 -2602 762
rect -2446 950 -2400 1015
rect -2440 758 -2406 950
rect -2250 950 -2204 1015
rect -2244 758 -2210 950
rect -2168 723 -2134 1023
rect -1990 1104 -1956 1312
rect -1794 1104 -1760 1312
rect -1598 1104 -1564 1312
rect -1402 1104 -1368 1312
rect -1990 758 -1956 966
rect -1794 758 -1760 966
rect -1598 758 -1564 966
rect -1402 758 -1368 966
rect -2168 689 -1874 723
rect -2042 649 -1874 689
rect 262 978 315 2542
rect 1034 2501 1111 2542
rect 738 2467 975 2497
rect 469 2428 975 2467
rect 469 1923 508 2428
rect 738 2401 975 2428
rect 1034 2405 2012 2501
rect 19892 3378 19926 3382
rect 19886 3125 19932 3378
rect 20088 3190 20122 3382
rect 20082 3125 20128 3190
rect 20284 3190 20318 3382
rect 20278 3125 20324 3190
rect 20742 3378 20776 3382
rect 19886 3117 20324 3125
rect 20736 3125 20782 3378
rect 20938 3190 20972 3382
rect 20932 3125 20978 3190
rect 21336 3451 21504 3491
rect 21210 3417 21504 3451
rect 21134 3190 21168 3382
rect 21128 3125 21174 3190
rect 20736 3117 21174 3125
rect 21210 3117 21244 3417
rect 19886 3102 20490 3117
rect 20532 3102 20700 3110
rect 19886 3079 20700 3102
rect 625 1923 659 2089
rect 895 2148 975 2222
rect 1026 2148 1104 2221
rect 871 1986 905 2114
rect 989 1986 1023 2114
rect 1107 1986 1141 2114
rect 1366 2148 1444 2222
rect 1313 1986 1347 2114
rect 465 1884 659 1923
rect 625 1649 659 1884
rect 693 1932 773 1950
rect 1401 1932 1435 2114
rect 1600 2215 1679 2234
rect 1600 2173 1794 2215
rect 1600 2154 1679 2173
rect 1603 1991 1637 2119
rect 1691 1991 1725 2119
rect 693 1884 1591 1932
rect 1759 1924 1794 2173
rect 1852 2160 2285 2238
rect 1829 1998 1863 2126
rect 1858 1924 2019 1957
rect 693 1859 860 1884
rect 777 1854 860 1859
rect 961 1695 995 1823
rect 1137 1695 1171 1884
rect 1117 1574 1189 1655
rect 1313 1695 1347 1884
rect 1431 1857 1591 1884
rect 1635 1857 1717 1923
rect 1759 1889 2019 1924
rect 1858 1857 2019 1889
rect 2065 1925 2099 2126
rect 2301 1925 2335 2126
rect 2474 1932 2554 1950
rect 2387 1925 2554 1932
rect 2065 1891 2554 1925
rect 1294 1573 1366 1654
rect 1514 1635 1548 1857
rect 1602 1635 1636 1823
rect 1954 1822 1988 1823
rect 2065 1822 2099 1891
rect 2387 1859 2554 1891
rect 2588 1932 2622 2089
rect 2783 1932 2863 1950
rect 2588 1884 2863 1932
rect 2387 1854 2470 1859
rect 1954 1785 2099 1822
rect 1954 1662 1988 1785
rect 2065 1662 2099 1785
rect 1954 1625 2099 1662
rect 2588 1649 2622 1884
rect 2696 1859 2863 1884
rect 2897 1923 2931 2089
rect 4613 2213 4647 2217
rect 4607 1960 4653 2213
rect 4809 2025 4843 2217
rect 4803 1960 4849 2025
rect 5005 2025 5039 2217
rect 4999 1960 5045 2025
rect 5463 2213 5497 2217
rect 4607 1952 5045 1960
rect 5457 1960 5503 2213
rect 5659 2025 5693 2217
rect 5653 1960 5699 2025
rect 6057 2286 6225 2326
rect 5931 2252 6225 2286
rect 5855 2025 5889 2217
rect 5849 1960 5895 2025
rect 5457 1952 5895 1960
rect 5931 1952 5965 2252
rect 2897 1884 4073 1923
rect 2696 1854 2779 1859
rect 2897 1649 2931 1884
rect 4034 1638 4073 1884
rect 4607 1937 5211 1952
rect 5253 1937 5421 1945
rect 4607 1914 5421 1937
rect 3990 1499 4106 1638
rect 625 978 659 1213
rect 961 1039 995 1167
rect 1117 1207 1189 1288
rect 777 1003 860 1008
rect 262 939 659 978
rect 262 925 508 939
rect 469 434 508 925
rect 625 773 659 939
rect 693 978 860 1003
rect 1137 978 1171 1167
rect 1294 1208 1366 1289
rect 1313 978 1347 1167
rect 1514 1005 1548 1227
rect 1602 1039 1636 1227
rect 1954 1200 2099 1237
rect 1954 1077 1988 1200
rect 2065 1077 2099 1200
rect 1954 1040 2099 1077
rect 1954 1039 1988 1040
rect 1431 978 1591 1005
rect 693 930 1591 978
rect 1635 939 1717 1005
rect 1858 973 2019 1005
rect 1759 938 2019 973
rect 693 912 773 930
rect 871 748 905 876
rect 989 748 1023 876
rect 1107 748 1141 876
rect 895 640 975 714
rect 1026 641 1104 714
rect 1313 748 1347 876
rect 1401 748 1435 930
rect 1366 640 1444 714
rect 1603 743 1637 871
rect 1691 743 1725 871
rect 1600 689 1679 708
rect 1759 689 1794 938
rect 1858 905 2019 938
rect 2065 971 2099 1040
rect 2387 1003 2470 1008
rect 2387 971 2554 1003
rect 2065 937 2554 971
rect 1829 736 1863 864
rect 2065 736 2099 937
rect 2301 736 2335 937
rect 2387 930 2554 937
rect 2474 912 2554 930
rect 2588 978 2622 1213
rect 2696 1003 2779 1008
rect 2696 978 2863 1003
rect 2588 930 2863 978
rect 1600 647 1794 689
rect 1600 628 1679 647
rect 1852 624 2285 702
rect 2588 773 2622 930
rect 2783 912 2863 930
rect 2897 978 2931 1213
rect 3563 978 3725 1039
rect 2897 939 3725 978
rect 2897 773 2931 939
rect 3563 885 3725 939
rect 4607 1821 4653 1914
rect 4613 1729 4647 1821
rect 4803 1821 4849 1914
rect 4999 1885 5421 1914
rect 4999 1882 5211 1885
rect 4809 1729 4843 1821
rect 4999 1821 5045 1882
rect 5253 1871 5421 1885
rect 5457 1914 5965 1952
rect 5005 1729 5039 1821
rect 5457 1821 5503 1914
rect 5463 1729 5497 1821
rect 5653 1821 5699 1914
rect 5849 1882 5965 1914
rect 6011 1960 6045 2217
rect 6109 2009 6143 2217
rect 6207 1960 6241 2217
rect 6305 2009 6339 2217
rect 6403 1960 6437 2217
rect 6501 2009 6535 2217
rect 6599 1960 6633 2217
rect 6697 2009 6731 2217
rect 6795 1960 6829 2217
rect 6011 1926 6829 1960
rect 5659 1729 5693 1821
rect 5849 1821 5895 1882
rect 5855 1729 5889 1821
rect 6011 1663 6045 1926
rect 6109 1663 6143 1871
rect 6207 1663 6241 1926
rect 6305 1663 6339 1871
rect 6403 1663 6437 1926
rect 6501 1663 6535 1871
rect 6599 1663 6633 1926
rect 6697 1663 6731 1871
rect 6795 1663 6829 1926
rect 5463 1330 5497 1422
rect 5457 1237 5503 1330
rect 5659 1330 5693 1422
rect 5653 1237 5699 1330
rect 5855 1330 5889 1422
rect 5849 1269 5895 1330
rect 5849 1237 5965 1269
rect 5457 1199 5965 1237
rect 5457 1191 5895 1199
rect 5457 938 5503 1191
rect 5463 934 5497 938
rect 5653 1126 5699 1191
rect 5659 934 5693 1126
rect 5849 1126 5895 1191
rect 5855 934 5889 1126
rect 5931 899 5965 1199
rect 6109 1280 6143 1488
rect 6305 1280 6339 1488
rect 6501 1280 6535 1488
rect 6697 1280 6731 1488
rect 6109 934 6143 1142
rect 6305 934 6339 1142
rect 6501 934 6535 1142
rect 6697 934 6731 1142
rect 5931 865 6225 899
rect 6057 825 6225 865
rect 7054 1845 7303 2079
rect 7736 1853 7770 2261
rect 7096 1568 7234 1845
rect 7972 1787 8006 2261
rect 8338 1853 8372 2261
rect 8574 1853 8608 2261
rect 8810 1853 8844 2261
rect 7972 1753 8180 1787
rect 7337 1634 7470 1680
rect 7947 1634 8023 1694
rect 7337 1573 8023 1634
rect 8146 1664 8180 1753
rect 8523 1664 8625 1712
rect 8146 1630 8625 1664
rect 9046 1667 9080 2261
rect 9412 1853 9446 2261
rect 9648 1853 9682 2261
rect 9884 1853 9918 2261
rect 10120 1853 10154 2261
rect 10356 1853 10390 2261
rect 10592 1853 10626 2261
rect 10828 1853 10862 2261
rect 9484 1667 9556 1741
rect 9046 1633 9556 1667
rect 7029 1334 7278 1568
rect 7337 1562 7470 1573
rect 7947 1517 8023 1573
rect 8523 1572 8625 1630
rect 9484 1585 9556 1633
rect 11064 1653 11098 2261
rect 11372 1653 11444 1707
rect 11064 1619 11444 1653
rect 11372 1551 11444 1619
rect 8028 1045 8062 1453
rect 8264 1045 8298 1453
rect 8500 1045 8534 1453
rect 8736 1045 8770 1453
rect 8972 1045 9006 1453
rect 9208 1045 9242 1453
rect 9444 1045 9478 1453
rect 19886 2986 19932 3079
rect 19892 2894 19926 2986
rect 20082 2986 20128 3079
rect 20278 3050 20700 3079
rect 20278 3047 20490 3050
rect 20088 2894 20122 2986
rect 20278 2986 20324 3047
rect 20532 3036 20700 3050
rect 20736 3079 21244 3117
rect 20284 2894 20318 2986
rect 20736 2986 20782 3079
rect 20742 2894 20776 2986
rect 20932 2986 20978 3079
rect 21128 3047 21244 3079
rect 21290 3125 21324 3382
rect 21388 3174 21422 3382
rect 21486 3125 21520 3382
rect 21584 3174 21618 3382
rect 21682 3125 21716 3382
rect 21780 3174 21814 3382
rect 21878 3125 21912 3382
rect 21976 3174 22010 3382
rect 22074 3125 22108 3382
rect 21290 3091 22108 3125
rect 20938 2894 20972 2986
rect 21128 2986 21174 3047
rect 21134 2894 21168 2986
rect 21290 2828 21324 3091
rect 21388 2828 21422 3036
rect 21486 2828 21520 3091
rect 21584 2828 21618 3036
rect 21682 2828 21716 3091
rect 21780 2828 21814 3036
rect 21878 2828 21912 3091
rect 21976 2828 22010 3036
rect 22074 2828 22108 3091
rect 20742 2495 20776 2587
rect 20736 2402 20782 2495
rect 20938 2495 20972 2587
rect 20932 2402 20978 2495
rect 21134 2495 21168 2587
rect 21128 2434 21174 2495
rect 21128 2402 21244 2434
rect 20736 2364 21244 2402
rect 20736 2356 21174 2364
rect 20736 2103 20782 2356
rect 20742 2099 20776 2103
rect 20932 2291 20978 2356
rect 20938 2099 20972 2291
rect 21128 2291 21174 2356
rect 21134 2099 21168 2291
rect 21210 2064 21244 2364
rect 21388 2445 21422 2653
rect 21584 2445 21618 2653
rect 21780 2445 21814 2653
rect 21976 2445 22010 2653
rect 21388 2099 21422 2307
rect 21584 2099 21618 2307
rect 21780 2099 21814 2307
rect 21976 2099 22010 2307
rect 21210 2030 21504 2064
rect 21336 1990 21504 2030
rect 22316 2711 22554 2900
rect 22376 2297 22532 2711
rect 25061 2297 25333 2372
rect 22376 2141 25333 2297
rect 25061 2085 25333 2141
rect 738 434 975 461
rect 469 395 975 434
rect 738 365 975 395
rect 1034 361 2012 457
rect -13197 -274 -7163 -135
rect -13197 -378 -5720 -274
rect -13197 -453 -7163 -378
rect -4954 -335 -4920 -331
rect -4960 -588 -4914 -335
rect -4758 -523 -4724 -331
rect -4764 -588 -4718 -523
rect -4562 -523 -4528 -331
rect -4568 -588 -4522 -523
rect -4104 -335 -4070 -331
rect -4960 -596 -4522 -588
rect -4110 -588 -4064 -335
rect -3908 -523 -3874 -331
rect -3914 -588 -3868 -523
rect -3510 -262 -3342 -222
rect -3636 -296 -3342 -262
rect -3712 -523 -3678 -331
rect -3718 -588 -3672 -523
rect -4110 -596 -3672 -588
rect -3636 -596 -3602 -296
rect -25553 -806 -25165 -654
rect -4960 -611 -4356 -596
rect -4314 -611 -4146 -603
rect -4960 -634 -4146 -611
rect -5976 -806 -5800 -784
rect -25553 -943 -5800 -806
rect -25553 -1050 -25165 -943
rect -5976 -1005 -5800 -943
rect -5052 -869 -5018 -711
rect -4960 -727 -4914 -634
rect -4954 -819 -4920 -727
rect -4856 -869 -4822 -711
rect -4764 -727 -4718 -634
rect -4568 -663 -4146 -634
rect -4568 -666 -4356 -663
rect -4758 -819 -4724 -727
rect -4660 -869 -4626 -711
rect -4568 -727 -4522 -666
rect -4314 -677 -4146 -663
rect -4110 -634 -3602 -596
rect -4562 -819 -4528 -727
rect -5052 -870 -4568 -869
rect -4202 -870 -4168 -711
rect -4110 -727 -4064 -634
rect -4104 -819 -4070 -727
rect -4006 -870 -3972 -711
rect -3914 -727 -3868 -634
rect -3718 -666 -3602 -634
rect -3556 -588 -3522 -331
rect -3458 -539 -3424 -331
rect -3360 -588 -3326 -331
rect -3262 -539 -3228 -331
rect -3164 -588 -3130 -331
rect -3066 -539 -3032 -331
rect -2968 -588 -2934 -331
rect -2870 -539 -2836 -331
rect -2772 -588 -2738 -331
rect -3556 -622 -2738 -588
rect -3908 -819 -3874 -727
rect -3810 -870 -3776 -711
rect -3718 -727 -3672 -666
rect -3712 -819 -3678 -727
rect -5061 -938 -3677 -870
rect -3556 -885 -3522 -622
rect -3458 -885 -3424 -677
rect -3360 -885 -3326 -622
rect -3262 -885 -3228 -677
rect -3164 -885 -3130 -622
rect -3066 -885 -3032 -677
rect -2968 -885 -2934 -622
rect -2870 -885 -2836 -677
rect -2772 -885 -2738 -622
rect -4211 -1075 -3677 -938
rect -4202 -1234 -4168 -1075
rect -4104 -1218 -4070 -1126
rect -4110 -1311 -4064 -1218
rect -4006 -1234 -3972 -1075
rect -3908 -1218 -3874 -1126
rect -3914 -1311 -3868 -1218
rect -3810 -1234 -3776 -1075
rect -3712 -1218 -3678 -1126
rect -3718 -1279 -3672 -1218
rect -3718 -1311 -3602 -1279
rect -4110 -1349 -3602 -1311
rect -4110 -1357 -3672 -1349
rect -4110 -1610 -4064 -1357
rect -4104 -1614 -4070 -1610
rect -3914 -1422 -3868 -1357
rect -3908 -1614 -3874 -1422
rect -3718 -1422 -3672 -1357
rect -3712 -1614 -3678 -1422
rect -3636 -1649 -3602 -1349
rect -3556 -1323 -3522 -1060
rect -3458 -1268 -3424 -1060
rect -3360 -1323 -3326 -1060
rect -3262 -1268 -3228 -1060
rect -3164 -1323 -3130 -1060
rect -3066 -1268 -3032 -1060
rect -2968 -1323 -2934 -1060
rect -2870 -1268 -2836 -1060
rect -2772 -1323 -2738 -1060
rect -3556 -1357 -2738 -1323
rect -3556 -1614 -3522 -1357
rect -3458 -1614 -3424 -1406
rect -3360 -1614 -3326 -1357
rect -3262 -1614 -3228 -1406
rect -3164 -1614 -3130 -1357
rect -3066 -1614 -3032 -1406
rect -2968 -1614 -2934 -1357
rect -2870 -1614 -2836 -1406
rect -2772 -1614 -2738 -1357
rect -3636 -1683 -3342 -1649
rect -3510 -1723 -3342 -1683
rect 25955 2273 26111 2333
rect 25955 2145 27588 2273
rect 25955 2116 26111 2145
rect 27791 2209 27952 2240
rect 27791 2179 28006 2209
rect 28063 2179 28219 2202
rect 27791 2161 28219 2179
rect 27913 2140 28219 2161
rect 28063 2125 28219 2140
rect 28109 1819 28143 2061
rect 28425 1853 28459 2061
rect 28741 1819 28775 2061
rect 28871 1858 28905 2066
rect 29101 2109 29269 2195
rect 29187 1819 29221 2066
rect 30488 2016 30522 2500
rect 30804 2016 30838 2500
rect 32647 2172 32812 2233
rect 32918 2172 33074 2195
rect 32647 2153 33074 2172
rect 32742 2133 33074 2153
rect 32918 2118 33074 2133
rect 29642 1922 30437 2004
rect 30488 1982 30838 2016
rect 29642 1819 29724 1922
rect 28000 1778 29803 1819
rect 28000 1290 28041 1778
rect 28109 1464 28143 1672
rect 28425 1464 28459 1778
rect 28741 1464 28775 1672
rect 28871 1464 28905 1778
rect 29075 1722 29803 1778
rect 29187 1464 29221 1672
rect 29806 1422 29847 1445
rect 29260 1356 29847 1422
rect 28000 1284 29070 1290
rect 30488 1436 30522 1982
rect 30804 1928 30838 1982
rect 30804 1894 31991 1928
rect 30804 1436 30838 1894
rect 31120 1436 31154 1894
rect 31436 1436 31470 1894
rect 27507 1246 29070 1284
rect 20064 28 20098 32
rect 20058 -225 20104 28
rect 20260 -160 20294 32
rect 20254 -225 20300 -160
rect 20456 -160 20490 32
rect 20450 -225 20496 -160
rect 20914 28 20948 32
rect 20058 -233 20496 -225
rect 20908 -225 20954 28
rect 21110 -160 21144 32
rect 21104 -225 21150 -160
rect 21508 101 21676 141
rect 21382 67 21676 101
rect 21306 -160 21340 32
rect 21300 -225 21346 -160
rect 20908 -233 21346 -225
rect 21382 -233 21416 67
rect 4628 -477 4662 -473
rect 4622 -730 4668 -477
rect 4824 -665 4858 -473
rect 4818 -730 4864 -665
rect 5020 -665 5054 -473
rect 5014 -730 5060 -665
rect 5478 -477 5512 -473
rect 4622 -738 5060 -730
rect 5472 -730 5518 -477
rect 5674 -665 5708 -473
rect 5668 -730 5714 -665
rect 6072 -404 6240 -364
rect 5946 -438 6240 -404
rect 5870 -665 5904 -473
rect 5864 -730 5910 -665
rect 5472 -738 5910 -730
rect 5946 -738 5980 -438
rect 4622 -753 5226 -738
rect 5268 -753 5436 -745
rect 4622 -776 5436 -753
rect 4622 -869 4668 -776
rect 4628 -961 4662 -869
rect 4818 -869 4864 -776
rect 5014 -805 5436 -776
rect 5014 -808 5226 -805
rect 4824 -961 4858 -869
rect 5014 -869 5060 -808
rect 5268 -819 5436 -805
rect 5472 -776 5980 -738
rect 5020 -961 5054 -869
rect 5472 -869 5518 -776
rect 5478 -961 5512 -869
rect 5668 -869 5714 -776
rect 5864 -808 5980 -776
rect 6026 -730 6060 -473
rect 6124 -681 6158 -473
rect 6222 -730 6256 -473
rect 6320 -681 6354 -473
rect 6418 -730 6452 -473
rect 6516 -681 6550 -473
rect 6614 -730 6648 -473
rect 6712 -681 6746 -473
rect 6810 -730 6844 -473
rect 6026 -764 6844 -730
rect 5674 -961 5708 -869
rect 5864 -869 5910 -808
rect 5870 -961 5904 -869
rect 6026 -1027 6060 -764
rect 6124 -1027 6158 -819
rect 6222 -1027 6256 -764
rect 6320 -1027 6354 -819
rect 6418 -1027 6452 -764
rect 6516 -1027 6550 -819
rect 6614 -1027 6648 -764
rect 6712 -1027 6746 -819
rect 6810 -1027 6844 -764
rect 5478 -1360 5512 -1268
rect 5472 -1453 5518 -1360
rect 5674 -1360 5708 -1268
rect 5668 -1453 5714 -1360
rect 5870 -1360 5904 -1268
rect 5864 -1421 5910 -1360
rect 5864 -1453 5980 -1421
rect 5472 -1491 5980 -1453
rect 5472 -1499 5910 -1491
rect 5472 -1752 5518 -1499
rect 5478 -1756 5512 -1752
rect 5668 -1564 5714 -1499
rect 5674 -1756 5708 -1564
rect 5864 -1564 5910 -1499
rect 5870 -1756 5904 -1564
rect 5946 -1791 5980 -1491
rect 6124 -1410 6158 -1202
rect 6320 -1410 6354 -1202
rect 6516 -1410 6550 -1202
rect 6712 -1410 6746 -1202
rect 6124 -1756 6158 -1548
rect 6320 -1756 6354 -1548
rect 6516 -1756 6550 -1548
rect 6712 -1756 6746 -1548
rect 5946 -1825 6240 -1791
rect 6072 -1865 6240 -1825
rect 20058 -248 20662 -233
rect 20704 -248 20872 -240
rect 20058 -271 20872 -248
rect 7695 -903 7729 -495
rect 7931 -969 7965 -495
rect 8297 -903 8331 -495
rect 8533 -903 8567 -495
rect 8769 -903 8803 -495
rect 7931 -1003 8139 -969
rect 7334 -1122 7443 -1093
rect 7906 -1122 7982 -1062
rect 7334 -1183 7982 -1122
rect 8105 -1092 8139 -1003
rect 8482 -1092 8584 -1044
rect 8105 -1126 8584 -1092
rect 9005 -1089 9039 -495
rect 9371 -903 9405 -495
rect 9607 -903 9641 -495
rect 9843 -903 9877 -495
rect 10079 -903 10113 -495
rect 10315 -903 10349 -495
rect 10551 -903 10585 -495
rect 10787 -903 10821 -495
rect 9443 -1089 9515 -1015
rect 9005 -1123 9515 -1089
rect 7334 -1207 7443 -1183
rect 7906 -1239 7982 -1183
rect 8482 -1184 8584 -1126
rect 9443 -1171 9515 -1123
rect 11023 -1103 11057 -495
rect 20058 -364 20104 -271
rect 20064 -456 20098 -364
rect 20254 -364 20300 -271
rect 20450 -300 20872 -271
rect 20450 -303 20662 -300
rect 20260 -456 20294 -364
rect 20450 -364 20496 -303
rect 20704 -314 20872 -300
rect 20908 -271 21416 -233
rect 20456 -456 20490 -364
rect 20908 -364 20954 -271
rect 20914 -456 20948 -364
rect 21104 -364 21150 -271
rect 21300 -303 21416 -271
rect 21462 -225 21496 32
rect 21560 -176 21594 32
rect 21658 -225 21692 32
rect 21756 -176 21790 32
rect 21854 -225 21888 32
rect 21952 -176 21986 32
rect 22050 -225 22084 32
rect 22148 -176 22182 32
rect 22246 -225 22280 32
rect 21462 -259 22280 -225
rect 21110 -456 21144 -364
rect 21300 -364 21346 -303
rect 21306 -456 21340 -364
rect 21462 -522 21496 -259
rect 21560 -522 21594 -314
rect 21658 -522 21692 -259
rect 21756 -522 21790 -314
rect 21854 -522 21888 -259
rect 21952 -522 21986 -314
rect 22050 -522 22084 -259
rect 22148 -522 22182 -314
rect 22246 -522 22280 -259
rect 20914 -855 20948 -763
rect 11331 -1103 11403 -1049
rect 11023 -1137 11403 -1103
rect 11331 -1205 11403 -1137
rect 20908 -948 20954 -855
rect 21110 -855 21144 -763
rect 21104 -948 21150 -855
rect 21306 -855 21340 -763
rect 21300 -916 21346 -855
rect 21300 -948 21416 -916
rect 20908 -986 21416 -948
rect 20908 -994 21346 -986
rect 7987 -1711 8021 -1303
rect 8223 -1711 8257 -1303
rect 8459 -1711 8493 -1303
rect 8695 -1711 8729 -1303
rect 8931 -1711 8965 -1303
rect 9167 -1711 9201 -1303
rect 9403 -1711 9437 -1303
rect 20908 -1247 20954 -994
rect 20914 -1251 20948 -1247
rect 21104 -1059 21150 -994
rect 21110 -1251 21144 -1059
rect 21300 -1059 21346 -994
rect 21306 -1251 21340 -1059
rect 21382 -1286 21416 -986
rect 21560 -905 21594 -697
rect 21756 -905 21790 -697
rect 21952 -905 21986 -697
rect 22148 -905 22182 -697
rect 21560 -1251 21594 -1043
rect 21756 -1251 21790 -1043
rect 21952 -1251 21986 -1043
rect 22148 -1251 22182 -1043
rect 21382 -1320 21676 -1286
rect 21508 -1360 21676 -1320
rect 26278 988 26470 1094
rect 27132 988 27450 1006
rect 26278 923 27450 988
rect 26278 836 26470 923
rect 27132 906 27450 923
rect 27507 772 27545 1246
rect 28000 1215 29070 1246
rect 28000 1199 28130 1215
rect 27655 885 27727 1035
rect 28096 935 28130 1199
rect 28254 935 28288 1143
rect 28412 935 28446 1143
rect 28570 935 28604 1143
rect 28728 935 28762 1215
rect 28846 935 28880 1143
rect 29004 935 29038 1143
rect 28159 885 28230 895
rect 28619 885 28697 896
rect 27655 818 29033 885
rect 27507 735 28880 772
rect 26241 367 26433 546
rect 28096 450 28130 693
rect 28254 485 28288 693
rect 28412 485 28446 735
rect 28570 485 28604 693
rect 28728 450 28762 693
rect 28846 485 28880 735
rect 28916 724 28985 818
rect 29004 485 29038 693
rect 29371 721 29446 869
rect 29390 575 29427 721
rect 29390 493 29797 575
rect 29390 450 29427 493
rect 28069 413 29427 450
rect 28049 367 28213 379
rect 26241 326 28213 367
rect 26241 288 26433 326
rect 28049 309 28213 326
rect 29715 358 29797 493
rect 29715 276 30437 358
rect 30488 298 30522 844
rect 30804 386 30838 844
rect 31120 386 31154 844
rect 31436 386 31470 844
rect 31930 999 31991 1894
rect 32964 1812 32998 2054
rect 33280 1846 33314 2054
rect 33596 1812 33630 2054
rect 33726 1851 33760 2059
rect 33956 2102 34124 2188
rect 34042 1812 34076 2059
rect 35223 2038 35257 2522
rect 35539 2038 35573 2522
rect 39284 2935 39318 2939
rect 39278 2682 39324 2935
rect 39480 2747 39514 2939
rect 39474 2682 39520 2747
rect 39676 2747 39710 2939
rect 39945 2753 40002 2917
rect 39670 2682 39716 2747
rect 40166 2935 40200 2939
rect 39278 2674 39716 2682
rect 40160 2682 40206 2935
rect 40362 2747 40396 2939
rect 40356 2682 40402 2747
rect 40776 2958 41404 2992
rect 40558 2747 40592 2939
rect 40776 2913 40812 2958
rect 40552 2682 40598 2747
rect 40160 2674 40598 2682
rect 40653 2698 40727 2866
rect 40777 2839 40811 2913
rect 40653 2674 40726 2698
rect 34534 1944 35172 2026
rect 35223 2004 35573 2038
rect 34534 1812 34616 1944
rect 32855 1771 34658 1812
rect 32855 1283 32896 1771
rect 32964 1457 32998 1665
rect 33280 1457 33314 1771
rect 33596 1457 33630 1665
rect 33726 1457 33760 1771
rect 33930 1715 34658 1771
rect 34042 1457 34076 1665
rect 34661 1415 34702 1438
rect 34115 1349 34702 1415
rect 35223 1458 35257 2004
rect 35539 1950 35573 2004
rect 36944 1995 36978 2479
rect 37260 1995 37294 2479
rect 39074 2593 39242 2667
rect 39278 2652 39746 2674
rect 39956 2656 40124 2667
rect 39804 2652 39864 2656
rect 39921 2652 40124 2656
rect 39278 2636 40124 2652
rect 39094 2199 39133 2593
rect 39278 2543 39324 2636
rect 39284 2451 39318 2543
rect 39474 2543 39520 2636
rect 39670 2610 40124 2636
rect 39670 2604 39746 2610
rect 39480 2451 39514 2543
rect 39670 2543 39716 2604
rect 39676 2451 39710 2543
rect 39804 2524 39864 2610
rect 39921 2598 40124 2610
rect 39956 2593 40124 2598
rect 40160 2636 40726 2674
rect 40160 2543 40206 2636
rect 40166 2451 40200 2543
rect 40356 2543 40402 2636
rect 40552 2604 40726 2636
rect 40771 2692 40818 2839
rect 40875 2832 40909 2924
rect 40972 2903 41014 2958
rect 40874 2780 40910 2832
rect 40973 2816 41007 2903
rect 41071 2834 41105 2924
rect 41166 2902 41208 2958
rect 41071 2816 41108 2834
rect 41169 2816 41203 2902
rect 41267 2834 41301 2924
rect 41362 2907 41404 2958
rect 41072 2780 41108 2816
rect 41266 2780 41302 2834
rect 41365 2816 41399 2907
rect 41463 2824 41497 2924
rect 41460 2780 41502 2824
rect 40874 2746 41502 2780
rect 40771 2618 40943 2692
rect 41327 2658 41502 2746
rect 41909 2935 41943 2939
rect 41903 2682 41949 2935
rect 42105 2747 42139 2939
rect 42099 2682 42145 2747
rect 42301 2747 42335 2939
rect 42645 2839 42702 2917
rect 42441 2794 42702 2839
rect 42295 2682 42341 2747
rect 41903 2674 42341 2682
rect 41699 2658 41867 2667
rect 40362 2451 40396 2543
rect 40552 2543 40598 2604
rect 40558 2451 40592 2543
rect 40771 2483 40818 2618
rect 41327 2601 41867 2658
rect 41327 2579 41502 2601
rect 41699 2593 41867 2601
rect 41903 2660 42371 2674
rect 42441 2660 42486 2794
rect 42645 2753 42702 2794
rect 42866 2935 42900 2939
rect 42860 2682 42906 2935
rect 43062 2747 43096 2939
rect 43056 2682 43102 2747
rect 43476 2958 44104 2992
rect 43258 2747 43292 2939
rect 43476 2913 43512 2958
rect 43252 2682 43298 2747
rect 42860 2674 43298 2682
rect 43353 2698 43427 2866
rect 43477 2839 43511 2913
rect 43353 2674 43426 2698
rect 41903 2636 42486 2660
rect 40871 2545 41502 2579
rect 40871 2504 40912 2545
rect 40777 2413 40811 2483
rect 40772 2355 40816 2413
rect 40875 2401 40909 2504
rect 40973 2424 41007 2509
rect 41069 2496 41110 2545
rect 40968 2355 41012 2424
rect 41071 2401 41105 2496
rect 41169 2424 41203 2509
rect 41263 2496 41304 2545
rect 41460 2538 41502 2545
rect 41164 2355 41208 2424
rect 41267 2401 41301 2496
rect 41365 2413 41399 2509
rect 41460 2505 41501 2538
rect 41454 2495 41501 2505
rect 41361 2355 41405 2413
rect 41454 2373 41500 2495
rect 41903 2543 41949 2636
rect 41909 2451 41943 2543
rect 42099 2543 42145 2636
rect 42295 2615 42486 2636
rect 42536 2656 42596 2657
rect 42656 2656 42824 2667
rect 42295 2604 42371 2615
rect 42105 2451 42139 2543
rect 42295 2543 42341 2604
rect 42301 2451 42335 2543
rect 42421 2500 42481 2615
rect 42536 2598 42824 2656
rect 42536 2525 42596 2598
rect 42656 2593 42824 2598
rect 42860 2636 43426 2674
rect 42860 2543 42906 2636
rect 42866 2451 42900 2543
rect 43056 2543 43102 2636
rect 43252 2604 43426 2636
rect 43471 2692 43518 2839
rect 43575 2832 43609 2924
rect 43672 2903 43714 2958
rect 43574 2780 43610 2832
rect 43673 2816 43707 2903
rect 43771 2834 43805 2924
rect 43866 2902 43908 2958
rect 43771 2816 43808 2834
rect 43869 2816 43903 2902
rect 43967 2834 44001 2924
rect 44062 2907 44104 2958
rect 43772 2780 43808 2816
rect 43966 2780 44002 2834
rect 44065 2816 44099 2907
rect 44163 2824 44197 2924
rect 44160 2780 44202 2824
rect 43574 2746 44202 2780
rect 43471 2618 43643 2692
rect 44027 2661 44202 2746
rect 44609 2935 44643 2939
rect 44603 2682 44649 2935
rect 44805 2747 44839 2939
rect 44799 2682 44845 2747
rect 45001 2747 45035 2939
rect 44995 2682 45041 2747
rect 44603 2674 45041 2682
rect 44399 2661 44567 2667
rect 43062 2451 43096 2543
rect 43252 2543 43298 2604
rect 43258 2451 43292 2543
rect 43471 2483 43518 2618
rect 44027 2608 44567 2661
rect 44027 2579 44202 2608
rect 44399 2593 44567 2608
rect 44603 2665 45071 2674
rect 44603 2663 45153 2665
rect 44603 2636 45154 2663
rect 43571 2545 44202 2579
rect 43571 2504 43612 2545
rect 43477 2413 43511 2483
rect 40772 2321 41405 2355
rect 43472 2355 43516 2413
rect 43575 2401 43609 2504
rect 43673 2424 43707 2509
rect 43769 2496 43810 2545
rect 43668 2355 43712 2424
rect 43771 2401 43805 2496
rect 43869 2424 43903 2509
rect 43963 2496 44004 2545
rect 44160 2538 44202 2545
rect 43864 2355 43908 2424
rect 43967 2401 44001 2496
rect 44065 2413 44099 2509
rect 44160 2495 44201 2538
rect 44061 2355 44105 2413
rect 44163 2401 44197 2495
rect 44603 2543 44649 2636
rect 44609 2451 44643 2543
rect 44799 2543 44845 2636
rect 44995 2626 45154 2636
rect 44995 2604 45071 2626
rect 44805 2451 44839 2543
rect 44995 2543 45041 2604
rect 45001 2451 45035 2543
rect 43472 2321 44105 2355
rect 39763 2285 39895 2296
rect 44286 2285 44418 2298
rect 39763 2246 44824 2285
rect 45106 2268 45154 2626
rect 39763 2236 39895 2246
rect 44286 2238 44418 2246
rect 41567 2199 41699 2210
rect 42508 2199 42645 2209
rect 39094 2160 44824 2199
rect 36596 1950 36893 1983
rect 35539 1916 36893 1950
rect 35539 1458 35573 1916
rect 35855 1458 35889 1916
rect 36171 1458 36205 1916
rect 36596 1901 36893 1916
rect 36944 1961 37294 1995
rect 36944 1415 36978 1961
rect 37260 1907 37294 1961
rect 38429 1942 38621 2013
rect 39153 1942 39245 2160
rect 41567 2150 41699 2160
rect 42508 2149 42645 2160
rect 45095 2131 45155 2268
rect 40161 1997 40794 2031
rect 38429 1907 39245 1942
rect 37260 1873 39245 1907
rect 32855 1277 33925 1283
rect 32362 1239 33925 1277
rect 31930 981 32305 999
rect 31922 916 32305 981
rect 31987 899 32305 916
rect 32362 765 32400 1239
rect 32855 1208 33925 1239
rect 32855 1192 32985 1208
rect 32510 878 32582 1028
rect 32951 928 32985 1192
rect 33109 928 33143 1136
rect 33267 928 33301 1136
rect 33425 928 33459 1136
rect 33583 928 33617 1208
rect 37260 1415 37294 1873
rect 37576 1415 37610 1873
rect 37892 1415 37926 1873
rect 38429 1850 39245 1873
rect 40069 1857 40103 1951
rect 40161 1939 40205 1997
rect 38429 1755 38621 1850
rect 40065 1814 40106 1857
rect 40167 1843 40201 1939
rect 40265 1856 40299 1951
rect 40358 1928 40402 1997
rect 40064 1807 40106 1814
rect 40262 1807 40303 1856
rect 40363 1843 40397 1928
rect 40461 1856 40495 1951
rect 40554 1928 40598 1997
rect 40456 1807 40497 1856
rect 40559 1843 40593 1928
rect 40657 1848 40691 1951
rect 40750 1939 40794 1997
rect 42861 1997 43494 2031
rect 40755 1869 40789 1939
rect 40654 1807 40695 1848
rect 40064 1775 40695 1807
rect 39989 1773 40695 1775
rect 39989 1715 40239 1773
rect 40748 1734 40795 1869
rect 40974 1809 41008 1901
rect 40968 1748 41014 1809
rect 41170 1809 41204 1901
rect 40064 1606 40239 1715
rect 40623 1660 40795 1734
rect 40064 1572 40692 1606
rect 40064 1528 40106 1572
rect 40069 1428 40103 1528
rect 40167 1445 40201 1536
rect 40264 1518 40300 1572
rect 40458 1536 40494 1572
rect 40162 1394 40204 1445
rect 40265 1428 40299 1518
rect 40363 1450 40397 1536
rect 40458 1518 40495 1536
rect 40358 1394 40400 1450
rect 40461 1428 40495 1518
rect 40559 1449 40593 1536
rect 40656 1520 40692 1572
rect 40552 1394 40594 1449
rect 40657 1428 40691 1520
rect 40748 1513 40795 1660
rect 40840 1716 41014 1748
rect 41164 1716 41210 1809
rect 41366 1809 41400 1901
rect 41360 1716 41406 1809
rect 41610 1759 41670 1918
rect 41811 1809 41845 1901
rect 40840 1678 41406 1716
rect 41442 1696 41670 1759
rect 41805 1748 41851 1809
rect 42007 1809 42041 1901
rect 41707 1716 41851 1748
rect 42001 1716 42047 1809
rect 42203 1809 42237 1901
rect 42197 1716 42243 1809
rect 42769 1857 42803 1951
rect 42861 1939 42905 1997
rect 42765 1814 42806 1857
rect 42867 1843 42901 1939
rect 42965 1856 42999 1951
rect 43058 1928 43102 1997
rect 42764 1807 42806 1814
rect 42962 1807 43003 1856
rect 43063 1843 43097 1928
rect 43161 1856 43195 1951
rect 43254 1928 43298 1997
rect 43156 1807 43197 1856
rect 43259 1843 43293 1928
rect 43357 1848 43391 1951
rect 43450 1939 43494 1997
rect 43455 1869 43489 1939
rect 43354 1807 43395 1848
rect 42764 1773 43395 1807
rect 41442 1685 41610 1696
rect 40840 1654 40913 1678
rect 40755 1439 40789 1513
rect 40839 1486 40913 1654
rect 40968 1670 41406 1678
rect 40968 1605 41014 1670
rect 40754 1394 40790 1439
rect 40974 1413 41008 1605
rect 40162 1360 40790 1394
rect 41164 1605 41210 1670
rect 41170 1413 41204 1605
rect 41360 1417 41406 1670
rect 41707 1678 42243 1716
rect 42279 1752 42447 1759
rect 42279 1692 42469 1752
rect 42673 1713 42939 1773
rect 43448 1734 43495 1869
rect 43674 1809 43708 1901
rect 43668 1748 43714 1809
rect 43870 1809 43904 1901
rect 42279 1685 42447 1692
rect 41366 1413 41400 1417
rect 41564 1549 41621 1599
rect 41707 1549 41769 1678
rect 41805 1670 42243 1678
rect 41805 1605 41851 1670
rect 41564 1487 41769 1549
rect 41564 1435 41621 1487
rect 41811 1413 41845 1605
rect 42001 1605 42047 1670
rect 42007 1413 42041 1605
rect 42197 1417 42243 1670
rect 42203 1413 42237 1417
rect 42764 1606 42939 1713
rect 43323 1660 43495 1734
rect 42764 1572 43392 1606
rect 42764 1528 42806 1572
rect 42769 1428 42803 1528
rect 42867 1445 42901 1536
rect 42964 1518 43000 1572
rect 43158 1536 43194 1572
rect 42862 1394 42904 1445
rect 42965 1428 42999 1518
rect 43063 1450 43097 1536
rect 43158 1518 43195 1536
rect 43058 1394 43100 1450
rect 43161 1428 43195 1518
rect 43259 1449 43293 1536
rect 43356 1520 43392 1572
rect 43252 1394 43294 1449
rect 43357 1428 43391 1520
rect 43448 1513 43495 1660
rect 43540 1716 43714 1748
rect 43864 1716 43910 1809
rect 44066 1809 44100 1901
rect 44060 1716 44106 1809
rect 44322 1759 44382 1903
rect 44511 1809 44545 1901
rect 43540 1678 44106 1716
rect 44142 1697 44382 1759
rect 44505 1748 44551 1809
rect 44707 1809 44741 1901
rect 44418 1716 44551 1748
rect 44701 1716 44747 1809
rect 44903 1809 44937 1901
rect 44897 1716 44943 1809
rect 45106 1759 45154 2131
rect 44142 1696 44345 1697
rect 44142 1685 44310 1696
rect 43540 1654 43613 1678
rect 43455 1439 43489 1513
rect 43539 1486 43613 1654
rect 43668 1670 44106 1678
rect 43668 1605 43714 1670
rect 43454 1394 43490 1439
rect 43674 1413 43708 1605
rect 42862 1360 43490 1394
rect 43864 1605 43910 1670
rect 43870 1413 43904 1605
rect 44060 1417 44106 1670
rect 44418 1678 44943 1716
rect 44979 1715 45154 1759
rect 44979 1685 45147 1715
rect 44066 1413 44100 1417
rect 44264 1548 44321 1599
rect 44418 1548 44464 1678
rect 44505 1670 44943 1678
rect 44505 1605 44551 1670
rect 44264 1499 44464 1548
rect 44264 1435 44321 1499
rect 44511 1413 44545 1605
rect 44701 1605 44747 1670
rect 44707 1413 44741 1605
rect 44897 1417 44943 1670
rect 44903 1413 44937 1417
rect 45351 1935 45497 2121
rect 45400 1852 45444 1935
rect 45677 1899 45711 1991
rect 45400 1849 45565 1852
rect 45400 1798 45635 1849
rect 45467 1775 45635 1798
rect 45671 1806 45717 1899
rect 45873 1899 45907 1991
rect 45867 1806 45913 1899
rect 46069 1899 46103 1991
rect 46063 1838 46109 1899
rect 46637 1838 46961 1997
rect 46063 1806 46961 1838
rect 45671 1768 46961 1806
rect 45671 1760 46109 1768
rect 45671 1507 45717 1760
rect 45677 1503 45711 1507
rect 45867 1695 45913 1760
rect 45873 1503 45907 1695
rect 46063 1695 46109 1760
rect 46069 1503 46103 1695
rect 46637 1686 46961 1768
rect 33701 928 33735 1136
rect 33859 928 33893 1136
rect 33014 878 33085 888
rect 33474 878 33552 889
rect 32510 811 33888 878
rect 46361 1295 46507 1357
rect 46361 1229 46864 1295
rect 46361 1171 46507 1229
rect 32362 728 33735 765
rect 32951 443 32985 686
rect 33109 478 33143 686
rect 33267 478 33301 728
rect 33425 478 33459 686
rect 33583 443 33617 686
rect 33701 478 33735 728
rect 33771 717 33840 811
rect 33859 478 33893 686
rect 34226 714 34301 862
rect 34245 547 34282 714
rect 34245 465 34616 547
rect 34245 443 34282 465
rect 32924 406 34282 443
rect 30804 360 31717 386
rect 34534 381 34616 465
rect 32904 360 33068 372
rect 30804 352 33068 360
rect 30804 298 30838 352
rect 31655 319 33068 352
rect 32904 302 33068 319
rect 34534 299 35172 381
rect 35223 321 35257 867
rect 35539 409 35573 867
rect 35855 409 35889 867
rect 36171 409 36205 867
rect 36596 409 36893 424
rect 35539 375 36893 409
rect 35539 321 35573 375
rect 36596 342 36893 375
rect 36944 364 36978 910
rect 37260 452 37294 910
rect 37576 452 37610 910
rect 37892 452 37926 910
rect 51014 2630 51048 3038
rect 51250 2564 51284 3038
rect 51616 2630 51650 3038
rect 51852 2630 51886 3038
rect 52088 2630 52122 3038
rect 51250 2530 51458 2564
rect 50510 2411 50749 2467
rect 51225 2411 51301 2471
rect 50510 2350 51301 2411
rect 51424 2441 51458 2530
rect 51801 2441 51903 2489
rect 51424 2407 51903 2441
rect 52324 2444 52358 3038
rect 52690 2630 52724 3038
rect 52926 2630 52960 3038
rect 53162 2630 53196 3038
rect 53398 2630 53432 3038
rect 53634 2630 53668 3038
rect 53870 2630 53904 3038
rect 54106 2630 54140 3038
rect 52762 2444 52834 2518
rect 52324 2410 52834 2444
rect 50510 2215 50749 2350
rect 51225 2294 51301 2350
rect 51801 2349 51903 2407
rect 52762 2362 52834 2410
rect 54342 2430 54376 3038
rect 54650 2430 54722 2484
rect 54342 2396 54722 2430
rect 54650 2328 54722 2396
rect 47896 1900 48216 1992
rect 50541 1900 50720 2215
rect 47896 1721 50720 1900
rect 51306 1822 51340 2230
rect 51542 1822 51576 2230
rect 51778 1822 51812 2230
rect 52014 1822 52048 2230
rect 52250 1822 52284 2230
rect 52486 1822 52520 2230
rect 52722 1822 52756 2230
rect 47896 1636 48216 1721
rect 38451 483 38643 565
rect 38451 452 38657 483
rect 37260 418 38657 452
rect 37260 364 37294 418
rect 30488 264 30838 298
rect 27809 -25 27843 183
rect 28125 -25 28159 183
rect 28441 -25 28475 183
rect 28757 -25 28791 183
rect 29073 -25 29107 183
rect 29389 -25 29423 183
rect 30488 -220 30522 264
rect 30804 -220 30838 264
rect 35223 287 35573 321
rect 36944 330 37294 364
rect 38451 380 38657 418
rect 32664 -32 32698 176
rect 32980 -32 33014 176
rect 33296 -32 33330 176
rect 33612 -32 33646 176
rect 33928 -32 33962 176
rect 34244 -32 34278 176
rect 35223 -197 35257 287
rect 35539 -197 35573 287
rect 36944 -154 36978 330
rect 37260 -154 37294 330
rect 38451 307 38643 380
rect 50811 -281 50845 127
rect 51047 -347 51081 127
rect 51413 -281 51447 127
rect 51649 -281 51683 127
rect 51885 -281 51919 127
rect 51047 -381 51255 -347
rect 50434 -500 50725 -478
rect 51022 -500 51098 -440
rect 50434 -561 51098 -500
rect 51221 -470 51255 -381
rect 51598 -470 51700 -422
rect 51221 -504 51700 -470
rect 52121 -467 52155 127
rect 52487 -281 52521 127
rect 52723 -281 52757 127
rect 52959 -281 52993 127
rect 53195 -281 53229 127
rect 53431 -281 53465 127
rect 53667 -281 53701 127
rect 53903 -281 53937 127
rect 52559 -467 52631 -393
rect 52121 -501 52631 -467
rect 50434 -572 50725 -561
rect 47758 -632 50725 -572
rect 51022 -617 51098 -561
rect 51598 -562 51700 -504
rect 52559 -549 52631 -501
rect 54139 -481 54173 127
rect 54447 -481 54519 -427
rect 54139 -515 54519 -481
rect 54447 -583 54519 -515
rect 47758 -726 50588 -632
rect 47758 -752 47953 -726
rect 51103 -1089 51137 -681
rect 51339 -1089 51373 -681
rect 51575 -1089 51609 -681
rect 51811 -1089 51845 -681
rect 52047 -1089 52081 -681
rect 52283 -1089 52317 -681
rect 52519 -1089 52553 -681
rect 50811 -3328 50845 -2920
rect 48966 -3547 49277 -3371
rect 51047 -3394 51081 -2920
rect 51413 -3328 51447 -2920
rect 51649 -3328 51683 -2920
rect 51885 -3328 51919 -2920
rect 51047 -3428 51255 -3394
rect 51022 -3547 51098 -3487
rect 48966 -3608 51098 -3547
rect 51221 -3517 51255 -3428
rect 51598 -3517 51700 -3469
rect 51221 -3551 51700 -3517
rect 52121 -3514 52155 -2920
rect 52487 -3328 52521 -2920
rect 52723 -3328 52757 -2920
rect 52959 -3328 52993 -2920
rect 53195 -3328 53229 -2920
rect 53431 -3328 53465 -2920
rect 53667 -3328 53701 -2920
rect 53903 -3328 53937 -2920
rect 52559 -3514 52631 -3440
rect 52121 -3548 52631 -3514
rect 48966 -3697 49277 -3608
rect 51022 -3664 51098 -3608
rect 51598 -3609 51700 -3551
rect 52559 -3596 52631 -3548
rect 54139 -3528 54173 -2920
rect 54387 -3328 54421 -2920
rect 54623 -3328 54657 -2920
rect 54859 -3328 54893 -2920
rect 55095 -3328 55129 -2920
rect 55331 -3328 55365 -2920
rect 55567 -3328 55601 -2920
rect 55803 -3328 55837 -2920
rect 56039 -3328 56073 -2920
rect 56275 -3328 56309 -2920
rect 56511 -3328 56545 -2920
rect 56747 -3328 56781 -2920
rect 56983 -3328 57017 -2920
rect 57219 -3328 57253 -2920
rect 57455 -3328 57489 -2920
rect 57691 -3328 57725 -2920
rect 57927 -3328 57961 -2920
rect 58163 -3432 58197 -2920
rect 62491 -2838 62525 -2834
rect 62485 -3091 62531 -2838
rect 62687 -3026 62721 -2834
rect 62681 -3091 62727 -3026
rect 62883 -3026 62917 -2834
rect 62877 -3091 62923 -3026
rect 63341 -2838 63375 -2834
rect 62485 -3099 62923 -3091
rect 63335 -3091 63381 -2838
rect 63537 -3026 63571 -2834
rect 63531 -3091 63577 -3026
rect 63935 -2765 64103 -2725
rect 63809 -2799 64103 -2765
rect 63733 -3026 63767 -2834
rect 63727 -3091 63773 -3026
rect 63335 -3099 63773 -3091
rect 63809 -3099 63843 -2799
rect 62485 -3114 63089 -3099
rect 63131 -3114 63299 -3106
rect 62485 -3137 63299 -3114
rect 61873 -3432 62067 -3407
rect 58163 -3474 62067 -3432
rect 54447 -3528 54519 -3474
rect 58163 -3508 62096 -3474
rect 61873 -3516 62067 -3508
rect 54139 -3562 54519 -3528
rect 54447 -3630 54519 -3562
rect 51103 -4136 51137 -3728
rect 51339 -4136 51373 -3728
rect 51575 -4136 51609 -3728
rect 51811 -4136 51845 -3728
rect 52047 -4136 52081 -3728
rect 52283 -4136 52317 -3728
rect 52519 -4136 52553 -3728
rect 52755 -4136 52789 -3728
rect 52991 -4136 53025 -3728
rect 53227 -4136 53261 -3728
rect 53463 -4136 53497 -3728
rect 53699 -4136 53733 -3728
rect 53935 -4136 53969 -3728
rect 54171 -4136 54205 -3728
rect 54407 -4136 54441 -3728
rect 62485 -3230 62531 -3137
rect 62491 -3322 62525 -3230
rect 62681 -3230 62727 -3137
rect 62877 -3166 63299 -3137
rect 62877 -3169 63089 -3166
rect 62687 -3322 62721 -3230
rect 62877 -3230 62923 -3169
rect 63131 -3180 63299 -3166
rect 63335 -3137 63843 -3099
rect 62883 -3322 62917 -3230
rect 63335 -3230 63381 -3137
rect 63341 -3322 63375 -3230
rect 63531 -3230 63577 -3137
rect 63727 -3169 63843 -3137
rect 63889 -3091 63923 -2834
rect 63987 -3042 64021 -2834
rect 64085 -3091 64119 -2834
rect 64183 -3042 64217 -2834
rect 64281 -3091 64315 -2834
rect 64379 -3042 64413 -2834
rect 64477 -3091 64511 -2834
rect 64575 -3042 64609 -2834
rect 64673 -3091 64707 -2834
rect 63889 -3125 64707 -3091
rect 63537 -3322 63571 -3230
rect 63727 -3230 63773 -3169
rect 63733 -3322 63767 -3230
rect 63889 -3388 63923 -3125
rect 63987 -3388 64021 -3180
rect 64085 -3388 64119 -3125
rect 64183 -3388 64217 -3180
rect 64281 -3388 64315 -3125
rect 64379 -3388 64413 -3180
rect 64477 -3388 64511 -3125
rect 64575 -3388 64609 -3180
rect 64673 -3388 64707 -3125
rect 63341 -3721 63375 -3629
rect 63335 -3814 63381 -3721
rect 63537 -3721 63571 -3629
rect 63531 -3814 63577 -3721
rect 63733 -3721 63767 -3629
rect 63727 -3782 63773 -3721
rect 63727 -3814 63843 -3782
rect 63335 -3852 63843 -3814
rect 63335 -3860 63773 -3852
rect 63335 -4113 63381 -3860
rect 63341 -4117 63375 -4113
rect 63531 -3925 63577 -3860
rect 63537 -4117 63571 -3925
rect 63727 -3925 63773 -3860
rect 63733 -4117 63767 -3925
rect 63809 -4152 63843 -3852
rect 63987 -3771 64021 -3563
rect 64183 -3771 64217 -3563
rect 64379 -3771 64413 -3563
rect 64575 -3771 64609 -3563
rect 63987 -4117 64021 -3909
rect 64183 -4117 64217 -3909
rect 64379 -4117 64413 -3909
rect 64575 -4117 64609 -3909
rect 63809 -4186 64103 -4152
rect 63935 -4226 64103 -4186
rect 87785 -3288 88210 -3189
rect 65127 -3507 88210 -3288
rect 87785 -3581 88210 -3507
rect -26907 -11088 -25983 -10980
rect -24373 -11088 -23278 -10959
rect -26907 -11732 -23278 -11088
rect -26907 -11904 -25983 -11732
rect -24373 -11840 -23278 -11732
rect -25931 -14188 -24870 -14108
rect -25931 -14808 -7185 -14188
rect -25931 -14876 -24870 -14808
rect -12874 -15119 -7870 -14969
rect -14982 -15239 -7795 -15119
rect -14951 -15732 -14917 -15324
rect -14833 -15732 -14799 -15324
rect -14715 -15732 -14681 -15324
rect -14597 -15732 -14563 -15324
rect -14479 -15732 -14445 -15324
rect -14361 -15732 -14327 -15324
rect -14243 -15732 -14209 -15324
rect -14125 -15732 -14091 -15324
rect -14007 -15732 -13973 -15324
rect -13889 -15732 -13855 -15324
rect -13771 -15732 -13737 -15324
rect -13653 -15732 -13619 -15324
rect -13535 -15732 -13501 -15324
rect -13417 -15732 -13383 -15324
rect -13299 -15732 -13265 -15324
rect -13181 -15732 -13147 -15324
rect -13063 -15732 -13029 -15324
rect -12945 -15732 -12911 -15324
rect -12827 -15732 -12793 -15324
rect -12709 -15732 -12675 -15324
rect -12591 -15732 -12557 -15324
rect -12473 -15732 -12439 -15324
rect -12355 -15732 -12321 -15324
rect -12237 -15732 -12203 -15324
rect -12119 -15732 -12085 -15324
rect -12001 -15732 -11967 -15324
rect -11883 -15732 -11849 -15324
rect -11765 -15732 -11731 -15324
rect -11647 -15732 -11613 -15324
rect -11529 -15732 -11495 -15324
rect -11411 -15732 -11377 -15239
rect -11175 -15732 -11141 -15239
rect -10939 -15732 -10905 -15239
rect -10703 -15732 -10669 -15239
rect -10467 -15732 -10433 -15239
rect -10231 -15732 -10197 -15239
rect -9995 -15732 -9961 -15239
rect -9759 -15732 -9725 -15239
rect -9523 -15732 -9489 -15239
rect -9405 -15732 -9371 -15324
rect -9287 -15732 -9253 -15239
rect -9169 -15732 -9135 -15324
rect -9051 -15732 -9017 -15239
rect -8933 -15732 -8899 -15324
rect -8815 -15732 -8781 -15239
rect -8697 -15732 -8663 -15324
rect -8579 -15732 -8545 -15239
rect -8461 -15732 -8427 -15324
rect -8343 -15732 -8309 -15239
rect -8225 -15732 -8191 -15324
rect -8107 -15732 -8073 -15239
rect -7989 -15732 -7955 -15324
rect -7871 -15732 -7837 -15239
rect -14977 -15796 -11347 -15732
rect -14977 -15824 -11495 -15796
rect -11371 -15898 -11299 -15830
rect -11371 -15932 -10991 -15898
rect -11371 -15986 -11299 -15932
rect -11025 -16540 -10991 -15932
rect -9483 -15912 -9411 -15864
rect -8552 -15909 -8450 -15851
rect -7950 -15852 -7874 -15796
rect -7536 -15852 -7185 -14808
rect -9483 -15946 -8973 -15912
rect -9483 -16020 -9411 -15946
rect -10789 -16540 -10755 -16132
rect -10553 -16540 -10519 -16132
rect -10317 -16540 -10283 -16132
rect -10081 -16540 -10047 -16132
rect -9845 -16540 -9811 -16132
rect -9609 -16540 -9575 -16132
rect -9373 -16540 -9339 -16132
rect -9007 -16540 -8973 -15946
rect -8552 -15943 -8073 -15909
rect -8552 -15991 -8450 -15943
rect -8107 -16032 -8073 -15943
rect -7950 -15913 -7185 -15852
rect -7950 -15973 -7874 -15913
rect -8107 -16066 -7899 -16032
rect -8771 -16540 -8737 -16132
rect -8535 -16540 -8501 -16132
rect -8299 -16540 -8265 -16132
rect -7933 -16540 -7899 -16066
rect -7697 -16540 -7663 -16132
rect 7543 -17611 18811 -17278
rect -15041 -18397 -15007 -18393
rect -15047 -18650 -15001 -18397
rect -14845 -18585 -14811 -18393
rect -14851 -18650 -14805 -18585
rect -14649 -18585 -14615 -18393
rect -14425 -18479 -14368 -18415
rect -14568 -18528 -14368 -18479
rect -14655 -18650 -14609 -18585
rect -15047 -18658 -14609 -18650
rect -14568 -18658 -14522 -18528
rect -14425 -18579 -14368 -18528
rect -14204 -18397 -14170 -18393
rect -15251 -18695 -15083 -18665
rect -22640 -19424 -22606 -19180
rect -22444 -19424 -22410 -19180
rect -22248 -19424 -22214 -19180
rect -22640 -19461 -22085 -19424
rect -22122 -19599 -22085 -19461
rect -21680 -19599 -21545 -19589
rect -22122 -19636 -21545 -19599
rect -22122 -19690 -22085 -19636
rect -21680 -19643 -21545 -19636
rect -22738 -19724 -22295 -19690
rect -22122 -19724 -21889 -19690
rect -22738 -20095 -22704 -19724
rect -22542 -19725 -22295 -19724
rect -22640 -20284 -22606 -19787
rect -22542 -20095 -22508 -19725
rect -22330 -19788 -22295 -19725
rect -22428 -20087 -22394 -19788
rect -22428 -20191 -22393 -20087
rect -22330 -20096 -22296 -19788
rect -22232 -20085 -22198 -19788
rect -22232 -20191 -22197 -20085
rect -22119 -20096 -22085 -19724
rect -22428 -20194 -22197 -20191
rect -22021 -20194 -21987 -19788
rect -21923 -20096 -21889 -19724
rect -22428 -20228 -21987 -20194
rect -21608 -20195 -21574 -19888
rect -21510 -20096 -21476 -19180
rect -20641 -19646 -20607 -19302
rect -20445 -19646 -20411 -19302
rect -20032 -19409 -19998 -19301
rect -19836 -19409 -19802 -19301
rect -20150 -19456 -20077 -19443
rect -20250 -19484 -20077 -19456
rect -20272 -19497 -20077 -19484
rect -20272 -19646 -20211 -19497
rect -20150 -19503 -20077 -19497
rect -19640 -19473 -19606 -19301
rect -18292 -19337 -16815 -19224
rect -19640 -19474 -19236 -19473
rect -19640 -19532 -19172 -19474
rect -20641 -19676 -20211 -19646
rect -20641 -19684 -20222 -19676
rect -20032 -19688 -19998 -19532
rect -19934 -19640 -19900 -19532
rect -19836 -19688 -19802 -19532
rect -19738 -19640 -19704 -19532
rect -19640 -19543 -19236 -19532
rect -19123 -19632 -18674 -19614
rect -18292 -19632 -18231 -19337
rect -17565 -19455 -17518 -19337
rect -19599 -19688 -18231 -19632
rect -20172 -19693 -18231 -19688
rect -20172 -19774 -19538 -19693
rect -19006 -19727 -18971 -19693
rect -20739 -20147 -20705 -19839
rect -20641 -20147 -20607 -19839
rect -20543 -20147 -20509 -19839
rect -20445 -20147 -20411 -19839
rect -20347 -20147 -20313 -19839
rect -20642 -20195 -20607 -20147
rect -19928 -20181 -19867 -19774
rect -19599 -19776 -19538 -19774
rect -19103 -20035 -19069 -19727
rect -19005 -20035 -18971 -19727
rect -18907 -20035 -18873 -19727
rect -18809 -20035 -18775 -19727
rect -18711 -20035 -18677 -19727
rect -19135 -20078 -19064 -20077
rect -18723 -20078 -18649 -20072
rect -19135 -20079 -18649 -20078
rect -19361 -20117 -18649 -20079
rect -18292 -20100 -18231 -19693
rect -17558 -19749 -17524 -19455
rect -17460 -19733 -17426 -19441
rect -17369 -19456 -17322 -19337
rect -17667 -19795 -17512 -19783
rect -17704 -19829 -17512 -19795
rect -17667 -19838 -17512 -19829
rect -17466 -19803 -17421 -19733
rect -17362 -19749 -17328 -19456
rect -17127 -19466 -17080 -19337
rect -17120 -19749 -17086 -19466
rect -17022 -19740 -16988 -19441
rect -17026 -19780 -16982 -19740
rect -17026 -19783 -15886 -19780
rect -17466 -19843 -17112 -19803
rect -17074 -19823 -15886 -19783
rect -17802 -19900 -17732 -19898
rect -17397 -19900 -17242 -19891
rect -17802 -19936 -17242 -19900
rect -19361 -20119 -19134 -20117
rect -18723 -20143 -18649 -20117
rect -19188 -20175 -19053 -20167
rect -19208 -20177 -19053 -20175
rect -20317 -20195 -19867 -20181
rect -21793 -20284 -19837 -20195
rect -19599 -20213 -19053 -20177
rect -18536 -20186 -17921 -20100
rect -22738 -20347 -19837 -20284
rect -22738 -20349 -21464 -20347
rect -24032 -20729 -23931 -20556
rect -19522 -20729 -19465 -20213
rect -19208 -20215 -19053 -20213
rect -19188 -20221 -19053 -20215
rect -19005 -20198 -18586 -20190
rect -19005 -20228 -18575 -20198
rect -19005 -20572 -18971 -20228
rect -18809 -20572 -18775 -20228
rect -18636 -20377 -18575 -20228
rect -18396 -20342 -18362 -20186
rect -18298 -20342 -18264 -20234
rect -18200 -20342 -18166 -20186
rect -18102 -20342 -18068 -20234
rect -17802 -20331 -17732 -19936
rect -17397 -19946 -17242 -19936
rect -17155 -19913 -17112 -19843
rect -17155 -19968 -16974 -19913
rect -17155 -19980 -17112 -19968
rect -17562 -20018 -17308 -19982
rect -18514 -20377 -18441 -20371
rect -18636 -20390 -18441 -20377
rect -18614 -20418 -18441 -20390
rect -18514 -20431 -18441 -20418
rect -18004 -20401 -17726 -20331
rect -18396 -20573 -18362 -20465
rect -18200 -20573 -18166 -20465
rect -18004 -20573 -17970 -20401
rect -17562 -20077 -17520 -20018
rect -24032 -20792 -19465 -20729
rect -17558 -20661 -17524 -20077
rect -17350 -20071 -17308 -20018
rect -17253 -20019 -17112 -19980
rect -17347 -20653 -17313 -20071
rect -17253 -20073 -17211 -20019
rect -17351 -20695 -17309 -20653
rect -17249 -20661 -17215 -20073
rect -17151 -20651 -17117 -20053
rect -16940 -20067 -16897 -19823
rect -16714 -19998 -16609 -19926
rect -17153 -20695 -17111 -20651
rect -17351 -20729 -17111 -20695
rect -16939 -20661 -16905 -20067
rect -24032 -20799 -23931 -20792
rect -22583 -21555 -22549 -21211
rect -22387 -21555 -22353 -21211
rect -21974 -21318 -21940 -21210
rect -21778 -21318 -21744 -21210
rect -22092 -21365 -22019 -21352
rect -22192 -21393 -22019 -21365
rect -22214 -21406 -22019 -21393
rect -22214 -21555 -22153 -21406
rect -22092 -21412 -22019 -21406
rect -21582 -21382 -21548 -21210
rect -20810 -21360 -20776 -21116
rect -20614 -21360 -20580 -21116
rect -20418 -21360 -20384 -21116
rect -20985 -21371 -20850 -21363
rect -21345 -21382 -20850 -21371
rect -21582 -21406 -20850 -21382
rect -20810 -21397 -20255 -21360
rect -22583 -21585 -22153 -21555
rect -22583 -21593 -22164 -21585
rect -21974 -21597 -21940 -21441
rect -21876 -21549 -21842 -21441
rect -21778 -21597 -21744 -21441
rect -21680 -21549 -21646 -21441
rect -21582 -21452 -21304 -21406
rect -21004 -21408 -20850 -21406
rect -20985 -21417 -20850 -21408
rect -21100 -21454 -21042 -21446
rect -20649 -21454 -20514 -21445
rect -21126 -21492 -20514 -21454
rect -22114 -21683 -21499 -21597
rect -22681 -22056 -22647 -21748
rect -22583 -22056 -22549 -21748
rect -22485 -22056 -22451 -21748
rect -22387 -22056 -22353 -21748
rect -22289 -22056 -22255 -21748
rect -22584 -22108 -22549 -22056
rect -21870 -22090 -21809 -21683
rect -21411 -21811 -21353 -21674
rect -21197 -21677 -21139 -21577
rect -21100 -21583 -21042 -21492
rect -20649 -21499 -20514 -21492
rect -20461 -21536 -20326 -21523
rect -21002 -21570 -20326 -21536
rect -21002 -21677 -20968 -21570
rect -20461 -21577 -20326 -21570
rect -20292 -21535 -20255 -21397
rect -19850 -21535 -19715 -21525
rect -20292 -21572 -19715 -21535
rect -20292 -21626 -20255 -21572
rect -19850 -21579 -19715 -21572
rect -19680 -21597 -19646 -21116
rect -18979 -21501 -18945 -21293
rect -18783 -21501 -18749 -21293
rect -18587 -21501 -18553 -21293
rect -18006 -21508 -17972 -21164
rect -17810 -21508 -17776 -21164
rect -17397 -21271 -17363 -21163
rect -17201 -21271 -17167 -21163
rect -17515 -21318 -17442 -21305
rect -17615 -21346 -17442 -21318
rect -17637 -21359 -17442 -21346
rect -17637 -21508 -17576 -21359
rect -17515 -21365 -17442 -21359
rect -17005 -21335 -16971 -21163
rect -16703 -21335 -16633 -19998
rect -18189 -21521 -18054 -21515
rect -18209 -21523 -18054 -21521
rect -19271 -21548 -19141 -21531
rect -19097 -21548 -19024 -21535
rect -19271 -21589 -19024 -21548
rect -18416 -21559 -18054 -21523
rect -18006 -21538 -17576 -21508
rect -18006 -21546 -17587 -21538
rect -17397 -21550 -17363 -21394
rect -17299 -21502 -17265 -21394
rect -17201 -21550 -17167 -21394
rect -17103 -21502 -17069 -21394
rect -17005 -21405 -16633 -21335
rect -18209 -21561 -18054 -21559
rect -18189 -21569 -18054 -21561
rect -19271 -21597 -19141 -21589
rect -19097 -21595 -19024 -21589
rect -21197 -21711 -20968 -21677
rect -20908 -21660 -20465 -21626
rect -20292 -21660 -20059 -21626
rect -21197 -21714 -21139 -21711
rect -20908 -22031 -20874 -21660
rect -20712 -21661 -20465 -21660
rect -22259 -22108 -21090 -22090
rect -22701 -22169 -21090 -22108
rect -22260 -22205 -21090 -22169
rect -21205 -22223 -21090 -22205
rect -20810 -22220 -20776 -21723
rect -20712 -22031 -20678 -21661
rect -20500 -21724 -20465 -21661
rect -20598 -22023 -20564 -21724
rect -20598 -22127 -20563 -22023
rect -20500 -22032 -20466 -21724
rect -20402 -22021 -20368 -21724
rect -20402 -22127 -20367 -22021
rect -20289 -22032 -20255 -21660
rect -20598 -22130 -20367 -22127
rect -20191 -22130 -20157 -21724
rect -20093 -22032 -20059 -21660
rect -19680 -21631 -19141 -21597
rect -18684 -21619 -18135 -21617
rect -17724 -21619 -17650 -21593
rect -18684 -21623 -17650 -21619
rect -20598 -22164 -20157 -22130
rect -19778 -22193 -19744 -21824
rect -19680 -22032 -19646 -21631
rect -19271 -21681 -19141 -21631
rect -18979 -21879 -18945 -21623
rect -18881 -21831 -18847 -21623
rect -18783 -21879 -18749 -21623
rect -18685 -21657 -17650 -21623
rect -17537 -21636 -16752 -21550
rect -18685 -21831 -18651 -21657
rect -18136 -21658 -17650 -21657
rect -18136 -21659 -18065 -21658
rect -17724 -21664 -17650 -21658
rect -19119 -21965 -18181 -21879
rect -18267 -22046 -18181 -21965
rect -18104 -22009 -18070 -21701
rect -18006 -22009 -17972 -21701
rect -17908 -22009 -17874 -21701
rect -17810 -22009 -17776 -21701
rect -17712 -22009 -17678 -21701
rect -18007 -22046 -17972 -22009
rect -17293 -22043 -17232 -21636
rect -17682 -22046 -17232 -22043
rect -18267 -22104 -17232 -22046
rect -18267 -22132 -17602 -22104
rect -18231 -22193 -18021 -22132
rect -19979 -22220 -18021 -22193
rect -20908 -22223 -18021 -22220
rect -21205 -22348 -18021 -22223
rect -17099 -22182 -16831 -22132
rect -16069 -22182 -15886 -19823
rect -15258 -18739 -15083 -18695
rect -15047 -18696 -14522 -18658
rect -14210 -18650 -14164 -18397
rect -14008 -18585 -13974 -18393
rect -14014 -18650 -13968 -18585
rect -13594 -18374 -12966 -18340
rect -13812 -18585 -13778 -18393
rect -13594 -18419 -13558 -18374
rect -13818 -18650 -13772 -18585
rect -14210 -18658 -13772 -18650
rect -13717 -18634 -13643 -18466
rect -13593 -18493 -13559 -18419
rect -13717 -18658 -13644 -18634
rect -14414 -18676 -14246 -18665
rect -14449 -18677 -14246 -18676
rect -15258 -19111 -15210 -18739
rect -15139 -18932 -15105 -18773
rect -15047 -18789 -15001 -18696
rect -15041 -18881 -15007 -18789
rect -14943 -18932 -14909 -18773
rect -14851 -18789 -14805 -18696
rect -14655 -18728 -14522 -18696
rect -14845 -18881 -14811 -18789
rect -14747 -18932 -14713 -18773
rect -14655 -18789 -14609 -18728
rect -14486 -18739 -14246 -18677
rect -14210 -18696 -13644 -18658
rect -14649 -18881 -14615 -18789
rect -14486 -18883 -14426 -18739
rect -14302 -18932 -14268 -18773
rect -14210 -18789 -14164 -18696
rect -14204 -18881 -14170 -18789
rect -14106 -18932 -14072 -18773
rect -14014 -18789 -13968 -18696
rect -13818 -18728 -13644 -18696
rect -13599 -18640 -13552 -18493
rect -13495 -18500 -13461 -18408
rect -13398 -18429 -13356 -18374
rect -13496 -18552 -13460 -18500
rect -13397 -18516 -13363 -18429
rect -13299 -18498 -13265 -18408
rect -13204 -18430 -13162 -18374
rect -13299 -18516 -13262 -18498
rect -13201 -18516 -13167 -18430
rect -13103 -18498 -13069 -18408
rect -13008 -18425 -12966 -18374
rect -13298 -18552 -13262 -18516
rect -13104 -18552 -13068 -18498
rect -13005 -18516 -12971 -18425
rect -12907 -18508 -12873 -18408
rect -12910 -18552 -12868 -18508
rect -13496 -18586 -12868 -18552
rect -13599 -18714 -13427 -18640
rect -13043 -18693 -12868 -18586
rect -12341 -18397 -12307 -18393
rect -12347 -18650 -12301 -18397
rect -12145 -18585 -12111 -18393
rect -12151 -18650 -12105 -18585
rect -11949 -18585 -11915 -18393
rect -11725 -18467 -11668 -18415
rect -11873 -18529 -11668 -18467
rect -11955 -18650 -11909 -18585
rect -12347 -18658 -11909 -18650
rect -11873 -18658 -11811 -18529
rect -11725 -18579 -11668 -18529
rect -11504 -18397 -11470 -18393
rect -12551 -18672 -12383 -18665
rect -14008 -18881 -13974 -18789
rect -13910 -18932 -13876 -18773
rect -13818 -18789 -13772 -18728
rect -13812 -18881 -13778 -18789
rect -13599 -18849 -13552 -18714
rect -13043 -18753 -12777 -18693
rect -12573 -18732 -12383 -18672
rect -12551 -18739 -12383 -18732
rect -12347 -18696 -11811 -18658
rect -11510 -18650 -11464 -18397
rect -11308 -18585 -11274 -18393
rect -11314 -18650 -11268 -18585
rect -10894 -18374 -10266 -18340
rect -11112 -18585 -11078 -18393
rect -10894 -18419 -10858 -18374
rect -11118 -18650 -11072 -18585
rect -11510 -18658 -11072 -18650
rect -11017 -18634 -10943 -18466
rect -10893 -18493 -10859 -18419
rect -11017 -18658 -10944 -18634
rect -11714 -18676 -11546 -18665
rect -13499 -18787 -12868 -18753
rect -13499 -18828 -13458 -18787
rect -13593 -18919 -13559 -18849
rect -15148 -19000 -13777 -18932
rect -13598 -18977 -13554 -18919
rect -13495 -18931 -13461 -18828
rect -13397 -18908 -13363 -18823
rect -13301 -18836 -13260 -18787
rect -13402 -18977 -13358 -18908
rect -13299 -18931 -13265 -18836
rect -13201 -18908 -13167 -18823
rect -13107 -18836 -13066 -18787
rect -12910 -18794 -12868 -18787
rect -13206 -18977 -13162 -18908
rect -13103 -18931 -13069 -18836
rect -13005 -18919 -12971 -18823
rect -12910 -18837 -12869 -18794
rect -13009 -18977 -12965 -18919
rect -12907 -18931 -12873 -18837
rect -12439 -18932 -12405 -18773
rect -12347 -18789 -12301 -18696
rect -12341 -18881 -12307 -18789
rect -12243 -18932 -12209 -18773
rect -12151 -18789 -12105 -18696
rect -11955 -18728 -11811 -18696
rect -12145 -18881 -12111 -18789
rect -12047 -18932 -12013 -18773
rect -11955 -18789 -11909 -18728
rect -11774 -18739 -11546 -18676
rect -11510 -18696 -10944 -18658
rect -11949 -18881 -11915 -18789
rect -11774 -18898 -11714 -18739
rect -11602 -18932 -11568 -18773
rect -11510 -18789 -11464 -18696
rect -11504 -18881 -11470 -18789
rect -11406 -18932 -11372 -18773
rect -11314 -18789 -11268 -18696
rect -11118 -18728 -10944 -18696
rect -10899 -18640 -10852 -18493
rect -10795 -18500 -10761 -18408
rect -10698 -18429 -10656 -18374
rect -10796 -18552 -10760 -18500
rect -10697 -18516 -10663 -18429
rect -10599 -18498 -10565 -18408
rect -10504 -18430 -10462 -18374
rect -10599 -18516 -10562 -18498
rect -10501 -18516 -10467 -18430
rect -10403 -18498 -10369 -18408
rect -10308 -18425 -10266 -18374
rect -10598 -18552 -10562 -18516
rect -10404 -18552 -10368 -18498
rect -10305 -18516 -10271 -18425
rect -10207 -18508 -10173 -18408
rect -10210 -18552 -10168 -18508
rect -10796 -18586 -10168 -18552
rect -10899 -18714 -10727 -18640
rect -10343 -18695 -10168 -18586
rect -11308 -18881 -11274 -18789
rect -11210 -18932 -11176 -18773
rect -11118 -18789 -11072 -18728
rect -11112 -18881 -11078 -18789
rect -10899 -18849 -10852 -18714
rect -10343 -18753 -10093 -18695
rect -10799 -18755 -10093 -18753
rect -10799 -18787 -10168 -18755
rect -10799 -18828 -10758 -18787
rect -10893 -18919 -10859 -18849
rect -14900 -19040 -14789 -19000
rect -14911 -19048 -14774 -19040
rect -14089 -19048 -13978 -19000
rect -13598 -19011 -12965 -18977
rect -12448 -18934 -11914 -18932
rect -11611 -18934 -11077 -18932
rect -12448 -19000 -11077 -18934
rect -10898 -18977 -10854 -18919
rect -10795 -18931 -10761 -18828
rect -10697 -18908 -10663 -18823
rect -10601 -18836 -10560 -18787
rect -10702 -18977 -10658 -18908
rect -10599 -18931 -10565 -18836
rect -10501 -18908 -10467 -18823
rect -10407 -18836 -10366 -18787
rect -10210 -18794 -10168 -18787
rect -10506 -18977 -10462 -18908
rect -10403 -18931 -10369 -18836
rect -10305 -18919 -10271 -18823
rect -10210 -18837 -10169 -18794
rect -10309 -18977 -10265 -18919
rect -10207 -18931 -10173 -18837
rect -12291 -19046 -12180 -19000
rect -12108 -19002 -11588 -19000
rect -12314 -19048 -12177 -19046
rect -11413 -19048 -11302 -19000
rect -10898 -19011 -10265 -18977
rect -8875 -18997 -8841 -18403
rect -8669 -18369 -8429 -18335
rect -8669 -18413 -8627 -18369
rect -9676 -19048 -9544 -19046
rect -14928 -19087 -9543 -19048
rect -14911 -19100 -14774 -19087
rect -12314 -19106 -12177 -19087
rect -9676 -19106 -9544 -19087
rect -15259 -19248 -15199 -19111
rect -12749 -19140 -12612 -19129
rect -11803 -19140 -11671 -19130
rect -14928 -19179 -9198 -19140
rect -12749 -19189 -12612 -19179
rect -11803 -19190 -11671 -19179
rect -14522 -19226 -14390 -19218
rect -9999 -19226 -9867 -19216
rect -15258 -19606 -15210 -19248
rect -14928 -19265 -9867 -19226
rect -9237 -19241 -9198 -19179
rect -8883 -19241 -8840 -18997
rect -8663 -19011 -8629 -18413
rect -8565 -18991 -8531 -18403
rect -8471 -18411 -8429 -18369
rect -8569 -19045 -8527 -18991
rect -8467 -18993 -8433 -18411
rect -8668 -19084 -8527 -19045
rect -8472 -19046 -8430 -18993
rect -8256 -18987 -8222 -18403
rect -8260 -19046 -8218 -18987
rect -7445 -18495 -6717 -18461
rect -7445 -18807 -7411 -18495
rect -7347 -18843 -7313 -18599
rect -7249 -18807 -7215 -18495
rect -7129 -18564 -6787 -18530
rect -7129 -18807 -7095 -18564
rect -7031 -18843 -6997 -18599
rect -6933 -18807 -6899 -18564
rect -7556 -18877 -6882 -18843
rect -8472 -19082 -8218 -19046
rect -8668 -19096 -8625 -19084
rect -8806 -19151 -8625 -19096
rect -8668 -19221 -8625 -19151
rect -8538 -19128 -8383 -19118
rect -7998 -19128 -7866 -19057
rect -8538 -19164 -7866 -19128
rect -8538 -19173 -8383 -19164
rect -14522 -19278 -14390 -19265
rect -9999 -19276 -9867 -19265
rect -9241 -19281 -8706 -19241
rect -8668 -19261 -8314 -19221
rect -9241 -19284 -8754 -19281
rect -15140 -19380 -14606 -19312
rect -14209 -19335 -13576 -19301
rect -15139 -19523 -15105 -19431
rect -15145 -19584 -15099 -19523
rect -15041 -19539 -15007 -19380
rect -14943 -19523 -14909 -19431
rect -15175 -19606 -15099 -19584
rect -15258 -19616 -15099 -19606
rect -14949 -19616 -14903 -19523
rect -14845 -19539 -14811 -19380
rect -14747 -19523 -14713 -19431
rect -14753 -19616 -14707 -19523
rect -14649 -19539 -14615 -19380
rect -14301 -19475 -14267 -19381
rect -14209 -19393 -14165 -19335
rect -14305 -19518 -14264 -19475
rect -14203 -19489 -14169 -19393
rect -14105 -19476 -14071 -19381
rect -14012 -19404 -13968 -19335
rect -14306 -19525 -14264 -19518
rect -14108 -19525 -14067 -19476
rect -14007 -19489 -13973 -19404
rect -13909 -19476 -13875 -19381
rect -13816 -19404 -13772 -19335
rect -13914 -19525 -13873 -19476
rect -13811 -19489 -13777 -19404
rect -13713 -19484 -13679 -19381
rect -13620 -19393 -13576 -19335
rect -13397 -19380 -11906 -19312
rect -11509 -19335 -10876 -19301
rect -13615 -19463 -13581 -19393
rect -13716 -19525 -13675 -19484
rect -14306 -19559 -13675 -19525
rect -15258 -19643 -14707 -19616
rect -15257 -19645 -14707 -19643
rect -15175 -19654 -14707 -19645
rect -14671 -19588 -14503 -19573
rect -14306 -19588 -14131 -19559
rect -14671 -19641 -14131 -19588
rect -13622 -19598 -13575 -19463
rect -13396 -19523 -13362 -19431
rect -13402 -19584 -13356 -19523
rect -13298 -19539 -13264 -19380
rect -13200 -19523 -13166 -19431
rect -14671 -19647 -14503 -19641
rect -15145 -19662 -14707 -19654
rect -15145 -19727 -15099 -19662
rect -15139 -19919 -15105 -19727
rect -14949 -19727 -14903 -19662
rect -14943 -19919 -14909 -19727
rect -14753 -19915 -14707 -19662
rect -14747 -19919 -14713 -19915
rect -14306 -19726 -14131 -19641
rect -13747 -19672 -13575 -19598
rect -14306 -19760 -13678 -19726
rect -14306 -19804 -14264 -19760
rect -14301 -19904 -14267 -19804
rect -14203 -19887 -14169 -19796
rect -14106 -19814 -14070 -19760
rect -13912 -19796 -13876 -19760
rect -14208 -19938 -14166 -19887
rect -14105 -19904 -14071 -19814
rect -14007 -19882 -13973 -19796
rect -13912 -19814 -13875 -19796
rect -14012 -19938 -13970 -19882
rect -13909 -19904 -13875 -19814
rect -13811 -19883 -13777 -19796
rect -13714 -19812 -13678 -19760
rect -13818 -19938 -13776 -19883
rect -13713 -19904 -13679 -19812
rect -13622 -19819 -13575 -19672
rect -13530 -19616 -13356 -19584
rect -13206 -19616 -13160 -19523
rect -13102 -19539 -13068 -19380
rect -13004 -19523 -12970 -19431
rect -13010 -19616 -12964 -19523
rect -12906 -19539 -12872 -19380
rect -13530 -19654 -12964 -19616
rect -12928 -19578 -12760 -19573
rect -12700 -19578 -12640 -19505
rect -12928 -19636 -12640 -19578
rect -12585 -19595 -12525 -19480
rect -12439 -19523 -12405 -19431
rect -12445 -19584 -12399 -19523
rect -12341 -19539 -12307 -19380
rect -12243 -19523 -12209 -19431
rect -12475 -19595 -12399 -19584
rect -12928 -19647 -12760 -19636
rect -12700 -19637 -12640 -19636
rect -12590 -19616 -12399 -19595
rect -12249 -19616 -12203 -19523
rect -12145 -19539 -12111 -19380
rect -12047 -19523 -12013 -19431
rect -12053 -19616 -12007 -19523
rect -11949 -19539 -11915 -19380
rect -11604 -19475 -11558 -19353
rect -11509 -19393 -11465 -19335
rect -11605 -19485 -11558 -19475
rect -11605 -19518 -11564 -19485
rect -11503 -19489 -11469 -19393
rect -11405 -19476 -11371 -19381
rect -11312 -19404 -11268 -19335
rect -11606 -19525 -11564 -19518
rect -11408 -19525 -11367 -19476
rect -11307 -19489 -11273 -19404
rect -11209 -19476 -11175 -19381
rect -11116 -19404 -11072 -19335
rect -11214 -19525 -11173 -19476
rect -11111 -19489 -11077 -19404
rect -11013 -19484 -10979 -19381
rect -10920 -19393 -10876 -19335
rect -10697 -19380 -9281 -19312
rect -10915 -19463 -10881 -19393
rect -11016 -19525 -10975 -19484
rect -11606 -19559 -10975 -19525
rect -12590 -19640 -12007 -19616
rect -13530 -19678 -13457 -19654
rect -13615 -19893 -13581 -19819
rect -13531 -19846 -13457 -19678
rect -13402 -19662 -12964 -19654
rect -13402 -19727 -13356 -19662
rect -13616 -19938 -13580 -19893
rect -13396 -19919 -13362 -19727
rect -14208 -19972 -13580 -19938
rect -13206 -19727 -13160 -19662
rect -13200 -19919 -13166 -19727
rect -13010 -19915 -12964 -19662
rect -13004 -19919 -12970 -19915
rect -12806 -19774 -12749 -19733
rect -12590 -19774 -12545 -19640
rect -12475 -19654 -12007 -19640
rect -11971 -19581 -11803 -19573
rect -11606 -19581 -11431 -19559
rect -11971 -19638 -11431 -19581
rect -10922 -19598 -10875 -19463
rect -10696 -19523 -10662 -19431
rect -10702 -19584 -10656 -19523
rect -10598 -19539 -10564 -19380
rect -10500 -19523 -10466 -19431
rect -11971 -19647 -11803 -19638
rect -12445 -19662 -12007 -19654
rect -12445 -19727 -12399 -19662
rect -12806 -19819 -12545 -19774
rect -12806 -19897 -12749 -19819
rect -12439 -19919 -12405 -19727
rect -12249 -19727 -12203 -19662
rect -12243 -19919 -12209 -19727
rect -12053 -19915 -12007 -19662
rect -12047 -19919 -12013 -19915
rect -11606 -19726 -11431 -19638
rect -11047 -19672 -10875 -19598
rect -11606 -19760 -10978 -19726
rect -11606 -19804 -11564 -19760
rect -11601 -19904 -11567 -19804
rect -11503 -19887 -11469 -19796
rect -11406 -19814 -11370 -19760
rect -11212 -19796 -11176 -19760
rect -11508 -19938 -11466 -19887
rect -11405 -19904 -11371 -19814
rect -11307 -19882 -11273 -19796
rect -11212 -19814 -11175 -19796
rect -11312 -19938 -11270 -19882
rect -11209 -19904 -11175 -19814
rect -11111 -19883 -11077 -19796
rect -11014 -19812 -10978 -19760
rect -11118 -19938 -11076 -19883
rect -11013 -19904 -10979 -19812
rect -10922 -19819 -10875 -19672
rect -10830 -19616 -10656 -19584
rect -10506 -19616 -10460 -19523
rect -10402 -19539 -10368 -19380
rect -10304 -19523 -10270 -19431
rect -10310 -19616 -10264 -19523
rect -10206 -19539 -10172 -19380
rect -10830 -19654 -10264 -19616
rect -10228 -19578 -10060 -19573
rect -10228 -19590 -10025 -19578
rect -9968 -19590 -9908 -19504
rect -9814 -19523 -9780 -19431
rect -9820 -19584 -9774 -19523
rect -9716 -19539 -9682 -19380
rect -9618 -19523 -9584 -19431
rect -9850 -19590 -9774 -19584
rect -10228 -19616 -9774 -19590
rect -9624 -19616 -9578 -19523
rect -9520 -19539 -9486 -19380
rect -9422 -19523 -9388 -19431
rect -9428 -19616 -9382 -19523
rect -9324 -19539 -9290 -19380
rect -9237 -19573 -9198 -19284
rect -8798 -19324 -8754 -19284
rect -10228 -19632 -9382 -19616
rect -10228 -19636 -10025 -19632
rect -9968 -19636 -9908 -19632
rect -10228 -19647 -10060 -19636
rect -9850 -19654 -9382 -19632
rect -9346 -19647 -9178 -19573
rect -8792 -19623 -8758 -19324
rect -8694 -19598 -8660 -19315
rect -10830 -19678 -10757 -19654
rect -10915 -19893 -10881 -19819
rect -10831 -19846 -10757 -19678
rect -10702 -19662 -10264 -19654
rect -10702 -19727 -10656 -19662
rect -10916 -19938 -10880 -19893
rect -10696 -19919 -10662 -19727
rect -11508 -19972 -10880 -19938
rect -10506 -19727 -10460 -19662
rect -10500 -19919 -10466 -19727
rect -10310 -19915 -10264 -19662
rect -9820 -19662 -9382 -19654
rect -10304 -19919 -10270 -19915
rect -9820 -19727 -9774 -19662
rect -10106 -19897 -10049 -19733
rect -9814 -19919 -9780 -19727
rect -9624 -19727 -9578 -19662
rect -9618 -19919 -9584 -19727
rect -9428 -19915 -9382 -19662
rect -9422 -19919 -9388 -19915
rect -9124 -19728 -8846 -19727
rect -8700 -19728 -8653 -19598
rect -8452 -19608 -8418 -19315
rect -8359 -19331 -8314 -19261
rect -8268 -19235 -8113 -19226
rect -8268 -19269 -7706 -19235
rect -8268 -19281 -8113 -19269
rect -8458 -19728 -8411 -19608
rect -8354 -19623 -8320 -19331
rect -8256 -19609 -8222 -19315
rect -8262 -19728 -8215 -19609
rect -9124 -19810 -8133 -19728
rect -17099 -22365 -15886 -22182
rect -13303 -20313 -11826 -20200
rect -14134 -20608 -13685 -20590
rect -13303 -20608 -13242 -20313
rect -12576 -20431 -12529 -20313
rect -14134 -20651 -13242 -20608
rect -14017 -20703 -13982 -20651
rect -13692 -20669 -13242 -20651
rect -14114 -21011 -14080 -20703
rect -14016 -21011 -13982 -20703
rect -13918 -21011 -13884 -20703
rect -13820 -21011 -13786 -20703
rect -13722 -21011 -13688 -20703
rect -13303 -21076 -13242 -20669
rect -12569 -20725 -12535 -20431
rect -12471 -20709 -12437 -20417
rect -12380 -20432 -12333 -20313
rect -12678 -20771 -12523 -20759
rect -12715 -20805 -12523 -20771
rect -12678 -20814 -12523 -20805
rect -12477 -20779 -12432 -20709
rect -12373 -20725 -12339 -20432
rect -12138 -20442 -12091 -20313
rect -12131 -20725 -12097 -20442
rect -12033 -20716 -11999 -20417
rect -12037 -20756 -11993 -20716
rect -12037 -20759 -8957 -20756
rect -12477 -20819 -12123 -20779
rect -12085 -20799 -8957 -20759
rect -12813 -20876 -12743 -20874
rect -12408 -20876 -12253 -20867
rect -12813 -20912 -12253 -20876
rect -14659 -21153 -14473 -21096
rect -14199 -21151 -14064 -21143
rect -14219 -21153 -14064 -21151
rect -14659 -21189 -14064 -21153
rect -13547 -21162 -12932 -21076
rect -14659 -21250 -14473 -21189
rect -14219 -21191 -14064 -21189
rect -14199 -21197 -14064 -21191
rect -14016 -21174 -13597 -21166
rect -14016 -21204 -13586 -21174
rect -14016 -21548 -13982 -21204
rect -13820 -21548 -13786 -21204
rect -13647 -21353 -13586 -21204
rect -13407 -21318 -13373 -21162
rect -13309 -21318 -13275 -21210
rect -13211 -21318 -13177 -21162
rect -13113 -21318 -13079 -21210
rect -12813 -21307 -12743 -20912
rect -12408 -20922 -12253 -20912
rect -12166 -20889 -12123 -20819
rect -12166 -20944 -11985 -20889
rect -12166 -20956 -12123 -20944
rect -12573 -20994 -12319 -20958
rect -13525 -21353 -13452 -21347
rect -13647 -21366 -13452 -21353
rect -13625 -21394 -13452 -21366
rect -13525 -21407 -13452 -21394
rect -13015 -21377 -12737 -21307
rect -13407 -21549 -13373 -21441
rect -13211 -21549 -13177 -21441
rect -13015 -21549 -12981 -21377
rect -12573 -21053 -12531 -20994
rect -12569 -21637 -12535 -21053
rect -12361 -21047 -12319 -20994
rect -12264 -20995 -12123 -20956
rect -12358 -21629 -12324 -21047
rect -12264 -21049 -12222 -20995
rect -12362 -21671 -12320 -21629
rect -12260 -21637 -12226 -21049
rect -12162 -21627 -12128 -21029
rect -11951 -21043 -11908 -20799
rect -9133 -20878 -8957 -20799
rect -11725 -20974 -11620 -20902
rect -12164 -21671 -12122 -21627
rect -12362 -21705 -12122 -21671
rect -11950 -21637 -11916 -21043
rect -17099 -22397 -16831 -22365
rect -19485 -22739 -15947 -22533
rect -16155 -22741 -15947 -22739
rect -25664 -22999 -25039 -22779
rect -17094 -22999 -16826 -22952
rect -25664 -23185 -16826 -22999
rect -13990 -22477 -13956 -22269
rect -13794 -22477 -13760 -22269
rect -13598 -22477 -13564 -22269
rect -13017 -22484 -12983 -22140
rect -12821 -22484 -12787 -22140
rect -12408 -22247 -12374 -22139
rect -12212 -22247 -12178 -22139
rect -12526 -22294 -12453 -22281
rect -12626 -22322 -12453 -22294
rect -12648 -22335 -12453 -22322
rect -12648 -22484 -12587 -22335
rect -12526 -22341 -12453 -22335
rect -12016 -22311 -11982 -22139
rect -11714 -22311 -11644 -20974
rect -7740 -21528 -7706 -19269
rect -7556 -20417 -7522 -18877
rect -7446 -19011 -7307 -18957
rect -6916 -18992 -6882 -18877
rect -6821 -18916 -6787 -18564
rect -6751 -18842 -6717 -18495
rect -6571 -18842 -6537 -18599
rect -6751 -18876 -6537 -18842
rect -6375 -18916 -6341 -18599
rect -6065 -18792 -6031 -18599
rect -6821 -18950 -6341 -18916
rect -6288 -18967 -6149 -18913
rect -6916 -19026 -6770 -18992
rect -7447 -19129 -7116 -19092
rect -7064 -19115 -6925 -19061
rect -6804 -19088 -6770 -19026
rect -6697 -19041 -6558 -18987
rect -6804 -19122 -6243 -19088
rect -7447 -19212 -7410 -19129
rect -7153 -19153 -7116 -19129
rect -7153 -19190 -6997 -19153
rect -7445 -19401 -7411 -19212
rect -7449 -19524 -7410 -19401
rect -7347 -19450 -7313 -19205
rect -7034 -19211 -6997 -19190
rect -7031 -19413 -6997 -19211
rect -6935 -19214 -6635 -19175
rect -6933 -19413 -6899 -19214
rect -6669 -19413 -6635 -19214
rect -6571 -19413 -6537 -19122
rect -6375 -19396 -6341 -19205
rect -6375 -19450 -6339 -19396
rect -6277 -19413 -6243 -19122
rect -6070 -19131 -6027 -18792
rect -5756 -18790 -5722 -18599
rect -5760 -18987 -5717 -18790
rect -5673 -18973 -5534 -18919
rect -5860 -19033 -5717 -18987
rect -5986 -19121 -5847 -19067
rect -6166 -19177 -6027 -19131
rect -6070 -19222 -6027 -19177
rect -6065 -19413 -6031 -19222
rect -5967 -19406 -5933 -19205
rect -5760 -19224 -5717 -19033
rect -7347 -19486 -6339 -19450
rect -5972 -19490 -5929 -19406
rect -5756 -19413 -5722 -19224
rect -5658 -19404 -5624 -19205
rect -4945 -18495 -4217 -18461
rect -4945 -18807 -4911 -18495
rect -4847 -18843 -4813 -18599
rect -4749 -18807 -4715 -18495
rect -4629 -18564 -4287 -18530
rect -4629 -18807 -4595 -18564
rect -4531 -18843 -4497 -18599
rect -4433 -18807 -4399 -18564
rect -5113 -18877 -4382 -18843
rect -5113 -19240 -5079 -18877
rect -4946 -19011 -4807 -18957
rect -4416 -18992 -4382 -18877
rect -4321 -18916 -4287 -18564
rect -4251 -18842 -4217 -18495
rect -4071 -18842 -4037 -18599
rect -4251 -18876 -4037 -18842
rect -3875 -18916 -3841 -18599
rect -3565 -18792 -3531 -18599
rect -4321 -18950 -3841 -18916
rect -3788 -18967 -3649 -18913
rect -4416 -19026 -4270 -18992
rect -4947 -19129 -4616 -19092
rect -4304 -19088 -4270 -19026
rect -4197 -19041 -4058 -18987
rect -4304 -19122 -3743 -19088
rect -4947 -19212 -4910 -19129
rect -4653 -19153 -4616 -19129
rect -4653 -19190 -4497 -19153
rect -5119 -19376 -5073 -19240
rect -4945 -19401 -4911 -19212
rect -5663 -19489 -5620 -19404
rect -4949 -19489 -4910 -19401
rect -4847 -19450 -4813 -19205
rect -4534 -19211 -4497 -19190
rect -4531 -19413 -4497 -19211
rect -4435 -19214 -4135 -19175
rect -4433 -19413 -4399 -19214
rect -4169 -19413 -4135 -19214
rect -4071 -19413 -4037 -19122
rect -3875 -19396 -3841 -19205
rect -3875 -19450 -3839 -19396
rect -3777 -19413 -3743 -19122
rect -3570 -19131 -3527 -18792
rect -3256 -18790 -3222 -18599
rect -3260 -18987 -3217 -18790
rect -3173 -18973 -3034 -18919
rect -3360 -19033 -3217 -18987
rect -3666 -19177 -3527 -19131
rect -3570 -19222 -3527 -19177
rect -3565 -19413 -3531 -19222
rect -3467 -19406 -3433 -19205
rect -3260 -19224 -3217 -19033
rect -4847 -19486 -3839 -19450
rect -5737 -19490 -4910 -19489
rect -3472 -19490 -3429 -19406
rect -3256 -19413 -3222 -19224
rect -3158 -19404 -3124 -19205
rect -2445 -18495 -1717 -18461
rect -2445 -18807 -2411 -18495
rect -2347 -18843 -2313 -18599
rect -2249 -18807 -2215 -18495
rect -2129 -18564 -1787 -18530
rect -2129 -18807 -2095 -18564
rect -2031 -18843 -1997 -18599
rect -1933 -18807 -1899 -18564
rect -2565 -18877 -1882 -18843
rect -2565 -19244 -2531 -18877
rect -2446 -19011 -2307 -18957
rect -1916 -18992 -1882 -18877
rect -1821 -18916 -1787 -18564
rect -1751 -18842 -1717 -18495
rect -1571 -18842 -1537 -18599
rect -1751 -18876 -1537 -18842
rect -1375 -18916 -1341 -18599
rect -1065 -18792 -1031 -18599
rect -1821 -18950 -1341 -18916
rect -1288 -18967 -1149 -18913
rect -1916 -19026 -1770 -18992
rect -2447 -19129 -2116 -19092
rect -1804 -19088 -1770 -19026
rect -1697 -19041 -1558 -18987
rect -1804 -19122 -1243 -19088
rect -2447 -19212 -2410 -19129
rect -2153 -19153 -2116 -19129
rect -2153 -19190 -1997 -19153
rect -2571 -19380 -2525 -19244
rect -2445 -19401 -2411 -19212
rect -3163 -19490 -3120 -19404
rect -6248 -19524 -4910 -19490
rect -3748 -19524 -3116 -19490
rect -2449 -19524 -2410 -19401
rect -2347 -19450 -2313 -19205
rect -2034 -19211 -1997 -19190
rect -2031 -19413 -1997 -19211
rect -1935 -19214 -1635 -19175
rect -1933 -19413 -1899 -19214
rect -1669 -19413 -1635 -19214
rect -1571 -19413 -1537 -19122
rect -1375 -19396 -1341 -19205
rect -1375 -19450 -1339 -19396
rect -1277 -19413 -1243 -19122
rect -1070 -19131 -1027 -18792
rect -756 -18790 -722 -18599
rect -760 -18987 -717 -18790
rect -673 -18973 -534 -18919
rect -860 -19033 -717 -18987
rect -1166 -19177 -1027 -19131
rect -1070 -19222 -1027 -19177
rect -1065 -19413 -1031 -19222
rect -967 -19406 -933 -19205
rect -760 -19224 -717 -19033
rect -2347 -19486 -1339 -19450
rect -972 -19490 -929 -19406
rect -756 -19413 -722 -19224
rect -658 -19404 -624 -19205
rect 55 -18495 783 -18461
rect 55 -18807 89 -18495
rect -85 -18843 -51 -18842
rect 153 -18843 187 -18599
rect 251 -18807 285 -18495
rect 371 -18564 713 -18530
rect 371 -18807 405 -18564
rect 469 -18843 503 -18599
rect 567 -18807 601 -18564
rect -85 -18877 618 -18843
rect -85 -19244 -51 -18877
rect 54 -19011 193 -18957
rect 584 -18992 618 -18877
rect 679 -18916 713 -18564
rect 749 -18842 783 -18495
rect 929 -18842 963 -18599
rect 749 -18876 963 -18842
rect 1125 -18916 1159 -18599
rect 1435 -18792 1469 -18599
rect 679 -18950 1159 -18916
rect 1212 -18967 1351 -18913
rect 584 -19026 730 -18992
rect 53 -19129 384 -19092
rect 696 -19088 730 -19026
rect 803 -19041 942 -18987
rect 696 -19122 1257 -19088
rect 53 -19212 90 -19129
rect 347 -19153 384 -19129
rect 347 -19190 503 -19153
rect -91 -19380 -45 -19244
rect 55 -19401 89 -19212
rect -663 -19490 -620 -19404
rect -1248 -19524 -616 -19490
rect 51 -19524 90 -19401
rect 153 -19450 187 -19205
rect 466 -19211 503 -19190
rect 469 -19413 503 -19211
rect 565 -19214 865 -19175
rect 567 -19413 601 -19214
rect 831 -19413 865 -19214
rect 929 -19413 963 -19122
rect 1125 -19396 1159 -19205
rect 1125 -19450 1161 -19396
rect 1223 -19413 1257 -19122
rect 1430 -19131 1473 -18792
rect 1744 -18790 1778 -18599
rect 2555 -18495 3283 -18461
rect 1740 -18987 1783 -18790
rect 2555 -18807 2589 -18495
rect 2653 -18843 2687 -18599
rect 2751 -18807 2785 -18495
rect 2871 -18564 3213 -18530
rect 2871 -18807 2905 -18564
rect 2969 -18843 3003 -18599
rect 3067 -18807 3101 -18564
rect 2331 -18877 3118 -18843
rect 1827 -18973 1966 -18919
rect 1640 -19033 1783 -18987
rect 1334 -19177 1473 -19131
rect 1430 -19222 1473 -19177
rect 1435 -19413 1469 -19222
rect 1533 -19406 1567 -19205
rect 1740 -19224 1783 -19033
rect 153 -19486 1161 -19450
rect 1528 -19490 1571 -19406
rect 1744 -19413 1778 -19224
rect 1842 -19404 1876 -19205
rect 2331 -19243 2365 -18877
rect 2554 -19011 2693 -18957
rect 3084 -18992 3118 -18877
rect 3179 -18916 3213 -18564
rect 3249 -18842 3283 -18495
rect 3429 -18842 3463 -18599
rect 3249 -18876 3463 -18842
rect 3625 -18916 3659 -18599
rect 3935 -18792 3969 -18599
rect 3179 -18950 3659 -18916
rect 3712 -18967 3851 -18913
rect 3084 -19026 3230 -18992
rect 2553 -19129 2884 -19092
rect 3196 -19088 3230 -19026
rect 3303 -19041 3442 -18987
rect 3196 -19122 3757 -19088
rect 2553 -19212 2590 -19129
rect 2847 -19153 2884 -19129
rect 2847 -19190 3003 -19153
rect 2331 -19244 2366 -19243
rect 2326 -19380 2372 -19244
rect 2555 -19401 2589 -19212
rect 1837 -19490 1880 -19404
rect 1252 -19524 1884 -19490
rect 2551 -19524 2590 -19401
rect 2653 -19450 2687 -19205
rect 2966 -19211 3003 -19190
rect 2969 -19413 3003 -19211
rect 3065 -19214 3365 -19175
rect 3067 -19413 3101 -19214
rect 3331 -19413 3365 -19214
rect 3429 -19413 3463 -19122
rect 3625 -19396 3659 -19205
rect 3625 -19450 3661 -19396
rect 3723 -19413 3757 -19122
rect 3930 -19131 3973 -18792
rect 4244 -18790 4278 -18599
rect 5555 -18495 6283 -18461
rect 4240 -18987 4283 -18790
rect 5555 -18807 5589 -18495
rect 5653 -18843 5687 -18599
rect 5751 -18807 5785 -18495
rect 5871 -18564 6213 -18530
rect 5871 -18807 5905 -18564
rect 5969 -18843 6003 -18599
rect 6067 -18807 6101 -18564
rect 5237 -18877 6118 -18843
rect 4327 -18973 4466 -18919
rect 4140 -19033 4283 -18987
rect 3834 -19177 3973 -19131
rect 3930 -19222 3973 -19177
rect 3935 -19413 3969 -19222
rect 4033 -19406 4067 -19205
rect 4240 -19224 4283 -19033
rect 2653 -19486 3661 -19450
rect 4028 -19490 4071 -19406
rect 4244 -19413 4278 -19224
rect 4342 -19404 4376 -19205
rect 5237 -19244 5271 -18877
rect 5554 -19011 5693 -18957
rect 6084 -18992 6118 -18877
rect 6179 -18916 6213 -18564
rect 6249 -18842 6283 -18495
rect 6429 -18842 6463 -18599
rect 6249 -18876 6463 -18842
rect 6625 -18916 6659 -18599
rect 6935 -18792 6969 -18599
rect 6179 -18950 6659 -18916
rect 6712 -18967 6851 -18913
rect 6084 -19026 6230 -18992
rect 5553 -19129 5884 -19092
rect 6196 -19088 6230 -19026
rect 6303 -19041 6442 -18987
rect 6196 -19122 6757 -19088
rect 5553 -19212 5590 -19129
rect 5847 -19153 5884 -19129
rect 5847 -19190 6003 -19153
rect 5231 -19380 5277 -19244
rect 5555 -19401 5589 -19212
rect 4337 -19490 4380 -19404
rect 3752 -19524 4384 -19490
rect 5551 -19524 5590 -19401
rect 5653 -19450 5687 -19205
rect 5966 -19211 6003 -19190
rect 5969 -19413 6003 -19211
rect 6065 -19214 6365 -19175
rect 6067 -19413 6101 -19214
rect 6331 -19413 6365 -19214
rect 6429 -19413 6463 -19122
rect 6625 -19396 6659 -19205
rect 6625 -19450 6661 -19396
rect 6723 -19413 6757 -19122
rect 6930 -19131 6973 -18792
rect 7244 -18790 7278 -18599
rect 7240 -18987 7283 -18790
rect 7327 -18973 7466 -18919
rect 7140 -19033 7283 -18987
rect 6834 -19177 6973 -19131
rect 6930 -19222 6973 -19177
rect 6935 -19413 6969 -19222
rect 7033 -19406 7067 -19205
rect 7240 -19224 7283 -19033
rect 5653 -19486 6661 -19450
rect 7028 -19472 7071 -19406
rect 7244 -19413 7278 -19224
rect 7342 -19404 7376 -19205
rect 7337 -19472 7380 -19404
rect 7543 -19472 7804 -17611
rect 16158 -17935 16355 -17754
rect 15814 -18410 16095 -18201
rect 8028 -18613 8228 -18579
rect 15454 -18613 15816 -18567
rect 8028 -18785 15816 -18613
rect 8028 -18950 8228 -18785
rect 15454 -18838 15816 -18785
rect 6736 -19524 7804 -19472
rect 15214 -19511 15506 -19510
rect -7449 -19576 7804 -19524
rect -7449 -19577 -5616 -19576
rect -4949 -19577 7804 -19576
rect -7017 -19597 -6483 -19577
rect -6248 -19586 -5616 -19577
rect -3748 -19586 -3116 -19577
rect -1248 -19586 -616 -19577
rect 1252 -19586 1884 -19577
rect 3752 -19586 4384 -19577
rect -7008 -19756 -6974 -19597
rect -6910 -19740 -6876 -19648
rect -6916 -19833 -6870 -19740
rect -6812 -19756 -6778 -19597
rect -6714 -19740 -6680 -19648
rect -6720 -19833 -6674 -19740
rect -6616 -19756 -6582 -19597
rect 6736 -19599 7804 -19577
rect -6518 -19740 -6484 -19648
rect -2406 -19662 -2270 -19616
rect 91 -19632 227 -19629
rect -2319 -19710 -2270 -19662
rect 58 -19666 2229 -19632
rect 91 -19675 227 -19666
rect -6524 -19801 -6478 -19740
rect -5501 -19801 -5455 -19735
rect -2319 -19746 2133 -19710
rect -6524 -19833 -5455 -19801
rect -6916 -19871 -5455 -19833
rect -6916 -19879 -6478 -19871
rect -6916 -20132 -6870 -19879
rect -6910 -20136 -6876 -20132
rect -6720 -19944 -6674 -19879
rect -6714 -20136 -6680 -19944
rect -6524 -19944 -6478 -19879
rect -6518 -20136 -6484 -19944
rect -5119 -20082 -5073 -19946
rect 2097 -19858 2133 -19746
rect 2195 -19790 2229 -19666
rect 5179 -19682 5315 -19676
rect 2274 -19701 2410 -19692
rect 2274 -19735 5075 -19701
rect 5179 -19716 5451 -19682
rect 5179 -19722 5315 -19716
rect 2274 -19738 2410 -19735
rect 5041 -19774 5075 -19735
rect 2195 -19824 3697 -19790
rect 5041 -19808 5381 -19774
rect -7596 -20463 -7460 -20417
rect -5116 -20335 -5076 -20082
rect -5116 -20381 -4980 -20335
rect -1363 -20554 -1226 -20503
rect -7740 -21591 -7556 -21528
rect -7719 -21592 -7556 -21591
rect -13200 -22497 -13065 -22491
rect -13220 -22499 -13065 -22497
rect -13427 -22535 -13065 -22499
rect -13017 -22514 -12587 -22484
rect -13017 -22522 -12598 -22514
rect -12408 -22526 -12374 -22370
rect -12310 -22478 -12276 -22370
rect -12212 -22526 -12178 -22370
rect -12114 -22478 -12080 -22370
rect -12016 -22381 -11644 -22311
rect -7265 -21023 -7231 -20831
rect -7271 -21088 -7225 -21023
rect -7069 -21023 -7035 -20831
rect -7075 -21088 -7029 -21023
rect -6873 -20835 -6839 -20831
rect -6879 -21088 -6833 -20835
rect -6334 -20812 -5706 -20778
rect -6427 -20946 -6393 -20846
rect -6334 -20863 -6292 -20812
rect -6432 -20990 -6390 -20946
rect -6329 -20954 -6295 -20863
rect -6231 -20936 -6197 -20846
rect -6138 -20868 -6096 -20812
rect -6232 -20990 -6196 -20936
rect -6133 -20954 -6099 -20868
rect -6035 -20936 -6001 -20846
rect -5944 -20867 -5902 -20812
rect -6038 -20954 -6001 -20936
rect -5937 -20954 -5903 -20867
rect -5839 -20938 -5805 -20846
rect -5742 -20857 -5706 -20812
rect -5741 -20931 -5707 -20857
rect -6038 -20990 -6002 -20954
rect -5840 -20990 -5804 -20938
rect -6432 -21024 -5804 -20990
rect -7271 -21096 -6833 -21088
rect -7301 -21105 -6833 -21096
rect -7383 -21107 -6833 -21105
rect -7384 -21134 -6833 -21107
rect -7384 -21144 -7225 -21134
rect -7384 -21502 -7336 -21144
rect -7301 -21166 -7225 -21144
rect -7271 -21227 -7225 -21166
rect -7265 -21319 -7231 -21227
rect -7167 -21370 -7133 -21211
rect -7075 -21227 -7029 -21134
rect -7069 -21319 -7035 -21227
rect -6971 -21370 -6937 -21211
rect -6879 -21227 -6833 -21134
rect -6797 -21109 -6629 -21103
rect -6432 -21109 -6257 -21024
rect -5748 -21078 -5701 -20931
rect -5657 -21072 -5583 -20904
rect -5522 -21023 -5488 -20831
rect -6797 -21162 -6257 -21109
rect -5873 -21152 -5701 -21078
rect -6797 -21177 -6629 -21162
rect -6432 -21191 -6257 -21162
rect -6873 -21319 -6839 -21227
rect -6775 -21370 -6741 -21211
rect -6432 -21225 -5801 -21191
rect -6432 -21232 -6390 -21225
rect -6431 -21275 -6390 -21232
rect -6427 -21369 -6393 -21275
rect -6329 -21357 -6295 -21261
rect -6234 -21274 -6193 -21225
rect -7266 -21438 -6732 -21370
rect -6335 -21415 -6291 -21357
rect -6231 -21369 -6197 -21274
rect -6133 -21346 -6099 -21261
rect -6040 -21274 -5999 -21225
rect -6138 -21415 -6094 -21346
rect -6035 -21369 -6001 -21274
rect -5937 -21346 -5903 -21261
rect -5842 -21266 -5801 -21225
rect -5942 -21415 -5898 -21346
rect -5839 -21369 -5805 -21266
rect -5748 -21287 -5701 -21152
rect -5656 -21096 -5583 -21072
rect -5528 -21088 -5482 -21023
rect -5326 -21023 -5292 -20831
rect -5332 -21088 -5286 -21023
rect -5130 -20835 -5096 -20831
rect -5136 -21088 -5090 -20835
rect -4932 -20931 -4875 -20853
rect -4932 -20976 -4671 -20931
rect -4932 -21017 -4875 -20976
rect -5528 -21096 -5090 -21088
rect -5656 -21134 -5090 -21096
rect -5656 -21166 -5482 -21134
rect -5528 -21227 -5482 -21166
rect -5741 -21357 -5707 -21287
rect -5522 -21319 -5488 -21227
rect -5746 -21415 -5702 -21357
rect -5424 -21370 -5390 -21211
rect -5332 -21227 -5286 -21134
rect -5326 -21319 -5292 -21227
rect -5228 -21370 -5194 -21211
rect -5136 -21227 -5090 -21134
rect -5054 -21114 -4886 -21103
rect -4716 -21110 -4671 -20976
rect -4565 -21023 -4531 -20831
rect -4571 -21088 -4525 -21023
rect -4369 -21023 -4335 -20831
rect -4375 -21088 -4329 -21023
rect -4173 -20835 -4139 -20831
rect -4179 -21088 -4133 -20835
rect -3634 -20812 -3006 -20778
rect -3727 -20946 -3693 -20846
rect -3634 -20863 -3592 -20812
rect -3732 -20990 -3690 -20946
rect -3629 -20954 -3595 -20863
rect -3531 -20936 -3497 -20846
rect -3438 -20868 -3396 -20812
rect -3532 -20990 -3496 -20936
rect -3433 -20954 -3399 -20868
rect -3335 -20936 -3301 -20846
rect -3244 -20867 -3202 -20812
rect -3338 -20954 -3301 -20936
rect -3237 -20954 -3203 -20867
rect -3139 -20938 -3105 -20846
rect -3042 -20857 -3006 -20812
rect -3041 -20931 -3007 -20857
rect -3338 -20990 -3302 -20954
rect -3140 -20990 -3104 -20938
rect -3732 -21024 -3104 -20990
rect -4571 -21096 -4133 -21088
rect -4601 -21110 -4133 -21096
rect -4826 -21114 -4766 -21113
rect -5054 -21172 -4766 -21114
rect -4716 -21134 -4133 -21110
rect -4716 -21155 -4525 -21134
rect -5054 -21177 -4886 -21172
rect -5130 -21319 -5096 -21227
rect -5032 -21370 -4998 -21211
rect -4826 -21245 -4766 -21172
rect -4711 -21270 -4651 -21155
rect -4601 -21166 -4525 -21155
rect -4571 -21227 -4525 -21166
rect -4565 -21319 -4531 -21227
rect -4467 -21370 -4433 -21211
rect -4375 -21227 -4329 -21134
rect -4369 -21319 -4335 -21227
rect -4271 -21370 -4237 -21211
rect -4179 -21227 -4133 -21134
rect -4097 -21112 -3929 -21103
rect -3732 -21112 -3557 -21024
rect -3048 -21078 -3001 -20931
rect -2957 -21072 -2883 -20904
rect -2822 -21023 -2788 -20831
rect -4097 -21169 -3557 -21112
rect -3173 -21152 -3001 -21078
rect -4097 -21177 -3929 -21169
rect -3732 -21191 -3557 -21169
rect -4173 -21319 -4139 -21227
rect -4075 -21370 -4041 -21211
rect -3732 -21225 -3101 -21191
rect -3732 -21232 -3690 -21225
rect -3731 -21265 -3690 -21232
rect -3731 -21275 -3684 -21265
rect -6335 -21449 -5702 -21415
rect -5523 -21438 -4032 -21370
rect -3730 -21397 -3684 -21275
rect -3629 -21357 -3595 -21261
rect -3534 -21274 -3493 -21225
rect -3635 -21415 -3591 -21357
rect -3531 -21369 -3497 -21274
rect -3433 -21346 -3399 -21261
rect -3340 -21274 -3299 -21225
rect -3438 -21415 -3394 -21346
rect -3335 -21369 -3301 -21274
rect -3237 -21346 -3203 -21261
rect -3142 -21266 -3101 -21225
rect -3242 -21415 -3198 -21346
rect -3139 -21369 -3105 -21266
rect -3048 -21287 -3001 -21152
rect -2956 -21096 -2883 -21072
rect -2828 -21088 -2782 -21023
rect -2626 -21023 -2592 -20831
rect -2632 -21088 -2586 -21023
rect -2430 -20835 -2396 -20831
rect -2436 -21088 -2390 -20835
rect -2232 -21017 -2175 -20853
rect -1940 -21023 -1906 -20831
rect -2828 -21096 -2390 -21088
rect -1946 -21088 -1900 -21023
rect -1744 -21023 -1710 -20831
rect -1750 -21088 -1704 -21023
rect -1548 -20835 -1514 -20831
rect -1554 -21088 -1508 -20835
rect -1946 -21096 -1508 -21088
rect -2956 -21134 -2390 -21096
rect -2956 -21166 -2782 -21134
rect -3041 -21357 -3007 -21287
rect -3046 -21415 -3002 -21357
rect -3635 -21449 -3002 -21415
rect -2957 -21362 -2883 -21203
rect -2828 -21227 -2782 -21166
rect -2822 -21319 -2788 -21227
rect -6648 -21485 -6516 -21472
rect -2957 -21485 -2882 -21362
rect -2724 -21370 -2690 -21211
rect -2632 -21227 -2586 -21134
rect -2626 -21319 -2592 -21227
rect -2528 -21370 -2494 -21211
rect -2436 -21227 -2390 -21134
rect -2354 -21114 -2186 -21103
rect -2354 -21172 -2151 -21114
rect -2094 -21118 -2034 -21114
rect -1976 -21118 -1508 -21096
rect -1363 -21103 -1324 -20554
rect 2097 -19894 3618 -19858
rect 1933 -20379 2069 -20333
rect 1829 -20463 1984 -20417
rect -2094 -21134 -1508 -21118
rect -2094 -21160 -1900 -21134
rect -2354 -21177 -2186 -21172
rect -2430 -21319 -2396 -21227
rect -2332 -21370 -2298 -21211
rect -2094 -21246 -2034 -21160
rect -1976 -21166 -1900 -21160
rect -1946 -21227 -1900 -21166
rect -1940 -21319 -1906 -21227
rect -1842 -21370 -1808 -21211
rect -1750 -21227 -1704 -21134
rect -1744 -21319 -1710 -21227
rect -1646 -21370 -1612 -21211
rect -1554 -21227 -1508 -21134
rect -1472 -21177 -1304 -21103
rect -1548 -21319 -1514 -21227
rect -1450 -21370 -1416 -21211
rect -2823 -21438 -1407 -21370
rect -1363 -21485 -1324 -21177
rect -1010 -21258 -976 -20848
rect -272 -21092 -238 -20848
rect -76 -21092 -42 -20848
rect 120 -21092 154 -20848
rect -401 -21129 154 -21092
rect 340 -21095 386 -21011
rect 723 -21033 757 -20861
rect 919 -20969 953 -20861
rect 1115 -20969 1149 -20861
rect -1161 -21311 -976 -21258
rect -941 -21267 -806 -21257
rect -401 -21267 -364 -21129
rect 194 -21149 386 -21095
rect 586 -21103 757 -21033
rect 1194 -21016 1267 -21003
rect 1194 -21044 1367 -21016
rect 1194 -21057 1389 -21044
rect 1194 -21063 1267 -21057
rect -142 -21186 -7 -21177
rect 421 -21186 557 -21185
rect -142 -21224 557 -21186
rect -142 -21231 -7 -21224
rect 421 -21231 557 -21224
rect -941 -21304 -364 -21267
rect -941 -21311 -806 -21304
rect -7385 -21639 -7325 -21502
rect -7054 -21524 -1324 -21485
rect -6648 -21532 -6516 -21524
rect -4875 -21571 -4738 -21561
rect -3929 -21571 -3797 -21560
rect -1915 -21571 -1783 -21561
rect -7054 -21610 -1783 -21571
rect -4875 -21621 -4738 -21610
rect -3929 -21620 -3797 -21610
rect -1915 -21621 -1783 -21610
rect -7384 -22011 -7336 -21639
rect -7037 -21663 -6900 -21650
rect -4440 -21663 -4303 -21644
rect -1672 -21663 -1540 -21644
rect -7054 -21702 -1539 -21663
rect -7037 -21710 -6900 -21702
rect -7026 -21750 -6915 -21710
rect -6215 -21750 -6104 -21702
rect -4440 -21704 -4303 -21702
rect -7274 -21818 -5903 -21750
rect -5724 -21773 -5091 -21739
rect -4417 -21750 -4306 -21704
rect -4234 -21750 -3714 -21748
rect -3539 -21750 -3428 -21702
rect -7265 -21977 -7231 -21818
rect -7167 -21961 -7133 -21869
rect -7384 -22055 -7209 -22011
rect -7377 -22085 -7209 -22055
rect -7173 -22054 -7127 -21961
rect -7069 -21977 -7035 -21818
rect -6971 -21961 -6937 -21869
rect -6977 -22054 -6931 -21961
rect -6873 -21977 -6839 -21818
rect -6775 -21961 -6741 -21869
rect -6781 -22022 -6735 -21961
rect -6612 -22011 -6552 -21867
rect -6428 -21977 -6394 -21818
rect -6330 -21961 -6296 -21869
rect -6781 -22054 -6648 -22022
rect -7173 -22092 -6648 -22054
rect -6612 -22073 -6372 -22011
rect -6575 -22074 -6372 -22073
rect -6540 -22085 -6372 -22074
rect -6336 -22054 -6290 -21961
rect -6232 -21977 -6198 -21818
rect -6134 -21961 -6100 -21869
rect -6140 -22054 -6094 -21961
rect -6036 -21977 -6002 -21818
rect -5724 -21831 -5680 -21773
rect -5938 -21961 -5904 -21869
rect -5719 -21901 -5685 -21831
rect -5944 -22022 -5898 -21961
rect -5944 -22054 -5770 -22022
rect -7173 -22100 -6735 -22092
rect -7173 -22353 -7127 -22100
rect -7167 -22357 -7133 -22353
rect -6977 -22165 -6931 -22100
rect -6971 -22357 -6937 -22165
rect -6781 -22165 -6735 -22100
rect -6775 -22357 -6741 -22165
rect -6694 -22222 -6648 -22092
rect -6336 -22092 -5770 -22054
rect -6336 -22100 -5898 -22092
rect -6551 -22222 -6494 -22171
rect -6694 -22271 -6494 -22222
rect -6551 -22335 -6494 -22271
rect -6336 -22353 -6290 -22100
rect -6330 -22357 -6296 -22353
rect -6140 -22165 -6094 -22100
rect -6134 -22357 -6100 -22165
rect -5944 -22165 -5898 -22100
rect -5843 -22116 -5770 -22092
rect -5725 -22036 -5678 -21901
rect -5621 -21922 -5587 -21819
rect -5528 -21842 -5484 -21773
rect -5625 -21963 -5584 -21922
rect -5523 -21927 -5489 -21842
rect -5425 -21914 -5391 -21819
rect -5332 -21842 -5288 -21773
rect -5427 -21963 -5386 -21914
rect -5327 -21927 -5293 -21842
rect -5229 -21914 -5195 -21819
rect -5135 -21831 -5091 -21773
rect -4574 -21816 -3203 -21750
rect -4574 -21818 -4040 -21816
rect -3737 -21818 -3203 -21816
rect -3024 -21773 -2391 -21739
rect -5233 -21963 -5192 -21914
rect -5131 -21927 -5097 -21831
rect -5033 -21913 -4999 -21819
rect -5036 -21956 -4995 -21913
rect -5036 -21963 -4994 -21956
rect -5625 -21997 -4994 -21963
rect -4565 -21977 -4531 -21818
rect -4467 -21961 -4433 -21869
rect -5725 -22110 -5553 -22036
rect -5169 -22057 -4903 -21997
rect -4677 -22018 -4509 -22011
rect -5938 -22357 -5904 -22165
rect -5843 -22284 -5769 -22116
rect -5725 -22257 -5678 -22110
rect -5169 -22164 -4994 -22057
rect -4699 -22078 -4509 -22018
rect -4677 -22085 -4509 -22078
rect -4473 -22054 -4427 -21961
rect -4369 -21977 -4335 -21818
rect -4271 -21961 -4237 -21869
rect -4277 -22054 -4231 -21961
rect -4173 -21977 -4139 -21818
rect -4075 -21961 -4041 -21869
rect -4081 -22022 -4035 -21961
rect -3900 -22011 -3840 -21852
rect -3728 -21977 -3694 -21818
rect -3630 -21961 -3596 -21869
rect -4081 -22054 -3937 -22022
rect -4473 -22092 -3937 -22054
rect -3900 -22074 -3672 -22011
rect -3840 -22085 -3672 -22074
rect -3636 -22054 -3590 -21961
rect -3532 -21977 -3498 -21818
rect -3434 -21961 -3400 -21869
rect -3440 -22054 -3394 -21961
rect -3336 -21977 -3302 -21818
rect -3024 -21831 -2980 -21773
rect -3238 -21961 -3204 -21869
rect -3019 -21901 -2985 -21831
rect -3244 -22022 -3198 -21961
rect -3244 -22054 -3070 -22022
rect -4473 -22100 -4035 -22092
rect -5622 -22198 -4994 -22164
rect -5622 -22250 -5586 -22198
rect -5424 -22234 -5388 -22198
rect -5719 -22331 -5685 -22257
rect -5720 -22376 -5684 -22331
rect -5621 -22342 -5587 -22250
rect -5523 -22321 -5489 -22234
rect -5425 -22252 -5388 -22234
rect -5524 -22376 -5482 -22321
rect -5425 -22342 -5391 -22252
rect -5327 -22320 -5293 -22234
rect -5230 -22252 -5194 -22198
rect -5330 -22376 -5288 -22320
rect -5229 -22342 -5195 -22252
rect -5131 -22325 -5097 -22234
rect -5036 -22242 -4994 -22198
rect -5134 -22376 -5092 -22325
rect -5033 -22342 -4999 -22242
rect -5720 -22410 -5092 -22376
rect -4473 -22353 -4427 -22100
rect -4467 -22357 -4433 -22353
rect -4277 -22165 -4231 -22100
rect -4271 -22357 -4237 -22165
rect -4081 -22165 -4035 -22100
rect -4075 -22357 -4041 -22165
rect -3999 -22221 -3937 -22092
rect -3636 -22092 -3070 -22054
rect -3636 -22100 -3198 -22092
rect -3851 -22221 -3794 -22171
rect -3999 -22283 -3794 -22221
rect -3851 -22335 -3794 -22283
rect -3636 -22353 -3590 -22100
rect -3630 -22357 -3596 -22353
rect -3440 -22165 -3394 -22100
rect -3434 -22357 -3400 -22165
rect -3244 -22165 -3198 -22100
rect -3143 -22116 -3070 -22092
rect -3025 -22036 -2978 -21901
rect -2921 -21922 -2887 -21819
rect -2828 -21842 -2784 -21773
rect -2925 -21963 -2884 -21922
rect -2823 -21927 -2789 -21842
rect -2725 -21914 -2691 -21819
rect -2632 -21842 -2588 -21773
rect -2727 -21963 -2686 -21914
rect -2627 -21927 -2593 -21842
rect -2529 -21914 -2495 -21819
rect -2435 -21831 -2391 -21773
rect -2533 -21963 -2492 -21914
rect -2431 -21927 -2397 -21831
rect -2333 -21913 -2299 -21819
rect -2336 -21956 -2295 -21913
rect -2336 -21963 -2294 -21956
rect -2925 -21995 -2294 -21963
rect -2925 -21997 -2219 -21995
rect -3025 -22110 -2853 -22036
rect -2469 -22055 -2219 -21997
rect -3238 -22357 -3204 -22165
rect -3143 -22284 -3069 -22116
rect -3025 -22257 -2978 -22110
rect -2469 -22164 -2294 -22055
rect -2922 -22198 -2294 -22164
rect -2922 -22250 -2886 -22198
rect -2724 -22234 -2688 -22198
rect -3019 -22331 -2985 -22257
rect -3020 -22376 -2984 -22331
rect -2921 -22342 -2887 -22250
rect -2823 -22321 -2789 -22234
rect -2725 -22252 -2688 -22234
rect -2824 -22376 -2782 -22321
rect -2725 -22342 -2691 -22252
rect -2627 -22320 -2593 -22234
rect -2530 -22252 -2494 -22198
rect -2630 -22376 -2588 -22320
rect -2529 -22342 -2495 -22252
rect -2431 -22325 -2397 -22234
rect -2336 -22242 -2294 -22198
rect -2434 -22376 -2392 -22325
rect -2333 -22342 -2299 -22242
rect -2055 -22282 -1757 -21702
rect -1672 -21704 -1540 -21702
rect -1010 -21764 -976 -21311
rect -401 -21358 -364 -21304
rect -330 -21268 -195 -21255
rect 592 -21268 626 -21103
rect 821 -21200 855 -21092
rect 919 -21248 953 -21092
rect 1017 -21200 1051 -21092
rect 1115 -21248 1149 -21092
rect 1328 -21206 1389 -21057
rect 1528 -21206 1562 -20862
rect 1724 -21206 1758 -20862
rect 1328 -21236 1758 -21206
rect 1948 -21213 1984 -20463
rect 1339 -21244 1758 -21236
rect 1806 -21221 1984 -21213
rect -330 -21302 626 -21268
rect -330 -21309 -195 -21302
rect 674 -21334 1289 -21248
rect 1806 -21257 1993 -21221
rect 1806 -21261 1971 -21257
rect 1806 -21267 1941 -21261
rect 1402 -21317 1476 -21291
rect 2029 -21315 2069 -20379
rect 2328 -21035 2362 -20863
rect 2524 -20971 2558 -20863
rect 2720 -20971 2754 -20863
rect 1887 -21317 2069 -21315
rect -597 -21392 -364 -21358
rect -191 -21392 252 -21358
rect -912 -21952 -878 -21556
rect -597 -21764 -563 -21392
rect -499 -21862 -465 -21456
rect -401 -21764 -367 -21392
rect -191 -21393 56 -21392
rect -191 -21456 -156 -21393
rect -288 -21753 -254 -21456
rect -289 -21859 -254 -21753
rect -190 -21764 -156 -21456
rect -92 -21755 -58 -21456
rect -93 -21859 -58 -21755
rect 22 -21763 56 -21393
rect -289 -21862 -58 -21859
rect -499 -21896 -58 -21862
rect 120 -21952 154 -21455
rect 218 -21763 252 -21392
rect 984 -21741 1045 -21334
rect 1402 -21355 2069 -21317
rect 2164 -21105 2362 -21035
rect 2799 -21018 2872 -21005
rect 2799 -21046 2972 -21018
rect 2799 -21059 2994 -21046
rect 2799 -21065 2872 -21059
rect 1402 -21356 1888 -21355
rect 1402 -21362 1476 -21356
rect 1817 -21357 1888 -21356
rect 1430 -21707 1464 -21399
rect 1528 -21707 1562 -21399
rect 1626 -21707 1660 -21399
rect 1724 -21707 1758 -21399
rect 1822 -21707 1856 -21399
rect 984 -21759 1434 -21741
rect 1724 -21759 1759 -21707
rect 984 -21802 1876 -21759
rect -1022 -22017 252 -21952
rect -1009 -22282 -879 -22017
rect -703 -22282 -573 -22017
rect -386 -22282 -256 -22017
rect 60 -22282 190 -22017
rect 984 -22282 1135 -21802
rect 1361 -21820 1876 -21802
rect 1361 -22282 1485 -21820
rect 1691 -22282 1815 -21820
rect 2164 -21840 2234 -21105
rect 2426 -21202 2460 -21094
rect 2524 -21250 2558 -21094
rect 2622 -21202 2656 -21094
rect 2720 -21250 2754 -21094
rect 2933 -21208 2994 -21059
rect 3133 -21208 3167 -20864
rect 3329 -21208 3363 -20864
rect 2933 -21238 3363 -21208
rect 2944 -21246 3363 -21238
rect 3411 -21221 3546 -21215
rect 3582 -21221 3618 -19894
rect 2279 -21336 2894 -21250
rect 3411 -21259 3618 -21221
rect 3411 -21261 3598 -21259
rect 3411 -21269 3546 -21261
rect 3007 -21319 3081 -21293
rect 3657 -21317 3697 -19824
rect 3492 -21319 3697 -21317
rect 2098 -21886 2234 -21840
rect 2589 -21743 2650 -21336
rect 3007 -21357 3697 -21319
rect 3007 -21358 3493 -21357
rect 3007 -21364 3081 -21358
rect 3422 -21359 3493 -21358
rect 3035 -21709 3069 -21401
rect 3133 -21709 3167 -21401
rect 3231 -21709 3265 -21401
rect 3329 -21709 3363 -21401
rect 3427 -21709 3461 -21401
rect 3952 -21439 3986 -20839
rect 4690 -21083 4724 -20839
rect 4886 -21083 4920 -20839
rect 5082 -21083 5116 -20839
rect 4561 -21120 5116 -21083
rect 5156 -21094 5291 -21086
rect 4021 -21258 4156 -21248
rect 4561 -21258 4598 -21120
rect 5155 -21131 5310 -21094
rect 5155 -21140 5291 -21131
rect 4820 -21177 4955 -21168
rect 5347 -21177 5381 -19808
rect 4820 -21215 5381 -21177
rect 4820 -21222 4955 -21215
rect 4021 -21295 4598 -21258
rect 4021 -21302 4156 -21295
rect 4561 -21349 4598 -21295
rect 4632 -21259 4767 -21246
rect 5417 -21259 5451 -19716
rect 5565 -20746 6293 -20712
rect 5565 -21058 5599 -20746
rect 5663 -21094 5697 -20850
rect 5761 -21058 5795 -20746
rect 5881 -20815 6223 -20781
rect 5881 -21058 5915 -20815
rect 5979 -21094 6013 -20850
rect 6077 -21058 6111 -20815
rect 5514 -21128 6128 -21094
rect 4632 -21293 5451 -21259
rect 5564 -21262 5703 -21208
rect 6094 -21243 6128 -21128
rect 6189 -21167 6223 -20815
rect 6259 -21093 6293 -20746
rect 6439 -21093 6473 -20850
rect 6259 -21127 6473 -21093
rect 6635 -21167 6669 -20850
rect 6945 -21043 6979 -20850
rect 6189 -21201 6669 -21167
rect 6722 -21218 6861 -21164
rect 6094 -21277 6240 -21243
rect 4632 -21300 4767 -21293
rect 3736 -21497 3986 -21439
rect 2589 -21761 3039 -21743
rect 3329 -21761 3364 -21709
rect 2589 -21804 3481 -21761
rect 2589 -22282 2740 -21804
rect 3031 -21822 3481 -21804
rect 3031 -22282 3182 -21822
rect 3324 -22282 3475 -21822
rect 3736 -21952 3801 -21497
rect 3952 -21755 3986 -21497
rect 4365 -21383 4598 -21349
rect 4771 -21383 5214 -21349
rect 4050 -21943 4084 -21547
rect 4365 -21755 4399 -21383
rect 4463 -21853 4497 -21447
rect 4561 -21755 4595 -21383
rect 4771 -21384 5018 -21383
rect 4771 -21447 4806 -21384
rect 4674 -21744 4708 -21447
rect 4673 -21850 4708 -21744
rect 4772 -21755 4806 -21447
rect 4870 -21746 4904 -21447
rect 4869 -21850 4904 -21746
rect 4984 -21754 5018 -21384
rect 4673 -21853 4904 -21850
rect 4463 -21887 4904 -21853
rect 5082 -21943 5116 -21446
rect 5180 -21754 5214 -21383
rect 5563 -21380 5894 -21343
rect 6206 -21339 6240 -21277
rect 6313 -21292 6452 -21238
rect 6206 -21373 6767 -21339
rect 5563 -21463 5600 -21380
rect 5857 -21404 5894 -21380
rect 5857 -21441 6013 -21404
rect 5565 -21652 5599 -21463
rect 5561 -21775 5600 -21652
rect 5663 -21701 5697 -21456
rect 5976 -21462 6013 -21441
rect 5979 -21664 6013 -21462
rect 6075 -21465 6375 -21426
rect 6077 -21664 6111 -21465
rect 6341 -21664 6375 -21465
rect 6439 -21664 6473 -21373
rect 6635 -21647 6669 -21456
rect 6635 -21701 6671 -21647
rect 6733 -21664 6767 -21373
rect 6940 -21382 6983 -21043
rect 7254 -21041 7288 -20850
rect 7250 -21238 7293 -21041
rect 7337 -21224 7476 -21170
rect 7150 -21284 7293 -21238
rect 6844 -21428 6983 -21382
rect 6940 -21473 6983 -21428
rect 6945 -21664 6979 -21473
rect 7043 -21657 7077 -21456
rect 7250 -21475 7293 -21284
rect 5663 -21737 6671 -21701
rect 7038 -21741 7081 -21657
rect 7254 -21664 7288 -21475
rect 7352 -21655 7386 -21456
rect 7347 -21741 7390 -21655
rect 6762 -21775 7394 -21741
rect 5561 -21828 7394 -21775
rect 3666 -21998 3802 -21952
rect 3940 -22008 5214 -21943
rect 3964 -22282 4110 -22008
rect 4409 -22282 4555 -22008
rect 4675 -22282 4821 -22008
rect 5035 -22282 5181 -22008
rect 5599 -22282 5796 -21828
rect 6132 -22282 6329 -21828
rect 6645 -21837 7394 -21828
rect 6645 -22282 6842 -21837
rect 7148 -22282 7345 -21837
rect 7543 -22282 7804 -19599
rect 8240 -19650 15506 -19511
rect 15267 -20114 15502 -20091
rect 9859 -20359 15502 -20114
rect 9859 -20361 15378 -20359
rect 15181 -20530 15448 -20494
rect 9836 -20765 15448 -20530
rect 15181 -20792 15448 -20765
rect 8268 -21124 8486 -21116
rect 15444 -21124 15597 -21085
rect 8268 -21199 15597 -21124
rect 8268 -21205 8486 -21199
rect 15444 -21236 15597 -21199
rect 9250 -21345 9300 -21339
rect 14762 -21345 14860 -21331
rect 9241 -21468 14860 -21345
rect 9250 -21472 9300 -21468
rect 14762 -21495 14860 -21468
rect 15679 -21750 15807 -18838
rect 15932 -21661 16064 -18410
rect 16174 -21085 16263 -17935
rect 18266 -19149 18811 -17611
rect 17683 -19655 83656 -19149
rect 17038 -20294 17256 -20048
rect 16174 -21236 16271 -21085
rect 17077 -21151 17219 -20294
rect 18266 -21119 18811 -19655
rect 25279 -20154 25609 -20071
rect 28012 -20116 28295 -19655
rect 27768 -20144 28433 -20116
rect 33380 -20131 33737 -20064
rect 34558 -20131 34915 -20098
rect 36411 -20127 36694 -19655
rect 25279 -20333 26458 -20154
rect 27768 -20202 28803 -20144
rect 27768 -20283 27854 -20202
rect 28028 -20239 28063 -20202
rect 28353 -20205 28803 -20202
rect 25279 -20365 25609 -20333
rect 26916 -20369 27854 -20283
rect 26764 -20659 26894 -20567
rect 27056 -20625 27090 -20369
rect 27154 -20625 27188 -20417
rect 27252 -20625 27286 -20369
rect 27350 -20591 27384 -20417
rect 27931 -20547 27965 -20239
rect 28029 -20547 28063 -20239
rect 28127 -20547 28161 -20239
rect 28225 -20547 28259 -20239
rect 28323 -20547 28357 -20239
rect 27899 -20590 27970 -20589
rect 28311 -20590 28385 -20584
rect 27899 -20591 28385 -20590
rect 27350 -20625 28385 -20591
rect 28742 -20612 28803 -20205
rect 33380 -20320 34915 -20131
rect 36208 -20155 36873 -20127
rect 36208 -20213 37243 -20155
rect 45323 -20166 45606 -19655
rect 54542 -20132 54825 -19655
rect 59891 -20100 60267 -20005
rect 63337 -20066 63644 -19655
rect 61492 -20100 61742 -20073
rect 36208 -20294 36294 -20213
rect 36468 -20250 36503 -20213
rect 36793 -20216 37243 -20213
rect 33380 -20331 33737 -20320
rect 34558 -20365 34915 -20320
rect 35356 -20380 36294 -20294
rect 27351 -20629 28385 -20625
rect 27351 -20631 27900 -20629
rect 26938 -20659 27011 -20653
rect 28311 -20655 28385 -20629
rect 26764 -20700 27011 -20659
rect 27846 -20687 27981 -20679
rect 27826 -20689 27981 -20687
rect 26764 -20717 26894 -20700
rect 26938 -20713 27011 -20700
rect 27619 -20725 27981 -20689
rect 28498 -20698 29283 -20612
rect 35204 -20670 35334 -20578
rect 35496 -20636 35530 -20380
rect 35594 -20636 35628 -20428
rect 35692 -20636 35726 -20380
rect 35790 -20602 35824 -20428
rect 36371 -20558 36405 -20250
rect 36469 -20558 36503 -20250
rect 36567 -20558 36601 -20250
rect 36665 -20558 36699 -20250
rect 36763 -20558 36797 -20250
rect 36339 -20601 36410 -20600
rect 36751 -20601 36825 -20595
rect 36339 -20602 36825 -20601
rect 35790 -20636 36825 -20602
rect 37182 -20623 37243 -20216
rect 41936 -20220 42201 -20189
rect 43462 -20220 43759 -20187
rect 41936 -20387 43759 -20220
rect 45071 -20194 45736 -20166
rect 45071 -20252 46106 -20194
rect 45071 -20333 45157 -20252
rect 45331 -20289 45366 -20252
rect 45656 -20255 46106 -20252
rect 41936 -20454 42201 -20387
rect 43462 -20409 43759 -20387
rect 44219 -20419 45157 -20333
rect 35791 -20640 36825 -20636
rect 35791 -20642 36340 -20640
rect 35378 -20670 35451 -20664
rect 36751 -20666 36825 -20640
rect 27826 -20727 27981 -20725
rect 27846 -20733 27981 -20727
rect 28029 -20710 28448 -20702
rect 28029 -20740 28459 -20710
rect 27056 -20955 27090 -20747
rect 27252 -20955 27286 -20747
rect 27448 -20955 27482 -20747
rect 19676 -21081 20304 -21047
rect 16174 -21569 16263 -21236
rect 17040 -21340 17219 -21151
rect 17368 -21225 19138 -21119
rect 19583 -21215 19617 -21115
rect 19676 -21132 19718 -21081
rect 17472 -21371 17520 -21225
rect 17477 -21542 17511 -21371
rect 17575 -21525 17609 -21334
rect 17666 -21374 17714 -21225
rect 17291 -21569 17436 -21562
rect 16174 -21610 17436 -21569
rect 17291 -21618 17436 -21610
rect 17571 -21576 17613 -21525
rect 17673 -21542 17707 -21374
rect 17771 -21525 17805 -21334
rect 17767 -21576 17809 -21525
rect 17571 -21618 18357 -21576
rect 18218 -21636 18357 -21618
rect 17620 -21661 17765 -21657
rect 15932 -21702 17765 -21661
rect 17620 -21713 17765 -21702
rect 17940 -21745 18085 -21689
rect 17940 -21750 18000 -21745
rect 15679 -21791 18000 -21750
rect 18218 -21818 18260 -21636
rect 17473 -21864 17922 -21827
rect -3020 -22410 -2392 -22376
rect -13220 -22537 -13065 -22535
rect -13200 -22545 -13065 -22537
rect -13695 -22595 -13146 -22593
rect -12735 -22595 -12661 -22569
rect -13695 -22599 -12661 -22595
rect -13990 -22855 -13956 -22599
rect -13892 -22807 -13858 -22599
rect -13794 -22855 -13760 -22599
rect -13696 -22633 -12661 -22599
rect -12548 -22612 -11763 -22526
rect -13696 -22807 -13662 -22633
rect -13147 -22634 -12661 -22633
rect -13147 -22635 -13076 -22634
rect -12735 -22640 -12661 -22634
rect -14130 -22941 -13192 -22855
rect -13278 -23022 -13192 -22941
rect -13115 -22985 -13081 -22677
rect -13017 -22985 -12983 -22677
rect -12919 -22985 -12885 -22677
rect -12821 -22985 -12787 -22677
rect -12723 -22985 -12689 -22677
rect -13018 -23022 -12983 -22985
rect -12304 -23019 -12243 -22612
rect -12693 -23022 -12243 -23019
rect -13278 -23080 -12243 -23022
rect -13278 -23108 -12613 -23080
rect -25664 -23404 -25039 -23185
rect -17094 -23217 -16826 -23185
rect -15041 -23324 -15007 -23320
rect -15047 -23577 -15001 -23324
rect -14845 -23512 -14811 -23320
rect -14851 -23577 -14805 -23512
rect -14649 -23512 -14615 -23320
rect -14425 -23406 -14368 -23342
rect -14568 -23455 -14368 -23406
rect -14655 -23577 -14609 -23512
rect -15047 -23585 -14609 -23577
rect -14568 -23585 -14522 -23455
rect -14425 -23506 -14368 -23455
rect -14204 -23324 -14170 -23320
rect -15251 -23622 -15083 -23592
rect -15258 -23666 -15083 -23622
rect -15047 -23623 -14522 -23585
rect -14210 -23577 -14164 -23324
rect -14008 -23512 -13974 -23320
rect -14014 -23577 -13968 -23512
rect -13594 -23301 -12966 -23267
rect -13812 -23512 -13778 -23320
rect -13594 -23346 -13558 -23301
rect -13818 -23577 -13772 -23512
rect -14210 -23585 -13772 -23577
rect -13717 -23561 -13643 -23393
rect -13593 -23420 -13559 -23346
rect -13717 -23585 -13644 -23561
rect -14414 -23603 -14246 -23592
rect -14449 -23604 -14246 -23603
rect -22518 -24996 -22484 -24405
rect -22218 -24369 -21755 -24335
rect -22522 -25047 -22481 -24996
rect -22306 -25003 -22272 -24405
rect -22218 -24411 -22165 -24369
rect -22311 -25047 -22269 -25003
rect -22208 -25013 -22174 -24411
rect -22110 -25002 -22076 -24405
rect -22009 -24411 -21953 -24369
rect -22115 -25047 -22073 -25002
rect -21997 -25013 -21963 -24411
rect -21899 -24995 -21865 -24405
rect -21811 -24411 -21755 -24369
rect -22522 -25084 -22073 -25047
rect -21903 -25051 -21861 -24995
rect -21801 -25013 -21767 -24411
rect -21312 -24737 -21278 -24334
rect -21108 -24298 -20864 -24260
rect -21313 -24776 -21277 -24737
rect -21108 -24362 -21062 -24298
rect -21101 -24742 -21067 -24362
rect -21003 -24732 -20969 -24334
rect -20910 -24362 -20864 -24298
rect -20905 -24696 -20871 -24362
rect -21010 -24776 -20965 -24732
rect -21313 -24812 -20965 -24776
rect -20908 -24928 -20858 -24696
rect -20407 -24738 -20373 -24335
rect -20203 -24299 -19959 -24261
rect -20408 -24777 -20372 -24738
rect -20203 -24363 -20157 -24299
rect -20196 -24743 -20162 -24363
rect -20098 -24733 -20064 -24335
rect -20005 -24363 -19959 -24299
rect -18292 -24337 -16815 -24224
rect -20000 -24697 -19966 -24363
rect -19123 -24632 -18674 -24614
rect -18292 -24632 -18231 -24337
rect -17565 -24455 -17518 -24337
rect -19635 -24693 -18231 -24632
rect -20105 -24777 -20060 -24733
rect -20408 -24813 -20060 -24777
rect -20908 -24941 -20762 -24928
rect -20003 -24929 -19953 -24697
rect -20964 -24950 -20762 -24941
rect -21903 -25093 -21735 -25051
rect -21219 -24986 -20762 -24950
rect -20003 -24942 -19831 -24929
rect -20059 -24951 -19831 -24942
rect -21777 -25277 -21735 -25093
rect -21312 -25185 -21278 -25026
rect -21219 -25035 -21174 -24986
rect -21786 -25293 -21649 -25277
rect -22424 -25335 -21649 -25293
rect -22518 -25540 -22484 -25369
rect -22424 -25386 -22382 -25335
rect -22523 -25669 -22475 -25540
rect -22420 -25577 -22386 -25386
rect -22322 -25537 -22288 -25369
rect -22228 -25386 -22186 -25335
rect -21316 -25337 -21272 -25185
rect -21214 -25234 -21180 -25035
rect -21116 -25186 -21082 -25026
rect -20314 -24987 -19831 -24951
rect -20407 -25186 -20373 -25027
rect -20314 -25036 -20269 -24987
rect -21122 -25337 -21078 -25186
rect -21445 -25372 -20848 -25337
rect -20411 -25338 -20367 -25186
rect -20309 -25235 -20275 -25036
rect -20211 -25187 -20177 -25027
rect -19635 -25051 -19574 -24693
rect -19006 -24727 -18971 -24693
rect -19103 -25035 -19069 -24727
rect -19005 -25035 -18971 -24727
rect -18907 -25035 -18873 -24727
rect -18809 -25035 -18775 -24727
rect -18711 -25035 -18677 -24727
rect -20022 -25112 -19574 -25051
rect -19135 -25078 -19064 -25077
rect -18723 -25078 -18649 -25072
rect -19135 -25079 -18649 -25078
rect -20217 -25338 -20173 -25187
rect -20022 -25338 -19961 -25112
rect -19361 -25117 -18649 -25079
rect -18292 -25100 -18231 -24693
rect -17558 -24749 -17524 -24455
rect -17460 -24733 -17426 -24441
rect -17369 -24456 -17322 -24337
rect -17667 -24795 -17512 -24783
rect -17704 -24829 -17512 -24795
rect -17667 -24838 -17512 -24829
rect -17466 -24803 -17421 -24733
rect -17362 -24749 -17328 -24456
rect -17127 -24466 -17080 -24337
rect -17120 -24749 -17086 -24466
rect -17022 -24740 -16988 -24441
rect -17026 -24780 -16982 -24740
rect -16134 -24780 -15997 -24710
rect -17026 -24783 -15997 -24780
rect -17466 -24843 -17112 -24803
rect -17074 -24823 -15997 -24783
rect -17802 -24900 -17732 -24898
rect -17397 -24900 -17242 -24891
rect -17802 -24936 -17242 -24900
rect -19361 -25119 -19134 -25117
rect -18723 -25143 -18649 -25117
rect -19707 -25177 -19590 -25162
rect -19188 -25175 -19053 -25167
rect -19208 -25177 -19053 -25175
rect -19707 -25213 -19053 -25177
rect -18536 -25186 -17921 -25100
rect -19707 -25285 -19590 -25213
rect -19208 -25215 -19053 -25213
rect -19188 -25221 -19053 -25215
rect -19005 -25198 -18586 -25190
rect -19005 -25228 -18575 -25198
rect -20540 -25372 -19943 -25338
rect -22329 -25669 -22281 -25537
rect -22224 -25577 -22190 -25386
rect -22000 -25427 -19943 -25372
rect -22000 -25488 -20159 -25427
rect -22000 -25669 -21884 -25488
rect -22658 -25686 -21854 -25669
rect -19005 -25572 -18971 -25228
rect -18809 -25572 -18775 -25228
rect -18636 -25377 -18575 -25228
rect -18396 -25342 -18362 -25186
rect -18298 -25342 -18264 -25234
rect -18200 -25342 -18166 -25186
rect -18102 -25342 -18068 -25234
rect -17802 -25331 -17732 -24936
rect -17397 -24946 -17242 -24936
rect -17155 -24913 -17112 -24843
rect -17155 -24968 -16974 -24913
rect -17155 -24980 -17112 -24968
rect -17562 -25018 -17308 -24982
rect -18514 -25377 -18441 -25371
rect -18636 -25390 -18441 -25377
rect -18614 -25418 -18441 -25390
rect -18514 -25431 -18441 -25418
rect -18004 -25401 -17726 -25331
rect -18396 -25573 -18362 -25465
rect -18200 -25573 -18166 -25465
rect -18004 -25573 -17970 -25401
rect -17562 -25077 -17520 -25018
rect -22658 -25792 -21770 -25686
rect -17558 -25661 -17524 -25077
rect -17350 -25071 -17308 -25018
rect -17253 -25019 -17112 -24980
rect -17347 -25653 -17313 -25071
rect -17253 -25073 -17211 -25019
rect -17351 -25695 -17309 -25653
rect -17249 -25661 -17215 -25073
rect -17151 -25651 -17117 -25053
rect -16940 -25067 -16897 -24823
rect -16134 -24876 -15997 -24823
rect -16714 -24998 -16609 -24926
rect -15258 -24038 -15210 -23666
rect -15139 -23859 -15105 -23700
rect -15047 -23716 -15001 -23623
rect -15041 -23808 -15007 -23716
rect -14943 -23859 -14909 -23700
rect -14851 -23716 -14805 -23623
rect -14655 -23655 -14522 -23623
rect -14845 -23808 -14811 -23716
rect -14747 -23859 -14713 -23700
rect -14655 -23716 -14609 -23655
rect -14486 -23666 -14246 -23604
rect -14210 -23623 -13644 -23585
rect -14649 -23808 -14615 -23716
rect -14486 -23810 -14426 -23666
rect -14302 -23859 -14268 -23700
rect -14210 -23716 -14164 -23623
rect -14204 -23808 -14170 -23716
rect -14106 -23859 -14072 -23700
rect -14014 -23716 -13968 -23623
rect -13818 -23655 -13644 -23623
rect -13599 -23567 -13552 -23420
rect -13495 -23427 -13461 -23335
rect -13398 -23356 -13356 -23301
rect -13496 -23479 -13460 -23427
rect -13397 -23443 -13363 -23356
rect -13299 -23425 -13265 -23335
rect -13204 -23357 -13162 -23301
rect -13299 -23443 -13262 -23425
rect -13201 -23443 -13167 -23357
rect -13103 -23425 -13069 -23335
rect -13008 -23352 -12966 -23301
rect -13298 -23479 -13262 -23443
rect -13104 -23479 -13068 -23425
rect -13005 -23443 -12971 -23352
rect -12907 -23435 -12873 -23335
rect -12910 -23479 -12868 -23435
rect -13496 -23513 -12868 -23479
rect -13599 -23641 -13427 -23567
rect -13043 -23620 -12868 -23513
rect -12341 -23324 -12307 -23320
rect -12347 -23577 -12301 -23324
rect -12145 -23512 -12111 -23320
rect -12151 -23577 -12105 -23512
rect -11949 -23512 -11915 -23320
rect -11725 -23394 -11668 -23342
rect -11873 -23456 -11668 -23394
rect -11955 -23577 -11909 -23512
rect -12347 -23585 -11909 -23577
rect -11873 -23585 -11811 -23456
rect -11725 -23506 -11668 -23456
rect -11504 -23324 -11470 -23320
rect -12551 -23599 -12383 -23592
rect -14008 -23808 -13974 -23716
rect -13910 -23859 -13876 -23700
rect -13818 -23716 -13772 -23655
rect -13812 -23808 -13778 -23716
rect -13599 -23776 -13552 -23641
rect -13043 -23680 -12777 -23620
rect -12573 -23659 -12383 -23599
rect -12551 -23666 -12383 -23659
rect -12347 -23623 -11811 -23585
rect -11510 -23577 -11464 -23324
rect -11308 -23512 -11274 -23320
rect -11314 -23577 -11268 -23512
rect -10894 -23301 -10266 -23267
rect -11112 -23512 -11078 -23320
rect -10894 -23346 -10858 -23301
rect -11118 -23577 -11072 -23512
rect -11510 -23585 -11072 -23577
rect -11017 -23561 -10943 -23393
rect -10893 -23420 -10859 -23346
rect -11017 -23585 -10944 -23561
rect -11714 -23603 -11546 -23592
rect -13499 -23714 -12868 -23680
rect -13499 -23755 -13458 -23714
rect -13593 -23846 -13559 -23776
rect -15148 -23927 -13777 -23859
rect -13598 -23904 -13554 -23846
rect -13495 -23858 -13461 -23755
rect -13397 -23835 -13363 -23750
rect -13301 -23763 -13260 -23714
rect -13402 -23904 -13358 -23835
rect -13299 -23858 -13265 -23763
rect -13201 -23835 -13167 -23750
rect -13107 -23763 -13066 -23714
rect -12910 -23721 -12868 -23714
rect -13206 -23904 -13162 -23835
rect -13103 -23858 -13069 -23763
rect -13005 -23846 -12971 -23750
rect -12910 -23764 -12869 -23721
rect -13009 -23904 -12965 -23846
rect -12907 -23858 -12873 -23764
rect -12439 -23859 -12405 -23700
rect -12347 -23716 -12301 -23623
rect -12341 -23808 -12307 -23716
rect -12243 -23859 -12209 -23700
rect -12151 -23716 -12105 -23623
rect -11955 -23655 -11811 -23623
rect -12145 -23808 -12111 -23716
rect -12047 -23859 -12013 -23700
rect -11955 -23716 -11909 -23655
rect -11774 -23666 -11546 -23603
rect -11510 -23623 -10944 -23585
rect -11949 -23808 -11915 -23716
rect -11774 -23825 -11714 -23666
rect -11602 -23859 -11568 -23700
rect -11510 -23716 -11464 -23623
rect -11504 -23808 -11470 -23716
rect -11406 -23859 -11372 -23700
rect -11314 -23716 -11268 -23623
rect -11118 -23655 -10944 -23623
rect -10899 -23567 -10852 -23420
rect -10795 -23427 -10761 -23335
rect -10698 -23356 -10656 -23301
rect -10796 -23479 -10760 -23427
rect -10697 -23443 -10663 -23356
rect -10599 -23425 -10565 -23335
rect -10504 -23357 -10462 -23301
rect -10599 -23443 -10562 -23425
rect -10501 -23443 -10467 -23357
rect -10403 -23425 -10369 -23335
rect -10308 -23352 -10266 -23301
rect -10598 -23479 -10562 -23443
rect -10404 -23479 -10368 -23425
rect -10305 -23443 -10271 -23352
rect -10207 -23435 -10173 -23335
rect -10210 -23479 -10168 -23435
rect -10796 -23513 -10168 -23479
rect -10899 -23641 -10727 -23567
rect -10343 -23622 -10168 -23513
rect -11308 -23808 -11274 -23716
rect -11210 -23859 -11176 -23700
rect -11118 -23716 -11072 -23655
rect -11112 -23808 -11078 -23716
rect -10899 -23776 -10852 -23641
rect -10343 -23680 -10093 -23622
rect -10799 -23682 -10093 -23680
rect -10799 -23714 -10168 -23682
rect -10799 -23755 -10758 -23714
rect -10893 -23846 -10859 -23776
rect -14900 -23967 -14789 -23927
rect -14911 -23975 -14774 -23967
rect -14089 -23975 -13978 -23927
rect -13598 -23938 -12965 -23904
rect -12448 -23861 -11914 -23859
rect -11611 -23861 -11077 -23859
rect -12448 -23927 -11077 -23861
rect -10898 -23904 -10854 -23846
rect -10795 -23858 -10761 -23755
rect -10697 -23835 -10663 -23750
rect -10601 -23763 -10560 -23714
rect -10702 -23904 -10658 -23835
rect -10599 -23858 -10565 -23763
rect -10501 -23835 -10467 -23750
rect -10407 -23763 -10366 -23714
rect -10210 -23721 -10168 -23714
rect -10506 -23904 -10462 -23835
rect -10403 -23858 -10369 -23763
rect -10305 -23846 -10271 -23750
rect -10210 -23764 -10169 -23721
rect -10309 -23904 -10265 -23846
rect -10207 -23858 -10173 -23764
rect -12291 -23973 -12180 -23927
rect -12108 -23929 -11588 -23927
rect -12314 -23975 -12177 -23973
rect -11413 -23975 -11302 -23927
rect -10898 -23938 -10265 -23904
rect -8848 -23931 -8814 -23337
rect -8642 -23303 -8402 -23269
rect -8642 -23347 -8600 -23303
rect -9676 -23975 -9544 -23973
rect -14928 -24014 -9543 -23975
rect -14911 -24027 -14774 -24014
rect -12314 -24033 -12177 -24014
rect -9676 -24033 -9544 -24014
rect -15259 -24175 -15199 -24038
rect -12749 -24067 -12612 -24056
rect -11803 -24067 -11671 -24057
rect -14928 -24106 -9198 -24067
rect -12749 -24116 -12612 -24106
rect -11803 -24117 -11671 -24106
rect -14522 -24153 -14390 -24145
rect -9999 -24153 -9867 -24143
rect -15258 -24533 -15210 -24175
rect -14928 -24192 -9867 -24153
rect -14522 -24205 -14390 -24192
rect -9999 -24203 -9867 -24192
rect -9237 -24175 -9198 -24106
rect -8856 -24175 -8813 -23931
rect -8636 -23945 -8602 -23347
rect -8538 -23925 -8504 -23337
rect -8444 -23345 -8402 -23303
rect -8542 -23979 -8500 -23925
rect -8440 -23927 -8406 -23345
rect -8641 -24018 -8500 -23979
rect -8445 -23980 -8403 -23927
rect -8229 -23921 -8195 -23337
rect -8233 -23980 -8191 -23921
rect -2055 -22543 7804 -22282
rect 17473 -21915 17514 -21864
rect -2055 -23401 -1757 -22543
rect -446 -23401 -185 -22543
rect 391 -23401 652 -22543
rect 1431 -23401 1692 -22543
rect 2889 -23401 3150 -22543
rect 4103 -23401 4364 -22543
rect 6049 -23401 6310 -22543
rect 7543 -23401 7804 -22543
rect 17477 -22506 17511 -21915
rect 17684 -21908 17726 -21864
rect 17689 -22506 17723 -21908
rect 17787 -22500 17821 -21898
rect 17880 -21909 17922 -21864
rect 18092 -21860 18260 -21818
rect 17777 -22542 17830 -22500
rect 17885 -22506 17919 -21909
rect 17998 -22500 18032 -21898
rect 18092 -21916 18134 -21860
rect 17986 -22542 18042 -22500
rect 18096 -22506 18130 -21916
rect 18194 -22500 18228 -21898
rect 18184 -22542 18240 -22500
rect 17777 -22576 18240 -22542
rect -8445 -24016 -8191 -23980
rect -8641 -24030 -8598 -24018
rect -8779 -24085 -8598 -24030
rect -8641 -24155 -8598 -24085
rect -8511 -24062 -8356 -24052
rect -7998 -24062 -7866 -24010
rect -8511 -24098 -7866 -24062
rect -8511 -24107 -8356 -24098
rect -9237 -24215 -8679 -24175
rect -8641 -24195 -8287 -24155
rect -9237 -24218 -8727 -24215
rect -15140 -24307 -14606 -24239
rect -14209 -24262 -13576 -24228
rect -15139 -24450 -15105 -24358
rect -15145 -24511 -15099 -24450
rect -15041 -24466 -15007 -24307
rect -14943 -24450 -14909 -24358
rect -15175 -24533 -15099 -24511
rect -15258 -24543 -15099 -24533
rect -14949 -24543 -14903 -24450
rect -14845 -24466 -14811 -24307
rect -14747 -24450 -14713 -24358
rect -14753 -24543 -14707 -24450
rect -14649 -24466 -14615 -24307
rect -14301 -24402 -14267 -24308
rect -14209 -24320 -14165 -24262
rect -14305 -24445 -14264 -24402
rect -14203 -24416 -14169 -24320
rect -14105 -24403 -14071 -24308
rect -14012 -24331 -13968 -24262
rect -14306 -24452 -14264 -24445
rect -14108 -24452 -14067 -24403
rect -14007 -24416 -13973 -24331
rect -13909 -24403 -13875 -24308
rect -13816 -24331 -13772 -24262
rect -13914 -24452 -13873 -24403
rect -13811 -24416 -13777 -24331
rect -13713 -24411 -13679 -24308
rect -13620 -24320 -13576 -24262
rect -13397 -24307 -11906 -24239
rect -11509 -24262 -10876 -24228
rect -13615 -24390 -13581 -24320
rect -13716 -24452 -13675 -24411
rect -14306 -24486 -13675 -24452
rect -15258 -24570 -14707 -24543
rect -15257 -24572 -14707 -24570
rect -15175 -24581 -14707 -24572
rect -14671 -24515 -14503 -24500
rect -14306 -24515 -14131 -24486
rect -14671 -24568 -14131 -24515
rect -13622 -24525 -13575 -24390
rect -13396 -24450 -13362 -24358
rect -13402 -24511 -13356 -24450
rect -13298 -24466 -13264 -24307
rect -13200 -24450 -13166 -24358
rect -14671 -24574 -14503 -24568
rect -15145 -24589 -14707 -24581
rect -15145 -24654 -15099 -24589
rect -15139 -24846 -15105 -24654
rect -14949 -24654 -14903 -24589
rect -14943 -24846 -14909 -24654
rect -14753 -24842 -14707 -24589
rect -14747 -24846 -14713 -24842
rect -14306 -24653 -14131 -24568
rect -13747 -24599 -13575 -24525
rect -14306 -24687 -13678 -24653
rect -14306 -24731 -14264 -24687
rect -14301 -24831 -14267 -24731
rect -14203 -24814 -14169 -24723
rect -14106 -24741 -14070 -24687
rect -13912 -24723 -13876 -24687
rect -14208 -24865 -14166 -24814
rect -14105 -24831 -14071 -24741
rect -14007 -24809 -13973 -24723
rect -13912 -24741 -13875 -24723
rect -14012 -24865 -13970 -24809
rect -13909 -24831 -13875 -24741
rect -13811 -24810 -13777 -24723
rect -13714 -24739 -13678 -24687
rect -13818 -24865 -13776 -24810
rect -13713 -24831 -13679 -24739
rect -13622 -24746 -13575 -24599
rect -13530 -24543 -13356 -24511
rect -13206 -24543 -13160 -24450
rect -13102 -24466 -13068 -24307
rect -13004 -24450 -12970 -24358
rect -13010 -24543 -12964 -24450
rect -12906 -24466 -12872 -24307
rect -13530 -24581 -12964 -24543
rect -12928 -24505 -12760 -24500
rect -12700 -24505 -12640 -24432
rect -12928 -24563 -12640 -24505
rect -12585 -24522 -12525 -24407
rect -12439 -24450 -12405 -24358
rect -12445 -24511 -12399 -24450
rect -12341 -24466 -12307 -24307
rect -12243 -24450 -12209 -24358
rect -12475 -24522 -12399 -24511
rect -12928 -24574 -12760 -24563
rect -12700 -24564 -12640 -24563
rect -12590 -24543 -12399 -24522
rect -12249 -24543 -12203 -24450
rect -12145 -24466 -12111 -24307
rect -12047 -24450 -12013 -24358
rect -12053 -24543 -12007 -24450
rect -11949 -24466 -11915 -24307
rect -11604 -24402 -11558 -24280
rect -11509 -24320 -11465 -24262
rect -11605 -24412 -11558 -24402
rect -11605 -24445 -11564 -24412
rect -11503 -24416 -11469 -24320
rect -11405 -24403 -11371 -24308
rect -11312 -24331 -11268 -24262
rect -11606 -24452 -11564 -24445
rect -11408 -24452 -11367 -24403
rect -11307 -24416 -11273 -24331
rect -11209 -24403 -11175 -24308
rect -11116 -24331 -11072 -24262
rect -11214 -24452 -11173 -24403
rect -11111 -24416 -11077 -24331
rect -11013 -24411 -10979 -24308
rect -10920 -24320 -10876 -24262
rect -10697 -24307 -9281 -24239
rect -10915 -24390 -10881 -24320
rect -11016 -24452 -10975 -24411
rect -11606 -24486 -10975 -24452
rect -12590 -24567 -12007 -24543
rect -13530 -24605 -13457 -24581
rect -13615 -24820 -13581 -24746
rect -13531 -24773 -13457 -24605
rect -13402 -24589 -12964 -24581
rect -13402 -24654 -13356 -24589
rect -13616 -24865 -13580 -24820
rect -13396 -24846 -13362 -24654
rect -14208 -24899 -13580 -24865
rect -13206 -24654 -13160 -24589
rect -13200 -24846 -13166 -24654
rect -13010 -24842 -12964 -24589
rect -13004 -24846 -12970 -24842
rect -12806 -24701 -12749 -24660
rect -12590 -24701 -12545 -24567
rect -12475 -24581 -12007 -24567
rect -11971 -24508 -11803 -24500
rect -11606 -24508 -11431 -24486
rect -11971 -24565 -11431 -24508
rect -10922 -24525 -10875 -24390
rect -10696 -24450 -10662 -24358
rect -10702 -24511 -10656 -24450
rect -10598 -24466 -10564 -24307
rect -10500 -24450 -10466 -24358
rect -11971 -24574 -11803 -24565
rect -12445 -24589 -12007 -24581
rect -12445 -24654 -12399 -24589
rect -12806 -24746 -12545 -24701
rect -12806 -24824 -12749 -24746
rect -12439 -24846 -12405 -24654
rect -12249 -24654 -12203 -24589
rect -12243 -24846 -12209 -24654
rect -12053 -24842 -12007 -24589
rect -12047 -24846 -12013 -24842
rect -11606 -24653 -11431 -24565
rect -11047 -24599 -10875 -24525
rect -11606 -24687 -10978 -24653
rect -11606 -24731 -11564 -24687
rect -11601 -24831 -11567 -24731
rect -11503 -24814 -11469 -24723
rect -11406 -24741 -11370 -24687
rect -11212 -24723 -11176 -24687
rect -11508 -24865 -11466 -24814
rect -11405 -24831 -11371 -24741
rect -11307 -24809 -11273 -24723
rect -11212 -24741 -11175 -24723
rect -11312 -24865 -11270 -24809
rect -11209 -24831 -11175 -24741
rect -11111 -24810 -11077 -24723
rect -11014 -24739 -10978 -24687
rect -11118 -24865 -11076 -24810
rect -11013 -24831 -10979 -24739
rect -10922 -24746 -10875 -24599
rect -10830 -24543 -10656 -24511
rect -10506 -24543 -10460 -24450
rect -10402 -24466 -10368 -24307
rect -10304 -24450 -10270 -24358
rect -10310 -24543 -10264 -24450
rect -10206 -24466 -10172 -24307
rect -10830 -24581 -10264 -24543
rect -10228 -24505 -10060 -24500
rect -10228 -24517 -10025 -24505
rect -9968 -24517 -9908 -24431
rect -9814 -24450 -9780 -24358
rect -9820 -24511 -9774 -24450
rect -9716 -24466 -9682 -24307
rect -9618 -24450 -9584 -24358
rect -9850 -24517 -9774 -24511
rect -10228 -24543 -9774 -24517
rect -9624 -24543 -9578 -24450
rect -9520 -24466 -9486 -24307
rect -9422 -24450 -9388 -24358
rect -9428 -24543 -9382 -24450
rect -9324 -24466 -9290 -24307
rect -9237 -24500 -9198 -24218
rect -8771 -24258 -8727 -24218
rect -10228 -24559 -9382 -24543
rect -10228 -24563 -10025 -24559
rect -9968 -24563 -9908 -24559
rect -10228 -24574 -10060 -24563
rect -9850 -24581 -9382 -24559
rect -9346 -24574 -9178 -24500
rect -8765 -24557 -8731 -24258
rect -8667 -24532 -8633 -24249
rect -10830 -24605 -10757 -24581
rect -10915 -24820 -10881 -24746
rect -10831 -24773 -10757 -24605
rect -10702 -24589 -10264 -24581
rect -10702 -24654 -10656 -24589
rect -10916 -24865 -10880 -24820
rect -10696 -24846 -10662 -24654
rect -11508 -24899 -10880 -24865
rect -10506 -24654 -10460 -24589
rect -10500 -24846 -10466 -24654
rect -10310 -24842 -10264 -24589
rect -9820 -24589 -9382 -24581
rect -10304 -24846 -10270 -24842
rect -9820 -24654 -9774 -24589
rect -10106 -24824 -10049 -24660
rect -9814 -24846 -9780 -24654
rect -9624 -24654 -9578 -24589
rect -9618 -24846 -9584 -24654
rect -9428 -24842 -9382 -24589
rect -9422 -24846 -9388 -24842
rect -8673 -24662 -8626 -24532
rect -8425 -24542 -8391 -24249
rect -8332 -24265 -8287 -24195
rect -8241 -24169 -8086 -24160
rect -7723 -24169 -7581 -24152
rect -8241 -24203 -7581 -24169
rect -8241 -24215 -8086 -24203
rect -7723 -24216 -7581 -24203
rect -8431 -24662 -8384 -24542
rect -8327 -24557 -8293 -24265
rect -8229 -24543 -8195 -24249
rect -8235 -24662 -8188 -24543
rect -7724 -24662 -7619 -24656
rect -8853 -24744 -7619 -24662
rect -7724 -24751 -7619 -24744
rect -17153 -25695 -17111 -25651
rect -17351 -25729 -17111 -25695
rect -16939 -25661 -16905 -25067
rect -22658 -25819 -21854 -25792
rect -22871 -26262 -21888 -26231
rect -22871 -26327 -21593 -26262
rect -22871 -26346 -21888 -26327
rect -22855 -27431 -22821 -26515
rect -22757 -26723 -22723 -26346
rect -22344 -26417 -21903 -26383
rect -22442 -26887 -22408 -26515
rect -22344 -26823 -22310 -26417
rect -22134 -26420 -21903 -26417
rect -22246 -26887 -22212 -26515
rect -22134 -26526 -22099 -26420
rect -22133 -26823 -22099 -26526
rect -22035 -26823 -22001 -26515
rect -21938 -26524 -21903 -26420
rect -21937 -26823 -21903 -26524
rect -22036 -26886 -22001 -26823
rect -21823 -26886 -21789 -26516
rect -21725 -26824 -21691 -26327
rect -22036 -26887 -21789 -26886
rect -21627 -26887 -21593 -26516
rect -22442 -26921 -22209 -26887
rect -22036 -26921 -21593 -26887
rect -22786 -26975 -22651 -26968
rect -22246 -26975 -22209 -26921
rect -22786 -27012 -22209 -26975
rect -22786 -27022 -22651 -27012
rect -22246 -27150 -22209 -27012
rect -22175 -26977 -22040 -26970
rect -21546 -26977 -21488 -26874
rect -22175 -27011 -21488 -26977
rect -22175 -27024 -22040 -27011
rect -21987 -27055 -21852 -27048
rect -20816 -27055 -20758 -26956
rect -18979 -26501 -18945 -26293
rect -18783 -26501 -18749 -26293
rect -18587 -26501 -18553 -26293
rect -18006 -26508 -17972 -26164
rect -17810 -26508 -17776 -26164
rect -17397 -26271 -17363 -26163
rect -17201 -26271 -17167 -26163
rect -17515 -26318 -17442 -26305
rect -17615 -26346 -17442 -26318
rect -17637 -26359 -17442 -26346
rect -17637 -26508 -17576 -26359
rect -17515 -26365 -17442 -26359
rect -17005 -26335 -16971 -26163
rect -16703 -26335 -16633 -24998
rect -7167 -23591 -7133 -23587
rect -7173 -23844 -7127 -23591
rect -6971 -23779 -6937 -23587
rect -6977 -23844 -6931 -23779
rect -6775 -23779 -6741 -23587
rect -6551 -23673 -6494 -23609
rect -6694 -23722 -6494 -23673
rect -6781 -23844 -6735 -23779
rect -7173 -23852 -6735 -23844
rect -6694 -23852 -6648 -23722
rect -6551 -23773 -6494 -23722
rect -6330 -23591 -6296 -23587
rect -7377 -23889 -7209 -23859
rect -7384 -23933 -7209 -23889
rect -7173 -23890 -6648 -23852
rect -6336 -23844 -6290 -23591
rect -6134 -23779 -6100 -23587
rect -6140 -23844 -6094 -23779
rect -5720 -23568 -5092 -23534
rect -5938 -23779 -5904 -23587
rect -5720 -23613 -5684 -23568
rect -5944 -23844 -5898 -23779
rect -6336 -23852 -5898 -23844
rect -5843 -23828 -5769 -23660
rect -5719 -23687 -5685 -23613
rect -5843 -23852 -5770 -23828
rect -6540 -23870 -6372 -23859
rect -6575 -23871 -6372 -23870
rect -7384 -24305 -7336 -23933
rect -7265 -24126 -7231 -23967
rect -7173 -23983 -7127 -23890
rect -7167 -24075 -7133 -23983
rect -7069 -24126 -7035 -23967
rect -6977 -23983 -6931 -23890
rect -6781 -23922 -6648 -23890
rect -6971 -24075 -6937 -23983
rect -6873 -24126 -6839 -23967
rect -6781 -23983 -6735 -23922
rect -6612 -23933 -6372 -23871
rect -6336 -23890 -5770 -23852
rect -6775 -24075 -6741 -23983
rect -6612 -24077 -6552 -23933
rect -6428 -24126 -6394 -23967
rect -6336 -23983 -6290 -23890
rect -6330 -24075 -6296 -23983
rect -6232 -24126 -6198 -23967
rect -6140 -23983 -6094 -23890
rect -5944 -23922 -5770 -23890
rect -5725 -23834 -5678 -23687
rect -5621 -23694 -5587 -23602
rect -5524 -23623 -5482 -23568
rect -5622 -23746 -5586 -23694
rect -5523 -23710 -5489 -23623
rect -5425 -23692 -5391 -23602
rect -5330 -23624 -5288 -23568
rect -5425 -23710 -5388 -23692
rect -5327 -23710 -5293 -23624
rect -5229 -23692 -5195 -23602
rect -5134 -23619 -5092 -23568
rect -5424 -23746 -5388 -23710
rect -5230 -23746 -5194 -23692
rect -5131 -23710 -5097 -23619
rect -5033 -23702 -4999 -23602
rect -5036 -23746 -4994 -23702
rect -5622 -23780 -4994 -23746
rect -5725 -23908 -5553 -23834
rect -5169 -23887 -4994 -23780
rect -4467 -23591 -4433 -23587
rect -4473 -23844 -4427 -23591
rect -4271 -23779 -4237 -23587
rect -4277 -23844 -4231 -23779
rect -4075 -23779 -4041 -23587
rect -3851 -23661 -3794 -23609
rect -3999 -23723 -3794 -23661
rect -4081 -23844 -4035 -23779
rect -4473 -23852 -4035 -23844
rect -3999 -23852 -3937 -23723
rect -3851 -23773 -3794 -23723
rect -3630 -23591 -3596 -23587
rect -4677 -23866 -4509 -23859
rect -6134 -24075 -6100 -23983
rect -6036 -24126 -6002 -23967
rect -5944 -23983 -5898 -23922
rect -5938 -24075 -5904 -23983
rect -5725 -24043 -5678 -23908
rect -5169 -23947 -4903 -23887
rect -4699 -23926 -4509 -23866
rect -4677 -23933 -4509 -23926
rect -4473 -23890 -3937 -23852
rect -3636 -23844 -3590 -23591
rect -3434 -23779 -3400 -23587
rect -3440 -23844 -3394 -23779
rect -3020 -23568 -2392 -23534
rect -3238 -23779 -3204 -23587
rect -3020 -23613 -2984 -23568
rect -3244 -23844 -3198 -23779
rect -3636 -23852 -3198 -23844
rect -3143 -23828 -3069 -23660
rect -3019 -23687 -2985 -23613
rect -3143 -23852 -3070 -23828
rect -3840 -23870 -3672 -23859
rect -5625 -23981 -4994 -23947
rect -5625 -24022 -5584 -23981
rect -5719 -24113 -5685 -24043
rect -7274 -24194 -5903 -24126
rect -5724 -24171 -5680 -24113
rect -5621 -24125 -5587 -24022
rect -5523 -24102 -5489 -24017
rect -5427 -24030 -5386 -23981
rect -5528 -24171 -5484 -24102
rect -5425 -24125 -5391 -24030
rect -5327 -24102 -5293 -24017
rect -5233 -24030 -5192 -23981
rect -5036 -23988 -4994 -23981
rect -5332 -24171 -5288 -24102
rect -5229 -24125 -5195 -24030
rect -5131 -24113 -5097 -24017
rect -5036 -24031 -4995 -23988
rect -5135 -24171 -5091 -24113
rect -5033 -24125 -4999 -24031
rect -4565 -24126 -4531 -23967
rect -4473 -23983 -4427 -23890
rect -4467 -24075 -4433 -23983
rect -4369 -24126 -4335 -23967
rect -4277 -23983 -4231 -23890
rect -4081 -23922 -3937 -23890
rect -4271 -24075 -4237 -23983
rect -4173 -24126 -4139 -23967
rect -4081 -23983 -4035 -23922
rect -3900 -23933 -3672 -23870
rect -3636 -23890 -3070 -23852
rect -4075 -24075 -4041 -23983
rect -3900 -24092 -3840 -23933
rect -3728 -24126 -3694 -23967
rect -3636 -23983 -3590 -23890
rect -3630 -24075 -3596 -23983
rect -3532 -24126 -3498 -23967
rect -3440 -23983 -3394 -23890
rect -3244 -23922 -3070 -23890
rect -3025 -23834 -2978 -23687
rect -2921 -23694 -2887 -23602
rect -2824 -23623 -2782 -23568
rect -2922 -23746 -2886 -23694
rect -2823 -23710 -2789 -23623
rect -2725 -23692 -2691 -23602
rect -2630 -23624 -2588 -23568
rect -2725 -23710 -2688 -23692
rect -2627 -23710 -2593 -23624
rect -2529 -23692 -2495 -23602
rect -2434 -23619 -2392 -23568
rect -2724 -23746 -2688 -23710
rect -2530 -23746 -2494 -23692
rect -2431 -23710 -2397 -23619
rect -2333 -23702 -2299 -23602
rect -2055 -23662 7804 -23401
rect 13550 -23274 14064 -23111
rect 15310 -23274 15531 -23246
rect 13550 -23404 15531 -23274
rect 13550 -23536 14064 -23404
rect -2336 -23746 -2294 -23702
rect -2922 -23780 -2294 -23746
rect -3025 -23908 -2853 -23834
rect -2469 -23889 -2294 -23780
rect -3434 -24075 -3400 -23983
rect -3336 -24126 -3302 -23967
rect -3244 -23983 -3198 -23922
rect -3238 -24075 -3204 -23983
rect -3025 -24043 -2978 -23908
rect -2469 -23947 -2219 -23889
rect -2925 -23949 -2219 -23947
rect -2925 -23981 -2294 -23949
rect -2925 -24022 -2884 -23981
rect -3019 -24113 -2985 -24043
rect -7026 -24234 -6915 -24194
rect -7037 -24242 -6900 -24234
rect -6215 -24242 -6104 -24194
rect -5724 -24205 -5091 -24171
rect -4574 -24128 -4040 -24126
rect -3737 -24128 -3203 -24126
rect -4574 -24194 -3203 -24128
rect -3024 -24171 -2980 -24113
rect -2921 -24125 -2887 -24022
rect -2823 -24102 -2789 -24017
rect -2727 -24030 -2686 -23981
rect -2828 -24171 -2784 -24102
rect -2725 -24125 -2691 -24030
rect -2627 -24102 -2593 -24017
rect -2533 -24030 -2492 -23981
rect -2336 -23988 -2294 -23981
rect -2632 -24171 -2588 -24102
rect -2529 -24125 -2495 -24030
rect -2431 -24113 -2397 -24017
rect -2336 -24031 -2295 -23988
rect -2435 -24171 -2391 -24113
rect -2333 -24125 -2299 -24031
rect -4417 -24240 -4306 -24194
rect -4234 -24196 -3714 -24194
rect -4440 -24242 -4303 -24240
rect -3539 -24242 -3428 -24194
rect -3024 -24205 -2391 -24171
rect -2055 -24240 -1757 -23662
rect -1009 -23927 -879 -23662
rect -703 -23927 -573 -23662
rect -386 -23927 -256 -23662
rect 60 -23927 190 -23662
rect -1022 -23992 252 -23927
rect -2055 -24242 -1670 -24240
rect -7054 -24281 -1669 -24242
rect -7037 -24294 -6900 -24281
rect -4440 -24300 -4303 -24281
rect -1802 -24300 -1670 -24281
rect -7385 -24442 -7325 -24305
rect -4875 -24334 -4738 -24323
rect -3929 -24334 -3797 -24324
rect -7054 -24373 -1324 -24334
rect -4875 -24383 -4738 -24373
rect -3929 -24384 -3797 -24373
rect -6648 -24420 -6516 -24412
rect -2125 -24420 -1993 -24410
rect -7384 -24800 -7336 -24442
rect -7054 -24459 -1993 -24420
rect -6648 -24472 -6516 -24459
rect -2125 -24470 -1993 -24459
rect -7266 -24574 -6732 -24506
rect -6335 -24529 -5702 -24495
rect -7265 -24717 -7231 -24625
rect -7271 -24778 -7225 -24717
rect -7167 -24733 -7133 -24574
rect -7069 -24717 -7035 -24625
rect -7301 -24800 -7225 -24778
rect -7384 -24810 -7225 -24800
rect -7075 -24810 -7029 -24717
rect -6971 -24733 -6937 -24574
rect -6873 -24717 -6839 -24625
rect -6879 -24810 -6833 -24717
rect -6775 -24733 -6741 -24574
rect -6427 -24669 -6393 -24575
rect -6335 -24587 -6291 -24529
rect -6431 -24712 -6390 -24669
rect -6329 -24683 -6295 -24587
rect -6231 -24670 -6197 -24575
rect -6138 -24598 -6094 -24529
rect -6432 -24719 -6390 -24712
rect -6234 -24719 -6193 -24670
rect -6133 -24683 -6099 -24598
rect -6035 -24670 -6001 -24575
rect -5942 -24598 -5898 -24529
rect -6040 -24719 -5999 -24670
rect -5937 -24683 -5903 -24598
rect -5839 -24678 -5805 -24575
rect -5746 -24587 -5702 -24529
rect -5523 -24574 -4032 -24506
rect -3635 -24529 -3002 -24495
rect -5741 -24657 -5707 -24587
rect -5842 -24719 -5801 -24678
rect -6432 -24753 -5801 -24719
rect -7384 -24837 -6833 -24810
rect -7383 -24839 -6833 -24837
rect -7301 -24848 -6833 -24839
rect -6797 -24782 -6629 -24767
rect -6432 -24782 -6257 -24753
rect -6797 -24835 -6257 -24782
rect -5748 -24792 -5701 -24657
rect -5522 -24717 -5488 -24625
rect -5528 -24778 -5482 -24717
rect -5424 -24733 -5390 -24574
rect -5326 -24717 -5292 -24625
rect -6797 -24841 -6629 -24835
rect -7271 -24856 -6833 -24848
rect -7271 -24921 -7225 -24856
rect -7265 -25113 -7231 -24921
rect -7075 -24921 -7029 -24856
rect -7069 -25113 -7035 -24921
rect -6879 -25109 -6833 -24856
rect -6873 -25113 -6839 -25109
rect -6432 -24920 -6257 -24835
rect -5873 -24866 -5701 -24792
rect -6432 -24954 -5804 -24920
rect -6432 -24998 -6390 -24954
rect -6427 -25098 -6393 -24998
rect -6329 -25081 -6295 -24990
rect -6232 -25008 -6196 -24954
rect -6038 -24990 -6002 -24954
rect -6334 -25132 -6292 -25081
rect -6231 -25098 -6197 -25008
rect -6133 -25076 -6099 -24990
rect -6038 -25008 -6001 -24990
rect -6138 -25132 -6096 -25076
rect -6035 -25098 -6001 -25008
rect -5937 -25077 -5903 -24990
rect -5840 -25006 -5804 -24954
rect -5944 -25132 -5902 -25077
rect -5839 -25098 -5805 -25006
rect -5748 -25013 -5701 -24866
rect -5656 -24810 -5482 -24778
rect -5332 -24810 -5286 -24717
rect -5228 -24733 -5194 -24574
rect -5130 -24717 -5096 -24625
rect -5136 -24810 -5090 -24717
rect -5032 -24733 -4998 -24574
rect -5656 -24848 -5090 -24810
rect -5054 -24772 -4886 -24767
rect -4826 -24772 -4766 -24699
rect -5054 -24830 -4766 -24772
rect -4711 -24789 -4651 -24674
rect -4565 -24717 -4531 -24625
rect -4571 -24778 -4525 -24717
rect -4467 -24733 -4433 -24574
rect -4369 -24717 -4335 -24625
rect -4601 -24789 -4525 -24778
rect -5054 -24841 -4886 -24830
rect -4826 -24831 -4766 -24830
rect -4716 -24810 -4525 -24789
rect -4375 -24810 -4329 -24717
rect -4271 -24733 -4237 -24574
rect -4173 -24717 -4139 -24625
rect -4179 -24810 -4133 -24717
rect -4075 -24733 -4041 -24574
rect -3730 -24669 -3684 -24547
rect -3635 -24587 -3591 -24529
rect -3731 -24679 -3684 -24669
rect -3731 -24712 -3690 -24679
rect -3629 -24683 -3595 -24587
rect -3531 -24670 -3497 -24575
rect -3438 -24598 -3394 -24529
rect -3732 -24719 -3690 -24712
rect -3534 -24719 -3493 -24670
rect -3433 -24683 -3399 -24598
rect -3335 -24670 -3301 -24575
rect -3242 -24598 -3198 -24529
rect -3340 -24719 -3299 -24670
rect -3237 -24683 -3203 -24598
rect -3139 -24678 -3105 -24575
rect -3046 -24587 -3002 -24529
rect -2823 -24574 -1407 -24506
rect -3041 -24657 -3007 -24587
rect -3142 -24719 -3101 -24678
rect -3732 -24753 -3101 -24719
rect -4716 -24834 -4133 -24810
rect -5656 -24872 -5583 -24848
rect -5741 -25087 -5707 -25013
rect -5657 -25040 -5583 -24872
rect -5528 -24856 -5090 -24848
rect -5528 -24921 -5482 -24856
rect -5742 -25132 -5706 -25087
rect -5522 -25113 -5488 -24921
rect -6334 -25166 -5706 -25132
rect -5332 -24921 -5286 -24856
rect -5326 -25113 -5292 -24921
rect -5136 -25109 -5090 -24856
rect -5130 -25113 -5096 -25109
rect -4932 -24968 -4875 -24927
rect -4716 -24968 -4671 -24834
rect -4601 -24848 -4133 -24834
rect -4097 -24775 -3929 -24767
rect -3732 -24775 -3557 -24753
rect -4097 -24832 -3557 -24775
rect -3048 -24792 -3001 -24657
rect -2822 -24717 -2788 -24625
rect -2828 -24778 -2782 -24717
rect -2724 -24733 -2690 -24574
rect -2626 -24717 -2592 -24625
rect -4097 -24841 -3929 -24832
rect -4571 -24856 -4133 -24848
rect -4571 -24921 -4525 -24856
rect -4932 -25013 -4671 -24968
rect -4932 -25091 -4875 -25013
rect -4565 -25113 -4531 -24921
rect -4375 -24921 -4329 -24856
rect -4369 -25113 -4335 -24921
rect -4179 -25109 -4133 -24856
rect -4173 -25113 -4139 -25109
rect -3732 -24920 -3557 -24832
rect -3173 -24866 -3001 -24792
rect -3732 -24954 -3104 -24920
rect -3732 -24998 -3690 -24954
rect -3727 -25098 -3693 -24998
rect -3629 -25081 -3595 -24990
rect -3532 -25008 -3496 -24954
rect -3338 -24990 -3302 -24954
rect -3634 -25132 -3592 -25081
rect -3531 -25098 -3497 -25008
rect -3433 -25076 -3399 -24990
rect -3338 -25008 -3301 -24990
rect -3438 -25132 -3396 -25076
rect -3335 -25098 -3301 -25008
rect -3237 -25077 -3203 -24990
rect -3140 -25006 -3104 -24954
rect -3244 -25132 -3202 -25077
rect -3139 -25098 -3105 -25006
rect -3048 -25013 -3001 -24866
rect -2956 -24810 -2782 -24778
rect -2632 -24810 -2586 -24717
rect -2528 -24733 -2494 -24574
rect -2430 -24717 -2396 -24625
rect -2436 -24810 -2390 -24717
rect -2332 -24733 -2298 -24574
rect -2956 -24848 -2390 -24810
rect -2354 -24772 -2186 -24767
rect -2354 -24784 -2151 -24772
rect -2094 -24784 -2034 -24698
rect -1940 -24717 -1906 -24625
rect -1946 -24778 -1900 -24717
rect -1842 -24733 -1808 -24574
rect -1744 -24717 -1710 -24625
rect -1976 -24784 -1900 -24778
rect -2354 -24810 -1900 -24784
rect -1750 -24810 -1704 -24717
rect -1646 -24733 -1612 -24574
rect -1548 -24717 -1514 -24625
rect -1554 -24810 -1508 -24717
rect -1450 -24733 -1416 -24574
rect -1363 -24767 -1324 -24373
rect -1010 -24633 -976 -24180
rect -912 -24388 -878 -23992
rect -499 -24082 -58 -24048
rect -597 -24552 -563 -24180
rect -499 -24488 -465 -24082
rect -289 -24085 -58 -24082
rect -401 -24552 -367 -24180
rect -289 -24191 -254 -24085
rect -288 -24488 -254 -24191
rect -190 -24488 -156 -24180
rect -93 -24189 -58 -24085
rect -92 -24488 -58 -24189
rect -191 -24551 -156 -24488
rect 22 -24551 56 -24181
rect 120 -24489 154 -23992
rect 984 -24142 1135 -23662
rect 1361 -24124 1485 -23662
rect 1691 -24124 1815 -23662
rect 2098 -24104 2234 -24058
rect 1361 -24142 1876 -24124
rect -191 -24552 56 -24551
rect 218 -24552 252 -24181
rect -597 -24586 -364 -24552
rect -191 -24586 252 -24552
rect 984 -24185 1876 -24142
rect 984 -24203 1434 -24185
rect -1161 -24686 -976 -24633
rect -2354 -24826 -1508 -24810
rect -2354 -24830 -2151 -24826
rect -2094 -24830 -2034 -24826
rect -2354 -24841 -2186 -24830
rect -1976 -24848 -1508 -24826
rect -1472 -24841 -1304 -24767
rect -2956 -24872 -2883 -24848
rect -3041 -25087 -3007 -25013
rect -2957 -25040 -2883 -24872
rect -2828 -24856 -2390 -24848
rect -2828 -24921 -2782 -24856
rect -3042 -25132 -3006 -25087
rect -2822 -25113 -2788 -24921
rect -3634 -25166 -3006 -25132
rect -2632 -24921 -2586 -24856
rect -2626 -25113 -2592 -24921
rect -2436 -25109 -2390 -24856
rect -1946 -24856 -1508 -24848
rect -2430 -25113 -2396 -25109
rect -1946 -24921 -1900 -24856
rect -2232 -25091 -2175 -24927
rect -1940 -25113 -1906 -24921
rect -1750 -24921 -1704 -24856
rect -1744 -25113 -1710 -24921
rect -1554 -25109 -1508 -24856
rect -1548 -25113 -1514 -25109
rect -7596 -25536 -7460 -25490
rect -18189 -26521 -18054 -26515
rect -18209 -26523 -18054 -26521
rect -19271 -26548 -19141 -26531
rect -19097 -26548 -19024 -26535
rect -19806 -26554 -19748 -26553
rect -19271 -26554 -19024 -26548
rect -19806 -26589 -19024 -26554
rect -18416 -26559 -18054 -26523
rect -18006 -26538 -17576 -26508
rect -18006 -26546 -17587 -26538
rect -17397 -26550 -17363 -26394
rect -17299 -26502 -17265 -26394
rect -17201 -26550 -17167 -26394
rect -17103 -26502 -17069 -26394
rect -17005 -26405 -16633 -26335
rect -18209 -26561 -18054 -26559
rect -18189 -26569 -18054 -26561
rect -19806 -26622 -19141 -26589
rect -19097 -26595 -19024 -26589
rect -19806 -26690 -19748 -26622
rect -19271 -26681 -19141 -26622
rect -18684 -26619 -18135 -26617
rect -17724 -26619 -17650 -26593
rect -18684 -26623 -17650 -26619
rect -18979 -26879 -18945 -26623
rect -18881 -26831 -18847 -26623
rect -18783 -26879 -18749 -26623
rect -18685 -26657 -17650 -26623
rect -17537 -26636 -16752 -26550
rect -18685 -26831 -18651 -26657
rect -18136 -26658 -17650 -26657
rect -18136 -26659 -18065 -26658
rect -17724 -26664 -17650 -26658
rect -19119 -26965 -18181 -26879
rect -21987 -27093 -20758 -27055
rect -21987 -27102 -21852 -27093
rect -21651 -27139 -21516 -27130
rect -19891 -27139 -19833 -27042
rect -18267 -27046 -18181 -26965
rect -18104 -27009 -18070 -26701
rect -18006 -27009 -17972 -26701
rect -17908 -27009 -17874 -26701
rect -17810 -27009 -17776 -26701
rect -17712 -27009 -17678 -26701
rect -18007 -27046 -17972 -27009
rect -17293 -27043 -17232 -26636
rect -17682 -27046 -17232 -27043
rect -18267 -27104 -17232 -27046
rect -7556 -27067 -7522 -25536
rect -5116 -25609 -4980 -25563
rect -5116 -25862 -5076 -25609
rect -5119 -25998 -5073 -25862
rect -1363 -25390 -1324 -24841
rect -1010 -25096 -976 -24686
rect -941 -24640 -806 -24633
rect -401 -24640 -364 -24586
rect 984 -24610 1045 -24203
rect 1724 -24237 1759 -24185
rect 1430 -24545 1464 -24237
rect 1528 -24545 1562 -24237
rect 1626 -24545 1660 -24237
rect 1724 -24545 1758 -24237
rect 1822 -24545 1856 -24237
rect 1402 -24588 1476 -24582
rect 1817 -24588 1888 -24587
rect 1402 -24589 1888 -24588
rect -941 -24677 -364 -24640
rect -941 -24687 -806 -24677
rect -401 -24815 -364 -24677
rect -330 -24642 -195 -24635
rect -330 -24676 626 -24642
rect -330 -24689 -195 -24676
rect -142 -24720 -7 -24713
rect 421 -24720 557 -24713
rect -142 -24758 557 -24720
rect -142 -24767 -7 -24758
rect 421 -24759 557 -24758
rect -401 -24852 154 -24815
rect 194 -24849 386 -24795
rect 592 -24841 626 -24676
rect 674 -24696 1289 -24610
rect 1402 -24627 2069 -24589
rect 1402 -24653 1476 -24627
rect 1887 -24629 2069 -24627
rect 1806 -24683 1941 -24677
rect 1806 -24687 1971 -24683
rect -272 -25096 -238 -24852
rect -76 -25096 -42 -24852
rect 120 -25096 154 -24852
rect 340 -24933 386 -24849
rect 586 -24911 757 -24841
rect 821 -24852 855 -24744
rect 919 -24852 953 -24696
rect 1017 -24852 1051 -24744
rect 1115 -24852 1149 -24696
rect 1339 -24708 1758 -24700
rect 1328 -24738 1758 -24708
rect 1806 -24723 1993 -24687
rect 1806 -24731 1984 -24723
rect 723 -25083 757 -24911
rect 1194 -24887 1267 -24881
rect 1328 -24887 1389 -24738
rect 1194 -24900 1389 -24887
rect 1194 -24928 1367 -24900
rect 1194 -24941 1267 -24928
rect 919 -25083 953 -24975
rect 1115 -25083 1149 -24975
rect 1528 -25082 1562 -24738
rect 1724 -25082 1758 -24738
rect -1363 -25441 -1226 -25390
rect 1948 -25481 1984 -24731
rect 1829 -25527 1984 -25481
rect 2029 -25565 2069 -24629
rect 2164 -24839 2234 -24104
rect 2589 -24140 2740 -23662
rect 3031 -24122 3182 -23662
rect 3324 -24122 3475 -23662
rect 3964 -23936 4110 -23662
rect 4409 -23936 4555 -23662
rect 4675 -23936 4821 -23662
rect 5035 -23936 5181 -23662
rect 3666 -23992 3802 -23946
rect 3031 -24140 3481 -24122
rect 2589 -24183 3481 -24140
rect 2589 -24201 3039 -24183
rect 2589 -24608 2650 -24201
rect 3329 -24235 3364 -24183
rect 3035 -24543 3069 -24235
rect 3133 -24543 3167 -24235
rect 3231 -24543 3265 -24235
rect 3329 -24543 3363 -24235
rect 3427 -24543 3461 -24235
rect 3736 -24447 3801 -23992
rect 3940 -24001 5214 -23936
rect 3952 -24447 3986 -24189
rect 4050 -24397 4084 -24001
rect 4463 -24091 4904 -24057
rect 3736 -24505 3986 -24447
rect 3007 -24586 3081 -24580
rect 3422 -24586 3493 -24585
rect 3007 -24587 3493 -24586
rect 2279 -24694 2894 -24608
rect 3007 -24625 3697 -24587
rect 3007 -24651 3081 -24625
rect 3492 -24627 3697 -24625
rect 3411 -24683 3546 -24675
rect 3411 -24685 3598 -24683
rect 2164 -24909 2362 -24839
rect 2426 -24850 2460 -24742
rect 2524 -24850 2558 -24694
rect 2622 -24850 2656 -24742
rect 2720 -24850 2754 -24694
rect 2944 -24706 3363 -24698
rect 2933 -24736 3363 -24706
rect 3411 -24723 3618 -24685
rect 3411 -24729 3546 -24723
rect 2328 -25081 2362 -24909
rect 2799 -24885 2872 -24879
rect 2933 -24885 2994 -24736
rect 2799 -24898 2994 -24885
rect 2799 -24926 2972 -24898
rect 2799 -24939 2872 -24926
rect 2524 -25081 2558 -24973
rect 2720 -25081 2754 -24973
rect 3133 -25080 3167 -24736
rect 3329 -25080 3363 -24736
rect 1933 -25611 2069 -25565
rect 3582 -26050 3618 -24723
rect 2097 -26086 3618 -26050
rect 2097 -26198 2133 -26086
rect 3657 -26120 3697 -24627
rect 3952 -25105 3986 -24505
rect 4365 -24561 4399 -24189
rect 4463 -24497 4497 -24091
rect 4673 -24094 4904 -24091
rect 4561 -24561 4595 -24189
rect 4673 -24200 4708 -24094
rect 4674 -24497 4708 -24200
rect 4772 -24497 4806 -24189
rect 4869 -24198 4904 -24094
rect 4870 -24497 4904 -24198
rect 4771 -24560 4806 -24497
rect 4984 -24560 5018 -24190
rect 5082 -24498 5116 -24001
rect 5599 -24116 5796 -23662
rect 6132 -24116 6329 -23662
rect 6645 -24107 6842 -23662
rect 7148 -24107 7345 -23662
rect 7543 -24089 7804 -23662
rect 9088 -23599 9152 -23576
rect 14453 -23599 14536 -23404
rect 15310 -23426 15531 -23404
rect 9088 -23682 14536 -23599
rect 9088 -23694 9152 -23682
rect 18393 -23760 18542 -21225
rect 18608 -21512 18740 -21377
rect 18608 -21847 18714 -21512
rect 18954 -21755 19138 -21225
rect 19578 -21259 19620 -21215
rect 19681 -21223 19715 -21132
rect 19779 -21205 19813 -21115
rect 19872 -21137 19914 -21081
rect 19778 -21259 19814 -21205
rect 19877 -21223 19911 -21137
rect 19975 -21205 20009 -21115
rect 20066 -21136 20108 -21081
rect 19972 -21223 20009 -21205
rect 20073 -21223 20107 -21136
rect 20171 -21207 20205 -21115
rect 20268 -21126 20304 -21081
rect 20269 -21200 20303 -21126
rect 19972 -21259 20008 -21223
rect 20170 -21259 20206 -21207
rect 19578 -21293 20206 -21259
rect 19578 -21402 19753 -21293
rect 20262 -21347 20309 -21200
rect 20353 -21341 20427 -21173
rect 20488 -21292 20522 -21100
rect 19503 -21460 19753 -21402
rect 20137 -21421 20309 -21347
rect 19503 -21462 20209 -21460
rect 19578 -21494 20209 -21462
rect 19578 -21501 19620 -21494
rect 19579 -21544 19620 -21501
rect 19583 -21638 19617 -21544
rect 19681 -21626 19715 -21530
rect 19776 -21543 19817 -21494
rect 19675 -21684 19719 -21626
rect 19779 -21638 19813 -21543
rect 19877 -21615 19911 -21530
rect 19970 -21543 20011 -21494
rect 19872 -21684 19916 -21615
rect 19975 -21638 20009 -21543
rect 20073 -21615 20107 -21530
rect 20168 -21535 20209 -21494
rect 20068 -21684 20112 -21615
rect 20171 -21638 20205 -21535
rect 20262 -21556 20309 -21421
rect 20354 -21365 20427 -21341
rect 20482 -21357 20528 -21292
rect 20684 -21292 20718 -21100
rect 20678 -21357 20724 -21292
rect 20880 -21104 20914 -21100
rect 20874 -21357 20920 -21104
rect 21078 -21174 21135 -21122
rect 21078 -21236 21283 -21174
rect 21078 -21286 21135 -21236
rect 20482 -21365 20920 -21357
rect 20354 -21403 20920 -21365
rect 21221 -21365 21283 -21236
rect 21325 -21292 21359 -21100
rect 21319 -21357 21365 -21292
rect 21521 -21292 21555 -21100
rect 21515 -21357 21561 -21292
rect 21717 -21104 21751 -21100
rect 21711 -21357 21757 -21104
rect 22376 -21081 23004 -21047
rect 22283 -21215 22317 -21115
rect 22376 -21132 22418 -21081
rect 22278 -21259 22320 -21215
rect 22381 -21223 22415 -21132
rect 22479 -21205 22513 -21115
rect 22572 -21137 22614 -21081
rect 22478 -21259 22514 -21205
rect 22577 -21223 22611 -21137
rect 22675 -21205 22709 -21115
rect 22766 -21136 22808 -21081
rect 22672 -21223 22709 -21205
rect 22773 -21223 22807 -21136
rect 22871 -21207 22905 -21115
rect 22968 -21126 23004 -21081
rect 22969 -21200 23003 -21126
rect 22672 -21259 22708 -21223
rect 22870 -21259 22906 -21207
rect 22278 -21293 22906 -21259
rect 21319 -21365 21757 -21357
rect 20354 -21435 20528 -21403
rect 20482 -21496 20528 -21435
rect 20269 -21626 20303 -21556
rect 20488 -21588 20522 -21496
rect 20264 -21684 20308 -21626
rect 20586 -21639 20620 -21480
rect 20678 -21496 20724 -21403
rect 20684 -21588 20718 -21496
rect 20782 -21639 20816 -21480
rect 20874 -21496 20920 -21403
rect 20956 -21383 21124 -21372
rect 20956 -21446 21184 -21383
rect 21221 -21403 21757 -21365
rect 21221 -21435 21365 -21403
rect 20880 -21588 20914 -21496
rect 20978 -21639 21012 -21480
rect 21124 -21605 21184 -21446
rect 21319 -21496 21365 -21435
rect 21325 -21588 21359 -21496
rect 21423 -21639 21457 -21480
rect 21515 -21496 21561 -21403
rect 21521 -21588 21555 -21496
rect 21619 -21639 21653 -21480
rect 21711 -21496 21757 -21403
rect 21793 -21379 21961 -21372
rect 21793 -21439 21983 -21379
rect 22278 -21400 22453 -21293
rect 22962 -21347 23009 -21200
rect 23053 -21341 23127 -21173
rect 23188 -21292 23222 -21100
rect 21793 -21446 21961 -21439
rect 22187 -21460 22453 -21400
rect 22837 -21421 23009 -21347
rect 21717 -21588 21751 -21496
rect 21815 -21639 21849 -21480
rect 22278 -21494 22909 -21460
rect 22278 -21501 22320 -21494
rect 22279 -21544 22320 -21501
rect 22283 -21638 22317 -21544
rect 22381 -21626 22415 -21530
rect 22476 -21543 22517 -21494
rect 19675 -21718 20308 -21684
rect 20487 -21641 21021 -21639
rect 21324 -21641 21858 -21639
rect 20487 -21707 21858 -21641
rect 22375 -21684 22419 -21626
rect 22479 -21638 22513 -21543
rect 22577 -21615 22611 -21530
rect 22670 -21543 22711 -21494
rect 22572 -21684 22616 -21615
rect 22675 -21638 22709 -21543
rect 22773 -21615 22807 -21530
rect 22868 -21535 22909 -21494
rect 22768 -21684 22812 -21615
rect 22871 -21638 22905 -21535
rect 22962 -21556 23009 -21421
rect 23054 -21365 23127 -21341
rect 23182 -21357 23228 -21292
rect 23384 -21292 23418 -21100
rect 23378 -21357 23424 -21292
rect 23580 -21104 23614 -21100
rect 23574 -21357 23620 -21104
rect 23778 -21186 23835 -21122
rect 23778 -21235 23978 -21186
rect 23778 -21286 23835 -21235
rect 23182 -21365 23620 -21357
rect 23054 -21403 23620 -21365
rect 23932 -21365 23978 -21235
rect 24025 -21292 24059 -21100
rect 24019 -21357 24065 -21292
rect 24221 -21292 24255 -21100
rect 24215 -21357 24261 -21292
rect 24417 -21104 24451 -21100
rect 24411 -21357 24457 -21104
rect 28029 -21084 28063 -20740
rect 28225 -21084 28259 -20740
rect 28398 -20889 28459 -20740
rect 28638 -20854 28672 -20698
rect 28736 -20854 28770 -20746
rect 28834 -20854 28868 -20698
rect 35204 -20711 35451 -20670
rect 36286 -20698 36421 -20690
rect 36266 -20700 36421 -20698
rect 35204 -20728 35334 -20711
rect 35378 -20724 35451 -20711
rect 36059 -20736 36421 -20700
rect 36938 -20709 37723 -20623
rect 44067 -20709 44197 -20617
rect 44359 -20675 44393 -20419
rect 44457 -20675 44491 -20467
rect 44555 -20675 44589 -20419
rect 44653 -20641 44687 -20467
rect 45234 -20597 45268 -20289
rect 45332 -20597 45366 -20289
rect 45430 -20597 45464 -20289
rect 45528 -20597 45562 -20289
rect 45626 -20597 45660 -20289
rect 45202 -20640 45273 -20639
rect 45614 -20640 45688 -20634
rect 45202 -20641 45688 -20640
rect 44653 -20675 45688 -20641
rect 46045 -20662 46106 -20255
rect 50800 -20223 51026 -20214
rect 52453 -20223 52699 -20143
rect 50800 -20356 52699 -20223
rect 54269 -20160 54934 -20132
rect 54269 -20218 55304 -20160
rect 54269 -20299 54355 -20218
rect 54529 -20255 54564 -20218
rect 54854 -20221 55304 -20218
rect 50800 -20448 51026 -20356
rect 52453 -20363 52699 -20356
rect 53417 -20385 54355 -20299
rect 44654 -20679 45688 -20675
rect 44654 -20681 45203 -20679
rect 44241 -20709 44314 -20703
rect 45614 -20705 45688 -20679
rect 36266 -20738 36421 -20736
rect 36286 -20744 36421 -20738
rect 36469 -20721 36888 -20713
rect 28932 -20854 28966 -20746
rect 36469 -20751 36899 -20721
rect 28520 -20889 28593 -20883
rect 28398 -20902 28593 -20889
rect 28420 -20930 28593 -20902
rect 28520 -20943 28593 -20930
rect 29030 -20913 29402 -20843
rect 28638 -21085 28672 -20977
rect 28834 -21085 28868 -20977
rect 29030 -21085 29064 -20913
rect 24019 -21365 24457 -21357
rect 23054 -21435 23228 -21403
rect 23182 -21496 23228 -21435
rect 22969 -21626 23003 -21556
rect 23188 -21588 23222 -21496
rect 22964 -21684 23008 -21626
rect 23286 -21639 23320 -21480
rect 23378 -21496 23424 -21403
rect 23384 -21588 23418 -21496
rect 23482 -21639 23516 -21480
rect 23574 -21496 23620 -21403
rect 23656 -21383 23824 -21372
rect 23656 -21384 23859 -21383
rect 23656 -21446 23896 -21384
rect 23932 -21403 24457 -21365
rect 23932 -21435 24065 -21403
rect 23580 -21588 23614 -21496
rect 23678 -21639 23712 -21480
rect 23836 -21590 23896 -21446
rect 24019 -21496 24065 -21435
rect 24025 -21588 24059 -21496
rect 24123 -21639 24157 -21480
rect 24215 -21496 24261 -21403
rect 24221 -21588 24255 -21496
rect 24319 -21639 24353 -21480
rect 24411 -21496 24457 -21403
rect 24493 -21402 24661 -21372
rect 24493 -21446 24668 -21402
rect 24417 -21588 24451 -21496
rect 24515 -21639 24549 -21480
rect 20712 -21755 20823 -21707
rect 20998 -21709 21518 -21707
rect 21590 -21753 21701 -21707
rect 22375 -21718 23008 -21684
rect 23187 -21707 24558 -21639
rect 21587 -21755 21724 -21753
rect 23388 -21755 23499 -21707
rect 24199 -21747 24310 -21707
rect 24184 -21755 24321 -21747
rect 18953 -21794 24338 -21755
rect 18954 -21813 19086 -21794
rect 21587 -21813 21724 -21794
rect 24184 -21807 24321 -21794
rect 24620 -21818 24668 -21446
rect 21081 -21847 21213 -21837
rect 22022 -21847 22159 -21836
rect 18608 -21886 24338 -21847
rect 18608 -22280 18647 -21886
rect 21081 -21897 21213 -21886
rect 22022 -21896 22159 -21886
rect 19277 -21933 19409 -21923
rect 23800 -21933 23932 -21925
rect 19277 -21972 24338 -21933
rect 24609 -21955 24669 -21818
rect 19277 -21983 19409 -21972
rect 23800 -21985 23932 -21972
rect 18691 -22087 20107 -22019
rect 20286 -22042 20919 -22008
rect 18700 -22246 18734 -22087
rect 18798 -22230 18832 -22138
rect 18588 -22354 18756 -22280
rect 18792 -22323 18838 -22230
rect 18896 -22246 18930 -22087
rect 18994 -22230 19028 -22138
rect 18988 -22323 19034 -22230
rect 19092 -22246 19126 -22087
rect 19190 -22230 19224 -22138
rect 19184 -22291 19230 -22230
rect 19184 -22297 19260 -22291
rect 19318 -22297 19378 -22211
rect 19582 -22246 19616 -22087
rect 19680 -22230 19714 -22138
rect 19470 -22285 19638 -22280
rect 19435 -22297 19638 -22285
rect 19184 -22323 19638 -22297
rect 18792 -22339 19638 -22323
rect 18792 -22361 19260 -22339
rect 19318 -22343 19378 -22339
rect 19435 -22343 19638 -22339
rect 19470 -22354 19638 -22343
rect 19674 -22323 19720 -22230
rect 19778 -22246 19812 -22087
rect 19876 -22230 19910 -22138
rect 19870 -22323 19916 -22230
rect 19974 -22246 20008 -22087
rect 20286 -22100 20330 -22042
rect 20072 -22230 20106 -22138
rect 20291 -22170 20325 -22100
rect 20066 -22291 20112 -22230
rect 20066 -22323 20240 -22291
rect 19674 -22361 20240 -22323
rect 18792 -22369 19230 -22361
rect 18792 -22622 18838 -22369
rect 18798 -22626 18832 -22622
rect 18988 -22434 19034 -22369
rect 18994 -22626 19028 -22434
rect 19184 -22434 19230 -22369
rect 19674 -22369 20112 -22361
rect 19190 -22626 19224 -22434
rect 19459 -22604 19516 -22440
rect 19674 -22622 19720 -22369
rect 19680 -22626 19714 -22622
rect 19870 -22434 19916 -22369
rect 19876 -22626 19910 -22434
rect 20066 -22434 20112 -22369
rect 20167 -22385 20240 -22361
rect 20285 -22305 20332 -22170
rect 20389 -22191 20423 -22088
rect 20482 -22111 20526 -22042
rect 20385 -22232 20426 -22191
rect 20487 -22196 20521 -22111
rect 20585 -22183 20619 -22088
rect 20678 -22111 20722 -22042
rect 20583 -22232 20624 -22183
rect 20683 -22196 20717 -22111
rect 20781 -22183 20815 -22088
rect 20875 -22100 20919 -22042
rect 20777 -22232 20818 -22183
rect 20879 -22196 20913 -22100
rect 20968 -22182 21014 -22060
rect 21316 -22087 22807 -22019
rect 22986 -22042 23619 -22008
rect 20968 -22192 21015 -22182
rect 20974 -22225 21015 -22192
rect 20974 -22232 21016 -22225
rect 20385 -22266 21016 -22232
rect 21325 -22246 21359 -22087
rect 21423 -22230 21457 -22138
rect 20841 -22288 21016 -22266
rect 21213 -22288 21381 -22280
rect 20285 -22379 20457 -22305
rect 20841 -22345 21381 -22288
rect 20072 -22626 20106 -22434
rect 20167 -22553 20241 -22385
rect 20285 -22526 20332 -22379
rect 20841 -22433 21016 -22345
rect 21213 -22354 21381 -22345
rect 21417 -22323 21463 -22230
rect 21521 -22246 21555 -22087
rect 21619 -22230 21653 -22138
rect 21613 -22323 21659 -22230
rect 21717 -22246 21751 -22087
rect 21815 -22230 21849 -22138
rect 21809 -22291 21855 -22230
rect 21809 -22302 21885 -22291
rect 21935 -22302 21995 -22187
rect 22050 -22285 22110 -22212
rect 22282 -22246 22316 -22087
rect 22380 -22230 22414 -22138
rect 22170 -22285 22338 -22280
rect 21809 -22323 22000 -22302
rect 21417 -22347 22000 -22323
rect 22050 -22343 22338 -22285
rect 22050 -22344 22110 -22343
rect 21417 -22361 21885 -22347
rect 21417 -22369 21855 -22361
rect 20388 -22467 21016 -22433
rect 20388 -22519 20424 -22467
rect 20586 -22503 20622 -22467
rect 20291 -22600 20325 -22526
rect 20290 -22645 20326 -22600
rect 20389 -22611 20423 -22519
rect 20487 -22590 20521 -22503
rect 20585 -22521 20622 -22503
rect 20486 -22645 20528 -22590
rect 20585 -22611 20619 -22521
rect 20683 -22589 20717 -22503
rect 20780 -22521 20816 -22467
rect 20680 -22645 20722 -22589
rect 20781 -22611 20815 -22521
rect 20879 -22594 20913 -22503
rect 20974 -22511 21016 -22467
rect 20876 -22645 20918 -22594
rect 20977 -22611 21011 -22511
rect 20290 -22679 20918 -22645
rect 21417 -22622 21463 -22369
rect 21423 -22626 21457 -22622
rect 21613 -22434 21659 -22369
rect 21619 -22626 21653 -22434
rect 21809 -22434 21855 -22369
rect 21815 -22626 21849 -22434
rect 21955 -22481 22000 -22347
rect 22170 -22354 22338 -22343
rect 22374 -22323 22420 -22230
rect 22478 -22246 22512 -22087
rect 22576 -22230 22610 -22138
rect 22570 -22323 22616 -22230
rect 22674 -22246 22708 -22087
rect 22986 -22100 23030 -22042
rect 22772 -22230 22806 -22138
rect 22991 -22170 23025 -22100
rect 22766 -22291 22812 -22230
rect 22766 -22323 22940 -22291
rect 22374 -22361 22940 -22323
rect 22374 -22369 22812 -22361
rect 22159 -22481 22216 -22440
rect 21955 -22526 22216 -22481
rect 22159 -22604 22216 -22526
rect 22374 -22622 22420 -22369
rect 22380 -22626 22414 -22622
rect 22570 -22434 22616 -22369
rect 22576 -22626 22610 -22434
rect 22766 -22434 22812 -22369
rect 22867 -22385 22940 -22361
rect 22985 -22305 23032 -22170
rect 23089 -22191 23123 -22088
rect 23182 -22111 23226 -22042
rect 23085 -22232 23126 -22191
rect 23187 -22196 23221 -22111
rect 23285 -22183 23319 -22088
rect 23378 -22111 23422 -22042
rect 23283 -22232 23324 -22183
rect 23383 -22196 23417 -22111
rect 23481 -22183 23515 -22088
rect 23575 -22100 23619 -22042
rect 24016 -22087 24550 -22019
rect 23477 -22232 23518 -22183
rect 23579 -22196 23613 -22100
rect 23677 -22182 23711 -22088
rect 23674 -22225 23715 -22182
rect 23674 -22232 23716 -22225
rect 23085 -22266 23716 -22232
rect 24025 -22246 24059 -22087
rect 24123 -22230 24157 -22138
rect 23541 -22295 23716 -22266
rect 23913 -22295 24081 -22280
rect 22985 -22379 23157 -22305
rect 23541 -22348 24081 -22295
rect 22772 -22626 22806 -22434
rect 22867 -22553 22941 -22385
rect 22985 -22526 23032 -22379
rect 23541 -22433 23716 -22348
rect 23913 -22354 24081 -22348
rect 24117 -22323 24163 -22230
rect 24221 -22246 24255 -22087
rect 24319 -22230 24353 -22138
rect 24313 -22323 24359 -22230
rect 24417 -22246 24451 -22087
rect 24515 -22230 24549 -22138
rect 24509 -22291 24555 -22230
rect 24509 -22313 24585 -22291
rect 24620 -22313 24668 -21955
rect 24509 -22323 24668 -22313
rect 24117 -22350 24668 -22323
rect 24117 -22352 24667 -22350
rect 24117 -22361 24585 -22352
rect 24117 -22369 24555 -22361
rect 23088 -22467 23716 -22433
rect 23088 -22519 23124 -22467
rect 23286 -22503 23322 -22467
rect 22991 -22600 23025 -22526
rect 22990 -22645 23026 -22600
rect 23089 -22611 23123 -22519
rect 23187 -22590 23221 -22503
rect 23285 -22521 23322 -22503
rect 23186 -22645 23228 -22590
rect 23285 -22611 23319 -22521
rect 23383 -22589 23417 -22503
rect 23480 -22521 23516 -22467
rect 23380 -22645 23422 -22589
rect 23481 -22611 23515 -22521
rect 23579 -22594 23613 -22503
rect 23674 -22511 23716 -22467
rect 23576 -22645 23618 -22594
rect 23677 -22611 23711 -22511
rect 22990 -22679 23618 -22645
rect 24117 -22622 24163 -22369
rect 24123 -22626 24157 -22622
rect 24313 -22434 24359 -22369
rect 24319 -22626 24353 -22434
rect 24509 -22434 24555 -22369
rect 24515 -22626 24549 -22434
rect 26198 -21924 26457 -21881
rect 25332 -22035 26457 -21924
rect 27030 -22020 27064 -21676
rect 27226 -22020 27260 -21676
rect 27639 -21783 27673 -21675
rect 27835 -21783 27869 -21675
rect 27521 -21830 27594 -21817
rect 27421 -21858 27594 -21830
rect 27399 -21871 27594 -21858
rect 27399 -22020 27460 -21871
rect 27521 -21877 27594 -21871
rect 28031 -21847 28065 -21675
rect 26847 -22033 26982 -22027
rect 26827 -22035 26982 -22033
rect 25332 -22071 26982 -22035
rect 27030 -22050 27460 -22020
rect 27030 -22058 27449 -22050
rect 27639 -22062 27673 -21906
rect 27737 -22014 27771 -21906
rect 27835 -22062 27869 -21906
rect 27933 -22014 27967 -21906
rect 28031 -21917 28309 -21847
rect 25332 -22129 26457 -22071
rect 26827 -22073 26982 -22071
rect 26847 -22081 26982 -22073
rect 26198 -22144 26457 -22129
rect 26674 -22131 26901 -22129
rect 27312 -22131 27386 -22105
rect 26674 -22169 27386 -22131
rect 27499 -22148 28114 -22062
rect 20723 -22980 20883 -22848
rect 20730 -23163 20865 -22980
rect 20720 -23295 20880 -23163
rect 21243 -23614 21277 -23170
rect 21439 -23614 21473 -23170
rect 21681 -23102 24605 -23005
rect 21243 -23615 21473 -23614
rect 20617 -23628 20749 -23618
rect 21060 -23627 21195 -23621
rect 21040 -23628 21195 -23627
rect 20617 -23664 21195 -23628
rect 21243 -23652 21487 -23615
rect 20617 -23678 20749 -23664
rect 21040 -23667 21195 -23664
rect 21060 -23675 21195 -23667
rect 21453 -23687 21487 -23652
rect 21583 -23687 21643 -23627
rect 19188 -23760 20784 -23717
rect 17339 -23782 20784 -23760
rect 20970 -23720 21129 -23719
rect 20970 -23725 21130 -23720
rect 21278 -23725 21413 -23719
rect 20970 -23764 21413 -23725
rect 20970 -23765 21184 -23764
rect 20970 -23778 21130 -23765
rect 21278 -23773 21413 -23764
rect 21453 -23748 21643 -23687
rect 20970 -23779 21129 -23778
rect 17339 -23849 19368 -23782
rect 8767 -23903 8826 -23896
rect 8767 -23986 12743 -23903
rect 8767 -23991 8826 -23986
rect 6645 -24116 7394 -24107
rect 5561 -24169 7394 -24116
rect 4771 -24561 5018 -24560
rect 5180 -24561 5214 -24190
rect 5561 -24292 5600 -24169
rect 6762 -24203 7394 -24169
rect 5663 -24243 6671 -24207
rect 5565 -24481 5599 -24292
rect 4365 -24595 4598 -24561
rect 4771 -24595 5214 -24561
rect 5563 -24564 5600 -24481
rect 5663 -24488 5697 -24243
rect 5979 -24482 6013 -24280
rect 6077 -24479 6111 -24280
rect 6341 -24479 6375 -24280
rect 5976 -24503 6013 -24482
rect 5857 -24540 6013 -24503
rect 6075 -24518 6375 -24479
rect 5857 -24564 5894 -24540
rect 4021 -24649 4156 -24642
rect 4561 -24649 4598 -24595
rect 5563 -24601 5894 -24564
rect 6439 -24571 6473 -24280
rect 6635 -24297 6671 -24243
rect 6635 -24488 6669 -24297
rect 6733 -24571 6767 -24280
rect 6945 -24471 6979 -24280
rect 7038 -24287 7081 -24203
rect 6940 -24516 6983 -24471
rect 7043 -24488 7077 -24287
rect 7254 -24469 7288 -24280
rect 7347 -24289 7390 -24203
rect 6844 -24562 6983 -24516
rect 6206 -24605 6767 -24571
rect 4021 -24686 4598 -24649
rect 4021 -24696 4156 -24686
rect 4561 -24824 4598 -24686
rect 4632 -24651 4767 -24644
rect 4632 -24685 5451 -24651
rect 6206 -24667 6240 -24605
rect 4632 -24698 4767 -24685
rect 4820 -24729 4955 -24722
rect 4820 -24767 5381 -24729
rect 4820 -24776 4955 -24767
rect 5155 -24813 5291 -24804
rect 4561 -24861 5116 -24824
rect 5155 -24850 5310 -24813
rect 5156 -24858 5291 -24850
rect 4690 -25105 4724 -24861
rect 4886 -25105 4920 -24861
rect 5082 -25105 5116 -24861
rect -2319 -26234 2133 -26198
rect 2195 -26154 3697 -26120
rect 5347 -26136 5381 -24767
rect -2319 -26282 -2270 -26234
rect 91 -26278 227 -26269
rect 2195 -26278 2229 -26154
rect 5041 -26170 5381 -26136
rect 2274 -26209 2410 -26206
rect 5041 -26209 5075 -26170
rect 2274 -26243 5075 -26209
rect 5179 -26228 5315 -26222
rect 5417 -26228 5451 -24685
rect 5564 -24736 5703 -24682
rect 6094 -24701 6240 -24667
rect 6094 -24816 6128 -24701
rect 6313 -24706 6452 -24652
rect 5514 -24850 6128 -24816
rect 6189 -24777 6669 -24743
rect 5565 -25198 5599 -24886
rect 5663 -25094 5697 -24850
rect 5761 -25198 5795 -24886
rect 5881 -25129 5915 -24886
rect 5979 -25094 6013 -24850
rect 6077 -25129 6111 -24886
rect 6189 -25129 6223 -24777
rect 5881 -25163 6223 -25129
rect 6259 -24851 6473 -24817
rect 6259 -25198 6293 -24851
rect 6439 -25094 6473 -24851
rect 5565 -25232 6293 -25198
rect 6635 -25094 6669 -24777
rect 6722 -24780 6861 -24726
rect 6940 -24901 6983 -24562
rect 7250 -24660 7293 -24469
rect 7352 -24488 7386 -24289
rect 7543 -24350 8698 -24089
rect 12080 -24175 12365 -24117
rect 12660 -24175 12743 -23986
rect 17468 -24001 17512 -23849
rect 17472 -24160 17506 -24001
rect 17570 -24151 17604 -23952
rect 17662 -24000 17706 -23849
rect 12080 -24203 17040 -24175
rect 17378 -24203 17524 -24195
rect 12080 -24239 17524 -24203
rect 17565 -24200 17610 -24151
rect 17668 -24160 17702 -24000
rect 18414 -24001 18458 -23849
rect 18418 -24160 18452 -24001
rect 18516 -24151 18550 -23952
rect 18608 -24000 18652 -23849
rect 17565 -24201 17959 -24200
rect 17565 -24236 18008 -24201
rect 18324 -24203 18470 -24195
rect 12080 -24269 17040 -24239
rect 17378 -24255 17524 -24239
rect 17820 -24245 18008 -24236
rect 18265 -24239 18470 -24203
rect 18511 -24200 18556 -24151
rect 18614 -24160 18648 -24000
rect 18511 -24236 19181 -24200
rect 17876 -24261 18008 -24245
rect 18324 -24255 18470 -24239
rect 18766 -24245 19181 -24236
rect 12080 -24336 12365 -24269
rect 17601 -24292 17744 -24275
rect 17143 -24328 17744 -24292
rect 7150 -24706 7293 -24660
rect 6945 -25094 6979 -24901
rect 7250 -24903 7293 -24706
rect 7337 -24774 7476 -24720
rect 7254 -25094 7288 -24903
rect 2274 -26252 2410 -26243
rect 5179 -26262 5451 -26228
rect 5179 -26268 5315 -26262
rect -2406 -26328 -2270 -26282
rect 58 -26312 2229 -26278
rect 91 -26315 227 -26312
rect 7543 -26345 7804 -24350
rect -6248 -26367 -5616 -26358
rect -3748 -26367 -3116 -26358
rect -1248 -26367 -616 -26358
rect 1252 -26367 1884 -26358
rect 3752 -26367 4384 -26358
rect 6736 -26367 7804 -26345
rect -7449 -26368 -5616 -26367
rect -4949 -26368 7804 -26367
rect -7449 -26420 7804 -26368
rect -7449 -26543 -7410 -26420
rect -6248 -26454 -4910 -26420
rect -3748 -26454 -3116 -26420
rect -7347 -26494 -6339 -26458
rect -7445 -26732 -7411 -26543
rect -7447 -26815 -7410 -26732
rect -7347 -26739 -7313 -26494
rect -7031 -26733 -6997 -26531
rect -6933 -26730 -6899 -26531
rect -6669 -26730 -6635 -26531
rect -7034 -26754 -6997 -26733
rect -7153 -26791 -6997 -26754
rect -6935 -26769 -6635 -26730
rect -7153 -26815 -7116 -26791
rect -7447 -26852 -7116 -26815
rect -6571 -26822 -6537 -26531
rect -6375 -26548 -6339 -26494
rect -6375 -26739 -6341 -26548
rect -6277 -26822 -6243 -26531
rect -6065 -26722 -6031 -26531
rect -5972 -26538 -5929 -26454
rect -5737 -26455 -4910 -26454
rect -6070 -26767 -6027 -26722
rect -5967 -26739 -5933 -26538
rect -5756 -26720 -5722 -26531
rect -5663 -26540 -5620 -26455
rect -6166 -26813 -6027 -26767
rect -6804 -26856 -6243 -26822
rect -6804 -26918 -6770 -26856
rect -7446 -26987 -7307 -26933
rect -6916 -26952 -6770 -26918
rect -6916 -27067 -6882 -26952
rect -6697 -26957 -6558 -26903
rect -7556 -27101 -6882 -27067
rect -6821 -27028 -6341 -26994
rect -18267 -27132 -17602 -27104
rect -22246 -27187 -21691 -27150
rect -21651 -27174 -19833 -27139
rect -21651 -27176 -21497 -27174
rect -21651 -27184 -21516 -27176
rect -19891 -27179 -19833 -27174
rect -22117 -27431 -22083 -27187
rect -21921 -27431 -21887 -27187
rect -21725 -27431 -21691 -27187
rect -9146 -27295 -8946 -27271
rect -19527 -27431 -8946 -27295
rect -9146 -27442 -8946 -27431
rect -7445 -27449 -7411 -27137
rect -7347 -27345 -7313 -27101
rect -7249 -27449 -7215 -27137
rect -7129 -27380 -7095 -27137
rect -7031 -27345 -6997 -27101
rect -6933 -27380 -6899 -27137
rect -6821 -27380 -6787 -27028
rect -7129 -27414 -6787 -27380
rect -6751 -27102 -6537 -27068
rect -6751 -27449 -6717 -27102
rect -7445 -27483 -6717 -27449
rect -6571 -27345 -6537 -27102
rect -6375 -27345 -6341 -27028
rect -6288 -27031 -6149 -26977
rect -6070 -27152 -6027 -26813
rect -5760 -26911 -5717 -26720
rect -5658 -26739 -5624 -26540
rect -4949 -26543 -4910 -26455
rect -4847 -26494 -3839 -26458
rect -5119 -26704 -5073 -26568
rect -5860 -26957 -5717 -26911
rect -6065 -27345 -6031 -27152
rect -5760 -27154 -5717 -26957
rect -5673 -27025 -5534 -26971
rect -5756 -27345 -5722 -27154
rect -8009 -27549 -7846 -27529
rect -19704 -27685 -7846 -27549
rect -5113 -27067 -5079 -26704
rect -4945 -26732 -4911 -26543
rect -4947 -26815 -4910 -26732
rect -4847 -26739 -4813 -26494
rect -4531 -26733 -4497 -26531
rect -4433 -26730 -4399 -26531
rect -4169 -26730 -4135 -26531
rect -4534 -26754 -4497 -26733
rect -4653 -26791 -4497 -26754
rect -4435 -26769 -4135 -26730
rect -4653 -26815 -4616 -26791
rect -4947 -26852 -4616 -26815
rect -4071 -26822 -4037 -26531
rect -3875 -26548 -3839 -26494
rect -3875 -26739 -3841 -26548
rect -3777 -26822 -3743 -26531
rect -3565 -26722 -3531 -26531
rect -3472 -26538 -3429 -26454
rect -3570 -26767 -3527 -26722
rect -3467 -26739 -3433 -26538
rect -3256 -26720 -3222 -26531
rect -3163 -26540 -3120 -26454
rect -3666 -26813 -3527 -26767
rect -4304 -26856 -3743 -26822
rect -4304 -26918 -4270 -26856
rect -4946 -26987 -4807 -26933
rect -4416 -26952 -4270 -26918
rect -4416 -27067 -4382 -26952
rect -4197 -26957 -4058 -26903
rect -5113 -27101 -4382 -27067
rect -4321 -27028 -3841 -26994
rect -4945 -27449 -4911 -27137
rect -4847 -27345 -4813 -27101
rect -4749 -27449 -4715 -27137
rect -4629 -27380 -4595 -27137
rect -4531 -27345 -4497 -27101
rect -4433 -27380 -4399 -27137
rect -4321 -27380 -4287 -27028
rect -4629 -27414 -4287 -27380
rect -4251 -27102 -4037 -27068
rect -4251 -27449 -4217 -27102
rect -4945 -27483 -4217 -27449
rect -4071 -27345 -4037 -27102
rect -3875 -27345 -3841 -27028
rect -3788 -27031 -3649 -26977
rect -3570 -27152 -3527 -26813
rect -3260 -26911 -3217 -26720
rect -3158 -26739 -3124 -26540
rect -2449 -26543 -2410 -26420
rect -1248 -26454 -616 -26420
rect -2347 -26494 -1339 -26458
rect -3360 -26957 -3217 -26911
rect -3565 -27345 -3531 -27152
rect -3260 -27154 -3217 -26957
rect -3173 -27025 -3034 -26971
rect -3256 -27345 -3222 -27154
rect -2571 -26700 -2525 -26564
rect -2565 -27067 -2531 -26700
rect -2445 -26732 -2411 -26543
rect -2447 -26815 -2410 -26732
rect -2347 -26739 -2313 -26494
rect -2031 -26733 -1997 -26531
rect -1933 -26730 -1899 -26531
rect -1669 -26730 -1635 -26531
rect -2034 -26754 -1997 -26733
rect -2153 -26791 -1997 -26754
rect -1935 -26769 -1635 -26730
rect -2153 -26815 -2116 -26791
rect -2447 -26852 -2116 -26815
rect -1571 -26822 -1537 -26531
rect -1375 -26548 -1339 -26494
rect -1375 -26739 -1341 -26548
rect -1277 -26822 -1243 -26531
rect -1065 -26722 -1031 -26531
rect -972 -26538 -929 -26454
rect -1070 -26767 -1027 -26722
rect -967 -26739 -933 -26538
rect -756 -26720 -722 -26531
rect -663 -26540 -620 -26454
rect -1166 -26813 -1027 -26767
rect -1804 -26856 -1243 -26822
rect -1804 -26918 -1770 -26856
rect -2446 -26987 -2307 -26933
rect -1916 -26952 -1770 -26918
rect -1916 -27067 -1882 -26952
rect -1697 -26957 -1558 -26903
rect -2565 -27101 -1882 -27067
rect -1821 -27028 -1341 -26994
rect -2445 -27449 -2411 -27137
rect -2347 -27345 -2313 -27101
rect -2249 -27449 -2215 -27137
rect -2129 -27380 -2095 -27137
rect -2031 -27345 -1997 -27101
rect -1933 -27380 -1899 -27137
rect -1821 -27380 -1787 -27028
rect -2129 -27414 -1787 -27380
rect -1751 -27102 -1537 -27068
rect -1751 -27449 -1717 -27102
rect -2445 -27483 -1717 -27449
rect -1571 -27345 -1537 -27102
rect -1375 -27345 -1341 -27028
rect -1288 -27031 -1149 -26977
rect -1070 -27152 -1027 -26813
rect -760 -26911 -717 -26720
rect -658 -26739 -624 -26540
rect 51 -26543 90 -26420
rect 1252 -26454 1884 -26420
rect 153 -26494 1161 -26458
rect -860 -26957 -717 -26911
rect -1065 -27345 -1031 -27152
rect -760 -27154 -717 -26957
rect -673 -27025 -534 -26971
rect -756 -27345 -722 -27154
rect -91 -26700 -45 -26564
rect -85 -27067 -51 -26700
rect 55 -26732 89 -26543
rect 53 -26815 90 -26732
rect 153 -26739 187 -26494
rect 469 -26733 503 -26531
rect 567 -26730 601 -26531
rect 831 -26730 865 -26531
rect 466 -26754 503 -26733
rect 347 -26791 503 -26754
rect 565 -26769 865 -26730
rect 347 -26815 384 -26791
rect 53 -26852 384 -26815
rect 929 -26822 963 -26531
rect 1125 -26548 1161 -26494
rect 1125 -26739 1159 -26548
rect 1223 -26822 1257 -26531
rect 1435 -26722 1469 -26531
rect 1528 -26538 1571 -26454
rect 1430 -26767 1473 -26722
rect 1533 -26739 1567 -26538
rect 1744 -26720 1778 -26531
rect 1837 -26540 1880 -26454
rect 1334 -26813 1473 -26767
rect 696 -26856 1257 -26822
rect 696 -26918 730 -26856
rect 54 -26987 193 -26933
rect 584 -26952 730 -26918
rect 584 -27067 618 -26952
rect 803 -26957 942 -26903
rect -85 -27101 618 -27067
rect 679 -27028 1159 -26994
rect -85 -27102 -51 -27101
rect 55 -27449 89 -27137
rect 153 -27345 187 -27101
rect 251 -27449 285 -27137
rect 371 -27380 405 -27137
rect 469 -27345 503 -27101
rect 567 -27380 601 -27137
rect 679 -27380 713 -27028
rect 371 -27414 713 -27380
rect 749 -27102 963 -27068
rect 749 -27449 783 -27102
rect 55 -27483 783 -27449
rect 929 -27345 963 -27102
rect 1125 -27345 1159 -27028
rect 1212 -27031 1351 -26977
rect 1430 -27152 1473 -26813
rect 1740 -26911 1783 -26720
rect 1842 -26739 1876 -26540
rect 2551 -26543 2590 -26420
rect 3752 -26454 4384 -26420
rect 2653 -26494 3661 -26458
rect 2326 -26700 2372 -26564
rect 2331 -26701 2366 -26700
rect 1640 -26957 1783 -26911
rect 1435 -27345 1469 -27152
rect 1740 -27154 1783 -26957
rect 1827 -27025 1966 -26971
rect 2331 -27067 2365 -26701
rect 2555 -26732 2589 -26543
rect 2553 -26815 2590 -26732
rect 2653 -26739 2687 -26494
rect 2969 -26733 3003 -26531
rect 3067 -26730 3101 -26531
rect 3331 -26730 3365 -26531
rect 2966 -26754 3003 -26733
rect 2847 -26791 3003 -26754
rect 3065 -26769 3365 -26730
rect 2847 -26815 2884 -26791
rect 2553 -26852 2884 -26815
rect 3429 -26822 3463 -26531
rect 3625 -26548 3661 -26494
rect 3625 -26739 3659 -26548
rect 3723 -26822 3757 -26531
rect 3935 -26722 3969 -26531
rect 4028 -26538 4071 -26454
rect 3930 -26767 3973 -26722
rect 4033 -26739 4067 -26538
rect 4244 -26720 4278 -26531
rect 4337 -26540 4380 -26454
rect 3834 -26813 3973 -26767
rect 3196 -26856 3757 -26822
rect 3196 -26918 3230 -26856
rect 2554 -26987 2693 -26933
rect 3084 -26952 3230 -26918
rect 3084 -27067 3118 -26952
rect 3303 -26957 3442 -26903
rect 2331 -27101 3118 -27067
rect 3179 -27028 3659 -26994
rect 1744 -27345 1778 -27154
rect 2555 -27449 2589 -27137
rect 2653 -27345 2687 -27101
rect 2751 -27449 2785 -27137
rect 2871 -27380 2905 -27137
rect 2969 -27345 3003 -27101
rect 3067 -27380 3101 -27137
rect 3179 -27380 3213 -27028
rect 2871 -27414 3213 -27380
rect 3249 -27102 3463 -27068
rect 3249 -27449 3283 -27102
rect 2555 -27483 3283 -27449
rect 3429 -27345 3463 -27102
rect 3625 -27345 3659 -27028
rect 3712 -27031 3851 -26977
rect 3930 -27152 3973 -26813
rect 4240 -26911 4283 -26720
rect 4342 -26739 4376 -26540
rect 5551 -26543 5590 -26420
rect 5653 -26494 6661 -26458
rect 6736 -26472 7804 -26420
rect 5231 -26700 5277 -26564
rect 4140 -26957 4283 -26911
rect 3935 -27345 3969 -27152
rect 4240 -27154 4283 -26957
rect 4327 -27025 4466 -26971
rect 5237 -27067 5271 -26700
rect 5555 -26732 5589 -26543
rect 5553 -26815 5590 -26732
rect 5653 -26739 5687 -26494
rect 5969 -26733 6003 -26531
rect 6067 -26730 6101 -26531
rect 6331 -26730 6365 -26531
rect 5966 -26754 6003 -26733
rect 5847 -26791 6003 -26754
rect 6065 -26769 6365 -26730
rect 5847 -26815 5884 -26791
rect 5553 -26852 5884 -26815
rect 6429 -26822 6463 -26531
rect 6625 -26548 6661 -26494
rect 6625 -26739 6659 -26548
rect 6723 -26822 6757 -26531
rect 6935 -26722 6969 -26531
rect 7028 -26538 7071 -26472
rect 6930 -26767 6973 -26722
rect 7033 -26739 7067 -26538
rect 7244 -26720 7278 -26531
rect 7337 -26540 7380 -26472
rect 6834 -26813 6973 -26767
rect 6196 -26856 6757 -26822
rect 6196 -26918 6230 -26856
rect 5554 -26987 5693 -26933
rect 6084 -26952 6230 -26918
rect 6084 -27067 6118 -26952
rect 6303 -26957 6442 -26903
rect 5237 -27101 6118 -27067
rect 6179 -27028 6659 -26994
rect 4244 -27345 4278 -27154
rect 5555 -27449 5589 -27137
rect 5653 -27345 5687 -27101
rect 5751 -27449 5785 -27137
rect 5871 -27380 5905 -27137
rect 5969 -27345 6003 -27101
rect 6067 -27380 6101 -27137
rect 6179 -27380 6213 -27028
rect 5871 -27414 6213 -27380
rect 6249 -27102 6463 -27068
rect 6249 -27449 6283 -27102
rect 5555 -27483 6283 -27449
rect 6429 -27345 6463 -27102
rect 6625 -27345 6659 -27028
rect 6712 -27031 6851 -26977
rect 6930 -27152 6973 -26813
rect 7240 -26911 7283 -26720
rect 7342 -26739 7376 -26540
rect 7140 -26957 7283 -26911
rect 6935 -27345 6969 -27152
rect 7240 -27154 7283 -26957
rect 7327 -27025 7466 -26971
rect 7244 -27345 7278 -27154
rect -19704 -27686 -19566 -27685
rect -22910 -27731 -22752 -27698
rect -8009 -27704 -7846 -27685
rect -19842 -27731 -19705 -27726
rect -22910 -27783 -19705 -27731
rect -22910 -27814 -22752 -27783
rect -19842 -27784 -19705 -27783
rect 8437 -25144 8698 -24350
rect 17143 -24381 17179 -24328
rect 17601 -24335 17744 -24328
rect 13062 -24543 17179 -24381
rect 17471 -24410 17819 -24374
rect 8920 -24706 8989 -24688
rect 14133 -24706 14244 -24543
rect 8920 -24817 14244 -24706
rect 8920 -24827 8989 -24817
rect 17471 -24449 17507 -24410
rect 17472 -24852 17506 -24449
rect 17683 -24824 17717 -24444
rect 17774 -24454 17819 -24410
rect 17676 -24888 17722 -24824
rect 17781 -24852 17815 -24454
rect 17876 -24490 17926 -24261
rect 18547 -24292 18690 -24275
rect 18264 -24328 18690 -24292
rect 18547 -24335 18690 -24328
rect 18417 -24410 18765 -24374
rect 17879 -24824 17913 -24490
rect 17874 -24888 17920 -24824
rect 18417 -24449 18453 -24410
rect 17676 -24926 17920 -24888
rect 18418 -24852 18452 -24449
rect 18629 -24824 18663 -24444
rect 18720 -24454 18765 -24410
rect 18622 -24888 18668 -24824
rect 18727 -24852 18761 -24454
rect 18822 -24490 18872 -24245
rect 18825 -24824 18859 -24490
rect 18912 -24510 18972 -24344
rect 19147 -24432 19181 -24245
rect 19236 -24342 19270 -23971
rect 19334 -24279 19368 -23849
rect 19546 -23872 19987 -23838
rect 19546 -23875 19777 -23872
rect 19432 -24341 19466 -23971
rect 19546 -23979 19581 -23875
rect 19546 -24278 19580 -23979
rect 19644 -24278 19678 -23970
rect 19742 -23981 19777 -23875
rect 19742 -24278 19776 -23981
rect 19644 -24341 19679 -24278
rect 19432 -24342 19679 -24341
rect 19855 -24342 19889 -23970
rect 19953 -24278 19987 -23872
rect 20051 -24342 20085 -23970
rect 20366 -24178 20400 -23782
rect 20468 -23798 20784 -23782
rect 20468 -23833 20783 -23798
rect 19236 -24376 19679 -24342
rect 19852 -24376 20085 -24342
rect 20464 -24363 20498 -23970
rect 20702 -24139 20783 -23833
rect 21145 -24136 21179 -23824
rect 21243 -24052 21277 -23824
rect 21355 -24052 21389 -23824
rect 21453 -24032 21487 -23748
rect 21583 -23761 21643 -23748
rect 21243 -24087 21389 -24052
rect 21112 -24139 21591 -24136
rect 21681 -24139 21751 -23102
rect 20702 -24297 21751 -24139
rect 21086 -24340 21751 -24297
rect 21808 -23981 21878 -23247
rect 21975 -23923 22009 -23102
rect 22073 -23979 22107 -23215
rect 22375 -23923 22409 -23102
rect 22305 -23979 22439 -23966
rect 21808 -24035 22037 -23981
rect 22073 -24013 22439 -23979
rect 19683 -24432 19818 -24425
rect 19142 -24466 19818 -24432
rect 19683 -24479 19818 -24466
rect 19852 -24430 19889 -24376
rect 20464 -24399 20741 -24363
rect 20294 -24430 20429 -24423
rect 19852 -24467 20429 -24430
rect 19495 -24510 19630 -24503
rect 18912 -24548 19630 -24510
rect 19495 -24557 19630 -24548
rect 19159 -24594 19294 -24585
rect 19027 -24629 19294 -24594
rect 19852 -24605 19889 -24467
rect 20294 -24477 20429 -24467
rect 19027 -24726 19087 -24629
rect 19140 -24631 19294 -24629
rect 19159 -24639 19294 -24631
rect 19334 -24642 19889 -24605
rect 18820 -24888 18866 -24824
rect 18622 -24926 18866 -24888
rect 19334 -24886 19368 -24642
rect 19530 -24886 19564 -24642
rect 19726 -24886 19760 -24642
rect 20464 -24886 20498 -24399
rect 20610 -24423 20741 -24399
rect 21095 -24499 21129 -24340
rect 21193 -24483 21227 -24391
rect 20983 -24607 21151 -24533
rect 21187 -24576 21233 -24483
rect 21291 -24499 21325 -24340
rect 21389 -24483 21423 -24391
rect 21383 -24576 21429 -24483
rect 21487 -24499 21521 -24340
rect 21585 -24483 21619 -24391
rect 21579 -24544 21625 -24483
rect 21808 -24544 21878 -24035
rect 21579 -24576 21878 -24544
rect 21187 -24614 21878 -24576
rect 21187 -24622 21625 -24614
rect 21187 -24875 21233 -24622
rect 21193 -24879 21227 -24875
rect 21383 -24687 21429 -24622
rect 21389 -24879 21423 -24687
rect 21579 -24687 21625 -24622
rect 21585 -24879 21619 -24687
rect 22073 -24808 22107 -24013
rect 22305 -24020 22439 -24013
rect 22473 -23969 22507 -23215
rect 22581 -23969 22699 -23957
rect 22473 -24003 22699 -23969
rect 22473 -24808 22507 -24003
rect 22581 -24015 22699 -24003
rect 22852 -23979 22922 -23798
rect 22975 -23923 23009 -23102
rect 22852 -24033 23026 -23979
rect 23073 -23989 23107 -23215
rect 23375 -23923 23409 -23102
rect 23305 -23989 23439 -23981
rect 23073 -24028 23439 -23989
rect 23073 -24808 23107 -24028
rect 23305 -24035 23439 -24028
rect 23473 -23996 23507 -23215
rect 23658 -23996 23776 -23984
rect 23473 -24030 23776 -23996
rect 23473 -24808 23507 -24030
rect 23658 -24042 23776 -24030
rect 23843 -23986 23913 -23799
rect 23975 -23923 24009 -23102
rect 23843 -24040 24026 -23986
rect 24073 -23990 24107 -23215
rect 24375 -23923 24409 -23102
rect 24473 -23980 24507 -23215
rect 24554 -23980 24672 -23972
rect 24298 -23990 24432 -23983
rect 24073 -24029 24432 -23990
rect 24073 -24808 24107 -24029
rect 24298 -24037 24432 -24029
rect 24473 -24014 24675 -23980
rect 24473 -24808 24507 -24014
rect 24554 -24030 24672 -24014
rect 26685 -23241 26761 -22169
rect 26900 -22170 27386 -22169
rect 26900 -22171 26971 -22170
rect 27312 -22176 27386 -22170
rect 26932 -22521 26966 -22213
rect 27030 -22521 27064 -22213
rect 27128 -22521 27162 -22213
rect 27226 -22521 27260 -22213
rect 27324 -22521 27358 -22213
rect 27029 -22573 27064 -22521
rect 27743 -22555 27804 -22148
rect 28233 -22312 28303 -21917
rect 28477 -22171 28511 -21587
rect 28684 -21553 28924 -21519
rect 28684 -21595 28726 -21553
rect 28473 -22230 28515 -22171
rect 28688 -22177 28722 -21595
rect 28786 -22175 28820 -21587
rect 28882 -21597 28924 -21553
rect 28685 -22230 28727 -22177
rect 28473 -22266 28727 -22230
rect 28782 -22229 28824 -22175
rect 28884 -22195 28918 -21597
rect 29096 -22181 29130 -21587
rect 28782 -22268 28923 -22229
rect 28880 -22280 28923 -22268
rect 28638 -22312 28793 -22302
rect 28233 -22348 28793 -22312
rect 28233 -22350 28303 -22348
rect 28638 -22357 28793 -22348
rect 28880 -22335 29061 -22280
rect 28880 -22405 28923 -22335
rect 28368 -22419 28523 -22410
rect 28331 -22453 28523 -22419
rect 28368 -22465 28523 -22453
rect 28569 -22445 28923 -22405
rect 29095 -22425 29138 -22181
rect 29332 -22250 29402 -20913
rect 35496 -20966 35530 -20758
rect 35692 -20966 35726 -20758
rect 35888 -20966 35922 -20758
rect 30469 -21945 30503 -21445
rect 30648 -21409 30969 -21375
rect 30468 -21991 30503 -21945
rect 30648 -21991 30688 -21409
rect 30737 -21449 30772 -21409
rect 30738 -21953 30772 -21449
rect 30836 -21946 30870 -21445
rect 30934 -21448 30969 -21409
rect 30468 -22031 30688 -21991
rect 30833 -22066 30871 -21946
rect 30934 -21953 30968 -21448
rect 31064 -22029 31098 -21445
rect 31390 -21959 31424 -21445
rect 31618 -21735 31652 -21445
rect 36469 -21095 36503 -20751
rect 36665 -21095 36699 -20751
rect 36838 -20900 36899 -20751
rect 37078 -20865 37112 -20709
rect 37176 -20865 37210 -20757
rect 37274 -20865 37308 -20709
rect 44067 -20750 44314 -20709
rect 45149 -20737 45284 -20729
rect 45129 -20739 45284 -20737
rect 37372 -20865 37406 -20757
rect 44067 -20767 44197 -20750
rect 44241 -20763 44314 -20750
rect 44922 -20775 45284 -20739
rect 45801 -20748 46586 -20662
rect 53265 -20675 53395 -20583
rect 53557 -20641 53591 -20385
rect 53655 -20641 53689 -20433
rect 53753 -20641 53787 -20385
rect 53851 -20607 53885 -20433
rect 54432 -20563 54466 -20255
rect 54530 -20563 54564 -20255
rect 54628 -20563 54662 -20255
rect 54726 -20563 54760 -20255
rect 54824 -20563 54858 -20255
rect 54400 -20606 54471 -20605
rect 54812 -20606 54886 -20600
rect 54400 -20607 54886 -20606
rect 53851 -20641 54886 -20607
rect 55243 -20628 55304 -20221
rect 59891 -20251 61742 -20100
rect 63023 -20094 63688 -20066
rect 63023 -20152 64058 -20094
rect 63023 -20233 63109 -20152
rect 63283 -20189 63318 -20152
rect 63608 -20155 64058 -20152
rect 59891 -20319 60267 -20251
rect 61492 -20302 61742 -20251
rect 62171 -20319 63109 -20233
rect 62019 -20609 62149 -20517
rect 62311 -20575 62345 -20319
rect 62409 -20575 62443 -20367
rect 62507 -20575 62541 -20319
rect 62605 -20541 62639 -20367
rect 63186 -20497 63220 -20189
rect 63284 -20497 63318 -20189
rect 63382 -20497 63416 -20189
rect 63480 -20497 63514 -20189
rect 63578 -20497 63612 -20189
rect 63154 -20540 63225 -20539
rect 63566 -20540 63640 -20534
rect 63154 -20541 63640 -20540
rect 62605 -20575 63640 -20541
rect 63997 -20562 64058 -20155
rect 68667 -20106 69005 -20010
rect 72443 -20049 72783 -19655
rect 77897 -20045 78167 -19924
rect 79910 -20045 80205 -20003
rect 81779 -20011 81990 -19655
rect 70655 -20106 70923 -20065
rect 68667 -20237 70923 -20106
rect 72176 -20077 72841 -20049
rect 72176 -20135 73211 -20077
rect 72176 -20216 72262 -20135
rect 72436 -20172 72471 -20135
rect 72761 -20138 73211 -20135
rect 68667 -20301 69005 -20237
rect 70655 -20305 70923 -20237
rect 71324 -20302 72262 -20216
rect 62606 -20579 63640 -20575
rect 62606 -20581 63155 -20579
rect 62193 -20609 62266 -20603
rect 63566 -20605 63640 -20579
rect 53852 -20645 54886 -20641
rect 53852 -20647 54401 -20645
rect 53439 -20675 53512 -20669
rect 54812 -20671 54886 -20645
rect 53265 -20716 53512 -20675
rect 54347 -20703 54482 -20695
rect 54327 -20705 54482 -20703
rect 53265 -20733 53395 -20716
rect 53439 -20729 53512 -20716
rect 54120 -20741 54482 -20705
rect 54999 -20714 55784 -20628
rect 62019 -20650 62266 -20609
rect 63101 -20637 63236 -20629
rect 63081 -20639 63236 -20637
rect 62019 -20667 62149 -20650
rect 62193 -20663 62266 -20650
rect 62874 -20675 63236 -20639
rect 63753 -20648 64538 -20562
rect 71172 -20592 71302 -20500
rect 71464 -20558 71498 -20302
rect 71562 -20558 71596 -20350
rect 71660 -20558 71694 -20302
rect 71758 -20524 71792 -20350
rect 72339 -20480 72373 -20172
rect 72437 -20480 72471 -20172
rect 72535 -20480 72569 -20172
rect 72633 -20480 72667 -20172
rect 72731 -20480 72765 -20172
rect 72307 -20523 72378 -20522
rect 72719 -20523 72793 -20517
rect 72307 -20524 72793 -20523
rect 71758 -20558 72793 -20524
rect 73150 -20545 73211 -20138
rect 77897 -20184 80205 -20045
rect 81540 -20039 82205 -20011
rect 81540 -20097 82575 -20039
rect 81540 -20178 81626 -20097
rect 81800 -20134 81835 -20097
rect 82125 -20100 82575 -20097
rect 77897 -20209 78167 -20184
rect 79910 -20276 80205 -20184
rect 80688 -20264 81626 -20178
rect 71759 -20562 72793 -20558
rect 71759 -20564 72308 -20562
rect 71346 -20592 71419 -20586
rect 72719 -20588 72793 -20562
rect 71172 -20633 71419 -20592
rect 72254 -20620 72389 -20612
rect 72234 -20622 72389 -20620
rect 63081 -20677 63236 -20675
rect 63101 -20683 63236 -20677
rect 63284 -20660 63703 -20652
rect 63284 -20690 63714 -20660
rect 54327 -20743 54482 -20741
rect 45129 -20777 45284 -20775
rect 45149 -20783 45284 -20777
rect 45332 -20760 45751 -20752
rect 45332 -20790 45762 -20760
rect 36960 -20900 37033 -20894
rect 36838 -20913 37033 -20900
rect 36860 -20941 37033 -20913
rect 36960 -20954 37033 -20941
rect 37470 -20924 37842 -20854
rect 37078 -21096 37112 -20988
rect 37274 -21096 37308 -20988
rect 37470 -21096 37504 -20924
rect 31617 -21828 31654 -21735
rect 31617 -21865 31754 -21828
rect 31390 -21993 31549 -21959
rect 31213 -22029 31351 -22018
rect 30469 -22104 30871 -22066
rect 30938 -22063 31351 -22029
rect 30232 -22115 30370 -22105
rect 29842 -22149 30370 -22115
rect 29321 -22322 29426 -22250
rect 29842 -22425 29885 -22149
rect 30232 -22159 30370 -22149
rect 30288 -22250 30426 -22241
rect 30078 -22284 30426 -22250
rect 30078 -22411 30150 -22284
rect 30288 -22295 30426 -22284
rect 30078 -22420 30162 -22411
rect 27354 -22573 27804 -22555
rect 26912 -22616 27804 -22573
rect 26912 -22634 27361 -22616
rect 27743 -22911 27804 -22616
rect 28477 -22793 28511 -22499
rect 28569 -22515 28614 -22445
rect 28961 -22465 29885 -22425
rect 29009 -22468 29885 -22465
rect 28470 -22911 28517 -22793
rect 28575 -22807 28609 -22515
rect 28673 -22792 28707 -22499
rect 28915 -22782 28949 -22499
rect 29009 -22508 29053 -22468
rect 30083 -22490 30162 -22420
rect 28666 -22911 28713 -22792
rect 28908 -22911 28955 -22782
rect 29013 -22807 29047 -22508
rect 30371 -22732 30405 -22441
rect 30369 -22843 30406 -22732
rect 30469 -22749 30503 -22104
rect 30698 -22174 30736 -22104
rect 30938 -22142 30972 -22063
rect 31213 -22072 31351 -22063
rect 30688 -22312 30742 -22174
rect 30841 -22176 30972 -22142
rect 31038 -22159 31176 -22105
rect 31423 -22174 31477 -22036
rect 31515 -22037 31549 -21993
rect 31515 -22091 31681 -22037
rect 30841 -22749 30875 -22176
rect 31515 -22206 31549 -22091
rect 31601 -22206 31655 -22189
rect 30939 -22245 31098 -22210
rect 31515 -22211 31655 -22206
rect 31487 -22240 31655 -22211
rect 30939 -22749 30973 -22245
rect 31064 -22749 31098 -22245
rect 31162 -22732 31196 -22241
rect 31292 -22731 31326 -22241
rect 29832 -22847 30443 -22843
rect 31161 -22847 31198 -22732
rect 31289 -22847 31326 -22731
rect 31390 -22749 31424 -22241
rect 31487 -22245 31549 -22240
rect 31488 -22749 31522 -22245
rect 31601 -22248 31655 -22240
rect 31716 -22358 31754 -21865
rect 31716 -22396 32008 -22358
rect 31618 -22730 31652 -22441
rect 31716 -22446 31754 -22396
rect 31616 -22847 31653 -22730
rect 31716 -22749 31750 -22446
rect 29832 -22911 31766 -22847
rect 27743 -22956 31766 -22911
rect 27743 -23024 29945 -22956
rect 30293 -23008 31766 -22956
rect 8437 -25405 9407 -25144
rect 8429 -25518 8620 -25512
rect 8429 -25601 8992 -25518
rect 8429 -25619 8620 -25601
rect 8909 -27466 8992 -25601
rect 9146 -27185 9407 -25405
rect 25889 -23297 26761 -23241
rect 31970 -23291 32008 -22396
rect 25889 -23373 29995 -23297
rect 25889 -23387 26761 -23373
rect 10670 -25660 10704 -25656
rect 10664 -25913 10710 -25660
rect 10866 -25848 10900 -25656
rect 10860 -25913 10906 -25848
rect 11062 -25848 11096 -25656
rect 11331 -25842 11388 -25678
rect 11056 -25913 11102 -25848
rect 11552 -25660 11586 -25656
rect 10664 -25921 11102 -25913
rect 11546 -25913 11592 -25660
rect 11748 -25848 11782 -25656
rect 11742 -25913 11788 -25848
rect 12162 -25637 12790 -25603
rect 11944 -25848 11978 -25656
rect 12162 -25682 12198 -25637
rect 11938 -25913 11984 -25848
rect 11546 -25921 11984 -25913
rect 12039 -25897 12113 -25729
rect 12163 -25756 12197 -25682
rect 12039 -25921 12112 -25897
rect 10460 -26002 10628 -25928
rect 10664 -25943 11132 -25921
rect 11342 -25939 11510 -25928
rect 11190 -25943 11250 -25939
rect 11307 -25943 11510 -25939
rect 10664 -25959 11510 -25943
rect 9859 -26396 10154 -26298
rect 10480 -26396 10519 -26002
rect 10572 -26195 10606 -26036
rect 10664 -26052 10710 -25959
rect 10670 -26144 10704 -26052
rect 10768 -26195 10802 -26036
rect 10860 -26052 10906 -25959
rect 11056 -25985 11510 -25959
rect 11056 -25991 11132 -25985
rect 10866 -26144 10900 -26052
rect 10964 -26195 10998 -26036
rect 11056 -26052 11102 -25991
rect 11062 -26144 11096 -26052
rect 11190 -26071 11250 -25985
rect 11307 -25997 11510 -25985
rect 11342 -26002 11510 -25997
rect 11546 -25959 12112 -25921
rect 11454 -26195 11488 -26036
rect 11546 -26052 11592 -25959
rect 11552 -26144 11586 -26052
rect 11650 -26195 11684 -26036
rect 11742 -26052 11788 -25959
rect 11938 -25991 12112 -25959
rect 12157 -25903 12204 -25756
rect 12261 -25763 12295 -25671
rect 12358 -25692 12400 -25637
rect 12260 -25815 12296 -25763
rect 12359 -25779 12393 -25692
rect 12457 -25761 12491 -25671
rect 12552 -25693 12594 -25637
rect 12457 -25779 12494 -25761
rect 12555 -25779 12589 -25693
rect 12653 -25761 12687 -25671
rect 12748 -25688 12790 -25637
rect 12458 -25815 12494 -25779
rect 12652 -25815 12688 -25761
rect 12751 -25779 12785 -25688
rect 12849 -25771 12883 -25671
rect 12846 -25815 12888 -25771
rect 12260 -25849 12888 -25815
rect 12157 -25977 12329 -25903
rect 12713 -25937 12888 -25849
rect 13295 -25660 13329 -25656
rect 13289 -25913 13335 -25660
rect 13491 -25848 13525 -25656
rect 13485 -25913 13531 -25848
rect 13687 -25848 13721 -25656
rect 14031 -25756 14088 -25678
rect 13827 -25801 14088 -25756
rect 13681 -25913 13727 -25848
rect 13289 -25921 13727 -25913
rect 13085 -25937 13253 -25928
rect 11748 -26144 11782 -26052
rect 11846 -26195 11880 -26036
rect 11938 -26052 11984 -25991
rect 11944 -26144 11978 -26052
rect 12157 -26112 12204 -25977
rect 12713 -25994 13253 -25937
rect 12713 -26016 12888 -25994
rect 13085 -26002 13253 -25994
rect 13289 -25935 13757 -25921
rect 13827 -25935 13872 -25801
rect 14031 -25842 14088 -25801
rect 14252 -25660 14286 -25656
rect 14246 -25913 14292 -25660
rect 14448 -25848 14482 -25656
rect 14442 -25913 14488 -25848
rect 14862 -25637 15490 -25603
rect 14644 -25848 14678 -25656
rect 14862 -25682 14898 -25637
rect 14638 -25913 14684 -25848
rect 14246 -25921 14684 -25913
rect 14739 -25897 14813 -25729
rect 14863 -25756 14897 -25682
rect 14739 -25921 14812 -25897
rect 13289 -25959 13872 -25935
rect 12257 -26050 12888 -26016
rect 12257 -26091 12298 -26050
rect 12163 -26182 12197 -26112
rect 10563 -26263 11979 -26195
rect 12158 -26240 12202 -26182
rect 12261 -26194 12295 -26091
rect 12359 -26171 12393 -26086
rect 12455 -26099 12496 -26050
rect 12354 -26240 12398 -26171
rect 12457 -26194 12491 -26099
rect 12555 -26171 12589 -26086
rect 12649 -26099 12690 -26050
rect 12846 -26057 12888 -26050
rect 12550 -26240 12594 -26171
rect 12653 -26194 12687 -26099
rect 12751 -26182 12785 -26086
rect 12846 -26090 12887 -26057
rect 12840 -26100 12887 -26090
rect 12747 -26240 12791 -26182
rect 12840 -26222 12886 -26100
rect 13197 -26195 13231 -26036
rect 13289 -26052 13335 -25959
rect 13295 -26144 13329 -26052
rect 13393 -26195 13427 -26036
rect 13485 -26052 13531 -25959
rect 13681 -25980 13872 -25959
rect 13922 -25939 13982 -25938
rect 14042 -25939 14210 -25928
rect 13681 -25991 13757 -25980
rect 13491 -26144 13525 -26052
rect 13589 -26195 13623 -26036
rect 13681 -26052 13727 -25991
rect 13687 -26144 13721 -26052
rect 13807 -26095 13867 -25980
rect 13922 -25997 14210 -25939
rect 13922 -26070 13982 -25997
rect 14042 -26002 14210 -25997
rect 14246 -25959 14812 -25921
rect 14154 -26195 14188 -26036
rect 14246 -26052 14292 -25959
rect 14252 -26144 14286 -26052
rect 14350 -26195 14384 -26036
rect 14442 -26052 14488 -25959
rect 14638 -25991 14812 -25959
rect 14857 -25903 14904 -25756
rect 14961 -25763 14995 -25671
rect 15058 -25692 15100 -25637
rect 14960 -25815 14996 -25763
rect 15059 -25779 15093 -25692
rect 15157 -25761 15191 -25671
rect 15252 -25693 15294 -25637
rect 15157 -25779 15194 -25761
rect 15255 -25779 15289 -25693
rect 15353 -25761 15387 -25671
rect 15448 -25688 15490 -25637
rect 15158 -25815 15194 -25779
rect 15352 -25815 15388 -25761
rect 15451 -25779 15485 -25688
rect 15549 -25771 15583 -25671
rect 15546 -25815 15588 -25771
rect 14960 -25849 15588 -25815
rect 14857 -25977 15029 -25903
rect 15413 -25934 15588 -25849
rect 15995 -25660 16029 -25656
rect 15989 -25913 16035 -25660
rect 16191 -25848 16225 -25656
rect 16185 -25913 16231 -25848
rect 16387 -25848 16421 -25656
rect 16381 -25913 16427 -25848
rect 15989 -25921 16427 -25913
rect 15785 -25934 15953 -25928
rect 14448 -26144 14482 -26052
rect 14546 -26195 14580 -26036
rect 14638 -26052 14684 -25991
rect 14644 -26144 14678 -26052
rect 14857 -26112 14904 -25977
rect 15413 -25987 15953 -25934
rect 15413 -26016 15588 -25987
rect 15785 -26002 15953 -25987
rect 15989 -25930 16457 -25921
rect 15989 -25932 16539 -25930
rect 15989 -25959 16540 -25932
rect 14957 -26050 15588 -26016
rect 14957 -26091 14998 -26050
rect 14863 -26182 14897 -26112
rect 12158 -26274 12791 -26240
rect 13188 -26263 14679 -26195
rect 14858 -26240 14902 -26182
rect 14961 -26194 14995 -26091
rect 15059 -26171 15093 -26086
rect 15155 -26099 15196 -26050
rect 15054 -26240 15098 -26171
rect 15157 -26194 15191 -26099
rect 15255 -26171 15289 -26086
rect 15349 -26099 15390 -26050
rect 15546 -26057 15588 -26050
rect 15250 -26240 15294 -26171
rect 15353 -26194 15387 -26099
rect 15451 -26182 15485 -26086
rect 15546 -26100 15587 -26057
rect 15447 -26240 15491 -26182
rect 15549 -26194 15583 -26100
rect 15897 -26195 15931 -26036
rect 15989 -26052 16035 -25959
rect 15995 -26144 16029 -26052
rect 16093 -26195 16127 -26036
rect 16185 -26052 16231 -25959
rect 16381 -25969 16540 -25959
rect 16381 -25991 16457 -25969
rect 16191 -26144 16225 -26052
rect 16289 -26195 16323 -26036
rect 16381 -26052 16427 -25991
rect 16387 -26144 16421 -26052
rect 14858 -26274 15491 -26240
rect 15888 -26263 16422 -26195
rect 11149 -26310 11281 -26299
rect 15672 -26310 15804 -26297
rect 11149 -26349 16210 -26310
rect 16492 -26327 16540 -25969
rect 11149 -26359 11281 -26349
rect 15672 -26357 15804 -26349
rect 12953 -26396 13085 -26385
rect 13894 -26396 14031 -26386
rect 9859 -26435 16210 -26396
rect 9859 -26501 10154 -26435
rect 12953 -26445 13085 -26435
rect 13894 -26446 14031 -26435
rect 16481 -26464 16541 -26327
rect 10826 -26488 10958 -26469
rect 13459 -26488 13596 -26469
rect 16056 -26488 16193 -26475
rect 10825 -26527 16210 -26488
rect 10826 -26529 11191 -26527
rect 10930 -27185 11191 -26529
rect 11547 -26598 12180 -26564
rect 12584 -26575 12695 -26527
rect 13459 -26529 13596 -26527
rect 12870 -26575 13390 -26573
rect 13462 -26575 13573 -26529
rect 11455 -26738 11489 -26644
rect 11547 -26656 11591 -26598
rect 11451 -26781 11492 -26738
rect 11553 -26752 11587 -26656
rect 11651 -26739 11685 -26644
rect 11744 -26667 11788 -26598
rect 11450 -26788 11492 -26781
rect 11648 -26788 11689 -26739
rect 11749 -26752 11783 -26667
rect 11847 -26739 11881 -26644
rect 11940 -26667 11984 -26598
rect 11842 -26788 11883 -26739
rect 11945 -26752 11979 -26667
rect 12043 -26747 12077 -26644
rect 12136 -26656 12180 -26598
rect 12359 -26641 13730 -26575
rect 12359 -26643 12893 -26641
rect 13196 -26643 13730 -26641
rect 14247 -26598 14880 -26564
rect 15260 -26575 15371 -26527
rect 16056 -26535 16193 -26527
rect 16071 -26575 16182 -26535
rect 12141 -26726 12175 -26656
rect 12040 -26788 12081 -26747
rect 11450 -26820 12081 -26788
rect 11375 -26822 12081 -26820
rect 11375 -26880 11625 -26822
rect 12134 -26861 12181 -26726
rect 12360 -26786 12394 -26694
rect 12354 -26847 12400 -26786
rect 12458 -26802 12492 -26643
rect 12556 -26786 12590 -26694
rect 11450 -26989 11625 -26880
rect 12009 -26935 12181 -26861
rect 11450 -27023 12078 -26989
rect 11450 -27067 11492 -27023
rect 11455 -27167 11489 -27067
rect 11553 -27150 11587 -27059
rect 11650 -27077 11686 -27023
rect 11844 -27059 11880 -27023
rect 9146 -27446 11191 -27185
rect 11548 -27201 11590 -27150
rect 11651 -27167 11685 -27077
rect 11749 -27145 11783 -27059
rect 11844 -27077 11881 -27059
rect 11744 -27201 11786 -27145
rect 11847 -27167 11881 -27077
rect 11945 -27146 11979 -27059
rect 12042 -27075 12078 -27023
rect 11938 -27201 11980 -27146
rect 12043 -27167 12077 -27075
rect 12134 -27082 12181 -26935
rect 12226 -26879 12400 -26847
rect 12550 -26879 12596 -26786
rect 12654 -26802 12688 -26643
rect 12752 -26786 12786 -26694
rect 12746 -26879 12792 -26786
rect 12850 -26802 12884 -26643
rect 12996 -26836 13056 -26677
rect 13197 -26786 13231 -26694
rect 12226 -26917 12792 -26879
rect 12828 -26899 13056 -26836
rect 13191 -26847 13237 -26786
rect 13295 -26802 13329 -26643
rect 13393 -26786 13427 -26694
rect 13093 -26879 13237 -26847
rect 13387 -26879 13433 -26786
rect 13491 -26802 13525 -26643
rect 13589 -26786 13623 -26694
rect 13583 -26879 13629 -26786
rect 13687 -26802 13721 -26643
rect 14155 -26738 14189 -26644
rect 14247 -26656 14291 -26598
rect 14151 -26781 14192 -26738
rect 14253 -26752 14287 -26656
rect 14351 -26739 14385 -26644
rect 14444 -26667 14488 -26598
rect 14150 -26788 14192 -26781
rect 14348 -26788 14389 -26739
rect 14449 -26752 14483 -26667
rect 14547 -26739 14581 -26644
rect 14640 -26667 14684 -26598
rect 14542 -26788 14583 -26739
rect 14645 -26752 14679 -26667
rect 14743 -26747 14777 -26644
rect 14836 -26656 14880 -26598
rect 15059 -26643 16430 -26575
rect 14841 -26726 14875 -26656
rect 14740 -26788 14781 -26747
rect 14150 -26822 14781 -26788
rect 12828 -26910 12996 -26899
rect 12226 -26941 12299 -26917
rect 12141 -27156 12175 -27082
rect 12225 -27109 12299 -26941
rect 12354 -26925 12792 -26917
rect 12354 -26990 12400 -26925
rect 12140 -27201 12176 -27156
rect 12360 -27182 12394 -26990
rect 11548 -27235 12176 -27201
rect 12550 -26990 12596 -26925
rect 12556 -27182 12590 -26990
rect 12746 -27178 12792 -26925
rect 13093 -26917 13629 -26879
rect 13665 -26843 13833 -26836
rect 13665 -26903 13855 -26843
rect 14059 -26882 14325 -26822
rect 14834 -26861 14881 -26726
rect 15060 -26786 15094 -26694
rect 15054 -26847 15100 -26786
rect 15158 -26802 15192 -26643
rect 15256 -26786 15290 -26694
rect 13665 -26910 13833 -26903
rect 12752 -27182 12786 -27178
rect 12950 -27046 13007 -26996
rect 13093 -27046 13155 -26917
rect 13191 -26925 13629 -26917
rect 13191 -26990 13237 -26925
rect 12950 -27108 13155 -27046
rect 12950 -27160 13007 -27108
rect 13197 -27182 13231 -26990
rect 13387 -26990 13433 -26925
rect 13393 -27182 13427 -26990
rect 13583 -27178 13629 -26925
rect 13589 -27182 13623 -27178
rect 14150 -26989 14325 -26882
rect 14709 -26935 14881 -26861
rect 14150 -27023 14778 -26989
rect 14150 -27067 14192 -27023
rect 14155 -27167 14189 -27067
rect 14253 -27150 14287 -27059
rect 14350 -27077 14386 -27023
rect 14544 -27059 14580 -27023
rect 14248 -27201 14290 -27150
rect 14351 -27167 14385 -27077
rect 14449 -27145 14483 -27059
rect 14544 -27077 14581 -27059
rect 14444 -27201 14486 -27145
rect 14547 -27167 14581 -27077
rect 14645 -27146 14679 -27059
rect 14742 -27075 14778 -27023
rect 14638 -27201 14680 -27146
rect 14743 -27167 14777 -27075
rect 14834 -27082 14881 -26935
rect 14926 -26879 15100 -26847
rect 15250 -26879 15296 -26786
rect 15354 -26802 15388 -26643
rect 15452 -26786 15486 -26694
rect 15446 -26879 15492 -26786
rect 15550 -26802 15584 -26643
rect 15708 -26836 15768 -26692
rect 15897 -26786 15931 -26694
rect 14926 -26917 15492 -26879
rect 15528 -26898 15768 -26836
rect 15891 -26847 15937 -26786
rect 15995 -26802 16029 -26643
rect 16093 -26786 16127 -26694
rect 15804 -26879 15937 -26847
rect 16087 -26879 16133 -26786
rect 16191 -26802 16225 -26643
rect 16289 -26786 16323 -26694
rect 16283 -26879 16329 -26786
rect 16387 -26802 16421 -26643
rect 16492 -26836 16540 -26464
rect 15528 -26899 15731 -26898
rect 15528 -26910 15696 -26899
rect 14926 -26941 14999 -26917
rect 14841 -27156 14875 -27082
rect 14925 -27109 14999 -26941
rect 15054 -26925 15492 -26917
rect 15054 -26990 15100 -26925
rect 14840 -27201 14876 -27156
rect 15060 -27182 15094 -26990
rect 14248 -27235 14876 -27201
rect 15250 -26990 15296 -26925
rect 15256 -27182 15290 -26990
rect 15446 -27178 15492 -26925
rect 15804 -26917 16329 -26879
rect 16365 -26880 16540 -26836
rect 16365 -26910 16533 -26880
rect 15452 -27182 15486 -27178
rect 15650 -27047 15707 -26996
rect 15804 -27047 15850 -26917
rect 15891 -26925 16329 -26917
rect 15891 -26990 15937 -26925
rect 15650 -27096 15850 -27047
rect 15650 -27160 15707 -27096
rect 15897 -27182 15931 -26990
rect 16087 -26990 16133 -26925
rect 16093 -27182 16127 -26990
rect 16283 -27178 16329 -26925
rect 16289 -27182 16323 -27178
rect 25889 -27137 26035 -23387
rect 26685 -23555 26761 -23387
rect 26685 -23631 26827 -23555
rect 26751 -24020 26827 -23631
rect 27760 -23597 28425 -23569
rect 27760 -23655 28795 -23597
rect 27760 -23736 27846 -23655
rect 28020 -23692 28055 -23655
rect 28345 -23658 28795 -23655
rect 26908 -23822 27846 -23736
rect 26751 -24112 26886 -24020
rect 27048 -24078 27082 -23822
rect 27146 -24078 27180 -23870
rect 27244 -24078 27278 -23822
rect 27342 -24044 27376 -23870
rect 27923 -24000 27957 -23692
rect 28021 -24000 28055 -23692
rect 28119 -24000 28153 -23692
rect 28217 -24000 28251 -23692
rect 28315 -24000 28349 -23692
rect 27891 -24043 27962 -24042
rect 28303 -24043 28377 -24037
rect 27891 -24044 28377 -24043
rect 27342 -24078 28377 -24044
rect 28734 -24065 28795 -23658
rect 27343 -24082 28377 -24078
rect 27343 -24084 27892 -24082
rect 26930 -24112 27003 -24106
rect 28303 -24108 28377 -24082
rect 26751 -24129 27003 -24112
rect 26756 -24153 27003 -24129
rect 27838 -24140 27973 -24132
rect 27818 -24142 27973 -24140
rect 26756 -24170 26886 -24153
rect 26930 -24166 27003 -24153
rect 27611 -24178 27973 -24142
rect 28490 -24151 29275 -24065
rect 27818 -24180 27973 -24178
rect 27838 -24186 27973 -24180
rect 28021 -24163 28440 -24155
rect 28021 -24193 28451 -24163
rect 27048 -24408 27082 -24200
rect 27244 -24408 27278 -24200
rect 27440 -24408 27474 -24200
rect 28021 -24537 28055 -24193
rect 28217 -24537 28251 -24193
rect 28390 -24342 28451 -24193
rect 28630 -24307 28664 -24151
rect 28728 -24307 28762 -24199
rect 28826 -24307 28860 -24151
rect 28924 -24307 28958 -24199
rect 28512 -24342 28585 -24336
rect 28390 -24355 28585 -24342
rect 28412 -24383 28585 -24355
rect 28512 -24396 28585 -24383
rect 29022 -24366 29394 -24296
rect 28630 -24538 28664 -24430
rect 28826 -24538 28860 -24430
rect 29022 -24538 29056 -24366
rect 27022 -25473 27056 -25129
rect 27218 -25473 27252 -25129
rect 27631 -25236 27665 -25128
rect 27827 -25236 27861 -25128
rect 27513 -25283 27586 -25270
rect 27413 -25311 27586 -25283
rect 27391 -25324 27586 -25311
rect 27391 -25473 27452 -25324
rect 27513 -25330 27586 -25324
rect 28023 -25300 28057 -25128
rect 27022 -25503 27452 -25473
rect 27022 -25511 27441 -25503
rect 27631 -25515 27665 -25359
rect 27729 -25467 27763 -25359
rect 27827 -25515 27861 -25359
rect 27925 -25467 27959 -25359
rect 28023 -25370 28301 -25300
rect 24023 -27139 26035 -27137
rect 26666 -25584 26893 -25582
rect 27304 -25584 27378 -25558
rect 26666 -25622 27378 -25584
rect 27491 -25601 28106 -25515
rect 26892 -25623 27378 -25622
rect 26892 -25624 26963 -25623
rect 27304 -25629 27378 -25623
rect 26924 -25974 26958 -25666
rect 27022 -25974 27056 -25666
rect 27120 -25974 27154 -25666
rect 27218 -25974 27252 -25666
rect 27316 -25974 27350 -25666
rect 27021 -26026 27056 -25974
rect 27735 -26008 27796 -25601
rect 28225 -25765 28295 -25370
rect 28469 -25624 28503 -25040
rect 28676 -25006 28916 -24972
rect 28676 -25048 28718 -25006
rect 28465 -25683 28507 -25624
rect 28680 -25630 28714 -25048
rect 28778 -25628 28812 -25040
rect 28874 -25050 28916 -25006
rect 28677 -25683 28719 -25630
rect 28465 -25719 28719 -25683
rect 28774 -25682 28816 -25628
rect 28876 -25648 28910 -25050
rect 29088 -25634 29122 -25040
rect 28774 -25721 28915 -25682
rect 28872 -25733 28915 -25721
rect 28630 -25765 28785 -25755
rect 28225 -25801 28785 -25765
rect 28225 -25803 28295 -25801
rect 28630 -25810 28785 -25801
rect 28872 -25788 29053 -25733
rect 28872 -25858 28915 -25788
rect 28360 -25872 28515 -25863
rect 28323 -25906 28515 -25872
rect 28360 -25918 28515 -25906
rect 28561 -25898 28915 -25858
rect 29087 -25878 29130 -25634
rect 29324 -25703 29394 -24366
rect 29569 -23654 29661 -23569
rect 29592 -25629 29635 -23654
rect 29919 -24077 29995 -23373
rect 30221 -23329 32008 -23291
rect 30221 -23707 30259 -23329
rect 31428 -23628 32093 -23600
rect 31428 -23686 32463 -23628
rect 30198 -23761 30271 -23707
rect 31428 -23767 31514 -23686
rect 31688 -23723 31723 -23686
rect 32013 -23689 32463 -23686
rect 30576 -23853 31514 -23767
rect 30424 -24077 30554 -24051
rect 29919 -24143 30554 -24077
rect 30716 -24109 30750 -23853
rect 30814 -24109 30848 -23901
rect 30912 -24109 30946 -23853
rect 31010 -24075 31044 -23901
rect 31591 -24031 31625 -23723
rect 31689 -24031 31723 -23723
rect 31787 -24031 31821 -23723
rect 31885 -24031 31919 -23723
rect 31983 -24031 32017 -23723
rect 31559 -24074 31630 -24073
rect 31971 -24074 32045 -24068
rect 31559 -24075 32045 -24074
rect 31010 -24109 32045 -24075
rect 32402 -24096 32463 -23689
rect 34199 -22046 34847 -21992
rect 35470 -22031 35504 -21687
rect 35666 -22031 35700 -21687
rect 36079 -21794 36113 -21686
rect 36275 -21794 36309 -21686
rect 35961 -21841 36034 -21828
rect 35861 -21869 36034 -21841
rect 35839 -21882 36034 -21869
rect 35839 -22031 35900 -21882
rect 35961 -21888 36034 -21882
rect 36471 -21858 36505 -21686
rect 35287 -22044 35422 -22038
rect 35267 -22046 35422 -22044
rect 34199 -22082 35422 -22046
rect 35470 -22061 35900 -22031
rect 35470 -22069 35889 -22061
rect 36079 -22073 36113 -21917
rect 36177 -22025 36211 -21917
rect 36275 -22073 36309 -21917
rect 36373 -22025 36407 -21917
rect 36471 -21928 36749 -21858
rect 34199 -22138 34847 -22082
rect 35267 -22084 35422 -22082
rect 35287 -22092 35422 -22084
rect 31011 -24113 32045 -24109
rect 31011 -24115 31560 -24113
rect 30598 -24143 30671 -24137
rect 31971 -24139 32045 -24113
rect 29919 -24153 30671 -24143
rect 30424 -24184 30671 -24153
rect 31506 -24171 31641 -24163
rect 31486 -24173 31641 -24171
rect 30424 -24201 30554 -24184
rect 30598 -24197 30671 -24184
rect 30451 -24251 30527 -24201
rect 31279 -24209 31641 -24173
rect 32158 -24182 32943 -24096
rect 31486 -24211 31641 -24209
rect 31506 -24217 31641 -24211
rect 31689 -24194 32108 -24186
rect 31689 -24224 32119 -24194
rect 30716 -24439 30750 -24231
rect 30912 -24439 30946 -24231
rect 31108 -24439 31142 -24231
rect 31689 -24568 31723 -24224
rect 31885 -24568 31919 -24224
rect 32058 -24373 32119 -24224
rect 32298 -24338 32332 -24182
rect 32396 -24338 32430 -24230
rect 32494 -24338 32528 -24182
rect 32592 -24338 32626 -24230
rect 32180 -24373 32253 -24367
rect 32058 -24386 32253 -24373
rect 32080 -24414 32253 -24386
rect 32180 -24427 32253 -24414
rect 32690 -24397 33062 -24327
rect 32298 -24569 32332 -24461
rect 32494 -24569 32528 -24461
rect 32690 -24569 32724 -24397
rect 30690 -25504 30724 -25160
rect 30886 -25504 30920 -25160
rect 31299 -25267 31333 -25159
rect 31495 -25267 31529 -25159
rect 31181 -25314 31254 -25301
rect 31081 -25342 31254 -25314
rect 31059 -25355 31254 -25342
rect 31059 -25504 31120 -25355
rect 31181 -25361 31254 -25355
rect 31691 -25331 31725 -25159
rect 30690 -25534 31120 -25504
rect 30690 -25542 31109 -25534
rect 31299 -25546 31333 -25390
rect 31397 -25498 31431 -25390
rect 31495 -25546 31529 -25390
rect 31593 -25498 31627 -25390
rect 31691 -25401 31969 -25331
rect 29592 -25672 29877 -25629
rect 29313 -25775 29418 -25703
rect 29834 -25878 29877 -25672
rect 27346 -26026 27796 -26008
rect 26904 -26069 27796 -26026
rect 26904 -26087 27353 -26069
rect 27735 -26364 27796 -26069
rect 28469 -26246 28503 -25952
rect 28561 -25968 28606 -25898
rect 28953 -25918 29877 -25878
rect 29001 -25921 29877 -25918
rect 28462 -26364 28509 -26246
rect 28567 -26260 28601 -25968
rect 28665 -26245 28699 -25952
rect 28907 -26235 28941 -25952
rect 29001 -25961 29045 -25921
rect 28658 -26364 28705 -26245
rect 28900 -26364 28947 -26235
rect 29005 -26260 29039 -25961
rect 27735 -26477 29212 -26364
rect 30334 -25615 30561 -25613
rect 30972 -25615 31046 -25589
rect 30334 -25653 31046 -25615
rect 31159 -25632 31774 -25546
rect 30560 -25654 31046 -25653
rect 30560 -25655 30631 -25654
rect 30972 -25660 31046 -25654
rect 30592 -26005 30626 -25697
rect 30690 -26005 30724 -25697
rect 30788 -26005 30822 -25697
rect 30886 -26005 30920 -25697
rect 30984 -26005 31018 -25697
rect 30689 -26057 30724 -26005
rect 31403 -26039 31464 -25632
rect 31893 -25796 31963 -25401
rect 32137 -25655 32171 -25071
rect 32344 -25037 32584 -25003
rect 32344 -25079 32386 -25037
rect 32133 -25714 32175 -25655
rect 32348 -25661 32382 -25079
rect 32446 -25659 32480 -25071
rect 32542 -25081 32584 -25037
rect 32345 -25714 32387 -25661
rect 32133 -25750 32387 -25714
rect 32442 -25713 32484 -25659
rect 32544 -25679 32578 -25081
rect 32756 -25665 32790 -25071
rect 32442 -25752 32583 -25713
rect 32540 -25764 32583 -25752
rect 32298 -25796 32453 -25786
rect 31893 -25832 32453 -25796
rect 31893 -25834 31963 -25832
rect 32298 -25841 32453 -25832
rect 32540 -25819 32721 -25764
rect 32540 -25889 32583 -25819
rect 32028 -25903 32183 -25894
rect 31991 -25937 32183 -25903
rect 32028 -25949 32183 -25937
rect 32229 -25929 32583 -25889
rect 32755 -25909 32798 -25665
rect 32992 -25734 33062 -24397
rect 32981 -25806 33086 -25734
rect 33487 -25909 33710 -25819
rect 31014 -26057 31464 -26039
rect 30572 -26100 31464 -26057
rect 30572 -26118 31021 -26100
rect 31403 -26395 31464 -26100
rect 32137 -26277 32171 -25983
rect 32229 -25999 32274 -25929
rect 32621 -25949 33823 -25909
rect 32669 -25952 33823 -25949
rect 32130 -26395 32177 -26277
rect 32235 -26291 32269 -25999
rect 32333 -26276 32367 -25983
rect 32575 -26266 32609 -25983
rect 32669 -25992 32713 -25952
rect 33487 -25989 33710 -25952
rect 32326 -26395 32373 -26276
rect 32568 -26395 32615 -26266
rect 32673 -26291 32707 -25992
rect 31403 -26508 32880 -26395
rect 24023 -27307 26054 -27139
rect 24023 -27308 25978 -27307
rect 8885 -27645 9013 -27466
rect 25904 -27701 26125 -27506
rect 34199 -27521 34345 -22138
rect 35114 -22142 35341 -22140
rect 35752 -22142 35826 -22116
rect 35114 -22180 35826 -22142
rect 35939 -22159 36554 -22073
rect 35125 -23030 35201 -22180
rect 35340 -22181 35826 -22180
rect 35340 -22182 35411 -22181
rect 35752 -22187 35826 -22181
rect 35372 -22532 35406 -22224
rect 35470 -22532 35504 -22224
rect 35568 -22532 35602 -22224
rect 35666 -22532 35700 -22224
rect 35764 -22532 35798 -22224
rect 35469 -22584 35504 -22532
rect 36183 -22566 36244 -22159
rect 36673 -22323 36743 -21928
rect 36917 -22182 36951 -21598
rect 37124 -21564 37364 -21530
rect 37124 -21606 37166 -21564
rect 36913 -22241 36955 -22182
rect 37128 -22188 37162 -21606
rect 37226 -22186 37260 -21598
rect 37322 -21608 37364 -21564
rect 37125 -22241 37167 -22188
rect 36913 -22277 37167 -22241
rect 37222 -22240 37264 -22186
rect 37324 -22206 37358 -21608
rect 37536 -22192 37570 -21598
rect 37222 -22279 37363 -22240
rect 37320 -22291 37363 -22279
rect 37078 -22323 37233 -22313
rect 36673 -22359 37233 -22323
rect 36673 -22361 36743 -22359
rect 37078 -22368 37233 -22359
rect 37320 -22346 37501 -22291
rect 37320 -22416 37363 -22346
rect 36808 -22430 36963 -22421
rect 36771 -22464 36963 -22430
rect 36808 -22476 36963 -22464
rect 37009 -22456 37363 -22416
rect 37535 -22436 37578 -22192
rect 37772 -22261 37842 -20924
rect 44359 -21005 44393 -20797
rect 44555 -21005 44589 -20797
rect 44751 -21005 44785 -20797
rect 45332 -21134 45366 -20790
rect 45528 -21134 45562 -20790
rect 45701 -20939 45762 -20790
rect 45941 -20904 45975 -20748
rect 46039 -20904 46073 -20796
rect 46137 -20904 46171 -20748
rect 54347 -20749 54482 -20743
rect 54530 -20726 54949 -20718
rect 54530 -20756 54960 -20726
rect 46235 -20904 46269 -20796
rect 45823 -20939 45896 -20933
rect 45701 -20952 45896 -20939
rect 45723 -20980 45896 -20952
rect 45823 -20993 45896 -20980
rect 46333 -20963 46705 -20893
rect 45941 -21135 45975 -21027
rect 46137 -21135 46171 -21027
rect 46333 -21135 46367 -20963
rect 38909 -21956 38943 -21456
rect 39088 -21420 39409 -21386
rect 38908 -22002 38943 -21956
rect 39088 -22002 39128 -21420
rect 39177 -21460 39212 -21420
rect 39178 -21964 39212 -21460
rect 39276 -21957 39310 -21456
rect 39374 -21459 39409 -21420
rect 38908 -22042 39128 -22002
rect 39273 -22077 39311 -21957
rect 39374 -21964 39408 -21459
rect 39504 -22040 39538 -21456
rect 39830 -21970 39864 -21456
rect 40058 -21746 40092 -21456
rect 40057 -21839 40094 -21746
rect 40057 -21876 40194 -21839
rect 39830 -22004 39989 -21970
rect 39653 -22040 39791 -22029
rect 38909 -22115 39311 -22077
rect 39378 -22074 39791 -22040
rect 38672 -22126 38810 -22116
rect 38282 -22160 38810 -22126
rect 37761 -22333 37866 -22261
rect 38282 -22436 38325 -22160
rect 38672 -22170 38810 -22160
rect 38728 -22261 38866 -22252
rect 38518 -22295 38866 -22261
rect 38518 -22422 38590 -22295
rect 38728 -22306 38866 -22295
rect 38518 -22431 38602 -22422
rect 35794 -22584 36244 -22566
rect 35352 -22627 36244 -22584
rect 35352 -22645 35801 -22627
rect 34469 -23176 35201 -23030
rect 36183 -22922 36244 -22627
rect 36917 -22804 36951 -22510
rect 37009 -22526 37054 -22456
rect 37401 -22476 38325 -22436
rect 37449 -22479 38325 -22476
rect 36910 -22922 36957 -22804
rect 37015 -22818 37049 -22526
rect 37113 -22803 37147 -22510
rect 37355 -22793 37389 -22510
rect 37449 -22519 37493 -22479
rect 38523 -22501 38602 -22431
rect 37106 -22922 37153 -22803
rect 37348 -22922 37395 -22793
rect 37453 -22818 37487 -22519
rect 38811 -22743 38845 -22452
rect 38809 -22854 38846 -22743
rect 38909 -22760 38943 -22115
rect 39138 -22185 39176 -22115
rect 39378 -22153 39412 -22074
rect 39653 -22083 39791 -22074
rect 39128 -22323 39182 -22185
rect 39281 -22187 39412 -22153
rect 39478 -22170 39616 -22116
rect 39863 -22185 39917 -22047
rect 39955 -22048 39989 -22004
rect 39955 -22102 40121 -22048
rect 39281 -22760 39315 -22187
rect 39955 -22217 39989 -22102
rect 40041 -22217 40095 -22200
rect 39379 -22256 39538 -22221
rect 39955 -22222 40095 -22217
rect 39927 -22251 40095 -22222
rect 39379 -22760 39413 -22256
rect 39504 -22760 39538 -22256
rect 39602 -22743 39636 -22252
rect 39732 -22742 39766 -22252
rect 38272 -22858 38883 -22854
rect 39601 -22858 39638 -22743
rect 39729 -22858 39766 -22742
rect 39830 -22760 39864 -22252
rect 39927 -22256 39989 -22251
rect 39928 -22760 39962 -22256
rect 40041 -22259 40095 -22251
rect 40156 -22369 40194 -21876
rect 40156 -22407 40448 -22369
rect 40058 -22741 40092 -22452
rect 40156 -22457 40194 -22407
rect 40056 -22858 40093 -22741
rect 40156 -22760 40190 -22457
rect 38272 -22922 40206 -22858
rect 36183 -22967 40206 -22922
rect 36183 -23035 38385 -22967
rect 38733 -23019 40206 -22967
rect 34469 -27159 34615 -23176
rect 35125 -23308 35201 -23176
rect 40410 -23302 40448 -22407
rect 35125 -23384 38435 -23308
rect 35125 -23566 35201 -23384
rect 35125 -23642 35267 -23566
rect 35191 -24031 35267 -23642
rect 36200 -23608 36865 -23580
rect 36200 -23666 37235 -23608
rect 36200 -23747 36286 -23666
rect 36460 -23703 36495 -23666
rect 36785 -23669 37235 -23666
rect 35348 -23833 36286 -23747
rect 35191 -24123 35326 -24031
rect 35488 -24089 35522 -23833
rect 35586 -24089 35620 -23881
rect 35684 -24089 35718 -23833
rect 35782 -24055 35816 -23881
rect 36363 -24011 36397 -23703
rect 36461 -24011 36495 -23703
rect 36559 -24011 36593 -23703
rect 36657 -24011 36691 -23703
rect 36755 -24011 36789 -23703
rect 36331 -24054 36402 -24053
rect 36743 -24054 36817 -24048
rect 36331 -24055 36817 -24054
rect 35782 -24089 36817 -24055
rect 37174 -24076 37235 -23669
rect 35783 -24093 36817 -24089
rect 35783 -24095 36332 -24093
rect 35370 -24123 35443 -24117
rect 36743 -24119 36817 -24093
rect 35191 -24140 35443 -24123
rect 35196 -24164 35443 -24140
rect 36278 -24151 36413 -24143
rect 36258 -24153 36413 -24151
rect 35196 -24181 35326 -24164
rect 35370 -24177 35443 -24164
rect 36051 -24189 36413 -24153
rect 36930 -24162 37715 -24076
rect 36258 -24191 36413 -24189
rect 36278 -24197 36413 -24191
rect 36461 -24174 36880 -24166
rect 36461 -24204 36891 -24174
rect 35488 -24419 35522 -24211
rect 35684 -24419 35718 -24211
rect 35880 -24419 35914 -24211
rect 36461 -24548 36495 -24204
rect 36657 -24548 36691 -24204
rect 36830 -24353 36891 -24204
rect 37070 -24318 37104 -24162
rect 37168 -24318 37202 -24210
rect 37266 -24318 37300 -24162
rect 37364 -24318 37398 -24210
rect 36952 -24353 37025 -24347
rect 36830 -24366 37025 -24353
rect 36852 -24394 37025 -24366
rect 36952 -24407 37025 -24394
rect 37462 -24377 37834 -24307
rect 37070 -24549 37104 -24441
rect 37266 -24549 37300 -24441
rect 37462 -24549 37496 -24377
rect 35462 -25484 35496 -25140
rect 35658 -25484 35692 -25140
rect 36071 -25247 36105 -25139
rect 36267 -25247 36301 -25139
rect 35953 -25294 36026 -25281
rect 35853 -25322 36026 -25294
rect 35831 -25335 36026 -25322
rect 35831 -25484 35892 -25335
rect 35953 -25341 36026 -25335
rect 36463 -25311 36497 -25139
rect 35462 -25514 35892 -25484
rect 35462 -25522 35881 -25514
rect 36071 -25526 36105 -25370
rect 36169 -25478 36203 -25370
rect 36267 -25526 36301 -25370
rect 36365 -25478 36399 -25370
rect 36463 -25381 36741 -25311
rect 35106 -25595 35333 -25593
rect 35744 -25595 35818 -25569
rect 35106 -25633 35818 -25595
rect 35931 -25612 36546 -25526
rect 35332 -25634 35818 -25633
rect 35332 -25635 35403 -25634
rect 35744 -25640 35818 -25634
rect 35364 -25985 35398 -25677
rect 35462 -25985 35496 -25677
rect 35560 -25985 35594 -25677
rect 35658 -25985 35692 -25677
rect 35756 -25985 35790 -25677
rect 35461 -26037 35496 -25985
rect 36175 -26019 36236 -25612
rect 36665 -25776 36735 -25381
rect 36909 -25635 36943 -25051
rect 37116 -25017 37356 -24983
rect 37116 -25059 37158 -25017
rect 36905 -25694 36947 -25635
rect 37120 -25641 37154 -25059
rect 37218 -25639 37252 -25051
rect 37314 -25061 37356 -25017
rect 37117 -25694 37159 -25641
rect 36905 -25730 37159 -25694
rect 37214 -25693 37256 -25639
rect 37316 -25659 37350 -25061
rect 37528 -25645 37562 -25051
rect 37214 -25732 37355 -25693
rect 37312 -25744 37355 -25732
rect 37070 -25776 37225 -25766
rect 36665 -25812 37225 -25776
rect 36665 -25814 36735 -25812
rect 37070 -25821 37225 -25812
rect 37312 -25799 37493 -25744
rect 37312 -25869 37355 -25799
rect 36800 -25883 36955 -25874
rect 36763 -25917 36955 -25883
rect 36800 -25929 36955 -25917
rect 37001 -25909 37355 -25869
rect 37527 -25889 37570 -25645
rect 37764 -25714 37834 -24377
rect 38009 -23665 38101 -23580
rect 38032 -25640 38075 -23665
rect 38359 -24088 38435 -23384
rect 38661 -23340 40448 -23302
rect 38661 -23718 38699 -23340
rect 39868 -23639 40533 -23611
rect 39868 -23697 40903 -23639
rect 38638 -23772 38711 -23718
rect 39868 -23778 39954 -23697
rect 40128 -23734 40163 -23697
rect 40453 -23700 40903 -23697
rect 39016 -23864 39954 -23778
rect 38864 -24088 38994 -24062
rect 38359 -24154 38994 -24088
rect 39156 -24120 39190 -23864
rect 39254 -24120 39288 -23912
rect 39352 -24120 39386 -23864
rect 39450 -24086 39484 -23912
rect 40031 -24042 40065 -23734
rect 40129 -24042 40163 -23734
rect 40227 -24042 40261 -23734
rect 40325 -24042 40359 -23734
rect 40423 -24042 40457 -23734
rect 39999 -24085 40070 -24084
rect 40411 -24085 40485 -24079
rect 39999 -24086 40485 -24085
rect 39450 -24120 40485 -24086
rect 40842 -24107 40903 -23700
rect 44333 -22070 44367 -21726
rect 44529 -22070 44563 -21726
rect 44942 -21833 44976 -21725
rect 45138 -21833 45172 -21725
rect 44824 -21880 44897 -21867
rect 44724 -21908 44897 -21880
rect 44702 -21921 44897 -21908
rect 44702 -22070 44763 -21921
rect 44824 -21927 44897 -21921
rect 45334 -21897 45368 -21725
rect 42881 -22085 43648 -22078
rect 44150 -22083 44285 -22077
rect 44130 -22085 44285 -22083
rect 42881 -22121 44285 -22085
rect 44333 -22100 44763 -22070
rect 44333 -22108 44752 -22100
rect 44942 -22112 44976 -21956
rect 45040 -22064 45074 -21956
rect 45138 -22112 45172 -21956
rect 45236 -22064 45270 -21956
rect 45334 -21967 45612 -21897
rect 42881 -22224 43648 -22121
rect 44130 -22123 44285 -22121
rect 44150 -22131 44285 -22123
rect 43977 -22181 44204 -22179
rect 44615 -22181 44689 -22155
rect 43977 -22219 44689 -22181
rect 44802 -22198 45417 -22112
rect 39451 -24124 40485 -24120
rect 39451 -24126 40000 -24124
rect 39038 -24154 39111 -24148
rect 40411 -24150 40485 -24124
rect 38359 -24164 39111 -24154
rect 38864 -24195 39111 -24164
rect 39946 -24182 40081 -24174
rect 39926 -24184 40081 -24182
rect 38864 -24212 38994 -24195
rect 39038 -24208 39111 -24195
rect 38891 -24262 38967 -24212
rect 39719 -24220 40081 -24184
rect 40598 -24193 41383 -24107
rect 39926 -24222 40081 -24220
rect 39946 -24228 40081 -24222
rect 40129 -24205 40548 -24197
rect 40129 -24235 40559 -24205
rect 39156 -24450 39190 -24242
rect 39352 -24450 39386 -24242
rect 39548 -24450 39582 -24242
rect 40129 -24579 40163 -24235
rect 40325 -24579 40359 -24235
rect 40498 -24384 40559 -24235
rect 40738 -24349 40772 -24193
rect 40836 -24349 40870 -24241
rect 40934 -24349 40968 -24193
rect 41032 -24349 41066 -24241
rect 40620 -24384 40693 -24378
rect 40498 -24397 40693 -24384
rect 40520 -24425 40693 -24397
rect 40620 -24438 40693 -24425
rect 41130 -24408 41502 -24338
rect 40738 -24580 40772 -24472
rect 40934 -24580 40968 -24472
rect 41130 -24580 41164 -24408
rect 39130 -25515 39164 -25171
rect 39326 -25515 39360 -25171
rect 39739 -25278 39773 -25170
rect 39935 -25278 39969 -25170
rect 39621 -25325 39694 -25312
rect 39521 -25353 39694 -25325
rect 39499 -25366 39694 -25353
rect 39499 -25515 39560 -25366
rect 39621 -25372 39694 -25366
rect 40131 -25342 40165 -25170
rect 39130 -25545 39560 -25515
rect 39130 -25553 39549 -25545
rect 39739 -25557 39773 -25401
rect 39837 -25509 39871 -25401
rect 39935 -25557 39969 -25401
rect 40033 -25509 40067 -25401
rect 40131 -25412 40409 -25342
rect 38032 -25683 38317 -25640
rect 37753 -25786 37858 -25714
rect 38274 -25889 38317 -25683
rect 35786 -26037 36236 -26019
rect 35344 -26080 36236 -26037
rect 35344 -26098 35793 -26080
rect 36175 -26375 36236 -26080
rect 36909 -26257 36943 -25963
rect 37001 -25979 37046 -25909
rect 37393 -25929 38317 -25889
rect 37441 -25932 38317 -25929
rect 36902 -26375 36949 -26257
rect 37007 -26271 37041 -25979
rect 37105 -26256 37139 -25963
rect 37347 -26246 37381 -25963
rect 37441 -25972 37485 -25932
rect 37098 -26375 37145 -26256
rect 37340 -26375 37387 -26246
rect 37445 -26271 37479 -25972
rect 36175 -26488 37652 -26375
rect 38774 -25626 39001 -25624
rect 39412 -25626 39486 -25600
rect 38774 -25664 39486 -25626
rect 39599 -25643 40214 -25557
rect 39000 -25665 39486 -25664
rect 39000 -25666 39071 -25665
rect 39412 -25671 39486 -25665
rect 39032 -26016 39066 -25708
rect 39130 -26016 39164 -25708
rect 39228 -26016 39262 -25708
rect 39326 -26016 39360 -25708
rect 39424 -26016 39458 -25708
rect 39129 -26068 39164 -26016
rect 39843 -26050 39904 -25643
rect 40333 -25807 40403 -25412
rect 40577 -25666 40611 -25082
rect 40784 -25048 41024 -25014
rect 40784 -25090 40826 -25048
rect 40573 -25725 40615 -25666
rect 40788 -25672 40822 -25090
rect 40886 -25670 40920 -25082
rect 40982 -25092 41024 -25048
rect 40785 -25725 40827 -25672
rect 40573 -25761 40827 -25725
rect 40882 -25724 40924 -25670
rect 40984 -25690 41018 -25092
rect 41196 -25676 41230 -25082
rect 40882 -25763 41023 -25724
rect 40980 -25775 41023 -25763
rect 40738 -25807 40893 -25797
rect 40333 -25843 40893 -25807
rect 40333 -25845 40403 -25843
rect 40738 -25852 40893 -25843
rect 40980 -25830 41161 -25775
rect 40980 -25900 41023 -25830
rect 40468 -25914 40623 -25905
rect 40431 -25948 40623 -25914
rect 40468 -25960 40623 -25948
rect 40669 -25940 41023 -25900
rect 41195 -25920 41238 -25676
rect 41432 -25745 41502 -24408
rect 41421 -25817 41526 -25745
rect 41936 -25920 42273 -25757
rect 39454 -26068 39904 -26050
rect 39012 -26111 39904 -26068
rect 39012 -26129 39461 -26111
rect 39843 -26406 39904 -26111
rect 40577 -26288 40611 -25994
rect 40669 -26010 40714 -25940
rect 41061 -25960 42273 -25920
rect 41109 -25963 42273 -25960
rect 40570 -26406 40617 -26288
rect 40675 -26302 40709 -26010
rect 40773 -26287 40807 -25994
rect 41015 -26277 41049 -25994
rect 41109 -26003 41153 -25963
rect 40766 -26406 40813 -26287
rect 41008 -26406 41055 -26277
rect 41113 -26302 41147 -26003
rect 41936 -26088 42273 -25963
rect 39843 -26519 41320 -26406
rect 34446 -27306 34649 -27159
rect 34130 -27724 34404 -27521
rect 41577 -27340 41894 -27049
rect 41594 -28120 41860 -27340
rect 42881 -27539 43027 -22224
rect 43988 -23157 44064 -22219
rect 44203 -22220 44689 -22219
rect 44203 -22221 44274 -22220
rect 44615 -22226 44689 -22220
rect 44235 -22571 44269 -22263
rect 44333 -22571 44367 -22263
rect 44431 -22571 44465 -22263
rect 44529 -22571 44563 -22263
rect 44627 -22571 44661 -22263
rect 44332 -22623 44367 -22571
rect 45046 -22605 45107 -22198
rect 45536 -22362 45606 -21967
rect 45780 -22221 45814 -21637
rect 45987 -21603 46227 -21569
rect 45987 -21645 46029 -21603
rect 45776 -22280 45818 -22221
rect 45991 -22227 46025 -21645
rect 46089 -22225 46123 -21637
rect 46185 -21647 46227 -21603
rect 45988 -22280 46030 -22227
rect 45776 -22316 46030 -22280
rect 46085 -22279 46127 -22225
rect 46187 -22245 46221 -21647
rect 46399 -22231 46433 -21637
rect 46085 -22318 46226 -22279
rect 46183 -22330 46226 -22318
rect 45941 -22362 46096 -22352
rect 45536 -22398 46096 -22362
rect 45536 -22400 45606 -22398
rect 45941 -22407 46096 -22398
rect 46183 -22385 46364 -22330
rect 46183 -22455 46226 -22385
rect 45671 -22469 45826 -22460
rect 45634 -22503 45826 -22469
rect 45671 -22515 45826 -22503
rect 45872 -22495 46226 -22455
rect 46398 -22475 46441 -22231
rect 46635 -22300 46705 -20963
rect 53557 -20971 53591 -20763
rect 53753 -20971 53787 -20763
rect 53949 -20971 53983 -20763
rect 54530 -21100 54564 -20756
rect 54726 -21100 54760 -20756
rect 54899 -20905 54960 -20756
rect 55139 -20870 55173 -20714
rect 55237 -20870 55271 -20762
rect 55335 -20870 55369 -20714
rect 55433 -20870 55467 -20762
rect 55021 -20905 55094 -20899
rect 54899 -20918 55094 -20905
rect 54921 -20946 55094 -20918
rect 55021 -20959 55094 -20946
rect 55531 -20929 55903 -20859
rect 55139 -21101 55173 -20993
rect 55335 -21101 55369 -20993
rect 55531 -21101 55565 -20929
rect 47772 -21995 47806 -21495
rect 47951 -21459 48272 -21425
rect 47771 -22041 47806 -21995
rect 47951 -22041 47991 -21459
rect 48040 -21499 48075 -21459
rect 48041 -22003 48075 -21499
rect 48139 -21996 48173 -21495
rect 48237 -21498 48272 -21459
rect 47771 -22081 47991 -22041
rect 48136 -22116 48174 -21996
rect 48237 -22003 48271 -21498
rect 48367 -22079 48401 -21495
rect 48693 -22009 48727 -21495
rect 48921 -21785 48955 -21495
rect 48920 -21878 48957 -21785
rect 48920 -21915 49057 -21878
rect 48693 -22043 48852 -22009
rect 48516 -22079 48654 -22068
rect 47772 -22154 48174 -22116
rect 48241 -22113 48654 -22079
rect 47535 -22165 47673 -22155
rect 47145 -22199 47673 -22165
rect 46624 -22372 46729 -22300
rect 47145 -22475 47188 -22199
rect 47535 -22209 47673 -22199
rect 47591 -22300 47729 -22291
rect 47381 -22334 47729 -22300
rect 47381 -22461 47453 -22334
rect 47591 -22345 47729 -22334
rect 47381 -22470 47465 -22461
rect 44657 -22623 45107 -22605
rect 44215 -22666 45107 -22623
rect 44215 -22684 44664 -22666
rect 45046 -22961 45107 -22666
rect 45780 -22843 45814 -22549
rect 45872 -22565 45917 -22495
rect 46264 -22515 47188 -22475
rect 46312 -22518 47188 -22515
rect 45773 -22961 45820 -22843
rect 45878 -22857 45912 -22565
rect 45976 -22842 46010 -22549
rect 46218 -22832 46252 -22549
rect 46312 -22558 46356 -22518
rect 47386 -22540 47465 -22470
rect 45969 -22961 46016 -22842
rect 46211 -22961 46258 -22832
rect 46316 -22857 46350 -22558
rect 47674 -22782 47708 -22491
rect 47672 -22893 47709 -22782
rect 47772 -22799 47806 -22154
rect 48001 -22224 48039 -22154
rect 48241 -22192 48275 -22113
rect 48516 -22122 48654 -22113
rect 47991 -22362 48045 -22224
rect 48144 -22226 48275 -22192
rect 48341 -22209 48479 -22155
rect 48726 -22224 48780 -22086
rect 48818 -22087 48852 -22043
rect 48818 -22141 48984 -22087
rect 48144 -22799 48178 -22226
rect 48818 -22256 48852 -22141
rect 48904 -22256 48958 -22239
rect 48242 -22295 48401 -22260
rect 48818 -22261 48958 -22256
rect 48790 -22290 48958 -22261
rect 48242 -22799 48276 -22295
rect 48367 -22799 48401 -22295
rect 48465 -22782 48499 -22291
rect 48595 -22781 48629 -22291
rect 47135 -22897 47746 -22893
rect 48464 -22897 48501 -22782
rect 48592 -22897 48629 -22781
rect 48693 -22799 48727 -22291
rect 48790 -22295 48852 -22290
rect 48791 -22799 48825 -22295
rect 48904 -22298 48958 -22290
rect 49019 -22408 49057 -21915
rect 49019 -22446 49311 -22408
rect 48921 -22780 48955 -22491
rect 49019 -22496 49057 -22446
rect 48919 -22897 48956 -22780
rect 49019 -22799 49053 -22496
rect 47135 -22961 49069 -22897
rect 45046 -23006 49069 -22961
rect 45046 -23074 47248 -23006
rect 47596 -23058 49069 -23006
rect 43338 -23303 44064 -23157
rect 43338 -27304 43484 -23303
rect 43988 -23347 44064 -23303
rect 49273 -23341 49311 -22446
rect 43988 -23423 47298 -23347
rect 43988 -23605 44064 -23423
rect 43988 -23681 44130 -23605
rect 44054 -24070 44130 -23681
rect 45063 -23647 45728 -23619
rect 45063 -23705 46098 -23647
rect 45063 -23786 45149 -23705
rect 45323 -23742 45358 -23705
rect 45648 -23708 46098 -23705
rect 44211 -23872 45149 -23786
rect 44054 -24162 44189 -24070
rect 44351 -24128 44385 -23872
rect 44449 -24128 44483 -23920
rect 44547 -24128 44581 -23872
rect 44645 -24094 44679 -23920
rect 45226 -24050 45260 -23742
rect 45324 -24050 45358 -23742
rect 45422 -24050 45456 -23742
rect 45520 -24050 45554 -23742
rect 45618 -24050 45652 -23742
rect 45194 -24093 45265 -24092
rect 45606 -24093 45680 -24087
rect 45194 -24094 45680 -24093
rect 44645 -24128 45680 -24094
rect 46037 -24115 46098 -23708
rect 44646 -24132 45680 -24128
rect 44646 -24134 45195 -24132
rect 44233 -24162 44306 -24156
rect 45606 -24158 45680 -24132
rect 44054 -24179 44306 -24162
rect 44059 -24203 44306 -24179
rect 45141 -24190 45276 -24182
rect 45121 -24192 45276 -24190
rect 44059 -24220 44189 -24203
rect 44233 -24216 44306 -24203
rect 44914 -24228 45276 -24192
rect 45793 -24201 46578 -24115
rect 45121 -24230 45276 -24228
rect 45141 -24236 45276 -24230
rect 45324 -24213 45743 -24205
rect 45324 -24243 45754 -24213
rect 44351 -24458 44385 -24250
rect 44547 -24458 44581 -24250
rect 44743 -24458 44777 -24250
rect 45324 -24587 45358 -24243
rect 45520 -24587 45554 -24243
rect 45693 -24392 45754 -24243
rect 45933 -24357 45967 -24201
rect 46031 -24357 46065 -24249
rect 46129 -24357 46163 -24201
rect 46227 -24357 46261 -24249
rect 45815 -24392 45888 -24386
rect 45693 -24405 45888 -24392
rect 45715 -24433 45888 -24405
rect 45815 -24446 45888 -24433
rect 46325 -24416 46697 -24346
rect 45933 -24588 45967 -24480
rect 46129 -24588 46163 -24480
rect 46325 -24588 46359 -24416
rect 44325 -25523 44359 -25179
rect 44521 -25523 44555 -25179
rect 44934 -25286 44968 -25178
rect 45130 -25286 45164 -25178
rect 44816 -25333 44889 -25320
rect 44716 -25361 44889 -25333
rect 44694 -25374 44889 -25361
rect 44694 -25523 44755 -25374
rect 44816 -25380 44889 -25374
rect 45326 -25350 45360 -25178
rect 44325 -25553 44755 -25523
rect 44325 -25561 44744 -25553
rect 44934 -25565 44968 -25409
rect 45032 -25517 45066 -25409
rect 45130 -25565 45164 -25409
rect 45228 -25517 45262 -25409
rect 45326 -25420 45604 -25350
rect 43969 -25634 44196 -25632
rect 44607 -25634 44681 -25608
rect 43969 -25672 44681 -25634
rect 44794 -25651 45409 -25565
rect 44195 -25673 44681 -25672
rect 44195 -25674 44266 -25673
rect 44607 -25679 44681 -25673
rect 44227 -26024 44261 -25716
rect 44325 -26024 44359 -25716
rect 44423 -26024 44457 -25716
rect 44521 -26024 44555 -25716
rect 44619 -26024 44653 -25716
rect 44324 -26076 44359 -26024
rect 45038 -26058 45099 -25651
rect 45528 -25815 45598 -25420
rect 45772 -25674 45806 -25090
rect 45979 -25056 46219 -25022
rect 45979 -25098 46021 -25056
rect 45768 -25733 45810 -25674
rect 45983 -25680 46017 -25098
rect 46081 -25678 46115 -25090
rect 46177 -25100 46219 -25056
rect 45980 -25733 46022 -25680
rect 45768 -25769 46022 -25733
rect 46077 -25732 46119 -25678
rect 46179 -25698 46213 -25100
rect 46391 -25684 46425 -25090
rect 46077 -25771 46218 -25732
rect 46175 -25783 46218 -25771
rect 45933 -25815 46088 -25805
rect 45528 -25851 46088 -25815
rect 45528 -25853 45598 -25851
rect 45933 -25860 46088 -25851
rect 46175 -25838 46356 -25783
rect 46175 -25908 46218 -25838
rect 45663 -25922 45818 -25913
rect 45626 -25956 45818 -25922
rect 45663 -25968 45818 -25956
rect 45864 -25948 46218 -25908
rect 46390 -25928 46433 -25684
rect 46627 -25753 46697 -24416
rect 46872 -23704 46964 -23619
rect 46895 -25679 46938 -23704
rect 47222 -24127 47298 -23423
rect 47524 -23379 49311 -23341
rect 47524 -23757 47562 -23379
rect 48731 -23678 49396 -23650
rect 48731 -23736 49766 -23678
rect 47501 -23811 47574 -23757
rect 48731 -23817 48817 -23736
rect 48991 -23773 49026 -23736
rect 49316 -23739 49766 -23736
rect 47879 -23903 48817 -23817
rect 47727 -24127 47857 -24101
rect 47222 -24193 47857 -24127
rect 48019 -24159 48053 -23903
rect 48117 -24159 48151 -23951
rect 48215 -24159 48249 -23903
rect 48313 -24125 48347 -23951
rect 48894 -24081 48928 -23773
rect 48992 -24081 49026 -23773
rect 49090 -24081 49124 -23773
rect 49188 -24081 49222 -23773
rect 49286 -24081 49320 -23773
rect 48862 -24124 48933 -24123
rect 49274 -24124 49348 -24118
rect 48862 -24125 49348 -24124
rect 48313 -24159 49348 -24125
rect 49705 -24146 49766 -23739
rect 52200 -22051 52929 -21986
rect 53531 -22036 53565 -21692
rect 53727 -22036 53761 -21692
rect 54140 -21799 54174 -21691
rect 54336 -21799 54370 -21691
rect 54022 -21846 54095 -21833
rect 53922 -21874 54095 -21846
rect 53900 -21887 54095 -21874
rect 53900 -22036 53961 -21887
rect 54022 -21893 54095 -21887
rect 54532 -21863 54566 -21691
rect 53348 -22049 53483 -22043
rect 53328 -22051 53483 -22049
rect 52200 -22087 53483 -22051
rect 53531 -22066 53961 -22036
rect 53531 -22074 53950 -22066
rect 54140 -22078 54174 -21922
rect 54238 -22030 54272 -21922
rect 54336 -22078 54370 -21922
rect 54434 -22030 54468 -21922
rect 54532 -21933 54810 -21863
rect 52200 -22132 52929 -22087
rect 53328 -22089 53483 -22087
rect 53348 -22097 53483 -22089
rect 48314 -24163 49348 -24159
rect 48314 -24165 48863 -24163
rect 47901 -24193 47974 -24187
rect 49274 -24189 49348 -24163
rect 47222 -24203 47974 -24193
rect 47727 -24234 47974 -24203
rect 48809 -24221 48944 -24213
rect 48789 -24223 48944 -24221
rect 47727 -24251 47857 -24234
rect 47901 -24247 47974 -24234
rect 47754 -24301 47830 -24251
rect 48582 -24259 48944 -24223
rect 49461 -24232 50246 -24146
rect 48789 -24261 48944 -24259
rect 48809 -24267 48944 -24261
rect 48992 -24244 49411 -24236
rect 48992 -24274 49422 -24244
rect 48019 -24489 48053 -24281
rect 48215 -24489 48249 -24281
rect 48411 -24489 48445 -24281
rect 48992 -24618 49026 -24274
rect 49188 -24618 49222 -24274
rect 49361 -24423 49422 -24274
rect 49601 -24388 49635 -24232
rect 49699 -24388 49733 -24280
rect 49797 -24388 49831 -24232
rect 49895 -24388 49929 -24280
rect 49483 -24423 49556 -24417
rect 49361 -24436 49556 -24423
rect 49383 -24464 49556 -24436
rect 49483 -24477 49556 -24464
rect 49993 -24447 50365 -24377
rect 49601 -24619 49635 -24511
rect 49797 -24619 49831 -24511
rect 49993 -24619 50027 -24447
rect 47993 -25554 48027 -25210
rect 48189 -25554 48223 -25210
rect 48602 -25317 48636 -25209
rect 48798 -25317 48832 -25209
rect 48484 -25364 48557 -25351
rect 48384 -25392 48557 -25364
rect 48362 -25405 48557 -25392
rect 48362 -25554 48423 -25405
rect 48484 -25411 48557 -25405
rect 48994 -25381 49028 -25209
rect 47993 -25584 48423 -25554
rect 47993 -25592 48412 -25584
rect 48602 -25596 48636 -25440
rect 48700 -25548 48734 -25440
rect 48798 -25596 48832 -25440
rect 48896 -25548 48930 -25440
rect 48994 -25451 49272 -25381
rect 46895 -25722 47180 -25679
rect 46616 -25825 46721 -25753
rect 47137 -25928 47180 -25722
rect 44649 -26076 45099 -26058
rect 44207 -26119 45099 -26076
rect 44207 -26137 44656 -26119
rect 45038 -26414 45099 -26119
rect 45772 -26296 45806 -26002
rect 45864 -26018 45909 -25948
rect 46256 -25968 47180 -25928
rect 46304 -25971 47180 -25968
rect 45765 -26414 45812 -26296
rect 45870 -26310 45904 -26018
rect 45968 -26295 46002 -26002
rect 46210 -26285 46244 -26002
rect 46304 -26011 46348 -25971
rect 45961 -26414 46008 -26295
rect 46203 -26414 46250 -26285
rect 46308 -26310 46342 -26011
rect 45038 -26527 46515 -26414
rect 47637 -25665 47864 -25663
rect 48275 -25665 48349 -25639
rect 47637 -25703 48349 -25665
rect 48462 -25682 49077 -25596
rect 47863 -25704 48349 -25703
rect 47863 -25705 47934 -25704
rect 48275 -25710 48349 -25704
rect 47895 -26055 47929 -25747
rect 47993 -26055 48027 -25747
rect 48091 -26055 48125 -25747
rect 48189 -26055 48223 -25747
rect 48287 -26055 48321 -25747
rect 47992 -26107 48027 -26055
rect 48706 -26089 48767 -25682
rect 49196 -25846 49266 -25451
rect 49440 -25705 49474 -25121
rect 49647 -25087 49887 -25053
rect 49647 -25129 49689 -25087
rect 49436 -25764 49478 -25705
rect 49651 -25711 49685 -25129
rect 49749 -25709 49783 -25121
rect 49845 -25131 49887 -25087
rect 49648 -25764 49690 -25711
rect 49436 -25800 49690 -25764
rect 49745 -25763 49787 -25709
rect 49847 -25729 49881 -25131
rect 50059 -25715 50093 -25121
rect 49745 -25802 49886 -25763
rect 49843 -25814 49886 -25802
rect 49601 -25846 49756 -25836
rect 49196 -25882 49756 -25846
rect 49196 -25884 49266 -25882
rect 49601 -25891 49756 -25882
rect 49843 -25869 50024 -25814
rect 49843 -25939 49886 -25869
rect 49331 -25953 49486 -25944
rect 49294 -25987 49486 -25953
rect 49331 -25999 49486 -25987
rect 49532 -25979 49886 -25939
rect 50058 -25959 50101 -25715
rect 50295 -25784 50365 -24447
rect 50284 -25856 50389 -25784
rect 50814 -25959 51028 -25844
rect 48317 -26107 48767 -26089
rect 47875 -26150 48767 -26107
rect 47875 -26168 48324 -26150
rect 48706 -26445 48767 -26150
rect 49440 -26327 49474 -26033
rect 49532 -26049 49577 -25979
rect 49924 -25999 51126 -25959
rect 49972 -26002 51126 -25999
rect 49433 -26445 49480 -26327
rect 49538 -26341 49572 -26049
rect 49636 -26326 49670 -26033
rect 49878 -26316 49912 -26033
rect 49972 -26042 50016 -26002
rect 49629 -26445 49676 -26326
rect 49871 -26445 49918 -26316
rect 49976 -26341 50010 -26042
rect 50814 -26064 51028 -26002
rect 48706 -26558 50183 -26445
rect 42827 -27678 43079 -27539
rect 41611 -28129 41851 -28120
rect 52200 -27500 52346 -22132
rect 53175 -22147 53402 -22145
rect 53813 -22147 53887 -22121
rect 53175 -22185 53887 -22147
rect 54000 -22164 54615 -22078
rect 53186 -23056 53262 -22185
rect 53401 -22186 53887 -22185
rect 53401 -22187 53472 -22186
rect 53813 -22192 53887 -22186
rect 53433 -22537 53467 -22229
rect 53531 -22537 53565 -22229
rect 53629 -22537 53663 -22229
rect 53727 -22537 53761 -22229
rect 53825 -22537 53859 -22229
rect 53530 -22589 53565 -22537
rect 54244 -22571 54305 -22164
rect 54734 -22328 54804 -21933
rect 54978 -22187 55012 -21603
rect 55185 -21569 55425 -21535
rect 55185 -21611 55227 -21569
rect 54974 -22246 55016 -22187
rect 55189 -22193 55223 -21611
rect 55287 -22191 55321 -21603
rect 55383 -21613 55425 -21569
rect 55186 -22246 55228 -22193
rect 54974 -22282 55228 -22246
rect 55283 -22245 55325 -22191
rect 55385 -22211 55419 -21613
rect 55597 -22197 55631 -21603
rect 55283 -22284 55424 -22245
rect 55381 -22296 55424 -22284
rect 55139 -22328 55294 -22318
rect 54734 -22364 55294 -22328
rect 54734 -22366 54804 -22364
rect 55139 -22373 55294 -22364
rect 55381 -22351 55562 -22296
rect 55381 -22421 55424 -22351
rect 54869 -22435 55024 -22426
rect 54832 -22469 55024 -22435
rect 54869 -22481 55024 -22469
rect 55070 -22461 55424 -22421
rect 55596 -22441 55639 -22197
rect 55833 -22266 55903 -20929
rect 62311 -20905 62345 -20697
rect 62507 -20905 62541 -20697
rect 62703 -20905 62737 -20697
rect 63284 -21034 63318 -20690
rect 63480 -21034 63514 -20690
rect 63653 -20839 63714 -20690
rect 63893 -20804 63927 -20648
rect 63991 -20804 64025 -20696
rect 64089 -20804 64123 -20648
rect 71172 -20650 71302 -20633
rect 71346 -20646 71419 -20633
rect 72027 -20658 72389 -20622
rect 72906 -20631 73691 -20545
rect 80536 -20554 80666 -20462
rect 80828 -20520 80862 -20264
rect 80926 -20520 80960 -20312
rect 81024 -20520 81058 -20264
rect 81122 -20486 81156 -20312
rect 81703 -20442 81737 -20134
rect 81801 -20442 81835 -20134
rect 81899 -20442 81933 -20134
rect 81997 -20442 82031 -20134
rect 82095 -20442 82129 -20134
rect 81671 -20485 81742 -20484
rect 82083 -20485 82157 -20479
rect 81671 -20486 82157 -20485
rect 81122 -20520 82157 -20486
rect 82514 -20507 82575 -20100
rect 81123 -20524 82157 -20520
rect 81123 -20526 81672 -20524
rect 80710 -20554 80783 -20548
rect 82083 -20550 82157 -20524
rect 80536 -20595 80783 -20554
rect 81618 -20582 81753 -20574
rect 81598 -20584 81753 -20582
rect 80536 -20612 80666 -20595
rect 80710 -20608 80783 -20595
rect 81391 -20620 81753 -20584
rect 82270 -20593 83055 -20507
rect 81598 -20622 81753 -20620
rect 81618 -20628 81753 -20622
rect 81801 -20605 82220 -20597
rect 72234 -20660 72389 -20658
rect 72254 -20666 72389 -20660
rect 72437 -20643 72856 -20635
rect 72437 -20673 72867 -20643
rect 64187 -20804 64221 -20696
rect 63775 -20839 63848 -20833
rect 63653 -20852 63848 -20839
rect 63675 -20880 63848 -20852
rect 63775 -20893 63848 -20880
rect 64285 -20863 64657 -20793
rect 63893 -21035 63927 -20927
rect 64089 -21035 64123 -20927
rect 64285 -21035 64319 -20863
rect 56970 -21961 57004 -21461
rect 57149 -21425 57470 -21391
rect 56969 -22007 57004 -21961
rect 57149 -22007 57189 -21425
rect 57238 -21465 57273 -21425
rect 57239 -21969 57273 -21465
rect 57337 -21962 57371 -21461
rect 57435 -21464 57470 -21425
rect 56969 -22047 57189 -22007
rect 57334 -22082 57372 -21962
rect 57435 -21969 57469 -21464
rect 57565 -22045 57599 -21461
rect 57891 -21975 57925 -21461
rect 58119 -21751 58153 -21461
rect 58118 -21844 58155 -21751
rect 58118 -21881 58255 -21844
rect 57891 -22009 58050 -21975
rect 57714 -22045 57852 -22034
rect 56970 -22120 57372 -22082
rect 57439 -22079 57852 -22045
rect 56733 -22131 56871 -22121
rect 56343 -22165 56871 -22131
rect 55822 -22338 55927 -22266
rect 56343 -22441 56386 -22165
rect 56733 -22175 56871 -22165
rect 56789 -22266 56927 -22257
rect 56579 -22300 56927 -22266
rect 56579 -22427 56651 -22300
rect 56789 -22311 56927 -22300
rect 56579 -22436 56663 -22427
rect 53855 -22589 54305 -22571
rect 53413 -22632 54305 -22589
rect 53413 -22650 53862 -22632
rect 54244 -22927 54305 -22632
rect 54978 -22809 55012 -22515
rect 55070 -22531 55115 -22461
rect 55462 -22481 56386 -22441
rect 55510 -22484 56386 -22481
rect 54971 -22927 55018 -22809
rect 55076 -22823 55110 -22531
rect 55174 -22808 55208 -22515
rect 55416 -22798 55450 -22515
rect 55510 -22524 55554 -22484
rect 56584 -22506 56663 -22436
rect 55167 -22927 55214 -22808
rect 55409 -22927 55456 -22798
rect 55514 -22823 55548 -22524
rect 56872 -22748 56906 -22457
rect 56870 -22859 56907 -22748
rect 56970 -22765 57004 -22120
rect 57199 -22190 57237 -22120
rect 57439 -22158 57473 -22079
rect 57714 -22088 57852 -22079
rect 57189 -22328 57243 -22190
rect 57342 -22192 57473 -22158
rect 57539 -22175 57677 -22121
rect 57924 -22190 57978 -22052
rect 58016 -22053 58050 -22009
rect 58016 -22107 58182 -22053
rect 57342 -22765 57376 -22192
rect 58016 -22222 58050 -22107
rect 58102 -22222 58156 -22205
rect 57440 -22261 57599 -22226
rect 58016 -22227 58156 -22222
rect 57988 -22256 58156 -22227
rect 57440 -22765 57474 -22261
rect 57565 -22765 57599 -22261
rect 57663 -22748 57697 -22257
rect 57793 -22747 57827 -22257
rect 56333 -22863 56944 -22859
rect 57662 -22863 57699 -22748
rect 57790 -22863 57827 -22747
rect 57891 -22765 57925 -22257
rect 57988 -22261 58050 -22256
rect 57989 -22765 58023 -22261
rect 58102 -22264 58156 -22256
rect 58217 -22374 58255 -21881
rect 58217 -22412 58509 -22374
rect 58119 -22746 58153 -22457
rect 58217 -22462 58255 -22412
rect 58117 -22863 58154 -22746
rect 58217 -22765 58251 -22462
rect 56333 -22927 58267 -22863
rect 54244 -22972 58267 -22927
rect 54244 -23040 56446 -22972
rect 56794 -23024 58267 -22972
rect 52475 -23217 53262 -23056
rect 52475 -27138 52636 -23217
rect 53186 -23313 53262 -23217
rect 58471 -23307 58509 -22412
rect 53186 -23389 56496 -23313
rect 53186 -23571 53262 -23389
rect 53186 -23647 53328 -23571
rect 53252 -24036 53328 -23647
rect 54261 -23613 54926 -23585
rect 54261 -23671 55296 -23613
rect 54261 -23752 54347 -23671
rect 54521 -23708 54556 -23671
rect 54846 -23674 55296 -23671
rect 53409 -23838 54347 -23752
rect 53252 -24128 53387 -24036
rect 53549 -24094 53583 -23838
rect 53647 -24094 53681 -23886
rect 53745 -24094 53779 -23838
rect 53843 -24060 53877 -23886
rect 54424 -24016 54458 -23708
rect 54522 -24016 54556 -23708
rect 54620 -24016 54654 -23708
rect 54718 -24016 54752 -23708
rect 54816 -24016 54850 -23708
rect 54392 -24059 54463 -24058
rect 54804 -24059 54878 -24053
rect 54392 -24060 54878 -24059
rect 53843 -24094 54878 -24060
rect 55235 -24081 55296 -23674
rect 53844 -24098 54878 -24094
rect 53844 -24100 54393 -24098
rect 53431 -24128 53504 -24122
rect 54804 -24124 54878 -24098
rect 53252 -24145 53504 -24128
rect 53257 -24169 53504 -24145
rect 54339 -24156 54474 -24148
rect 54319 -24158 54474 -24156
rect 53257 -24186 53387 -24169
rect 53431 -24182 53504 -24169
rect 54112 -24194 54474 -24158
rect 54991 -24167 55776 -24081
rect 54319 -24196 54474 -24194
rect 54339 -24202 54474 -24196
rect 54522 -24179 54941 -24171
rect 54522 -24209 54952 -24179
rect 53549 -24424 53583 -24216
rect 53745 -24424 53779 -24216
rect 53941 -24424 53975 -24216
rect 54522 -24553 54556 -24209
rect 54718 -24553 54752 -24209
rect 54891 -24358 54952 -24209
rect 55131 -24323 55165 -24167
rect 55229 -24323 55263 -24215
rect 55327 -24323 55361 -24167
rect 55425 -24323 55459 -24215
rect 55013 -24358 55086 -24352
rect 54891 -24371 55086 -24358
rect 54913 -24399 55086 -24371
rect 55013 -24412 55086 -24399
rect 55523 -24382 55895 -24312
rect 55131 -24554 55165 -24446
rect 55327 -24554 55361 -24446
rect 55523 -24554 55557 -24382
rect 53523 -25489 53557 -25145
rect 53719 -25489 53753 -25145
rect 54132 -25252 54166 -25144
rect 54328 -25252 54362 -25144
rect 54014 -25299 54087 -25286
rect 53914 -25327 54087 -25299
rect 53892 -25340 54087 -25327
rect 53892 -25489 53953 -25340
rect 54014 -25346 54087 -25340
rect 54524 -25316 54558 -25144
rect 53523 -25519 53953 -25489
rect 53523 -25527 53942 -25519
rect 54132 -25531 54166 -25375
rect 54230 -25483 54264 -25375
rect 54328 -25531 54362 -25375
rect 54426 -25483 54460 -25375
rect 54524 -25386 54802 -25316
rect 53167 -25600 53394 -25598
rect 53805 -25600 53879 -25574
rect 53167 -25638 53879 -25600
rect 53992 -25617 54607 -25531
rect 53393 -25639 53879 -25638
rect 53393 -25640 53464 -25639
rect 53805 -25645 53879 -25639
rect 53425 -25990 53459 -25682
rect 53523 -25990 53557 -25682
rect 53621 -25990 53655 -25682
rect 53719 -25990 53753 -25682
rect 53817 -25990 53851 -25682
rect 53522 -26042 53557 -25990
rect 54236 -26024 54297 -25617
rect 54726 -25781 54796 -25386
rect 54970 -25640 55004 -25056
rect 55177 -25022 55417 -24988
rect 55177 -25064 55219 -25022
rect 54966 -25699 55008 -25640
rect 55181 -25646 55215 -25064
rect 55279 -25644 55313 -25056
rect 55375 -25066 55417 -25022
rect 55178 -25699 55220 -25646
rect 54966 -25735 55220 -25699
rect 55275 -25698 55317 -25644
rect 55377 -25664 55411 -25066
rect 55589 -25650 55623 -25056
rect 55275 -25737 55416 -25698
rect 55373 -25749 55416 -25737
rect 55131 -25781 55286 -25771
rect 54726 -25817 55286 -25781
rect 54726 -25819 54796 -25817
rect 55131 -25826 55286 -25817
rect 55373 -25804 55554 -25749
rect 55373 -25874 55416 -25804
rect 54861 -25888 55016 -25879
rect 54824 -25922 55016 -25888
rect 54861 -25934 55016 -25922
rect 55062 -25914 55416 -25874
rect 55588 -25894 55631 -25650
rect 55825 -25719 55895 -24382
rect 56070 -23670 56162 -23585
rect 56093 -25645 56136 -23670
rect 56420 -24093 56496 -23389
rect 56722 -23345 58509 -23307
rect 56722 -23723 56760 -23345
rect 57929 -23644 58594 -23616
rect 57929 -23702 58964 -23644
rect 56699 -23777 56772 -23723
rect 57929 -23783 58015 -23702
rect 58189 -23739 58224 -23702
rect 58514 -23705 58964 -23702
rect 57077 -23869 58015 -23783
rect 56925 -24093 57055 -24067
rect 56420 -24159 57055 -24093
rect 57217 -24125 57251 -23869
rect 57315 -24125 57349 -23917
rect 57413 -24125 57447 -23869
rect 57511 -24091 57545 -23917
rect 58092 -24047 58126 -23739
rect 58190 -24047 58224 -23739
rect 58288 -24047 58322 -23739
rect 58386 -24047 58420 -23739
rect 58484 -24047 58518 -23739
rect 58060 -24090 58131 -24089
rect 58472 -24090 58546 -24084
rect 58060 -24091 58546 -24090
rect 57511 -24125 58546 -24091
rect 58903 -24112 58964 -23705
rect 60727 -21985 61653 -21861
rect 62285 -21970 62319 -21626
rect 62481 -21970 62515 -21626
rect 62894 -21733 62928 -21625
rect 63090 -21733 63124 -21625
rect 62776 -21780 62849 -21767
rect 62676 -21808 62849 -21780
rect 62654 -21821 62849 -21808
rect 62654 -21970 62715 -21821
rect 62776 -21827 62849 -21821
rect 63286 -21797 63320 -21625
rect 62102 -21983 62237 -21977
rect 62082 -21985 62237 -21983
rect 60727 -22021 62237 -21985
rect 62285 -22000 62715 -21970
rect 62285 -22008 62704 -22000
rect 62894 -22012 62928 -21856
rect 62992 -21964 63026 -21856
rect 63090 -22012 63124 -21856
rect 63188 -21964 63222 -21856
rect 63286 -21867 63564 -21797
rect 60727 -22100 61653 -22021
rect 62082 -22023 62237 -22021
rect 62102 -22031 62237 -22023
rect 61929 -22081 62156 -22079
rect 62567 -22081 62641 -22055
rect 57512 -24129 58546 -24125
rect 57512 -24131 58061 -24129
rect 57099 -24159 57172 -24153
rect 58472 -24155 58546 -24129
rect 56420 -24169 57172 -24159
rect 56925 -24200 57172 -24169
rect 58007 -24187 58142 -24179
rect 57987 -24189 58142 -24187
rect 56925 -24217 57055 -24200
rect 57099 -24213 57172 -24200
rect 56952 -24267 57028 -24217
rect 57780 -24225 58142 -24189
rect 58659 -24198 59444 -24112
rect 57987 -24227 58142 -24225
rect 58007 -24233 58142 -24227
rect 58190 -24210 58609 -24202
rect 58190 -24240 58620 -24210
rect 57217 -24455 57251 -24247
rect 57413 -24455 57447 -24247
rect 57609 -24455 57643 -24247
rect 58190 -24584 58224 -24240
rect 58386 -24584 58420 -24240
rect 58559 -24389 58620 -24240
rect 58799 -24354 58833 -24198
rect 58897 -24354 58931 -24246
rect 58995 -24354 59029 -24198
rect 59093 -24354 59127 -24246
rect 58681 -24389 58754 -24383
rect 58559 -24402 58754 -24389
rect 58581 -24430 58754 -24402
rect 58681 -24443 58754 -24430
rect 59191 -24413 59563 -24343
rect 58799 -24585 58833 -24477
rect 58995 -24585 59029 -24477
rect 59191 -24585 59225 -24413
rect 57191 -25520 57225 -25176
rect 57387 -25520 57421 -25176
rect 57800 -25283 57834 -25175
rect 57996 -25283 58030 -25175
rect 57682 -25330 57755 -25317
rect 57582 -25358 57755 -25330
rect 57560 -25371 57755 -25358
rect 57560 -25520 57621 -25371
rect 57682 -25377 57755 -25371
rect 58192 -25347 58226 -25175
rect 57191 -25550 57621 -25520
rect 57191 -25558 57610 -25550
rect 57800 -25562 57834 -25406
rect 57898 -25514 57932 -25406
rect 57996 -25562 58030 -25406
rect 58094 -25514 58128 -25406
rect 58192 -25417 58470 -25347
rect 56093 -25688 56378 -25645
rect 55814 -25791 55919 -25719
rect 56335 -25894 56378 -25688
rect 53847 -26042 54297 -26024
rect 53405 -26085 54297 -26042
rect 53405 -26103 53854 -26085
rect 54236 -26380 54297 -26085
rect 54970 -26262 55004 -25968
rect 55062 -25984 55107 -25914
rect 55454 -25934 56378 -25894
rect 55502 -25937 56378 -25934
rect 54963 -26380 55010 -26262
rect 55068 -26276 55102 -25984
rect 55166 -26261 55200 -25968
rect 55408 -26251 55442 -25968
rect 55502 -25977 55546 -25937
rect 55159 -26380 55206 -26261
rect 55401 -26380 55448 -26251
rect 55506 -26276 55540 -25977
rect 54236 -26493 55713 -26380
rect 56835 -25631 57062 -25629
rect 57473 -25631 57547 -25605
rect 56835 -25669 57547 -25631
rect 57660 -25648 58275 -25562
rect 57061 -25670 57547 -25669
rect 57061 -25671 57132 -25670
rect 57473 -25676 57547 -25670
rect 57093 -26021 57127 -25713
rect 57191 -26021 57225 -25713
rect 57289 -26021 57323 -25713
rect 57387 -26021 57421 -25713
rect 57485 -26021 57519 -25713
rect 57190 -26073 57225 -26021
rect 57904 -26055 57965 -25648
rect 58394 -25812 58464 -25417
rect 58638 -25671 58672 -25087
rect 58845 -25053 59085 -25019
rect 58845 -25095 58887 -25053
rect 58634 -25730 58676 -25671
rect 58849 -25677 58883 -25095
rect 58947 -25675 58981 -25087
rect 59043 -25097 59085 -25053
rect 58846 -25730 58888 -25677
rect 58634 -25766 58888 -25730
rect 58943 -25729 58985 -25675
rect 59045 -25695 59079 -25097
rect 59257 -25681 59291 -25087
rect 58943 -25768 59084 -25729
rect 59041 -25780 59084 -25768
rect 58799 -25812 58954 -25802
rect 58394 -25848 58954 -25812
rect 58394 -25850 58464 -25848
rect 58799 -25857 58954 -25848
rect 59041 -25835 59222 -25780
rect 59041 -25905 59084 -25835
rect 58529 -25919 58684 -25910
rect 58492 -25953 58684 -25919
rect 58529 -25965 58684 -25953
rect 58730 -25945 59084 -25905
rect 59256 -25925 59299 -25681
rect 59493 -25750 59563 -24413
rect 59482 -25822 59587 -25750
rect 59940 -25925 60232 -25756
rect 57515 -26073 57965 -26055
rect 57073 -26116 57965 -26073
rect 57073 -26134 57522 -26116
rect 57904 -26411 57965 -26116
rect 58638 -26293 58672 -25999
rect 58730 -26015 58775 -25945
rect 59122 -25965 60324 -25925
rect 59170 -25968 60324 -25965
rect 58631 -26411 58678 -26293
rect 58736 -26307 58770 -26015
rect 58834 -26292 58868 -25999
rect 59076 -26282 59110 -25999
rect 59170 -26008 59214 -25968
rect 58827 -26411 58874 -26292
rect 59069 -26411 59116 -26282
rect 59174 -26307 59208 -26008
rect 59940 -26055 60232 -25968
rect 57904 -26524 59381 -26411
rect 52457 -27305 52651 -27138
rect 52166 -27705 52398 -27500
rect 60727 -27485 60966 -22100
rect 61929 -22119 62641 -22081
rect 62754 -22098 63369 -22012
rect 61940 -23083 62016 -22119
rect 62155 -22120 62641 -22119
rect 62155 -22121 62226 -22120
rect 62567 -22126 62641 -22120
rect 62187 -22471 62221 -22163
rect 62285 -22471 62319 -22163
rect 62383 -22471 62417 -22163
rect 62481 -22471 62515 -22163
rect 62579 -22471 62613 -22163
rect 62284 -22523 62319 -22471
rect 62998 -22505 63059 -22098
rect 63488 -22262 63558 -21867
rect 63732 -22121 63766 -21537
rect 63939 -21503 64179 -21469
rect 63939 -21545 63981 -21503
rect 63728 -22180 63770 -22121
rect 63943 -22127 63977 -21545
rect 64041 -22125 64075 -21537
rect 64137 -21547 64179 -21503
rect 63940 -22180 63982 -22127
rect 63728 -22216 63982 -22180
rect 64037 -22179 64079 -22125
rect 64139 -22145 64173 -21547
rect 64351 -22131 64385 -21537
rect 64037 -22218 64178 -22179
rect 64135 -22230 64178 -22218
rect 63893 -22262 64048 -22252
rect 63488 -22298 64048 -22262
rect 63488 -22300 63558 -22298
rect 63893 -22307 64048 -22298
rect 64135 -22285 64316 -22230
rect 64135 -22355 64178 -22285
rect 63623 -22369 63778 -22360
rect 63586 -22403 63778 -22369
rect 63623 -22415 63778 -22403
rect 63824 -22395 64178 -22355
rect 64350 -22375 64393 -22131
rect 64587 -22200 64657 -20863
rect 71464 -20888 71498 -20680
rect 71660 -20888 71694 -20680
rect 71856 -20888 71890 -20680
rect 72437 -21017 72471 -20673
rect 72633 -21017 72667 -20673
rect 72806 -20822 72867 -20673
rect 73046 -20787 73080 -20631
rect 73144 -20787 73178 -20679
rect 73242 -20787 73276 -20631
rect 81801 -20635 82231 -20605
rect 73340 -20787 73374 -20679
rect 72928 -20822 73001 -20816
rect 72806 -20835 73001 -20822
rect 72828 -20863 73001 -20835
rect 72928 -20876 73001 -20863
rect 73438 -20846 73810 -20776
rect 73046 -21018 73080 -20910
rect 73242 -21018 73276 -20910
rect 73438 -21018 73472 -20846
rect 65724 -21895 65758 -21395
rect 65903 -21359 66224 -21325
rect 65723 -21941 65758 -21895
rect 65903 -21941 65943 -21359
rect 65992 -21399 66027 -21359
rect 65993 -21903 66027 -21399
rect 66091 -21896 66125 -21395
rect 66189 -21398 66224 -21359
rect 65723 -21981 65943 -21941
rect 66088 -22016 66126 -21896
rect 66189 -21903 66223 -21398
rect 66319 -21979 66353 -21395
rect 66645 -21909 66679 -21395
rect 66873 -21685 66907 -21395
rect 66872 -21778 66909 -21685
rect 66872 -21815 67009 -21778
rect 66645 -21943 66804 -21909
rect 66468 -21979 66606 -21968
rect 65724 -22054 66126 -22016
rect 66193 -22013 66606 -21979
rect 65487 -22065 65625 -22055
rect 65097 -22099 65625 -22065
rect 64576 -22272 64681 -22200
rect 65097 -22375 65140 -22099
rect 65487 -22109 65625 -22099
rect 65543 -22200 65681 -22191
rect 65333 -22234 65681 -22200
rect 65333 -22361 65405 -22234
rect 65543 -22245 65681 -22234
rect 65333 -22370 65417 -22361
rect 62609 -22523 63059 -22505
rect 62167 -22566 63059 -22523
rect 62167 -22584 62616 -22566
rect 62998 -22861 63059 -22566
rect 63732 -22743 63766 -22449
rect 63824 -22465 63869 -22395
rect 64216 -22415 65140 -22375
rect 64264 -22418 65140 -22415
rect 63725 -22861 63772 -22743
rect 63830 -22757 63864 -22465
rect 63928 -22742 63962 -22449
rect 64170 -22732 64204 -22449
rect 64264 -22458 64308 -22418
rect 65338 -22440 65417 -22370
rect 63921 -22861 63968 -22742
rect 64163 -22861 64210 -22732
rect 64268 -22757 64302 -22458
rect 65626 -22682 65660 -22391
rect 65624 -22793 65661 -22682
rect 65724 -22699 65758 -22054
rect 65953 -22124 65991 -22054
rect 66193 -22092 66227 -22013
rect 66468 -22022 66606 -22013
rect 65943 -22262 65997 -22124
rect 66096 -22126 66227 -22092
rect 66293 -22109 66431 -22055
rect 66678 -22124 66732 -21986
rect 66770 -21987 66804 -21943
rect 66770 -22041 66936 -21987
rect 66096 -22699 66130 -22126
rect 66770 -22156 66804 -22041
rect 66856 -22156 66910 -22139
rect 66194 -22195 66353 -22160
rect 66770 -22161 66910 -22156
rect 66742 -22190 66910 -22161
rect 66194 -22699 66228 -22195
rect 66319 -22699 66353 -22195
rect 66417 -22682 66451 -22191
rect 66547 -22681 66581 -22191
rect 65087 -22797 65698 -22793
rect 66416 -22797 66453 -22682
rect 66544 -22797 66581 -22681
rect 66645 -22699 66679 -22191
rect 66742 -22195 66804 -22190
rect 66743 -22699 66777 -22195
rect 66856 -22198 66910 -22190
rect 66971 -22308 67009 -21815
rect 66971 -22346 67263 -22308
rect 66873 -22680 66907 -22391
rect 66971 -22396 67009 -22346
rect 66871 -22797 66908 -22680
rect 66971 -22699 67005 -22396
rect 65087 -22861 67021 -22797
rect 62998 -22906 67021 -22861
rect 62998 -22974 65200 -22906
rect 65548 -22958 67021 -22906
rect 61227 -23247 62016 -23083
rect 67225 -23241 67263 -22346
rect 61227 -23300 65250 -23247
rect 60665 -27717 61013 -27485
rect 61227 -27870 61444 -23300
rect 61940 -23323 65250 -23300
rect 61940 -23505 62016 -23323
rect 61940 -23581 62082 -23505
rect 62006 -23970 62082 -23581
rect 63015 -23547 63680 -23519
rect 63015 -23605 64050 -23547
rect 63015 -23686 63101 -23605
rect 63275 -23642 63310 -23605
rect 63600 -23608 64050 -23605
rect 62163 -23772 63101 -23686
rect 62006 -24062 62141 -23970
rect 62303 -24028 62337 -23772
rect 62401 -24028 62435 -23820
rect 62499 -24028 62533 -23772
rect 62597 -23994 62631 -23820
rect 63178 -23950 63212 -23642
rect 63276 -23950 63310 -23642
rect 63374 -23950 63408 -23642
rect 63472 -23950 63506 -23642
rect 63570 -23950 63604 -23642
rect 63146 -23993 63217 -23992
rect 63558 -23993 63632 -23987
rect 63146 -23994 63632 -23993
rect 62597 -24028 63632 -23994
rect 63989 -24015 64050 -23608
rect 62598 -24032 63632 -24028
rect 62598 -24034 63147 -24032
rect 62185 -24062 62258 -24056
rect 63558 -24058 63632 -24032
rect 62006 -24079 62258 -24062
rect 62011 -24103 62258 -24079
rect 63093 -24090 63228 -24082
rect 63073 -24092 63228 -24090
rect 62011 -24120 62141 -24103
rect 62185 -24116 62258 -24103
rect 62866 -24128 63228 -24092
rect 63745 -24101 64530 -24015
rect 63073 -24130 63228 -24128
rect 63093 -24136 63228 -24130
rect 63276 -24113 63695 -24105
rect 63276 -24143 63706 -24113
rect 62303 -24358 62337 -24150
rect 62499 -24358 62533 -24150
rect 62695 -24358 62729 -24150
rect 63276 -24487 63310 -24143
rect 63472 -24487 63506 -24143
rect 63645 -24292 63706 -24143
rect 63885 -24257 63919 -24101
rect 63983 -24257 64017 -24149
rect 64081 -24257 64115 -24101
rect 64179 -24257 64213 -24149
rect 63767 -24292 63840 -24286
rect 63645 -24305 63840 -24292
rect 63667 -24333 63840 -24305
rect 63767 -24346 63840 -24333
rect 64277 -24316 64649 -24246
rect 63885 -24488 63919 -24380
rect 64081 -24488 64115 -24380
rect 64277 -24488 64311 -24316
rect 62277 -25423 62311 -25079
rect 62473 -25423 62507 -25079
rect 62886 -25186 62920 -25078
rect 63082 -25186 63116 -25078
rect 62768 -25233 62841 -25220
rect 62668 -25261 62841 -25233
rect 62646 -25274 62841 -25261
rect 62646 -25423 62707 -25274
rect 62768 -25280 62841 -25274
rect 63278 -25250 63312 -25078
rect 62277 -25453 62707 -25423
rect 62277 -25461 62696 -25453
rect 62886 -25465 62920 -25309
rect 62984 -25417 63018 -25309
rect 63082 -25465 63116 -25309
rect 63180 -25417 63214 -25309
rect 63278 -25320 63556 -25250
rect 61921 -25534 62148 -25532
rect 62559 -25534 62633 -25508
rect 61921 -25572 62633 -25534
rect 62746 -25551 63361 -25465
rect 62147 -25573 62633 -25572
rect 62147 -25574 62218 -25573
rect 62559 -25579 62633 -25573
rect 62179 -25924 62213 -25616
rect 62277 -25924 62311 -25616
rect 62375 -25924 62409 -25616
rect 62473 -25924 62507 -25616
rect 62571 -25924 62605 -25616
rect 62276 -25976 62311 -25924
rect 62990 -25958 63051 -25551
rect 63480 -25715 63550 -25320
rect 63724 -25574 63758 -24990
rect 63931 -24956 64171 -24922
rect 63931 -24998 63973 -24956
rect 63720 -25633 63762 -25574
rect 63935 -25580 63969 -24998
rect 64033 -25578 64067 -24990
rect 64129 -25000 64171 -24956
rect 63932 -25633 63974 -25580
rect 63720 -25669 63974 -25633
rect 64029 -25632 64071 -25578
rect 64131 -25598 64165 -25000
rect 64343 -25584 64377 -24990
rect 64029 -25671 64170 -25632
rect 64127 -25683 64170 -25671
rect 63885 -25715 64040 -25705
rect 63480 -25751 64040 -25715
rect 63480 -25753 63550 -25751
rect 63885 -25760 64040 -25751
rect 64127 -25738 64308 -25683
rect 64127 -25808 64170 -25738
rect 63615 -25822 63770 -25813
rect 63578 -25856 63770 -25822
rect 63615 -25868 63770 -25856
rect 63816 -25848 64170 -25808
rect 64342 -25828 64385 -25584
rect 64579 -25653 64649 -24316
rect 64824 -23604 64916 -23519
rect 64847 -25579 64890 -23604
rect 65174 -24027 65250 -23323
rect 65476 -23279 67263 -23241
rect 65476 -23657 65514 -23279
rect 66683 -23578 67348 -23550
rect 66683 -23636 67718 -23578
rect 65453 -23711 65526 -23657
rect 66683 -23717 66769 -23636
rect 66943 -23673 66978 -23636
rect 67268 -23639 67718 -23636
rect 65831 -23803 66769 -23717
rect 65679 -24027 65809 -24001
rect 65174 -24093 65809 -24027
rect 65971 -24059 66005 -23803
rect 66069 -24059 66103 -23851
rect 66167 -24059 66201 -23803
rect 66265 -24025 66299 -23851
rect 66846 -23981 66880 -23673
rect 66944 -23981 66978 -23673
rect 67042 -23981 67076 -23673
rect 67140 -23981 67174 -23673
rect 67238 -23981 67272 -23673
rect 66814 -24024 66885 -24023
rect 67226 -24024 67300 -24018
rect 66814 -24025 67300 -24024
rect 66265 -24059 67300 -24025
rect 67657 -24046 67718 -23639
rect 70055 -21968 70719 -21889
rect 71438 -21953 71472 -21609
rect 71634 -21953 71668 -21609
rect 72047 -21716 72081 -21608
rect 72243 -21716 72277 -21608
rect 71929 -21763 72002 -21750
rect 71829 -21791 72002 -21763
rect 71807 -21804 72002 -21791
rect 71807 -21953 71868 -21804
rect 71929 -21810 72002 -21804
rect 72439 -21780 72473 -21608
rect 71255 -21966 71390 -21960
rect 71235 -21968 71390 -21966
rect 70055 -22004 71390 -21968
rect 71438 -21983 71868 -21953
rect 71438 -21991 71857 -21983
rect 72047 -21995 72081 -21839
rect 72145 -21947 72179 -21839
rect 72243 -21995 72277 -21839
rect 72341 -21947 72375 -21839
rect 72439 -21850 72717 -21780
rect 70055 -22074 70719 -22004
rect 71235 -22006 71390 -22004
rect 71255 -22014 71390 -22006
rect 71082 -22064 71309 -22062
rect 71720 -22064 71794 -22038
rect 66266 -24063 67300 -24059
rect 66266 -24065 66815 -24063
rect 65853 -24093 65926 -24087
rect 67226 -24089 67300 -24063
rect 65174 -24103 65926 -24093
rect 65679 -24134 65926 -24103
rect 66761 -24121 66896 -24113
rect 66741 -24123 66896 -24121
rect 65679 -24151 65809 -24134
rect 65853 -24147 65926 -24134
rect 65706 -24201 65782 -24151
rect 66534 -24159 66896 -24123
rect 67413 -24132 68198 -24046
rect 66741 -24161 66896 -24159
rect 66761 -24167 66896 -24161
rect 66944 -24144 67363 -24136
rect 66944 -24174 67374 -24144
rect 65971 -24389 66005 -24181
rect 66167 -24389 66201 -24181
rect 66363 -24389 66397 -24181
rect 66944 -24518 66978 -24174
rect 67140 -24518 67174 -24174
rect 67313 -24323 67374 -24174
rect 67553 -24288 67587 -24132
rect 67651 -24288 67685 -24180
rect 67749 -24288 67783 -24132
rect 67847 -24288 67881 -24180
rect 67435 -24323 67508 -24317
rect 67313 -24336 67508 -24323
rect 67335 -24364 67508 -24336
rect 67435 -24377 67508 -24364
rect 67945 -24347 68317 -24277
rect 67553 -24519 67587 -24411
rect 67749 -24519 67783 -24411
rect 67945 -24519 67979 -24347
rect 65945 -25454 65979 -25110
rect 66141 -25454 66175 -25110
rect 66554 -25217 66588 -25109
rect 66750 -25217 66784 -25109
rect 66436 -25264 66509 -25251
rect 66336 -25292 66509 -25264
rect 66314 -25305 66509 -25292
rect 66314 -25454 66375 -25305
rect 66436 -25311 66509 -25305
rect 66946 -25281 66980 -25109
rect 65945 -25484 66375 -25454
rect 65945 -25492 66364 -25484
rect 66554 -25496 66588 -25340
rect 66652 -25448 66686 -25340
rect 66750 -25496 66784 -25340
rect 66848 -25448 66882 -25340
rect 66946 -25351 67224 -25281
rect 64847 -25622 65132 -25579
rect 64568 -25725 64673 -25653
rect 65089 -25828 65132 -25622
rect 62601 -25976 63051 -25958
rect 62159 -26019 63051 -25976
rect 62159 -26037 62608 -26019
rect 62990 -26314 63051 -26019
rect 63724 -26196 63758 -25902
rect 63816 -25918 63861 -25848
rect 64208 -25868 65132 -25828
rect 64256 -25871 65132 -25868
rect 63717 -26314 63764 -26196
rect 63822 -26210 63856 -25918
rect 63920 -26195 63954 -25902
rect 64162 -26185 64196 -25902
rect 64256 -25911 64300 -25871
rect 63913 -26314 63960 -26195
rect 64155 -26314 64202 -26185
rect 64260 -26210 64294 -25911
rect 62990 -26427 64467 -26314
rect 65589 -25565 65816 -25563
rect 66227 -25565 66301 -25539
rect 65589 -25603 66301 -25565
rect 66414 -25582 67029 -25496
rect 65815 -25604 66301 -25603
rect 65815 -25605 65886 -25604
rect 66227 -25610 66301 -25604
rect 65847 -25955 65881 -25647
rect 65945 -25955 65979 -25647
rect 66043 -25955 66077 -25647
rect 66141 -25955 66175 -25647
rect 66239 -25955 66273 -25647
rect 65944 -26007 65979 -25955
rect 66658 -25989 66719 -25582
rect 67148 -25746 67218 -25351
rect 67392 -25605 67426 -25021
rect 67599 -24987 67839 -24953
rect 67599 -25029 67641 -24987
rect 67388 -25664 67430 -25605
rect 67603 -25611 67637 -25029
rect 67701 -25609 67735 -25021
rect 67797 -25031 67839 -24987
rect 67600 -25664 67642 -25611
rect 67388 -25700 67642 -25664
rect 67697 -25663 67739 -25609
rect 67799 -25629 67833 -25031
rect 68011 -25615 68045 -25021
rect 67697 -25702 67838 -25663
rect 67795 -25714 67838 -25702
rect 67553 -25746 67708 -25736
rect 67148 -25782 67708 -25746
rect 67148 -25784 67218 -25782
rect 67553 -25791 67708 -25782
rect 67795 -25769 67976 -25714
rect 67795 -25839 67838 -25769
rect 67283 -25853 67438 -25844
rect 67246 -25887 67438 -25853
rect 67283 -25899 67438 -25887
rect 67484 -25879 67838 -25839
rect 68010 -25859 68053 -25615
rect 68247 -25684 68317 -24347
rect 68236 -25756 68341 -25684
rect 68705 -25859 68966 -25698
rect 66269 -26007 66719 -25989
rect 65827 -26050 66719 -26007
rect 65827 -26068 66276 -26050
rect 66658 -26345 66719 -26050
rect 67392 -26227 67426 -25933
rect 67484 -25949 67529 -25879
rect 67876 -25899 69078 -25859
rect 67924 -25902 69078 -25899
rect 67385 -26345 67432 -26227
rect 67490 -26241 67524 -25949
rect 67588 -26226 67622 -25933
rect 67830 -26216 67864 -25933
rect 67924 -25942 67968 -25902
rect 67581 -26345 67628 -26226
rect 67823 -26345 67870 -26216
rect 67928 -26241 67962 -25942
rect 68705 -26002 68966 -25902
rect 66658 -26458 68135 -26345
rect 61170 -28153 61514 -27870
rect 70055 -27482 70240 -22074
rect 71082 -22102 71794 -22064
rect 71907 -22081 72522 -21995
rect 71093 -23124 71169 -22102
rect 71308 -22103 71794 -22102
rect 71308 -22104 71379 -22103
rect 71720 -22109 71794 -22103
rect 71340 -22454 71374 -22146
rect 71438 -22454 71472 -22146
rect 71536 -22454 71570 -22146
rect 71634 -22454 71668 -22146
rect 71732 -22454 71766 -22146
rect 71437 -22506 71472 -22454
rect 72151 -22488 72212 -22081
rect 72641 -22245 72711 -21850
rect 72885 -22104 72919 -21520
rect 73092 -21486 73332 -21452
rect 73092 -21528 73134 -21486
rect 72881 -22163 72923 -22104
rect 73096 -22110 73130 -21528
rect 73194 -22108 73228 -21520
rect 73290 -21530 73332 -21486
rect 73093 -22163 73135 -22110
rect 72881 -22199 73135 -22163
rect 73190 -22162 73232 -22108
rect 73292 -22128 73326 -21530
rect 73504 -22114 73538 -21520
rect 73190 -22201 73331 -22162
rect 73288 -22213 73331 -22201
rect 73046 -22245 73201 -22235
rect 72641 -22281 73201 -22245
rect 72641 -22283 72711 -22281
rect 73046 -22290 73201 -22281
rect 73288 -22268 73469 -22213
rect 73288 -22338 73331 -22268
rect 72776 -22352 72931 -22343
rect 72739 -22386 72931 -22352
rect 72776 -22398 72931 -22386
rect 72977 -22378 73331 -22338
rect 73503 -22358 73546 -22114
rect 73740 -22183 73810 -20846
rect 80828 -20850 80862 -20642
rect 81024 -20850 81058 -20642
rect 81220 -20850 81254 -20642
rect 81801 -20979 81835 -20635
rect 81997 -20979 82031 -20635
rect 82170 -20784 82231 -20635
rect 82410 -20749 82444 -20593
rect 82508 -20749 82542 -20641
rect 82606 -20749 82640 -20593
rect 82704 -20749 82738 -20641
rect 82292 -20784 82365 -20778
rect 82170 -20797 82365 -20784
rect 82192 -20825 82365 -20797
rect 82292 -20838 82365 -20825
rect 82802 -20808 83174 -20738
rect 82410 -20980 82444 -20872
rect 82606 -20980 82640 -20872
rect 82802 -20980 82836 -20808
rect 74877 -21878 74911 -21378
rect 75056 -21342 75377 -21308
rect 74876 -21924 74911 -21878
rect 75056 -21924 75096 -21342
rect 75145 -21382 75180 -21342
rect 75146 -21886 75180 -21382
rect 75244 -21879 75278 -21378
rect 75342 -21381 75377 -21342
rect 74876 -21964 75096 -21924
rect 75241 -21999 75279 -21879
rect 75342 -21886 75376 -21381
rect 75472 -21962 75506 -21378
rect 75798 -21892 75832 -21378
rect 76026 -21668 76060 -21378
rect 76025 -21761 76062 -21668
rect 76025 -21798 76162 -21761
rect 75798 -21926 75957 -21892
rect 75621 -21962 75759 -21951
rect 74877 -22037 75279 -21999
rect 75346 -21996 75759 -21962
rect 74640 -22048 74778 -22038
rect 74250 -22082 74778 -22048
rect 73729 -22255 73834 -22183
rect 74250 -22358 74293 -22082
rect 74640 -22092 74778 -22082
rect 74696 -22183 74834 -22174
rect 74486 -22217 74834 -22183
rect 74486 -22344 74558 -22217
rect 74696 -22228 74834 -22217
rect 74486 -22353 74570 -22344
rect 71762 -22506 72212 -22488
rect 71320 -22549 72212 -22506
rect 71320 -22567 71769 -22549
rect 72151 -22844 72212 -22549
rect 72885 -22726 72919 -22432
rect 72977 -22448 73022 -22378
rect 73369 -22398 74293 -22358
rect 73417 -22401 74293 -22398
rect 72878 -22844 72925 -22726
rect 72983 -22740 73017 -22448
rect 73081 -22725 73115 -22432
rect 73323 -22715 73357 -22432
rect 73417 -22441 73461 -22401
rect 74491 -22423 74570 -22353
rect 73074 -22844 73121 -22725
rect 73316 -22844 73363 -22715
rect 73421 -22740 73455 -22441
rect 74779 -22665 74813 -22374
rect 74777 -22776 74814 -22665
rect 74877 -22682 74911 -22037
rect 75106 -22107 75144 -22037
rect 75346 -22075 75380 -21996
rect 75621 -22005 75759 -21996
rect 75096 -22245 75150 -22107
rect 75249 -22109 75380 -22075
rect 75446 -22092 75584 -22038
rect 75831 -22107 75885 -21969
rect 75923 -21970 75957 -21926
rect 75923 -22024 76089 -21970
rect 75249 -22682 75283 -22109
rect 75923 -22139 75957 -22024
rect 76009 -22139 76063 -22122
rect 75347 -22178 75506 -22143
rect 75923 -22144 76063 -22139
rect 75895 -22173 76063 -22144
rect 75347 -22682 75381 -22178
rect 75472 -22682 75506 -22178
rect 75570 -22665 75604 -22174
rect 75700 -22664 75734 -22174
rect 74240 -22780 74851 -22776
rect 75569 -22780 75606 -22665
rect 75697 -22780 75734 -22664
rect 75798 -22682 75832 -22174
rect 75895 -22178 75957 -22173
rect 75896 -22682 75930 -22178
rect 76009 -22181 76063 -22173
rect 76124 -22291 76162 -21798
rect 76124 -22329 76416 -22291
rect 76026 -22663 76060 -22374
rect 76124 -22379 76162 -22329
rect 76024 -22780 76061 -22663
rect 76124 -22682 76158 -22379
rect 74240 -22844 76174 -22780
rect 72151 -22889 76174 -22844
rect 72151 -22957 74353 -22889
rect 74701 -22941 76174 -22889
rect 70418 -23230 71169 -23124
rect 76378 -23224 76416 -22329
rect 70418 -23294 74403 -23230
rect 70418 -27130 70588 -23294
rect 71093 -23306 74403 -23294
rect 71093 -23488 71169 -23306
rect 71093 -23564 71235 -23488
rect 71159 -23953 71235 -23564
rect 72168 -23530 72833 -23502
rect 72168 -23588 73203 -23530
rect 72168 -23669 72254 -23588
rect 72428 -23625 72463 -23588
rect 72753 -23591 73203 -23588
rect 71316 -23755 72254 -23669
rect 71159 -24045 71294 -23953
rect 71456 -24011 71490 -23755
rect 71554 -24011 71588 -23803
rect 71652 -24011 71686 -23755
rect 71750 -23977 71784 -23803
rect 72331 -23933 72365 -23625
rect 72429 -23933 72463 -23625
rect 72527 -23933 72561 -23625
rect 72625 -23933 72659 -23625
rect 72723 -23933 72757 -23625
rect 72299 -23976 72370 -23975
rect 72711 -23976 72785 -23970
rect 72299 -23977 72785 -23976
rect 71750 -24011 72785 -23977
rect 73142 -23998 73203 -23591
rect 71751 -24015 72785 -24011
rect 71751 -24017 72300 -24015
rect 71338 -24045 71411 -24039
rect 72711 -24041 72785 -24015
rect 71159 -24062 71411 -24045
rect 71164 -24086 71411 -24062
rect 72246 -24073 72381 -24065
rect 72226 -24075 72381 -24073
rect 71164 -24103 71294 -24086
rect 71338 -24099 71411 -24086
rect 72019 -24111 72381 -24075
rect 72898 -24084 73683 -23998
rect 72226 -24113 72381 -24111
rect 72246 -24119 72381 -24113
rect 72429 -24096 72848 -24088
rect 72429 -24126 72859 -24096
rect 71456 -24341 71490 -24133
rect 71652 -24341 71686 -24133
rect 71848 -24341 71882 -24133
rect 72429 -24470 72463 -24126
rect 72625 -24470 72659 -24126
rect 72798 -24275 72859 -24126
rect 73038 -24240 73072 -24084
rect 73136 -24240 73170 -24132
rect 73234 -24240 73268 -24084
rect 73332 -24240 73366 -24132
rect 72920 -24275 72993 -24269
rect 72798 -24288 72993 -24275
rect 72820 -24316 72993 -24288
rect 72920 -24329 72993 -24316
rect 73430 -24299 73802 -24229
rect 73038 -24471 73072 -24363
rect 73234 -24471 73268 -24363
rect 73430 -24471 73464 -24299
rect 71430 -25406 71464 -25062
rect 71626 -25406 71660 -25062
rect 72039 -25169 72073 -25061
rect 72235 -25169 72269 -25061
rect 71921 -25216 71994 -25203
rect 71821 -25244 71994 -25216
rect 71799 -25257 71994 -25244
rect 71799 -25406 71860 -25257
rect 71921 -25263 71994 -25257
rect 72431 -25233 72465 -25061
rect 71430 -25436 71860 -25406
rect 71430 -25444 71849 -25436
rect 72039 -25448 72073 -25292
rect 72137 -25400 72171 -25292
rect 72235 -25448 72269 -25292
rect 72333 -25400 72367 -25292
rect 72431 -25303 72709 -25233
rect 71074 -25517 71301 -25515
rect 71712 -25517 71786 -25491
rect 71074 -25555 71786 -25517
rect 71899 -25534 72514 -25448
rect 71300 -25556 71786 -25555
rect 71300 -25557 71371 -25556
rect 71712 -25562 71786 -25556
rect 71332 -25907 71366 -25599
rect 71430 -25907 71464 -25599
rect 71528 -25907 71562 -25599
rect 71626 -25907 71660 -25599
rect 71724 -25907 71758 -25599
rect 71429 -25959 71464 -25907
rect 72143 -25941 72204 -25534
rect 72633 -25698 72703 -25303
rect 72877 -25557 72911 -24973
rect 73084 -24939 73324 -24905
rect 73084 -24981 73126 -24939
rect 72873 -25616 72915 -25557
rect 73088 -25563 73122 -24981
rect 73186 -25561 73220 -24973
rect 73282 -24983 73324 -24939
rect 73085 -25616 73127 -25563
rect 72873 -25652 73127 -25616
rect 73182 -25615 73224 -25561
rect 73284 -25581 73318 -24983
rect 73496 -25567 73530 -24973
rect 73182 -25654 73323 -25615
rect 73280 -25666 73323 -25654
rect 73038 -25698 73193 -25688
rect 72633 -25734 73193 -25698
rect 72633 -25736 72703 -25734
rect 73038 -25743 73193 -25734
rect 73280 -25721 73461 -25666
rect 73280 -25791 73323 -25721
rect 72768 -25805 72923 -25796
rect 72731 -25839 72923 -25805
rect 72768 -25851 72923 -25839
rect 72969 -25831 73323 -25791
rect 73495 -25811 73538 -25567
rect 73732 -25636 73802 -24299
rect 73977 -23587 74069 -23502
rect 74000 -25562 74043 -23587
rect 74327 -24010 74403 -23306
rect 74629 -23262 76416 -23224
rect 74629 -23640 74667 -23262
rect 75836 -23561 76501 -23533
rect 75836 -23619 76871 -23561
rect 74606 -23694 74679 -23640
rect 75836 -23700 75922 -23619
rect 76096 -23656 76131 -23619
rect 76421 -23622 76871 -23619
rect 74984 -23786 75922 -23700
rect 74832 -24010 74962 -23984
rect 74327 -24076 74962 -24010
rect 75124 -24042 75158 -23786
rect 75222 -24042 75256 -23834
rect 75320 -24042 75354 -23786
rect 75418 -24008 75452 -23834
rect 75999 -23964 76033 -23656
rect 76097 -23964 76131 -23656
rect 76195 -23964 76229 -23656
rect 76293 -23964 76327 -23656
rect 76391 -23964 76425 -23656
rect 75967 -24007 76038 -24006
rect 76379 -24007 76453 -24001
rect 75967 -24008 76453 -24007
rect 75418 -24042 76453 -24008
rect 76810 -24029 76871 -23622
rect 78972 -21930 80180 -21747
rect 80802 -21915 80836 -21571
rect 80998 -21915 81032 -21571
rect 81411 -21678 81445 -21570
rect 81607 -21678 81641 -21570
rect 81293 -21725 81366 -21712
rect 81193 -21753 81366 -21725
rect 81171 -21766 81366 -21753
rect 81171 -21915 81232 -21766
rect 81293 -21772 81366 -21766
rect 81803 -21742 81837 -21570
rect 80619 -21928 80754 -21922
rect 80599 -21930 80754 -21928
rect 78972 -21966 80754 -21930
rect 80802 -21945 81232 -21915
rect 80802 -21953 81221 -21945
rect 81411 -21957 81445 -21801
rect 81509 -21909 81543 -21801
rect 81607 -21957 81641 -21801
rect 81705 -21909 81739 -21801
rect 81803 -21812 82081 -21742
rect 78972 -22041 80180 -21966
rect 80599 -21968 80754 -21966
rect 80619 -21976 80754 -21968
rect 80446 -22026 80673 -22024
rect 81084 -22026 81158 -22000
rect 75419 -24046 76453 -24042
rect 75419 -24048 75968 -24046
rect 75006 -24076 75079 -24070
rect 76379 -24072 76453 -24046
rect 74327 -24086 75079 -24076
rect 74832 -24117 75079 -24086
rect 75914 -24104 76049 -24096
rect 75894 -24106 76049 -24104
rect 74832 -24134 74962 -24117
rect 75006 -24130 75079 -24117
rect 74859 -24184 74935 -24134
rect 75687 -24142 76049 -24106
rect 76566 -24115 77351 -24029
rect 75894 -24144 76049 -24142
rect 75914 -24150 76049 -24144
rect 76097 -24127 76516 -24119
rect 76097 -24157 76527 -24127
rect 75124 -24372 75158 -24164
rect 75320 -24372 75354 -24164
rect 75516 -24372 75550 -24164
rect 76097 -24501 76131 -24157
rect 76293 -24501 76327 -24157
rect 76466 -24306 76527 -24157
rect 76706 -24271 76740 -24115
rect 76804 -24271 76838 -24163
rect 76902 -24271 76936 -24115
rect 77000 -24271 77034 -24163
rect 76588 -24306 76661 -24300
rect 76466 -24319 76661 -24306
rect 76488 -24347 76661 -24319
rect 76588 -24360 76661 -24347
rect 77098 -24330 77470 -24260
rect 76706 -24502 76740 -24394
rect 76902 -24502 76936 -24394
rect 77098 -24502 77132 -24330
rect 75098 -25437 75132 -25093
rect 75294 -25437 75328 -25093
rect 75707 -25200 75741 -25092
rect 75903 -25200 75937 -25092
rect 75589 -25247 75662 -25234
rect 75489 -25275 75662 -25247
rect 75467 -25288 75662 -25275
rect 75467 -25437 75528 -25288
rect 75589 -25294 75662 -25288
rect 76099 -25264 76133 -25092
rect 75098 -25467 75528 -25437
rect 75098 -25475 75517 -25467
rect 75707 -25479 75741 -25323
rect 75805 -25431 75839 -25323
rect 75903 -25479 75937 -25323
rect 76001 -25431 76035 -25323
rect 76099 -25334 76377 -25264
rect 74000 -25605 74285 -25562
rect 73721 -25708 73826 -25636
rect 74242 -25811 74285 -25605
rect 71754 -25959 72204 -25941
rect 71312 -26002 72204 -25959
rect 71312 -26020 71761 -26002
rect 72143 -26297 72204 -26002
rect 72877 -26179 72911 -25885
rect 72969 -25901 73014 -25831
rect 73361 -25851 74285 -25811
rect 73409 -25854 74285 -25851
rect 72870 -26297 72917 -26179
rect 72975 -26193 73009 -25901
rect 73073 -26178 73107 -25885
rect 73315 -26168 73349 -25885
rect 73409 -25894 73453 -25854
rect 73066 -26297 73113 -26178
rect 73308 -26297 73355 -26168
rect 73413 -26193 73447 -25894
rect 72143 -26410 73620 -26297
rect 74742 -25548 74969 -25546
rect 75380 -25548 75454 -25522
rect 74742 -25586 75454 -25548
rect 75567 -25565 76182 -25479
rect 74968 -25587 75454 -25586
rect 74968 -25588 75039 -25587
rect 75380 -25593 75454 -25587
rect 75000 -25938 75034 -25630
rect 75098 -25938 75132 -25630
rect 75196 -25938 75230 -25630
rect 75294 -25938 75328 -25630
rect 75392 -25938 75426 -25630
rect 75097 -25990 75132 -25938
rect 75811 -25972 75872 -25565
rect 76301 -25729 76371 -25334
rect 76545 -25588 76579 -25004
rect 76752 -24970 76992 -24936
rect 76752 -25012 76794 -24970
rect 76541 -25647 76583 -25588
rect 76756 -25594 76790 -25012
rect 76854 -25592 76888 -25004
rect 76950 -25014 76992 -24970
rect 76753 -25647 76795 -25594
rect 76541 -25683 76795 -25647
rect 76850 -25646 76892 -25592
rect 76952 -25612 76986 -25014
rect 77164 -25598 77198 -25004
rect 76850 -25685 76991 -25646
rect 76948 -25697 76991 -25685
rect 76706 -25729 76861 -25719
rect 76301 -25765 76861 -25729
rect 76301 -25767 76371 -25765
rect 76706 -25774 76861 -25765
rect 76948 -25752 77129 -25697
rect 76948 -25822 76991 -25752
rect 76436 -25836 76591 -25827
rect 76399 -25870 76591 -25836
rect 76436 -25882 76591 -25870
rect 76637 -25862 76991 -25822
rect 77163 -25842 77206 -25598
rect 77400 -25667 77470 -24330
rect 77389 -25739 77494 -25667
rect 77991 -25842 78093 -25804
rect 75422 -25990 75872 -25972
rect 74980 -26033 75872 -25990
rect 74980 -26051 75429 -26033
rect 75811 -26328 75872 -26033
rect 76545 -26210 76579 -25916
rect 76637 -25932 76682 -25862
rect 77029 -25882 78231 -25842
rect 77077 -25885 78231 -25882
rect 76538 -26328 76585 -26210
rect 76643 -26224 76677 -25932
rect 76741 -26209 76775 -25916
rect 76983 -26199 77017 -25916
rect 77077 -25925 77121 -25885
rect 77991 -25915 78093 -25885
rect 76734 -26328 76781 -26209
rect 76976 -26328 77023 -26199
rect 77081 -26224 77115 -25925
rect 75811 -26441 77288 -26328
rect 70379 -27310 70625 -27130
rect 69970 -27727 70352 -27482
rect 78972 -27485 79266 -22041
rect 80446 -22064 81158 -22026
rect 81271 -22043 81886 -21957
rect 80457 -23045 80533 -22064
rect 80672 -22065 81158 -22064
rect 80672 -22066 80743 -22065
rect 81084 -22071 81158 -22065
rect 80704 -22416 80738 -22108
rect 80802 -22416 80836 -22108
rect 80900 -22416 80934 -22108
rect 80998 -22416 81032 -22108
rect 81096 -22416 81130 -22108
rect 80801 -22468 80836 -22416
rect 81515 -22450 81576 -22043
rect 82005 -22207 82075 -21812
rect 82249 -22066 82283 -21482
rect 82456 -21448 82696 -21414
rect 82456 -21490 82498 -21448
rect 82245 -22125 82287 -22066
rect 82460 -22072 82494 -21490
rect 82558 -22070 82592 -21482
rect 82654 -21492 82696 -21448
rect 82457 -22125 82499 -22072
rect 82245 -22161 82499 -22125
rect 82554 -22124 82596 -22070
rect 82656 -22090 82690 -21492
rect 82868 -22076 82902 -21482
rect 82554 -22163 82695 -22124
rect 82652 -22175 82695 -22163
rect 82410 -22207 82565 -22197
rect 82005 -22243 82565 -22207
rect 82005 -22245 82075 -22243
rect 82410 -22252 82565 -22243
rect 82652 -22230 82833 -22175
rect 82652 -22300 82695 -22230
rect 82140 -22314 82295 -22305
rect 82103 -22348 82295 -22314
rect 82140 -22360 82295 -22348
rect 82341 -22340 82695 -22300
rect 82867 -22320 82910 -22076
rect 83104 -22145 83174 -20808
rect 84241 -21840 84275 -21340
rect 84420 -21304 84741 -21270
rect 84240 -21886 84275 -21840
rect 84420 -21886 84460 -21304
rect 84509 -21344 84544 -21304
rect 84510 -21848 84544 -21344
rect 84608 -21841 84642 -21340
rect 84706 -21343 84741 -21304
rect 84240 -21926 84460 -21886
rect 84605 -21961 84643 -21841
rect 84706 -21848 84740 -21343
rect 84836 -21924 84870 -21340
rect 85162 -21854 85196 -21340
rect 85390 -21630 85424 -21340
rect 85389 -21723 85426 -21630
rect 85389 -21760 85526 -21723
rect 85162 -21888 85321 -21854
rect 84985 -21924 85123 -21913
rect 84241 -21999 84643 -21961
rect 84710 -21958 85123 -21924
rect 84004 -22010 84142 -22000
rect 83614 -22044 84142 -22010
rect 83093 -22217 83198 -22145
rect 83614 -22320 83657 -22044
rect 84004 -22054 84142 -22044
rect 84060 -22145 84198 -22136
rect 83850 -22179 84198 -22145
rect 83850 -22306 83922 -22179
rect 84060 -22190 84198 -22179
rect 83850 -22315 83934 -22306
rect 81126 -22468 81576 -22450
rect 80684 -22511 81576 -22468
rect 80684 -22529 81133 -22511
rect 81515 -22806 81576 -22511
rect 82249 -22688 82283 -22394
rect 82341 -22410 82386 -22340
rect 82733 -22360 83657 -22320
rect 82781 -22363 83657 -22360
rect 82242 -22806 82289 -22688
rect 82347 -22702 82381 -22410
rect 82445 -22687 82479 -22394
rect 82687 -22677 82721 -22394
rect 82781 -22403 82825 -22363
rect 83855 -22385 83934 -22315
rect 82438 -22806 82485 -22687
rect 82680 -22806 82727 -22677
rect 82785 -22702 82819 -22403
rect 84143 -22627 84177 -22336
rect 84141 -22738 84178 -22627
rect 84241 -22644 84275 -21999
rect 84470 -22069 84508 -21999
rect 84710 -22037 84744 -21958
rect 84985 -21967 85123 -21958
rect 84460 -22207 84514 -22069
rect 84613 -22071 84744 -22037
rect 84810 -22054 84948 -22000
rect 85195 -22069 85249 -21931
rect 85287 -21932 85321 -21888
rect 85287 -21986 85453 -21932
rect 84613 -22644 84647 -22071
rect 85287 -22101 85321 -21986
rect 85373 -22101 85427 -22084
rect 84711 -22140 84870 -22105
rect 85287 -22106 85427 -22101
rect 85259 -22135 85427 -22106
rect 84711 -22644 84745 -22140
rect 84836 -22644 84870 -22140
rect 84934 -22627 84968 -22136
rect 85064 -22626 85098 -22136
rect 83604 -22742 84215 -22738
rect 84933 -22742 84970 -22627
rect 85061 -22742 85098 -22626
rect 85162 -22644 85196 -22136
rect 85259 -22140 85321 -22135
rect 85260 -22644 85294 -22140
rect 85373 -22143 85427 -22135
rect 85488 -22253 85526 -21760
rect 85488 -22291 85780 -22253
rect 85390 -22625 85424 -22336
rect 85488 -22341 85526 -22291
rect 85388 -22742 85425 -22625
rect 85488 -22644 85522 -22341
rect 83604 -22806 85538 -22742
rect 81515 -22851 85538 -22806
rect 81515 -22919 83717 -22851
rect 84065 -22903 85538 -22851
rect 79694 -23192 80575 -23045
rect 85742 -23186 85780 -22291
rect 79694 -23268 83767 -23192
rect 79694 -23271 80575 -23268
rect 78923 -27723 79323 -27485
rect 79694 -27873 79920 -23271
rect 80457 -23450 80533 -23271
rect 80457 -23526 80599 -23450
rect 80523 -23915 80599 -23526
rect 81532 -23492 82197 -23464
rect 81532 -23550 82567 -23492
rect 81532 -23631 81618 -23550
rect 81792 -23587 81827 -23550
rect 82117 -23553 82567 -23550
rect 80680 -23717 81618 -23631
rect 80523 -24007 80658 -23915
rect 80820 -23973 80854 -23717
rect 80918 -23973 80952 -23765
rect 81016 -23973 81050 -23717
rect 81114 -23939 81148 -23765
rect 81695 -23895 81729 -23587
rect 81793 -23895 81827 -23587
rect 81891 -23895 81925 -23587
rect 81989 -23895 82023 -23587
rect 82087 -23895 82121 -23587
rect 81663 -23938 81734 -23937
rect 82075 -23938 82149 -23932
rect 81663 -23939 82149 -23938
rect 81114 -23973 82149 -23939
rect 82506 -23960 82567 -23553
rect 81115 -23977 82149 -23973
rect 81115 -23979 81664 -23977
rect 80702 -24007 80775 -24001
rect 82075 -24003 82149 -23977
rect 80523 -24024 80775 -24007
rect 80528 -24048 80775 -24024
rect 81610 -24035 81745 -24027
rect 81590 -24037 81745 -24035
rect 80528 -24065 80658 -24048
rect 80702 -24061 80775 -24048
rect 81383 -24073 81745 -24037
rect 82262 -24046 83047 -23960
rect 81590 -24075 81745 -24073
rect 81610 -24081 81745 -24075
rect 81793 -24058 82212 -24050
rect 81793 -24088 82223 -24058
rect 80820 -24303 80854 -24095
rect 81016 -24303 81050 -24095
rect 81212 -24303 81246 -24095
rect 81793 -24432 81827 -24088
rect 81989 -24432 82023 -24088
rect 82162 -24237 82223 -24088
rect 82402 -24202 82436 -24046
rect 82500 -24202 82534 -24094
rect 82598 -24202 82632 -24046
rect 82696 -24202 82730 -24094
rect 82284 -24237 82357 -24231
rect 82162 -24250 82357 -24237
rect 82184 -24278 82357 -24250
rect 82284 -24291 82357 -24278
rect 82794 -24261 83166 -24191
rect 82402 -24433 82436 -24325
rect 82598 -24433 82632 -24325
rect 82794 -24433 82828 -24261
rect 80794 -25368 80828 -25024
rect 80990 -25368 81024 -25024
rect 81403 -25131 81437 -25023
rect 81599 -25131 81633 -25023
rect 81285 -25178 81358 -25165
rect 81185 -25206 81358 -25178
rect 81163 -25219 81358 -25206
rect 81163 -25368 81224 -25219
rect 81285 -25225 81358 -25219
rect 81795 -25195 81829 -25023
rect 80794 -25398 81224 -25368
rect 80794 -25406 81213 -25398
rect 81403 -25410 81437 -25254
rect 81501 -25362 81535 -25254
rect 81599 -25410 81633 -25254
rect 81697 -25362 81731 -25254
rect 81795 -25265 82073 -25195
rect 80438 -25479 80665 -25477
rect 81076 -25479 81150 -25453
rect 80438 -25517 81150 -25479
rect 81263 -25496 81878 -25410
rect 80664 -25518 81150 -25517
rect 80664 -25519 80735 -25518
rect 81076 -25524 81150 -25518
rect 80696 -25869 80730 -25561
rect 80794 -25869 80828 -25561
rect 80892 -25869 80926 -25561
rect 80990 -25869 81024 -25561
rect 81088 -25869 81122 -25561
rect 80793 -25921 80828 -25869
rect 81507 -25903 81568 -25496
rect 81997 -25660 82067 -25265
rect 82241 -25519 82275 -24935
rect 82448 -24901 82688 -24867
rect 82448 -24943 82490 -24901
rect 82237 -25578 82279 -25519
rect 82452 -25525 82486 -24943
rect 82550 -25523 82584 -24935
rect 82646 -24945 82688 -24901
rect 82449 -25578 82491 -25525
rect 82237 -25614 82491 -25578
rect 82546 -25577 82588 -25523
rect 82648 -25543 82682 -24945
rect 82860 -25529 82894 -24935
rect 82546 -25616 82687 -25577
rect 82644 -25628 82687 -25616
rect 82402 -25660 82557 -25650
rect 81997 -25696 82557 -25660
rect 81997 -25698 82067 -25696
rect 82402 -25705 82557 -25696
rect 82644 -25683 82825 -25628
rect 82644 -25753 82687 -25683
rect 82132 -25767 82287 -25758
rect 82095 -25801 82287 -25767
rect 82132 -25813 82287 -25801
rect 82333 -25793 82687 -25753
rect 82859 -25773 82902 -25529
rect 83096 -25598 83166 -24261
rect 83341 -23549 83433 -23464
rect 83364 -25524 83407 -23549
rect 83691 -23972 83767 -23268
rect 83993 -23224 85780 -23186
rect 83993 -23602 84031 -23224
rect 85200 -23523 85865 -23495
rect 85200 -23581 86235 -23523
rect 83970 -23656 84043 -23602
rect 85200 -23662 85286 -23581
rect 85460 -23618 85495 -23581
rect 85785 -23584 86235 -23581
rect 84348 -23748 85286 -23662
rect 84196 -23972 84326 -23946
rect 83691 -24038 84326 -23972
rect 84488 -24004 84522 -23748
rect 84586 -24004 84620 -23796
rect 84684 -24004 84718 -23748
rect 84782 -23970 84816 -23796
rect 85363 -23926 85397 -23618
rect 85461 -23926 85495 -23618
rect 85559 -23926 85593 -23618
rect 85657 -23926 85691 -23618
rect 85755 -23926 85789 -23618
rect 85331 -23969 85402 -23968
rect 85743 -23969 85817 -23963
rect 85331 -23970 85817 -23969
rect 84782 -24004 85817 -23970
rect 86174 -23991 86235 -23584
rect 84783 -24008 85817 -24004
rect 84783 -24010 85332 -24008
rect 84370 -24038 84443 -24032
rect 85743 -24034 85817 -24008
rect 83691 -24048 84443 -24038
rect 84196 -24079 84443 -24048
rect 85278 -24066 85413 -24058
rect 85258 -24068 85413 -24066
rect 84196 -24096 84326 -24079
rect 84370 -24092 84443 -24079
rect 84223 -24146 84299 -24096
rect 85051 -24104 85413 -24068
rect 85930 -24077 86715 -23991
rect 85258 -24106 85413 -24104
rect 85278 -24112 85413 -24106
rect 85461 -24089 85880 -24081
rect 85461 -24119 85891 -24089
rect 84488 -24334 84522 -24126
rect 84684 -24334 84718 -24126
rect 84880 -24334 84914 -24126
rect 85461 -24463 85495 -24119
rect 85657 -24463 85691 -24119
rect 85830 -24268 85891 -24119
rect 86070 -24233 86104 -24077
rect 86168 -24233 86202 -24125
rect 86266 -24233 86300 -24077
rect 86364 -24233 86398 -24125
rect 85952 -24268 86025 -24262
rect 85830 -24281 86025 -24268
rect 85852 -24309 86025 -24281
rect 85952 -24322 86025 -24309
rect 86462 -24292 86834 -24222
rect 86070 -24464 86104 -24356
rect 86266 -24464 86300 -24356
rect 86462 -24464 86496 -24292
rect 84462 -25399 84496 -25055
rect 84658 -25399 84692 -25055
rect 85071 -25162 85105 -25054
rect 85267 -25162 85301 -25054
rect 84953 -25209 85026 -25196
rect 84853 -25237 85026 -25209
rect 84831 -25250 85026 -25237
rect 84831 -25399 84892 -25250
rect 84953 -25256 85026 -25250
rect 85463 -25226 85497 -25054
rect 84462 -25429 84892 -25399
rect 84462 -25437 84881 -25429
rect 85071 -25441 85105 -25285
rect 85169 -25393 85203 -25285
rect 85267 -25441 85301 -25285
rect 85365 -25393 85399 -25285
rect 85463 -25296 85741 -25226
rect 83364 -25567 83649 -25524
rect 83085 -25670 83190 -25598
rect 83606 -25773 83649 -25567
rect 81118 -25921 81568 -25903
rect 80676 -25964 81568 -25921
rect 80676 -25982 81125 -25964
rect 81507 -26259 81568 -25964
rect 82241 -26141 82275 -25847
rect 82333 -25863 82378 -25793
rect 82725 -25813 83649 -25773
rect 82773 -25816 83649 -25813
rect 82234 -26259 82281 -26141
rect 82339 -26155 82373 -25863
rect 82437 -26140 82471 -25847
rect 82679 -26130 82713 -25847
rect 82773 -25856 82817 -25816
rect 82430 -26259 82477 -26140
rect 82672 -26259 82719 -26130
rect 82777 -26155 82811 -25856
rect 81507 -26372 82984 -26259
rect 84106 -25510 84333 -25508
rect 84744 -25510 84818 -25484
rect 84106 -25548 84818 -25510
rect 84931 -25527 85546 -25441
rect 84332 -25549 84818 -25548
rect 84332 -25550 84403 -25549
rect 84744 -25555 84818 -25549
rect 84364 -25900 84398 -25592
rect 84462 -25900 84496 -25592
rect 84560 -25900 84594 -25592
rect 84658 -25900 84692 -25592
rect 84756 -25900 84790 -25592
rect 84461 -25952 84496 -25900
rect 85175 -25934 85236 -25527
rect 85665 -25691 85735 -25296
rect 85909 -25550 85943 -24966
rect 86116 -24932 86356 -24898
rect 86116 -24974 86158 -24932
rect 85905 -25609 85947 -25550
rect 86120 -25556 86154 -24974
rect 86218 -25554 86252 -24966
rect 86314 -24976 86356 -24932
rect 86117 -25609 86159 -25556
rect 85905 -25645 86159 -25609
rect 86214 -25608 86256 -25554
rect 86316 -25574 86350 -24976
rect 86528 -25560 86562 -24966
rect 86214 -25647 86355 -25608
rect 86312 -25659 86355 -25647
rect 86070 -25691 86225 -25681
rect 85665 -25727 86225 -25691
rect 85665 -25729 85735 -25727
rect 86070 -25736 86225 -25727
rect 86312 -25714 86493 -25659
rect 86312 -25784 86355 -25714
rect 85800 -25798 85955 -25789
rect 85763 -25832 85955 -25798
rect 85800 -25844 85955 -25832
rect 86001 -25824 86355 -25784
rect 86527 -25804 86570 -25560
rect 86764 -25629 86834 -24292
rect 86753 -25701 86858 -25629
rect 87382 -25804 87741 -25654
rect 84786 -25952 85236 -25934
rect 84344 -25995 85236 -25952
rect 84344 -26013 84793 -25995
rect 85175 -26290 85236 -25995
rect 85909 -26172 85943 -25878
rect 86001 -25894 86046 -25824
rect 86393 -25844 87741 -25804
rect 86441 -25847 87741 -25844
rect 85902 -26290 85949 -26172
rect 86007 -26186 86041 -25894
rect 86105 -26171 86139 -25878
rect 86347 -26161 86381 -25878
rect 86441 -25887 86485 -25847
rect 86098 -26290 86145 -26171
rect 86340 -26290 86387 -26161
rect 86445 -26186 86479 -25887
rect 87382 -25997 87741 -25847
rect 85175 -26403 86652 -26290
rect 79605 -28149 79992 -27873
rect -24201 -29799 -23988 -29767
rect -24757 -29935 10154 -29799
rect -24201 -29945 -23988 -29935
rect -8007 -30195 16937 -30059
rect -24757 -30432 10411 -30297
rect -27604 -37174 -27464 -37004
rect -27029 -37174 -26909 -34086
rect -26416 -34117 -26324 -34091
rect -26824 -34151 -26324 -34117
rect -26416 -34235 -26324 -34151
rect -26824 -34269 -26324 -34235
rect -26416 -34353 -26324 -34269
rect -26824 -34387 -26324 -34353
rect -26416 -34471 -26324 -34387
rect -26824 -34505 -26324 -34471
rect -26416 -34589 -26324 -34505
rect -26824 -34623 -26324 -34589
rect -26416 -34707 -26324 -34623
rect -26824 -34741 -26324 -34707
rect -26416 -34825 -26324 -34741
rect -26824 -34859 -26324 -34825
rect -26416 -34943 -26324 -34859
rect -26824 -34977 -26324 -34943
rect -26416 -35061 -26324 -34977
rect -26824 -35095 -26324 -35061
rect 8241 -34202 19509 -33869
rect -26416 -35179 -26324 -35095
rect -26824 -35213 -26324 -35179
rect -26416 -35297 -26324 -35213
rect -26824 -35331 -26324 -35297
rect -26416 -35415 -26324 -35331
rect -26824 -35449 -26324 -35415
rect -26416 -35533 -26324 -35449
rect -26824 -35567 -26324 -35533
rect -14343 -34988 -14309 -34984
rect -14349 -35241 -14303 -34988
rect -14147 -35176 -14113 -34984
rect -14153 -35241 -14107 -35176
rect -13951 -35176 -13917 -34984
rect -13727 -35070 -13670 -35006
rect -13870 -35119 -13670 -35070
rect -13957 -35241 -13911 -35176
rect -14349 -35249 -13911 -35241
rect -13870 -35249 -13824 -35119
rect -13727 -35170 -13670 -35119
rect -13506 -34988 -13472 -34984
rect -14553 -35286 -14385 -35256
rect -26416 -35651 -26324 -35567
rect -26824 -35685 -26324 -35651
rect -26416 -35769 -26324 -35685
rect -26824 -35803 -26324 -35769
rect -26416 -35887 -26324 -35803
rect -26824 -35921 -26324 -35887
rect -26416 -36005 -26324 -35921
rect -26824 -36039 -26324 -36005
rect -26416 -36123 -26324 -36039
rect -26824 -36157 -26324 -36123
rect -26416 -36241 -26324 -36157
rect -26824 -36275 -26324 -36241
rect -21942 -36015 -21908 -35771
rect -21746 -36015 -21712 -35771
rect -21550 -36015 -21516 -35771
rect -21942 -36052 -21387 -36015
rect -21424 -36190 -21387 -36052
rect -20982 -36190 -20847 -36180
rect -21424 -36227 -20847 -36190
rect -26416 -36359 -26324 -36275
rect -21424 -36281 -21387 -36227
rect -20982 -36234 -20847 -36227
rect -26824 -36393 -26324 -36359
rect -26416 -36477 -26324 -36393
rect -26824 -36511 -26324 -36477
rect -26416 -36595 -26324 -36511
rect -26824 -36629 -26324 -36595
rect -26416 -36713 -26324 -36629
rect -26824 -36747 -26324 -36713
rect -26416 -36831 -26324 -36747
rect -26824 -36865 -26324 -36831
rect -26416 -36949 -26324 -36865
rect -26824 -36983 -26324 -36949
rect -26416 -37067 -26324 -36983
rect -26824 -37101 -26324 -37067
rect -27604 -37351 -26909 -37174
rect -26416 -37185 -26324 -37101
rect -26824 -37219 -26324 -37185
rect -26416 -37303 -26324 -37219
rect -26824 -37337 -26324 -37303
rect -27604 -37685 -27464 -37351
rect -27029 -37657 -26909 -37351
rect -26416 -37421 -26324 -37337
rect -26824 -37455 -26324 -37421
rect -22040 -36315 -21597 -36281
rect -21424 -36315 -21191 -36281
rect -22040 -36686 -22006 -36315
rect -21844 -36316 -21597 -36315
rect -21942 -36875 -21908 -36378
rect -21844 -36686 -21810 -36316
rect -21632 -36379 -21597 -36316
rect -21730 -36678 -21696 -36379
rect -21730 -36782 -21695 -36678
rect -21632 -36687 -21598 -36379
rect -21534 -36676 -21500 -36379
rect -21534 -36782 -21499 -36676
rect -21421 -36687 -21387 -36315
rect -21730 -36785 -21499 -36782
rect -21323 -36785 -21289 -36379
rect -21225 -36687 -21191 -36315
rect -21730 -36819 -21289 -36785
rect -20910 -36786 -20876 -36479
rect -20812 -36687 -20778 -35771
rect -20356 -36252 -20219 -36235
rect -19943 -36237 -19909 -35893
rect -19747 -36237 -19713 -35893
rect -19334 -36000 -19300 -35892
rect -19138 -36000 -19104 -35892
rect -19452 -36047 -19379 -36034
rect -19552 -36075 -19379 -36047
rect -19574 -36088 -19379 -36075
rect -19574 -36237 -19513 -36088
rect -19452 -36094 -19379 -36088
rect -18942 -36064 -18908 -35892
rect -17594 -35928 -16117 -35815
rect -18942 -36065 -18538 -36064
rect -18942 -36123 -18474 -36065
rect -20126 -36250 -19991 -36244
rect -20146 -36252 -19991 -36250
rect -20356 -36288 -19991 -36252
rect -19943 -36267 -19513 -36237
rect -19943 -36275 -19524 -36267
rect -19334 -36279 -19300 -36123
rect -19236 -36231 -19202 -36123
rect -19138 -36279 -19104 -36123
rect -19040 -36231 -19006 -36123
rect -18942 -36134 -18538 -36123
rect -18425 -36223 -17976 -36205
rect -17594 -36223 -17533 -35928
rect -16867 -36046 -16820 -35928
rect -18901 -36279 -17533 -36223
rect -20356 -36293 -20219 -36288
rect -20146 -36290 -19991 -36288
rect -20126 -36298 -19991 -36290
rect -19474 -36284 -17533 -36279
rect -19474 -36365 -18840 -36284
rect -18308 -36318 -18273 -36284
rect -20041 -36738 -20007 -36430
rect -19943 -36738 -19909 -36430
rect -19845 -36738 -19811 -36430
rect -19747 -36738 -19713 -36430
rect -19649 -36738 -19615 -36430
rect -19944 -36786 -19909 -36738
rect -19230 -36772 -19169 -36365
rect -18901 -36367 -18840 -36365
rect -18405 -36626 -18371 -36318
rect -18307 -36626 -18273 -36318
rect -18209 -36626 -18175 -36318
rect -18111 -36626 -18077 -36318
rect -18013 -36626 -17979 -36318
rect -18437 -36669 -18366 -36668
rect -18025 -36669 -17951 -36663
rect -18437 -36670 -17951 -36669
rect -18663 -36708 -17951 -36670
rect -17594 -36691 -17533 -36284
rect -16860 -36340 -16826 -36046
rect -16762 -36324 -16728 -36032
rect -16671 -36047 -16624 -35928
rect -16969 -36386 -16814 -36374
rect -17006 -36420 -16814 -36386
rect -16969 -36429 -16814 -36420
rect -16768 -36394 -16723 -36324
rect -16664 -36340 -16630 -36047
rect -16429 -36057 -16382 -35928
rect -16422 -36340 -16388 -36057
rect -16324 -36331 -16290 -36032
rect -16328 -36371 -16284 -36331
rect -16328 -36374 -15188 -36371
rect -16768 -36434 -16414 -36394
rect -16376 -36414 -15188 -36374
rect -17104 -36491 -17034 -36489
rect -16699 -36491 -16544 -36482
rect -17104 -36527 -16544 -36491
rect -18663 -36710 -18436 -36708
rect -18025 -36734 -17951 -36708
rect -19619 -36786 -19169 -36772
rect -21095 -36875 -19139 -36786
rect -17838 -36777 -17223 -36691
rect -22674 -37099 -22613 -36921
rect -22040 -36938 -19139 -36875
rect -22040 -36940 -20766 -36938
rect -20386 -37099 -20333 -37003
rect -22674 -37135 -20333 -37099
rect -22674 -37137 -22613 -37135
rect -18307 -36789 -17888 -36781
rect -18307 -36819 -17877 -36789
rect -18307 -37163 -18273 -36819
rect -18111 -37163 -18077 -36819
rect -17938 -36968 -17877 -36819
rect -17698 -36933 -17664 -36777
rect -17600 -36933 -17566 -36825
rect -17502 -36933 -17468 -36777
rect -17404 -36933 -17370 -36825
rect -17104 -36922 -17034 -36527
rect -16699 -36537 -16544 -36527
rect -16457 -36504 -16414 -36434
rect -16457 -36559 -16276 -36504
rect -16457 -36571 -16414 -36559
rect -16864 -36609 -16610 -36573
rect -17816 -36968 -17743 -36962
rect -17938 -36981 -17743 -36968
rect -17916 -37009 -17743 -36981
rect -17816 -37022 -17743 -37009
rect -17306 -36992 -17028 -36922
rect -17698 -37164 -17664 -37056
rect -17502 -37164 -17468 -37056
rect -17306 -37164 -17272 -36992
rect -16864 -36668 -16822 -36609
rect -16860 -37252 -16826 -36668
rect -16652 -36662 -16610 -36609
rect -16555 -36610 -16414 -36571
rect -16649 -37244 -16615 -36662
rect -16555 -36664 -16513 -36610
rect -16653 -37286 -16611 -37244
rect -16551 -37252 -16517 -36664
rect -16453 -37242 -16419 -36644
rect -16242 -36658 -16199 -36414
rect -16016 -36589 -15911 -36517
rect -16455 -37286 -16413 -37242
rect -16653 -37320 -16413 -37286
rect -16241 -37252 -16207 -36658
rect -26416 -37539 -26324 -37455
rect -26824 -37573 -26324 -37539
rect -26416 -37657 -26352 -37573
rect -27029 -37685 -26352 -37657
rect -27604 -37691 -26352 -37685
rect -27604 -37862 -26909 -37691
rect -26416 -37721 -26352 -37691
rect -26318 -37769 -26162 -37697
rect -27604 -38300 -27464 -37862
rect -27029 -37893 -26909 -37862
rect -27029 -37927 -26416 -37893
rect -27029 -38129 -26909 -37927
rect -26250 -38043 -26216 -37769
rect -26250 -38077 -25608 -38043
rect -27029 -38163 -26416 -38129
rect -27029 -38300 -26909 -38163
rect -22415 -38161 -22355 -37962
rect -21885 -38146 -21851 -37802
rect -21689 -38146 -21655 -37802
rect -21276 -37909 -21242 -37801
rect -21080 -37909 -21046 -37801
rect -21394 -37956 -21321 -37943
rect -21494 -37984 -21321 -37956
rect -21516 -37997 -21321 -37984
rect -21516 -38146 -21455 -37997
rect -21394 -38003 -21321 -37997
rect -20884 -37973 -20850 -37801
rect -20112 -37951 -20078 -37707
rect -19916 -37951 -19882 -37707
rect -19720 -37951 -19686 -37707
rect -20287 -37962 -20152 -37954
rect -20647 -37973 -20152 -37962
rect -20884 -37997 -20152 -37973
rect -20112 -37988 -19557 -37951
rect -22068 -38159 -21933 -38153
rect -22088 -38161 -21933 -38159
rect -22415 -38197 -21933 -38161
rect -21885 -38176 -21455 -38146
rect -21885 -38184 -21466 -38176
rect -21276 -38188 -21242 -38032
rect -21178 -38140 -21144 -38032
rect -21080 -38188 -21046 -38032
rect -20982 -38140 -20948 -38032
rect -20884 -38043 -20606 -37997
rect -20306 -37999 -20152 -37997
rect -20287 -38008 -20152 -37999
rect -20402 -38045 -20344 -38037
rect -19951 -38045 -19816 -38036
rect -20428 -38083 -19816 -38045
rect -22415 -38199 -22355 -38197
rect -22088 -38199 -21933 -38197
rect -22068 -38207 -21933 -38199
rect -27604 -38365 -26909 -38300
rect -26016 -38313 -25608 -38279
rect -27604 -38399 -26416 -38365
rect -27604 -38477 -26909 -38399
rect -22541 -38257 -22014 -38255
rect -21603 -38257 -21529 -38231
rect -22541 -38295 -21529 -38257
rect -21416 -38274 -20801 -38188
rect -22541 -38400 -22501 -38295
rect -22015 -38296 -21529 -38295
rect -22015 -38297 -21944 -38296
rect -21603 -38302 -21529 -38296
rect -27604 -39092 -27464 -38477
rect -27029 -38601 -26909 -38477
rect -26016 -38549 -25608 -38515
rect -27029 -38635 -26416 -38601
rect -27029 -38837 -26909 -38635
rect -22558 -38637 -22498 -38400
rect -21983 -38647 -21949 -38339
rect -21885 -38647 -21851 -38339
rect -21787 -38647 -21753 -38339
rect -21689 -38647 -21655 -38339
rect -21591 -38647 -21557 -38339
rect -26016 -38785 -25608 -38751
rect -27029 -38871 -26416 -38837
rect -21886 -38699 -21851 -38647
rect -21172 -38681 -21111 -38274
rect -20713 -38402 -20655 -38265
rect -20499 -38268 -20441 -38168
rect -20402 -38174 -20344 -38083
rect -19951 -38090 -19816 -38083
rect -19763 -38127 -19628 -38114
rect -20304 -38161 -19628 -38127
rect -20304 -38268 -20270 -38161
rect -19763 -38168 -19628 -38161
rect -19594 -38126 -19557 -37988
rect -19152 -38126 -19017 -38116
rect -19594 -38163 -19017 -38126
rect -19594 -38217 -19557 -38163
rect -19152 -38170 -19017 -38163
rect -18982 -38188 -18948 -37707
rect -18281 -38092 -18247 -37884
rect -18085 -38092 -18051 -37884
rect -17889 -38092 -17855 -37884
rect -17308 -38099 -17274 -37755
rect -17112 -38099 -17078 -37755
rect -16699 -37862 -16665 -37754
rect -16503 -37862 -16469 -37754
rect -16817 -37909 -16744 -37896
rect -16917 -37937 -16744 -37909
rect -16939 -37950 -16744 -37937
rect -16939 -38099 -16878 -37950
rect -16817 -37956 -16744 -37950
rect -16307 -37926 -16273 -37754
rect -16005 -37926 -15935 -36589
rect -17491 -38112 -17356 -38106
rect -17511 -38114 -17356 -38112
rect -18573 -38139 -18443 -38122
rect -18399 -38139 -18326 -38126
rect -18573 -38180 -18326 -38139
rect -17718 -38150 -17356 -38114
rect -17308 -38129 -16878 -38099
rect -17308 -38137 -16889 -38129
rect -16699 -38141 -16665 -37985
rect -16601 -38093 -16567 -37985
rect -16503 -38141 -16469 -37985
rect -16405 -38093 -16371 -37985
rect -16307 -37996 -15935 -37926
rect -17511 -38152 -17356 -38150
rect -17491 -38160 -17356 -38152
rect -18573 -38188 -18443 -38180
rect -18399 -38186 -18326 -38180
rect -20499 -38302 -20270 -38268
rect -20210 -38251 -19767 -38217
rect -19594 -38251 -19361 -38217
rect -20499 -38305 -20441 -38302
rect -20210 -38622 -20176 -38251
rect -20014 -38252 -19767 -38251
rect -20537 -38681 -20422 -38680
rect -21561 -38699 -20392 -38681
rect -22003 -38760 -20392 -38699
rect -21562 -38796 -20392 -38760
rect -27029 -39073 -26909 -38871
rect -20537 -38814 -20392 -38796
rect -20112 -38811 -20078 -38314
rect -20014 -38622 -19980 -38252
rect -19802 -38315 -19767 -38252
rect -19900 -38614 -19866 -38315
rect -19900 -38718 -19865 -38614
rect -19802 -38623 -19768 -38315
rect -19704 -38612 -19670 -38315
rect -19704 -38718 -19669 -38612
rect -19591 -38623 -19557 -38251
rect -19900 -38721 -19669 -38718
rect -19493 -38721 -19459 -38315
rect -19395 -38623 -19361 -38251
rect -18982 -38222 -18443 -38188
rect -17986 -38210 -17437 -38208
rect -17026 -38210 -16952 -38184
rect -17986 -38214 -16952 -38210
rect -19900 -38755 -19459 -38721
rect -19080 -38784 -19046 -38415
rect -18982 -38623 -18948 -38222
rect -18573 -38272 -18443 -38222
rect -18281 -38470 -18247 -38214
rect -18183 -38422 -18149 -38214
rect -18085 -38470 -18051 -38214
rect -17987 -38248 -16952 -38214
rect -16839 -38227 -16054 -38141
rect -17987 -38422 -17953 -38248
rect -17438 -38249 -16952 -38248
rect -17438 -38250 -17367 -38249
rect -17026 -38255 -16952 -38249
rect -18421 -38556 -17483 -38470
rect -17569 -38637 -17483 -38556
rect -17406 -38600 -17372 -38292
rect -17308 -38600 -17274 -38292
rect -17210 -38600 -17176 -38292
rect -17112 -38600 -17078 -38292
rect -17014 -38600 -16980 -38292
rect -17309 -38637 -17274 -38600
rect -16595 -38634 -16534 -38227
rect -16984 -38637 -16534 -38634
rect -17569 -38695 -16534 -38637
rect -17569 -38723 -16904 -38695
rect -17533 -38784 -17323 -38723
rect -19281 -38811 -17323 -38784
rect -20210 -38814 -17323 -38811
rect -20537 -38893 -17323 -38814
rect -26016 -39021 -25608 -38987
rect -27029 -39092 -26416 -39073
rect -27604 -39107 -26416 -39092
rect -27604 -39269 -26909 -39107
rect -26016 -39257 -25608 -39223
rect -27604 -39973 -27464 -39269
rect -27029 -39309 -26909 -39269
rect -27029 -39343 -26416 -39309
rect -27029 -39545 -26909 -39343
rect -26016 -39493 -25608 -39459
rect -27029 -39579 -26416 -39545
rect -27029 -39781 -26909 -39579
rect -26284 -39657 -26128 -39585
rect -26824 -39697 -26416 -39663
rect -27029 -39815 -26416 -39781
rect -27029 -39973 -26909 -39815
rect -26824 -39933 -26416 -39899
rect -27604 -40017 -26909 -39973
rect -27604 -40051 -26416 -40017
rect -27604 -40150 -26909 -40051
rect -26236 -40061 -26202 -39657
rect -26016 -39729 -25608 -39695
rect -26236 -40095 -25608 -40061
rect -27604 -40795 -27464 -40150
rect -27029 -40253 -26909 -40150
rect -26824 -40169 -26416 -40135
rect -27029 -40287 -26416 -40253
rect -27029 -40489 -26909 -40287
rect -26016 -40331 -25608 -40297
rect -26824 -40405 -26416 -40371
rect -27029 -40523 -26416 -40489
rect -27029 -40725 -26909 -40523
rect -26824 -40641 -26416 -40607
rect -26297 -40618 -26157 -40516
rect -26016 -40567 -25608 -40533
rect -27029 -40759 -26416 -40725
rect -27029 -40795 -26909 -40759
rect -27604 -40961 -26909 -40795
rect -26824 -40877 -26416 -40843
rect -26239 -40961 -26205 -40618
rect -26016 -40803 -25608 -40769
rect -27604 -40972 -26416 -40961
rect -27604 -41184 -27464 -40972
rect -27029 -40995 -26416 -40972
rect -26239 -40995 -26082 -40961
rect -27029 -41197 -26909 -40995
rect -26824 -41113 -26416 -41079
rect -26352 -41194 -26175 -41118
rect -26116 -41135 -26082 -40995
rect -26116 -41169 -25608 -41135
rect -27029 -41231 -26416 -41197
rect -27029 -41273 -26909 -41231
rect -26296 -41401 -26235 -41194
rect -26388 -41420 -26202 -41401
rect -26016 -41405 -25608 -41371
rect -26388 -44174 -26195 -41420
rect -24450 -38939 -17323 -38893
rect -16401 -38773 -16133 -38723
rect -15371 -38773 -15188 -36414
rect -14560 -35330 -14385 -35286
rect -14349 -35287 -13824 -35249
rect -13512 -35241 -13466 -34988
rect -13310 -35176 -13276 -34984
rect -13316 -35241 -13270 -35176
rect -12896 -34965 -12268 -34931
rect -13114 -35176 -13080 -34984
rect -12896 -35010 -12860 -34965
rect -13120 -35241 -13074 -35176
rect -13512 -35249 -13074 -35241
rect -13019 -35225 -12945 -35057
rect -12895 -35084 -12861 -35010
rect -13019 -35249 -12946 -35225
rect -13716 -35267 -13548 -35256
rect -13751 -35268 -13548 -35267
rect -14560 -35702 -14512 -35330
rect -14441 -35523 -14407 -35364
rect -14349 -35380 -14303 -35287
rect -14343 -35472 -14309 -35380
rect -14245 -35523 -14211 -35364
rect -14153 -35380 -14107 -35287
rect -13957 -35319 -13824 -35287
rect -14147 -35472 -14113 -35380
rect -14049 -35523 -14015 -35364
rect -13957 -35380 -13911 -35319
rect -13788 -35330 -13548 -35268
rect -13512 -35287 -12946 -35249
rect -13951 -35472 -13917 -35380
rect -13788 -35474 -13728 -35330
rect -13604 -35523 -13570 -35364
rect -13512 -35380 -13466 -35287
rect -13506 -35472 -13472 -35380
rect -13408 -35523 -13374 -35364
rect -13316 -35380 -13270 -35287
rect -13120 -35319 -12946 -35287
rect -12901 -35231 -12854 -35084
rect -12797 -35091 -12763 -34999
rect -12700 -35020 -12658 -34965
rect -12798 -35143 -12762 -35091
rect -12699 -35107 -12665 -35020
rect -12601 -35089 -12567 -34999
rect -12506 -35021 -12464 -34965
rect -12601 -35107 -12564 -35089
rect -12503 -35107 -12469 -35021
rect -12405 -35089 -12371 -34999
rect -12310 -35016 -12268 -34965
rect -12600 -35143 -12564 -35107
rect -12406 -35143 -12370 -35089
rect -12307 -35107 -12273 -35016
rect -12209 -35099 -12175 -34999
rect -12212 -35143 -12170 -35099
rect -12798 -35177 -12170 -35143
rect -12901 -35305 -12729 -35231
rect -12345 -35284 -12170 -35177
rect -11643 -34988 -11609 -34984
rect -11649 -35241 -11603 -34988
rect -11447 -35176 -11413 -34984
rect -11453 -35241 -11407 -35176
rect -11251 -35176 -11217 -34984
rect -11027 -35058 -10970 -35006
rect -11175 -35120 -10970 -35058
rect -11257 -35241 -11211 -35176
rect -11649 -35249 -11211 -35241
rect -11175 -35249 -11113 -35120
rect -11027 -35170 -10970 -35120
rect -10806 -34988 -10772 -34984
rect -11853 -35263 -11685 -35256
rect -13310 -35472 -13276 -35380
rect -13212 -35523 -13178 -35364
rect -13120 -35380 -13074 -35319
rect -13114 -35472 -13080 -35380
rect -12901 -35440 -12854 -35305
rect -12345 -35344 -12079 -35284
rect -11875 -35323 -11685 -35263
rect -11853 -35330 -11685 -35323
rect -11649 -35287 -11113 -35249
rect -10812 -35241 -10766 -34988
rect -10610 -35176 -10576 -34984
rect -10616 -35241 -10570 -35176
rect -10196 -34965 -9568 -34931
rect -10414 -35176 -10380 -34984
rect -10196 -35010 -10160 -34965
rect -10420 -35241 -10374 -35176
rect -10812 -35249 -10374 -35241
rect -10319 -35225 -10245 -35057
rect -10195 -35084 -10161 -35010
rect -10319 -35249 -10246 -35225
rect -11016 -35267 -10848 -35256
rect -12801 -35378 -12170 -35344
rect -12801 -35419 -12760 -35378
rect -12895 -35510 -12861 -35440
rect -14450 -35591 -13079 -35523
rect -12900 -35568 -12856 -35510
rect -12797 -35522 -12763 -35419
rect -12699 -35499 -12665 -35414
rect -12603 -35427 -12562 -35378
rect -12704 -35568 -12660 -35499
rect -12601 -35522 -12567 -35427
rect -12503 -35499 -12469 -35414
rect -12409 -35427 -12368 -35378
rect -12212 -35385 -12170 -35378
rect -12508 -35568 -12464 -35499
rect -12405 -35522 -12371 -35427
rect -12307 -35510 -12273 -35414
rect -12212 -35428 -12171 -35385
rect -12311 -35568 -12267 -35510
rect -12209 -35522 -12175 -35428
rect -11741 -35523 -11707 -35364
rect -11649 -35380 -11603 -35287
rect -11643 -35472 -11609 -35380
rect -11545 -35523 -11511 -35364
rect -11453 -35380 -11407 -35287
rect -11257 -35319 -11113 -35287
rect -11447 -35472 -11413 -35380
rect -11349 -35523 -11315 -35364
rect -11257 -35380 -11211 -35319
rect -11076 -35330 -10848 -35267
rect -10812 -35287 -10246 -35249
rect -11251 -35472 -11217 -35380
rect -11076 -35489 -11016 -35330
rect -10904 -35523 -10870 -35364
rect -10812 -35380 -10766 -35287
rect -10806 -35472 -10772 -35380
rect -10708 -35523 -10674 -35364
rect -10616 -35380 -10570 -35287
rect -10420 -35319 -10246 -35287
rect -10201 -35231 -10154 -35084
rect -10097 -35091 -10063 -34999
rect -10000 -35020 -9958 -34965
rect -10098 -35143 -10062 -35091
rect -9999 -35107 -9965 -35020
rect -9901 -35089 -9867 -34999
rect -9806 -35021 -9764 -34965
rect -9901 -35107 -9864 -35089
rect -9803 -35107 -9769 -35021
rect -9705 -35089 -9671 -34999
rect -9610 -35016 -9568 -34965
rect -9900 -35143 -9864 -35107
rect -9706 -35143 -9670 -35089
rect -9607 -35107 -9573 -35016
rect -9509 -35099 -9475 -34999
rect -9512 -35143 -9470 -35099
rect -10098 -35177 -9470 -35143
rect -10201 -35305 -10029 -35231
rect -9645 -35286 -9470 -35177
rect -10610 -35472 -10576 -35380
rect -10512 -35523 -10478 -35364
rect -10420 -35380 -10374 -35319
rect -10414 -35472 -10380 -35380
rect -10201 -35440 -10154 -35305
rect -9645 -35344 -9395 -35286
rect -10101 -35346 -9395 -35344
rect -10101 -35378 -9470 -35346
rect -10101 -35419 -10060 -35378
rect -10195 -35510 -10161 -35440
rect -14202 -35631 -14091 -35591
rect -14213 -35639 -14076 -35631
rect -13391 -35639 -13280 -35591
rect -12900 -35602 -12267 -35568
rect -11750 -35525 -11216 -35523
rect -10913 -35525 -10379 -35523
rect -11750 -35591 -10379 -35525
rect -10200 -35568 -10156 -35510
rect -10097 -35522 -10063 -35419
rect -9999 -35499 -9965 -35414
rect -9903 -35427 -9862 -35378
rect -10004 -35568 -9960 -35499
rect -9901 -35522 -9867 -35427
rect -9803 -35499 -9769 -35414
rect -9709 -35427 -9668 -35378
rect -9512 -35385 -9470 -35378
rect -9808 -35568 -9764 -35499
rect -9705 -35522 -9671 -35427
rect -9607 -35510 -9573 -35414
rect -9512 -35428 -9471 -35385
rect -9611 -35568 -9567 -35510
rect -9509 -35522 -9475 -35428
rect -11593 -35637 -11482 -35591
rect -11410 -35593 -10890 -35591
rect -11616 -35639 -11479 -35637
rect -10715 -35639 -10604 -35591
rect -10200 -35602 -9567 -35568
rect -8177 -35588 -8143 -34994
rect -7971 -34960 -7731 -34926
rect -7971 -35004 -7929 -34960
rect -8978 -35639 -8846 -35637
rect -14230 -35678 -8845 -35639
rect -14213 -35691 -14076 -35678
rect -11616 -35697 -11479 -35678
rect -8978 -35697 -8846 -35678
rect -14561 -35839 -14501 -35702
rect -12051 -35731 -11914 -35720
rect -11105 -35731 -10973 -35721
rect -14230 -35770 -8500 -35731
rect -12051 -35780 -11914 -35770
rect -11105 -35781 -10973 -35770
rect -13824 -35817 -13692 -35809
rect -9301 -35817 -9169 -35807
rect -14560 -36197 -14512 -35839
rect -14230 -35856 -9169 -35817
rect -8539 -35832 -8500 -35770
rect -8185 -35832 -8142 -35588
rect -7965 -35602 -7931 -35004
rect -7867 -35582 -7833 -34994
rect -7773 -35002 -7731 -34960
rect -7871 -35636 -7829 -35582
rect -7769 -35584 -7735 -35002
rect -7970 -35675 -7829 -35636
rect -7774 -35637 -7732 -35584
rect -7558 -35578 -7524 -34994
rect -7562 -35637 -7520 -35578
rect -6747 -35086 -6019 -35052
rect -6747 -35398 -6713 -35086
rect -6649 -35434 -6615 -35190
rect -6551 -35398 -6517 -35086
rect -6431 -35155 -6089 -35121
rect -6431 -35398 -6397 -35155
rect -6333 -35434 -6299 -35190
rect -6235 -35398 -6201 -35155
rect -6858 -35468 -6184 -35434
rect -7774 -35673 -7520 -35637
rect -7970 -35687 -7927 -35675
rect -8108 -35742 -7927 -35687
rect -7970 -35812 -7927 -35742
rect -7840 -35719 -7685 -35709
rect -7300 -35719 -7168 -35648
rect -7840 -35755 -7168 -35719
rect -7840 -35764 -7685 -35755
rect -13824 -35869 -13692 -35856
rect -9301 -35867 -9169 -35856
rect -8543 -35872 -8008 -35832
rect -7970 -35852 -7616 -35812
rect -8543 -35875 -8056 -35872
rect -14442 -35971 -13908 -35903
rect -13511 -35926 -12878 -35892
rect -14441 -36114 -14407 -36022
rect -14447 -36175 -14401 -36114
rect -14343 -36130 -14309 -35971
rect -14245 -36114 -14211 -36022
rect -14477 -36197 -14401 -36175
rect -14560 -36207 -14401 -36197
rect -14251 -36207 -14205 -36114
rect -14147 -36130 -14113 -35971
rect -14049 -36114 -14015 -36022
rect -14055 -36207 -14009 -36114
rect -13951 -36130 -13917 -35971
rect -13603 -36066 -13569 -35972
rect -13511 -35984 -13467 -35926
rect -13607 -36109 -13566 -36066
rect -13505 -36080 -13471 -35984
rect -13407 -36067 -13373 -35972
rect -13314 -35995 -13270 -35926
rect -13608 -36116 -13566 -36109
rect -13410 -36116 -13369 -36067
rect -13309 -36080 -13275 -35995
rect -13211 -36067 -13177 -35972
rect -13118 -35995 -13074 -35926
rect -13216 -36116 -13175 -36067
rect -13113 -36080 -13079 -35995
rect -13015 -36075 -12981 -35972
rect -12922 -35984 -12878 -35926
rect -12699 -35971 -11208 -35903
rect -10811 -35926 -10178 -35892
rect -12917 -36054 -12883 -35984
rect -13018 -36116 -12977 -36075
rect -13608 -36150 -12977 -36116
rect -14560 -36234 -14009 -36207
rect -14559 -36236 -14009 -36234
rect -14477 -36245 -14009 -36236
rect -13973 -36179 -13805 -36164
rect -13608 -36179 -13433 -36150
rect -13973 -36232 -13433 -36179
rect -12924 -36189 -12877 -36054
rect -12698 -36114 -12664 -36022
rect -12704 -36175 -12658 -36114
rect -12600 -36130 -12566 -35971
rect -12502 -36114 -12468 -36022
rect -13973 -36238 -13805 -36232
rect -14447 -36253 -14009 -36245
rect -14447 -36318 -14401 -36253
rect -14441 -36510 -14407 -36318
rect -14251 -36318 -14205 -36253
rect -14245 -36510 -14211 -36318
rect -14055 -36506 -14009 -36253
rect -14049 -36510 -14015 -36506
rect -13608 -36317 -13433 -36232
rect -13049 -36263 -12877 -36189
rect -13608 -36351 -12980 -36317
rect -13608 -36395 -13566 -36351
rect -13603 -36495 -13569 -36395
rect -13505 -36478 -13471 -36387
rect -13408 -36405 -13372 -36351
rect -13214 -36387 -13178 -36351
rect -13510 -36529 -13468 -36478
rect -13407 -36495 -13373 -36405
rect -13309 -36473 -13275 -36387
rect -13214 -36405 -13177 -36387
rect -13314 -36529 -13272 -36473
rect -13211 -36495 -13177 -36405
rect -13113 -36474 -13079 -36387
rect -13016 -36403 -12980 -36351
rect -13120 -36529 -13078 -36474
rect -13015 -36495 -12981 -36403
rect -12924 -36410 -12877 -36263
rect -12832 -36207 -12658 -36175
rect -12508 -36207 -12462 -36114
rect -12404 -36130 -12370 -35971
rect -12306 -36114 -12272 -36022
rect -12312 -36207 -12266 -36114
rect -12208 -36130 -12174 -35971
rect -12832 -36245 -12266 -36207
rect -12230 -36169 -12062 -36164
rect -12002 -36169 -11942 -36096
rect -12230 -36227 -11942 -36169
rect -11887 -36186 -11827 -36071
rect -11741 -36114 -11707 -36022
rect -11747 -36175 -11701 -36114
rect -11643 -36130 -11609 -35971
rect -11545 -36114 -11511 -36022
rect -11777 -36186 -11701 -36175
rect -12230 -36238 -12062 -36227
rect -12002 -36228 -11942 -36227
rect -11892 -36207 -11701 -36186
rect -11551 -36207 -11505 -36114
rect -11447 -36130 -11413 -35971
rect -11349 -36114 -11315 -36022
rect -11355 -36207 -11309 -36114
rect -11251 -36130 -11217 -35971
rect -10906 -36066 -10860 -35944
rect -10811 -35984 -10767 -35926
rect -10907 -36076 -10860 -36066
rect -10907 -36109 -10866 -36076
rect -10805 -36080 -10771 -35984
rect -10707 -36067 -10673 -35972
rect -10614 -35995 -10570 -35926
rect -10908 -36116 -10866 -36109
rect -10710 -36116 -10669 -36067
rect -10609 -36080 -10575 -35995
rect -10511 -36067 -10477 -35972
rect -10418 -35995 -10374 -35926
rect -10516 -36116 -10475 -36067
rect -10413 -36080 -10379 -35995
rect -10315 -36075 -10281 -35972
rect -10222 -35984 -10178 -35926
rect -9999 -35971 -8583 -35903
rect -10217 -36054 -10183 -35984
rect -10318 -36116 -10277 -36075
rect -10908 -36150 -10277 -36116
rect -11892 -36231 -11309 -36207
rect -12832 -36269 -12759 -36245
rect -12917 -36484 -12883 -36410
rect -12833 -36437 -12759 -36269
rect -12704 -36253 -12266 -36245
rect -12704 -36318 -12658 -36253
rect -12918 -36529 -12882 -36484
rect -12698 -36510 -12664 -36318
rect -13510 -36563 -12882 -36529
rect -12508 -36318 -12462 -36253
rect -12502 -36510 -12468 -36318
rect -12312 -36506 -12266 -36253
rect -12306 -36510 -12272 -36506
rect -12108 -36365 -12051 -36324
rect -11892 -36365 -11847 -36231
rect -11777 -36245 -11309 -36231
rect -11273 -36172 -11105 -36164
rect -10908 -36172 -10733 -36150
rect -11273 -36229 -10733 -36172
rect -10224 -36189 -10177 -36054
rect -9998 -36114 -9964 -36022
rect -10004 -36175 -9958 -36114
rect -9900 -36130 -9866 -35971
rect -9802 -36114 -9768 -36022
rect -11273 -36238 -11105 -36229
rect -11747 -36253 -11309 -36245
rect -11747 -36318 -11701 -36253
rect -12108 -36410 -11847 -36365
rect -12108 -36488 -12051 -36410
rect -11741 -36510 -11707 -36318
rect -11551 -36318 -11505 -36253
rect -11545 -36510 -11511 -36318
rect -11355 -36506 -11309 -36253
rect -11349 -36510 -11315 -36506
rect -10908 -36317 -10733 -36229
rect -10349 -36263 -10177 -36189
rect -10908 -36351 -10280 -36317
rect -10908 -36395 -10866 -36351
rect -10903 -36495 -10869 -36395
rect -10805 -36478 -10771 -36387
rect -10708 -36405 -10672 -36351
rect -10514 -36387 -10478 -36351
rect -10810 -36529 -10768 -36478
rect -10707 -36495 -10673 -36405
rect -10609 -36473 -10575 -36387
rect -10514 -36405 -10477 -36387
rect -10614 -36529 -10572 -36473
rect -10511 -36495 -10477 -36405
rect -10413 -36474 -10379 -36387
rect -10316 -36403 -10280 -36351
rect -10420 -36529 -10378 -36474
rect -10315 -36495 -10281 -36403
rect -10224 -36410 -10177 -36263
rect -10132 -36207 -9958 -36175
rect -9808 -36207 -9762 -36114
rect -9704 -36130 -9670 -35971
rect -9606 -36114 -9572 -36022
rect -9612 -36207 -9566 -36114
rect -9508 -36130 -9474 -35971
rect -10132 -36245 -9566 -36207
rect -9530 -36169 -9362 -36164
rect -9530 -36181 -9327 -36169
rect -9270 -36181 -9210 -36095
rect -9116 -36114 -9082 -36022
rect -9122 -36175 -9076 -36114
rect -9018 -36130 -8984 -35971
rect -8920 -36114 -8886 -36022
rect -9152 -36181 -9076 -36175
rect -9530 -36207 -9076 -36181
rect -8926 -36207 -8880 -36114
rect -8822 -36130 -8788 -35971
rect -8724 -36114 -8690 -36022
rect -8730 -36207 -8684 -36114
rect -8626 -36130 -8592 -35971
rect -8539 -36164 -8500 -35875
rect -8100 -35915 -8056 -35875
rect -9530 -36223 -8684 -36207
rect -9530 -36227 -9327 -36223
rect -9270 -36227 -9210 -36223
rect -9530 -36238 -9362 -36227
rect -9152 -36245 -8684 -36223
rect -8648 -36238 -8480 -36164
rect -8094 -36214 -8060 -35915
rect -7996 -36189 -7962 -35906
rect -10132 -36269 -10059 -36245
rect -10217 -36484 -10183 -36410
rect -10133 -36437 -10059 -36269
rect -10004 -36253 -9566 -36245
rect -10004 -36318 -9958 -36253
rect -10218 -36529 -10182 -36484
rect -9998 -36510 -9964 -36318
rect -10810 -36563 -10182 -36529
rect -9808 -36318 -9762 -36253
rect -9802 -36510 -9768 -36318
rect -9612 -36506 -9566 -36253
rect -9122 -36253 -8684 -36245
rect -9606 -36510 -9572 -36506
rect -9122 -36318 -9076 -36253
rect -9408 -36488 -9351 -36324
rect -9116 -36510 -9082 -36318
rect -8926 -36318 -8880 -36253
rect -8920 -36510 -8886 -36318
rect -8730 -36506 -8684 -36253
rect -8724 -36510 -8690 -36506
rect -8426 -36319 -8148 -36318
rect -8002 -36319 -7955 -36189
rect -7754 -36199 -7720 -35906
rect -7661 -35922 -7616 -35852
rect -7570 -35826 -7415 -35817
rect -7570 -35860 -7008 -35826
rect -7570 -35872 -7415 -35860
rect -7760 -36319 -7713 -36199
rect -7656 -36214 -7622 -35922
rect -7558 -36200 -7524 -35906
rect -7564 -36319 -7517 -36200
rect -8426 -36401 -7435 -36319
rect -24450 -39008 -20422 -38939
rect -16401 -38956 -15188 -38773
rect -12605 -36904 -11128 -36791
rect -13436 -37199 -12987 -37181
rect -12605 -37199 -12544 -36904
rect -11878 -37022 -11831 -36904
rect -13436 -37242 -12544 -37199
rect -13319 -37294 -13284 -37242
rect -12994 -37260 -12544 -37242
rect -13416 -37602 -13382 -37294
rect -13318 -37602 -13284 -37294
rect -13220 -37602 -13186 -37294
rect -13122 -37602 -13088 -37294
rect -13024 -37602 -12990 -37294
rect -12605 -37667 -12544 -37260
rect -11871 -37316 -11837 -37022
rect -11773 -37300 -11739 -37008
rect -11682 -37023 -11635 -36904
rect -11980 -37362 -11825 -37350
rect -12017 -37396 -11825 -37362
rect -11980 -37405 -11825 -37396
rect -11779 -37370 -11734 -37300
rect -11675 -37316 -11641 -37023
rect -11440 -37033 -11393 -36904
rect -11433 -37316 -11399 -37033
rect -11335 -37307 -11301 -37008
rect -11339 -37347 -11295 -37307
rect -11339 -37350 -8259 -37347
rect -11779 -37410 -11425 -37370
rect -11387 -37390 -8259 -37350
rect -12115 -37467 -12045 -37465
rect -11710 -37467 -11555 -37458
rect -12115 -37503 -11555 -37467
rect -13961 -37744 -13775 -37687
rect -13501 -37742 -13366 -37734
rect -13521 -37744 -13366 -37742
rect -13961 -37780 -13366 -37744
rect -12849 -37753 -12234 -37667
rect -13961 -37841 -13775 -37780
rect -13521 -37782 -13366 -37780
rect -13501 -37788 -13366 -37782
rect -13318 -37765 -12899 -37757
rect -13318 -37795 -12888 -37765
rect -13318 -38139 -13284 -37795
rect -13122 -38139 -13088 -37795
rect -12949 -37944 -12888 -37795
rect -12709 -37909 -12675 -37753
rect -12611 -37909 -12577 -37801
rect -12513 -37909 -12479 -37753
rect -12415 -37909 -12381 -37801
rect -12115 -37898 -12045 -37503
rect -11710 -37513 -11555 -37503
rect -11468 -37480 -11425 -37410
rect -11468 -37535 -11287 -37480
rect -11468 -37547 -11425 -37535
rect -11875 -37585 -11621 -37549
rect -12827 -37944 -12754 -37938
rect -12949 -37957 -12754 -37944
rect -12927 -37985 -12754 -37957
rect -12827 -37998 -12754 -37985
rect -12317 -37968 -12039 -37898
rect -12709 -38140 -12675 -38032
rect -12513 -38140 -12479 -38032
rect -12317 -38140 -12283 -37968
rect -11875 -37644 -11833 -37585
rect -11871 -38228 -11837 -37644
rect -11663 -37638 -11621 -37585
rect -11566 -37586 -11425 -37547
rect -11660 -38220 -11626 -37638
rect -11566 -37640 -11524 -37586
rect -11664 -38262 -11622 -38220
rect -11562 -38228 -11528 -37640
rect -11464 -38218 -11430 -37620
rect -11253 -37634 -11210 -37390
rect -8435 -37469 -8259 -37390
rect -11027 -37565 -10922 -37493
rect -11466 -38262 -11424 -38218
rect -11664 -38296 -11424 -38262
rect -11252 -38228 -11218 -37634
rect -16401 -38988 -16133 -38956
rect -25977 -42872 -25639 -42789
rect -24450 -42872 -24335 -39008
rect -18787 -39330 -15249 -39124
rect -15457 -39332 -15249 -39330
rect -16396 -39590 -16128 -39543
rect -23799 -39776 -16128 -39590
rect -13292 -39068 -13258 -38860
rect -13096 -39068 -13062 -38860
rect -12900 -39068 -12866 -38860
rect -12319 -39075 -12285 -38731
rect -12123 -39075 -12089 -38731
rect -11710 -38838 -11676 -38730
rect -11514 -38838 -11480 -38730
rect -11828 -38885 -11755 -38872
rect -11928 -38913 -11755 -38885
rect -11950 -38926 -11755 -38913
rect -11950 -39075 -11889 -38926
rect -11828 -38932 -11755 -38926
rect -11318 -38902 -11284 -38730
rect -11016 -38902 -10946 -37565
rect -7042 -38119 -7008 -35860
rect -6858 -37008 -6824 -35468
rect -6748 -35602 -6609 -35548
rect -6218 -35583 -6184 -35468
rect -6123 -35507 -6089 -35155
rect -6053 -35433 -6019 -35086
rect -5873 -35433 -5839 -35190
rect -6053 -35467 -5839 -35433
rect -5677 -35507 -5643 -35190
rect -5367 -35383 -5333 -35190
rect -6123 -35541 -5643 -35507
rect -5590 -35558 -5451 -35504
rect -6218 -35617 -6072 -35583
rect -6749 -35720 -6418 -35683
rect -6366 -35706 -6227 -35652
rect -6106 -35679 -6072 -35617
rect -5999 -35632 -5860 -35578
rect -6106 -35713 -5545 -35679
rect -6749 -35803 -6712 -35720
rect -6455 -35744 -6418 -35720
rect -6455 -35781 -6299 -35744
rect -6747 -35992 -6713 -35803
rect -6751 -36115 -6712 -35992
rect -6649 -36041 -6615 -35796
rect -6336 -35802 -6299 -35781
rect -6333 -36004 -6299 -35802
rect -6237 -35805 -5937 -35766
rect -6235 -36004 -6201 -35805
rect -5971 -36004 -5937 -35805
rect -5873 -36004 -5839 -35713
rect -5677 -35987 -5643 -35796
rect -5677 -36041 -5641 -35987
rect -5579 -36004 -5545 -35713
rect -5372 -35722 -5329 -35383
rect -5058 -35381 -5024 -35190
rect -5062 -35578 -5019 -35381
rect -4975 -35564 -4836 -35510
rect -5162 -35624 -5019 -35578
rect -5288 -35712 -5149 -35658
rect -5468 -35768 -5329 -35722
rect -5372 -35813 -5329 -35768
rect -5367 -36004 -5333 -35813
rect -5269 -35997 -5235 -35796
rect -5062 -35815 -5019 -35624
rect -6649 -36077 -5641 -36041
rect -5274 -36081 -5231 -35997
rect -5058 -36004 -5024 -35815
rect -4960 -35995 -4926 -35796
rect -4247 -35086 -3519 -35052
rect -4247 -35398 -4213 -35086
rect -4149 -35434 -4115 -35190
rect -4051 -35398 -4017 -35086
rect -3931 -35155 -3589 -35121
rect -3931 -35398 -3897 -35155
rect -3833 -35434 -3799 -35190
rect -3735 -35398 -3701 -35155
rect -4415 -35468 -3684 -35434
rect -4415 -35831 -4381 -35468
rect -4248 -35602 -4109 -35548
rect -3718 -35583 -3684 -35468
rect -3623 -35507 -3589 -35155
rect -3553 -35433 -3519 -35086
rect -3373 -35433 -3339 -35190
rect -3553 -35467 -3339 -35433
rect -3177 -35507 -3143 -35190
rect -2867 -35383 -2833 -35190
rect -3623 -35541 -3143 -35507
rect -3090 -35558 -2951 -35504
rect -3718 -35617 -3572 -35583
rect -4249 -35720 -3918 -35683
rect -3866 -35706 -3727 -35652
rect -3606 -35679 -3572 -35617
rect -3499 -35632 -3360 -35578
rect -3606 -35713 -3045 -35679
rect -4249 -35803 -4212 -35720
rect -3955 -35744 -3918 -35720
rect -3955 -35781 -3799 -35744
rect -4421 -35967 -4375 -35831
rect -4247 -35992 -4213 -35803
rect -4965 -36080 -4922 -35995
rect -4251 -36080 -4212 -35992
rect -4149 -36041 -4115 -35796
rect -3836 -35802 -3799 -35781
rect -3833 -36004 -3799 -35802
rect -3737 -35805 -3437 -35766
rect -3735 -36004 -3701 -35805
rect -3471 -36004 -3437 -35805
rect -3373 -36004 -3339 -35713
rect -3177 -35987 -3143 -35796
rect -3177 -36041 -3141 -35987
rect -3079 -36004 -3045 -35713
rect -2872 -35722 -2829 -35383
rect -2558 -35381 -2524 -35190
rect -2562 -35578 -2519 -35381
rect -2475 -35564 -2336 -35510
rect -2662 -35624 -2519 -35578
rect -2788 -35712 -2649 -35658
rect -2968 -35768 -2829 -35722
rect -2872 -35813 -2829 -35768
rect -2867 -36004 -2833 -35813
rect -2769 -35997 -2735 -35796
rect -2562 -35815 -2519 -35624
rect -4149 -36077 -3141 -36041
rect -5039 -36081 -4212 -36080
rect -2774 -36081 -2731 -35997
rect -2558 -36004 -2524 -35815
rect -2460 -35995 -2426 -35796
rect -1747 -35086 -1019 -35052
rect -1747 -35398 -1713 -35086
rect -1649 -35434 -1615 -35190
rect -1551 -35398 -1517 -35086
rect -1431 -35155 -1089 -35121
rect -1431 -35398 -1397 -35155
rect -1333 -35434 -1299 -35190
rect -1235 -35398 -1201 -35155
rect -1867 -35468 -1184 -35434
rect -1867 -35835 -1833 -35468
rect -1748 -35602 -1609 -35548
rect -1218 -35583 -1184 -35468
rect -1123 -35507 -1089 -35155
rect -1053 -35433 -1019 -35086
rect -873 -35433 -839 -35190
rect -1053 -35467 -839 -35433
rect -677 -35507 -643 -35190
rect -367 -35383 -333 -35190
rect -1123 -35541 -643 -35507
rect -590 -35558 -451 -35504
rect -1218 -35617 -1072 -35583
rect -1749 -35720 -1418 -35683
rect -1366 -35706 -1227 -35652
rect -1106 -35679 -1072 -35617
rect -999 -35632 -860 -35578
rect -1106 -35713 -545 -35679
rect -1749 -35803 -1712 -35720
rect -1455 -35744 -1418 -35720
rect -1455 -35781 -1299 -35744
rect -1873 -35971 -1827 -35835
rect -1747 -35992 -1713 -35803
rect -2465 -36081 -2422 -35995
rect -5550 -36115 -4212 -36081
rect -3050 -36115 -2418 -36081
rect -1751 -36115 -1712 -35992
rect -1649 -36041 -1615 -35796
rect -1336 -35802 -1299 -35781
rect -1333 -36004 -1299 -35802
rect -1237 -35805 -937 -35766
rect -1235 -36004 -1201 -35805
rect -971 -36004 -937 -35805
rect -873 -36004 -839 -35713
rect -677 -35987 -643 -35796
rect -677 -36041 -641 -35987
rect -579 -36004 -545 -35713
rect -372 -35722 -329 -35383
rect -58 -35381 -24 -35190
rect -62 -35578 -19 -35381
rect 25 -35564 164 -35510
rect -162 -35624 -19 -35578
rect -288 -35712 -149 -35658
rect -468 -35768 -329 -35722
rect -372 -35813 -329 -35768
rect -367 -36004 -333 -35813
rect -269 -35997 -235 -35796
rect -62 -35815 -19 -35624
rect -1649 -36077 -641 -36041
rect -274 -36081 -231 -35997
rect -58 -36004 -24 -35815
rect 40 -35995 74 -35796
rect 753 -35086 1481 -35052
rect 753 -35398 787 -35086
rect 613 -35434 647 -35433
rect 851 -35434 885 -35190
rect 949 -35398 983 -35086
rect 1069 -35155 1411 -35121
rect 1069 -35398 1103 -35155
rect 1167 -35434 1201 -35190
rect 1265 -35398 1299 -35155
rect 613 -35468 1316 -35434
rect 613 -35835 647 -35468
rect 752 -35602 891 -35548
rect 1282 -35583 1316 -35468
rect 1377 -35507 1411 -35155
rect 1447 -35433 1481 -35086
rect 1627 -35433 1661 -35190
rect 1447 -35467 1661 -35433
rect 1823 -35507 1857 -35190
rect 2133 -35383 2167 -35190
rect 1377 -35541 1857 -35507
rect 1910 -35558 2049 -35504
rect 1282 -35617 1428 -35583
rect 751 -35720 1082 -35683
rect 1134 -35706 1273 -35652
rect 1394 -35679 1428 -35617
rect 1501 -35632 1640 -35578
rect 1394 -35713 1955 -35679
rect 751 -35803 788 -35720
rect 1045 -35744 1082 -35720
rect 1045 -35781 1201 -35744
rect 607 -35971 653 -35835
rect 753 -35992 787 -35803
rect 35 -36081 78 -35995
rect -550 -36115 82 -36081
rect 749 -36115 788 -35992
rect 851 -36041 885 -35796
rect 1164 -35802 1201 -35781
rect 1167 -36004 1201 -35802
rect 1263 -35805 1563 -35766
rect 1265 -36004 1299 -35805
rect 1529 -36004 1563 -35805
rect 1627 -36004 1661 -35713
rect 1823 -35987 1857 -35796
rect 1823 -36041 1859 -35987
rect 1921 -36004 1955 -35713
rect 2128 -35722 2171 -35383
rect 2442 -35381 2476 -35190
rect 3253 -35086 3981 -35052
rect 2438 -35578 2481 -35381
rect 3253 -35398 3287 -35086
rect 3351 -35434 3385 -35190
rect 3449 -35398 3483 -35086
rect 3569 -35155 3911 -35121
rect 3569 -35398 3603 -35155
rect 3667 -35434 3701 -35190
rect 3765 -35398 3799 -35155
rect 3029 -35468 3816 -35434
rect 2525 -35564 2664 -35510
rect 2338 -35624 2481 -35578
rect 2212 -35712 2351 -35658
rect 2032 -35768 2171 -35722
rect 2128 -35813 2171 -35768
rect 2133 -36004 2167 -35813
rect 2231 -35997 2265 -35796
rect 2438 -35815 2481 -35624
rect 851 -36077 1859 -36041
rect 2226 -36081 2269 -35997
rect 2442 -36004 2476 -35815
rect 2540 -35995 2574 -35796
rect 3029 -35834 3063 -35468
rect 3252 -35602 3391 -35548
rect 3782 -35583 3816 -35468
rect 3877 -35507 3911 -35155
rect 3947 -35433 3981 -35086
rect 4127 -35433 4161 -35190
rect 3947 -35467 4161 -35433
rect 4323 -35507 4357 -35190
rect 4633 -35383 4667 -35190
rect 3877 -35541 4357 -35507
rect 4410 -35558 4549 -35504
rect 3782 -35617 3928 -35583
rect 3251 -35720 3582 -35683
rect 3894 -35679 3928 -35617
rect 4001 -35632 4140 -35578
rect 3894 -35713 4455 -35679
rect 3251 -35803 3288 -35720
rect 3545 -35744 3582 -35720
rect 3545 -35781 3701 -35744
rect 3029 -35835 3064 -35834
rect 3024 -35971 3070 -35835
rect 3253 -35992 3287 -35803
rect 2535 -36081 2578 -35995
rect 1950 -36115 2582 -36081
rect 3249 -36115 3288 -35992
rect 3351 -36041 3385 -35796
rect 3664 -35802 3701 -35781
rect 3667 -36004 3701 -35802
rect 3763 -35805 4063 -35766
rect 3765 -36004 3799 -35805
rect 4029 -36004 4063 -35805
rect 4127 -36004 4161 -35713
rect 4323 -35987 4357 -35796
rect 4323 -36041 4359 -35987
rect 4421 -36004 4455 -35713
rect 4628 -35722 4671 -35383
rect 4942 -35381 4976 -35190
rect 6253 -35086 6981 -35052
rect 4938 -35578 4981 -35381
rect 6253 -35398 6287 -35086
rect 6351 -35434 6385 -35190
rect 6449 -35398 6483 -35086
rect 6569 -35155 6911 -35121
rect 6569 -35398 6603 -35155
rect 6667 -35434 6701 -35190
rect 6765 -35398 6799 -35155
rect 5935 -35468 6816 -35434
rect 5025 -35564 5164 -35510
rect 4838 -35624 4981 -35578
rect 4532 -35768 4671 -35722
rect 4628 -35813 4671 -35768
rect 4633 -36004 4667 -35813
rect 4731 -35997 4765 -35796
rect 4938 -35815 4981 -35624
rect 3351 -36077 4359 -36041
rect 4726 -36081 4769 -35997
rect 4942 -36004 4976 -35815
rect 5040 -35995 5074 -35796
rect 5935 -35835 5969 -35468
rect 6252 -35602 6391 -35548
rect 6782 -35583 6816 -35468
rect 6877 -35507 6911 -35155
rect 6947 -35433 6981 -35086
rect 7127 -35433 7161 -35190
rect 6947 -35467 7161 -35433
rect 7323 -35507 7357 -35190
rect 7633 -35383 7667 -35190
rect 6877 -35541 7357 -35507
rect 7410 -35558 7549 -35504
rect 6782 -35617 6928 -35583
rect 6251 -35720 6582 -35683
rect 6894 -35679 6928 -35617
rect 7001 -35632 7140 -35578
rect 6894 -35713 7455 -35679
rect 6251 -35803 6288 -35720
rect 6545 -35744 6582 -35720
rect 6545 -35781 6701 -35744
rect 5929 -35971 5975 -35835
rect 6253 -35992 6287 -35803
rect 5035 -36081 5078 -35995
rect 4450 -36115 5082 -36081
rect 6249 -36115 6288 -35992
rect 6351 -36041 6385 -35796
rect 6664 -35802 6701 -35781
rect 6667 -36004 6701 -35802
rect 6763 -35805 7063 -35766
rect 6765 -36004 6799 -35805
rect 7029 -36004 7063 -35805
rect 7127 -36004 7161 -35713
rect 7323 -35987 7357 -35796
rect 7323 -36041 7359 -35987
rect 7421 -36004 7455 -35713
rect 7628 -35722 7671 -35383
rect 7942 -35381 7976 -35190
rect 7938 -35578 7981 -35381
rect 8025 -35564 8164 -35510
rect 7838 -35624 7981 -35578
rect 7532 -35768 7671 -35722
rect 7628 -35813 7671 -35768
rect 7633 -36004 7667 -35813
rect 7731 -35997 7765 -35796
rect 7938 -35815 7981 -35624
rect 6351 -36077 7359 -36041
rect 7726 -36063 7769 -35997
rect 7942 -36004 7976 -35815
rect 8040 -35995 8074 -35796
rect 8035 -36063 8078 -35995
rect 8241 -36063 8502 -34202
rect 16856 -34526 17053 -34345
rect 16512 -35001 16793 -34792
rect 8726 -35204 8926 -35170
rect 16152 -35204 16514 -35158
rect 8726 -35376 16514 -35204
rect 8726 -35541 8926 -35376
rect 16152 -35429 16514 -35376
rect 7434 -36115 8502 -36063
rect 15912 -36102 16204 -36101
rect -6751 -36167 8502 -36115
rect -6751 -36168 -4918 -36167
rect -4251 -36168 8502 -36167
rect -6319 -36188 -5785 -36168
rect -5550 -36177 -4918 -36168
rect -3050 -36177 -2418 -36168
rect -550 -36177 82 -36168
rect 1950 -36177 2582 -36168
rect 4450 -36177 5082 -36168
rect -6310 -36347 -6276 -36188
rect -6212 -36331 -6178 -36239
rect -6218 -36424 -6172 -36331
rect -6114 -36347 -6080 -36188
rect -6016 -36331 -5982 -36239
rect -6022 -36424 -5976 -36331
rect -5918 -36347 -5884 -36188
rect 7434 -36190 8502 -36168
rect -5820 -36331 -5786 -36239
rect -1708 -36253 -1572 -36207
rect 789 -36223 925 -36220
rect -1621 -36301 -1572 -36253
rect 756 -36257 2927 -36223
rect 789 -36266 925 -36257
rect -5826 -36392 -5780 -36331
rect -4803 -36392 -4757 -36326
rect -1621 -36337 2831 -36301
rect -5826 -36424 -4757 -36392
rect -6218 -36462 -4757 -36424
rect -6218 -36470 -5780 -36462
rect -6218 -36723 -6172 -36470
rect -6212 -36727 -6178 -36723
rect -6022 -36535 -5976 -36470
rect -6016 -36727 -5982 -36535
rect -5826 -36535 -5780 -36470
rect -5820 -36727 -5786 -36535
rect -4421 -36673 -4375 -36537
rect 2795 -36449 2831 -36337
rect 2893 -36381 2927 -36257
rect 5877 -36273 6013 -36267
rect 2972 -36292 3108 -36283
rect 2972 -36326 5773 -36292
rect 5877 -36307 6149 -36273
rect 5877 -36313 6013 -36307
rect 2972 -36329 3108 -36326
rect 5739 -36365 5773 -36326
rect 2893 -36415 4395 -36381
rect 5739 -36399 6079 -36365
rect -6898 -37054 -6762 -37008
rect -4418 -36926 -4378 -36673
rect -4418 -36972 -4282 -36926
rect -7042 -38182 -6858 -38119
rect -7021 -38183 -6858 -38182
rect -12502 -39088 -12367 -39082
rect -12522 -39090 -12367 -39088
rect -12729 -39126 -12367 -39090
rect -12319 -39105 -11889 -39075
rect -12319 -39113 -11900 -39105
rect -11710 -39117 -11676 -38961
rect -11612 -39069 -11578 -38961
rect -11514 -39117 -11480 -38961
rect -11416 -39069 -11382 -38961
rect -11318 -38972 -10946 -38902
rect -6567 -37614 -6533 -37422
rect -6573 -37679 -6527 -37614
rect -6371 -37614 -6337 -37422
rect -6377 -37679 -6331 -37614
rect -6175 -37426 -6141 -37422
rect -6181 -37679 -6135 -37426
rect -5636 -37403 -5008 -37369
rect -5729 -37537 -5695 -37437
rect -5636 -37454 -5594 -37403
rect -5734 -37581 -5692 -37537
rect -5631 -37545 -5597 -37454
rect -5533 -37527 -5499 -37437
rect -5440 -37459 -5398 -37403
rect -5534 -37581 -5498 -37527
rect -5435 -37545 -5401 -37459
rect -5337 -37527 -5303 -37437
rect -5246 -37458 -5204 -37403
rect -5340 -37545 -5303 -37527
rect -5239 -37545 -5205 -37458
rect -5141 -37529 -5107 -37437
rect -5044 -37448 -5008 -37403
rect -5043 -37522 -5009 -37448
rect -5340 -37581 -5304 -37545
rect -5142 -37581 -5106 -37529
rect -5734 -37615 -5106 -37581
rect -6573 -37687 -6135 -37679
rect -6603 -37696 -6135 -37687
rect -6685 -37698 -6135 -37696
rect -6686 -37725 -6135 -37698
rect -6686 -37735 -6527 -37725
rect -6686 -38093 -6638 -37735
rect -6603 -37757 -6527 -37735
rect -6573 -37818 -6527 -37757
rect -6567 -37910 -6533 -37818
rect -6469 -37961 -6435 -37802
rect -6377 -37818 -6331 -37725
rect -6371 -37910 -6337 -37818
rect -6273 -37961 -6239 -37802
rect -6181 -37818 -6135 -37725
rect -6099 -37700 -5931 -37694
rect -5734 -37700 -5559 -37615
rect -5050 -37669 -5003 -37522
rect -4959 -37663 -4885 -37495
rect -4824 -37614 -4790 -37422
rect -6099 -37753 -5559 -37700
rect -5175 -37743 -5003 -37669
rect -6099 -37768 -5931 -37753
rect -5734 -37782 -5559 -37753
rect -6175 -37910 -6141 -37818
rect -6077 -37961 -6043 -37802
rect -5734 -37816 -5103 -37782
rect -5734 -37823 -5692 -37816
rect -5733 -37866 -5692 -37823
rect -5729 -37960 -5695 -37866
rect -5631 -37948 -5597 -37852
rect -5536 -37865 -5495 -37816
rect -6568 -38029 -6034 -37961
rect -5637 -38006 -5593 -37948
rect -5533 -37960 -5499 -37865
rect -5435 -37937 -5401 -37852
rect -5342 -37865 -5301 -37816
rect -5440 -38006 -5396 -37937
rect -5337 -37960 -5303 -37865
rect -5239 -37937 -5205 -37852
rect -5144 -37857 -5103 -37816
rect -5244 -38006 -5200 -37937
rect -5141 -37960 -5107 -37857
rect -5050 -37878 -5003 -37743
rect -4958 -37687 -4885 -37663
rect -4830 -37679 -4784 -37614
rect -4628 -37614 -4594 -37422
rect -4634 -37679 -4588 -37614
rect -4432 -37426 -4398 -37422
rect -4438 -37679 -4392 -37426
rect -4234 -37522 -4177 -37444
rect -4234 -37567 -3973 -37522
rect -4234 -37608 -4177 -37567
rect -4830 -37687 -4392 -37679
rect -4958 -37725 -4392 -37687
rect -4958 -37757 -4784 -37725
rect -4830 -37818 -4784 -37757
rect -5043 -37948 -5009 -37878
rect -4824 -37910 -4790 -37818
rect -5048 -38006 -5004 -37948
rect -4726 -37961 -4692 -37802
rect -4634 -37818 -4588 -37725
rect -4628 -37910 -4594 -37818
rect -4530 -37961 -4496 -37802
rect -4438 -37818 -4392 -37725
rect -4356 -37705 -4188 -37694
rect -4018 -37701 -3973 -37567
rect -3867 -37614 -3833 -37422
rect -3873 -37679 -3827 -37614
rect -3671 -37614 -3637 -37422
rect -3677 -37679 -3631 -37614
rect -3475 -37426 -3441 -37422
rect -3481 -37679 -3435 -37426
rect -2936 -37403 -2308 -37369
rect -3029 -37537 -2995 -37437
rect -2936 -37454 -2894 -37403
rect -3034 -37581 -2992 -37537
rect -2931 -37545 -2897 -37454
rect -2833 -37527 -2799 -37437
rect -2740 -37459 -2698 -37403
rect -2834 -37581 -2798 -37527
rect -2735 -37545 -2701 -37459
rect -2637 -37527 -2603 -37437
rect -2546 -37458 -2504 -37403
rect -2640 -37545 -2603 -37527
rect -2539 -37545 -2505 -37458
rect -2441 -37529 -2407 -37437
rect -2344 -37448 -2308 -37403
rect -2343 -37522 -2309 -37448
rect -2640 -37581 -2604 -37545
rect -2442 -37581 -2406 -37529
rect -3034 -37615 -2406 -37581
rect -3873 -37687 -3435 -37679
rect -3903 -37701 -3435 -37687
rect -4128 -37705 -4068 -37704
rect -4356 -37763 -4068 -37705
rect -4018 -37725 -3435 -37701
rect -4018 -37746 -3827 -37725
rect -4356 -37768 -4188 -37763
rect -4432 -37910 -4398 -37818
rect -4334 -37961 -4300 -37802
rect -4128 -37836 -4068 -37763
rect -4013 -37861 -3953 -37746
rect -3903 -37757 -3827 -37746
rect -3873 -37818 -3827 -37757
rect -3867 -37910 -3833 -37818
rect -3769 -37961 -3735 -37802
rect -3677 -37818 -3631 -37725
rect -3671 -37910 -3637 -37818
rect -3573 -37961 -3539 -37802
rect -3481 -37818 -3435 -37725
rect -3399 -37703 -3231 -37694
rect -3034 -37703 -2859 -37615
rect -2350 -37669 -2303 -37522
rect -2259 -37663 -2185 -37495
rect -2124 -37614 -2090 -37422
rect -3399 -37760 -2859 -37703
rect -2475 -37743 -2303 -37669
rect -3399 -37768 -3231 -37760
rect -3034 -37782 -2859 -37760
rect -3475 -37910 -3441 -37818
rect -3377 -37961 -3343 -37802
rect -3034 -37816 -2403 -37782
rect -3034 -37823 -2992 -37816
rect -3033 -37856 -2992 -37823
rect -3033 -37866 -2986 -37856
rect -5637 -38040 -5004 -38006
rect -4825 -38029 -3334 -37961
rect -3032 -37988 -2986 -37866
rect -2931 -37948 -2897 -37852
rect -2836 -37865 -2795 -37816
rect -2937 -38006 -2893 -37948
rect -2833 -37960 -2799 -37865
rect -2735 -37937 -2701 -37852
rect -2642 -37865 -2601 -37816
rect -2740 -38006 -2696 -37937
rect -2637 -37960 -2603 -37865
rect -2539 -37937 -2505 -37852
rect -2444 -37857 -2403 -37816
rect -2544 -38006 -2500 -37937
rect -2441 -37960 -2407 -37857
rect -2350 -37878 -2303 -37743
rect -2258 -37687 -2185 -37663
rect -2130 -37679 -2084 -37614
rect -1928 -37614 -1894 -37422
rect -1934 -37679 -1888 -37614
rect -1732 -37426 -1698 -37422
rect -1738 -37679 -1692 -37426
rect -1534 -37608 -1477 -37444
rect -1242 -37614 -1208 -37422
rect -2130 -37687 -1692 -37679
rect -1248 -37679 -1202 -37614
rect -1046 -37614 -1012 -37422
rect -1052 -37679 -1006 -37614
rect -850 -37426 -816 -37422
rect -856 -37679 -810 -37426
rect -1248 -37687 -810 -37679
rect -2258 -37725 -1692 -37687
rect -2258 -37757 -2084 -37725
rect -2343 -37948 -2309 -37878
rect -2348 -38006 -2304 -37948
rect -2937 -38040 -2304 -38006
rect -2130 -37818 -2084 -37757
rect -2124 -37910 -2090 -37818
rect -2026 -37961 -1992 -37802
rect -1934 -37818 -1888 -37725
rect -1928 -37910 -1894 -37818
rect -1830 -37961 -1796 -37802
rect -1738 -37818 -1692 -37725
rect -1396 -37709 -1336 -37705
rect -1278 -37709 -810 -37687
rect 2795 -36485 4316 -36449
rect 2631 -36970 2767 -36924
rect 2527 -37054 2682 -37008
rect -1396 -37725 -810 -37709
rect -1396 -37751 -1202 -37725
rect -1732 -37910 -1698 -37818
rect -1634 -37961 -1600 -37802
rect -1396 -37837 -1336 -37751
rect -1278 -37757 -1202 -37751
rect -1248 -37818 -1202 -37757
rect -1242 -37910 -1208 -37818
rect -1144 -37961 -1110 -37802
rect -1052 -37818 -1006 -37725
rect -1046 -37910 -1012 -37818
rect -948 -37961 -914 -37802
rect -856 -37818 -810 -37725
rect -850 -37910 -816 -37818
rect -752 -37961 -718 -37802
rect -2125 -38029 -709 -37961
rect -312 -37849 -278 -37439
rect 426 -37683 460 -37439
rect 622 -37683 656 -37439
rect 818 -37683 852 -37439
rect 297 -37720 852 -37683
rect 1038 -37686 1084 -37602
rect 1421 -37624 1455 -37452
rect 1617 -37560 1651 -37452
rect 1813 -37560 1847 -37452
rect -463 -37902 -278 -37849
rect -243 -37858 -108 -37848
rect 297 -37858 334 -37720
rect 892 -37740 1084 -37686
rect 1284 -37694 1455 -37624
rect 1892 -37607 1965 -37594
rect 1892 -37635 2065 -37607
rect 1892 -37648 2087 -37635
rect 1892 -37654 1965 -37648
rect 556 -37777 691 -37768
rect 1119 -37777 1255 -37776
rect 556 -37815 1255 -37777
rect 556 -37822 691 -37815
rect 1119 -37822 1255 -37815
rect -243 -37895 334 -37858
rect -243 -37902 -108 -37895
rect -6687 -38230 -6627 -38093
rect -4177 -38162 -4040 -38152
rect -3231 -38162 -3099 -38151
rect -1217 -38162 -1085 -38152
rect -6356 -38201 -1085 -38162
rect -4177 -38212 -4040 -38201
rect -3231 -38211 -3099 -38201
rect -1217 -38212 -1085 -38201
rect -6686 -38602 -6638 -38230
rect -6339 -38254 -6202 -38241
rect -3742 -38254 -3605 -38235
rect -974 -38254 -842 -38235
rect -6356 -38293 -841 -38254
rect -6339 -38301 -6202 -38293
rect -6328 -38341 -6217 -38301
rect -5517 -38341 -5406 -38293
rect -3742 -38295 -3605 -38293
rect -6576 -38409 -5205 -38341
rect -5026 -38364 -4393 -38330
rect -3719 -38341 -3608 -38295
rect -3536 -38341 -3016 -38339
rect -2841 -38341 -2730 -38293
rect -6567 -38568 -6533 -38409
rect -6469 -38552 -6435 -38460
rect -6686 -38646 -6511 -38602
rect -6679 -38676 -6511 -38646
rect -6475 -38645 -6429 -38552
rect -6371 -38568 -6337 -38409
rect -6273 -38552 -6239 -38460
rect -6279 -38645 -6233 -38552
rect -6175 -38568 -6141 -38409
rect -6077 -38552 -6043 -38460
rect -6083 -38613 -6037 -38552
rect -5730 -38568 -5696 -38409
rect -5632 -38552 -5598 -38460
rect -6083 -38645 -5950 -38613
rect -6475 -38683 -5950 -38645
rect -5638 -38645 -5592 -38552
rect -5534 -38568 -5500 -38409
rect -5436 -38552 -5402 -38460
rect -5442 -38645 -5396 -38552
rect -5338 -38568 -5304 -38409
rect -5026 -38422 -4982 -38364
rect -5240 -38552 -5206 -38460
rect -5021 -38492 -4987 -38422
rect -5246 -38613 -5200 -38552
rect -5246 -38645 -5072 -38613
rect -6475 -38691 -6037 -38683
rect -6475 -38944 -6429 -38691
rect -6469 -38948 -6435 -38944
rect -6279 -38756 -6233 -38691
rect -6273 -38948 -6239 -38756
rect -6083 -38756 -6037 -38691
rect -6077 -38948 -6043 -38756
rect -5996 -38813 -5950 -38683
rect -5638 -38683 -5072 -38645
rect -5638 -38691 -5200 -38683
rect -5853 -38813 -5796 -38762
rect -5996 -38862 -5796 -38813
rect -5853 -38926 -5796 -38862
rect -5638 -38944 -5592 -38691
rect -5632 -38948 -5598 -38944
rect -5442 -38756 -5396 -38691
rect -5436 -38948 -5402 -38756
rect -5246 -38756 -5200 -38691
rect -5145 -38707 -5072 -38683
rect -5027 -38627 -4980 -38492
rect -4923 -38513 -4889 -38410
rect -4830 -38433 -4786 -38364
rect -4927 -38554 -4886 -38513
rect -4825 -38518 -4791 -38433
rect -4727 -38505 -4693 -38410
rect -4634 -38433 -4590 -38364
rect -4729 -38554 -4688 -38505
rect -4629 -38518 -4595 -38433
rect -4531 -38505 -4497 -38410
rect -4437 -38422 -4393 -38364
rect -3876 -38407 -2505 -38341
rect -3876 -38409 -3342 -38407
rect -3039 -38409 -2505 -38407
rect -2326 -38364 -1693 -38330
rect -4535 -38554 -4494 -38505
rect -4433 -38518 -4399 -38422
rect -4335 -38504 -4301 -38410
rect -4338 -38547 -4297 -38504
rect -4338 -38554 -4296 -38547
rect -4927 -38588 -4296 -38554
rect -3867 -38568 -3833 -38409
rect -3769 -38552 -3735 -38460
rect -5027 -38701 -4855 -38627
rect -4471 -38648 -4205 -38588
rect -3979 -38609 -3811 -38602
rect -5240 -38948 -5206 -38756
rect -5145 -38875 -5071 -38707
rect -5027 -38848 -4980 -38701
rect -4471 -38755 -4296 -38648
rect -4001 -38669 -3811 -38609
rect -3979 -38676 -3811 -38669
rect -3775 -38645 -3729 -38552
rect -3671 -38568 -3637 -38409
rect -3573 -38552 -3539 -38460
rect -3579 -38645 -3533 -38552
rect -3475 -38568 -3441 -38409
rect -3377 -38552 -3343 -38460
rect -3383 -38613 -3337 -38552
rect -3202 -38602 -3142 -38443
rect -3030 -38568 -2996 -38409
rect -2932 -38552 -2898 -38460
rect -3383 -38645 -3239 -38613
rect -3775 -38683 -3239 -38645
rect -3202 -38665 -2974 -38602
rect -3142 -38676 -2974 -38665
rect -2938 -38645 -2892 -38552
rect -2834 -38568 -2800 -38409
rect -2736 -38552 -2702 -38460
rect -2742 -38645 -2696 -38552
rect -2638 -38568 -2604 -38409
rect -2326 -38422 -2282 -38364
rect -2540 -38552 -2506 -38460
rect -2321 -38492 -2287 -38422
rect -2546 -38613 -2500 -38552
rect -2546 -38645 -2372 -38613
rect -3775 -38691 -3337 -38683
rect -4924 -38789 -4296 -38755
rect -4924 -38841 -4888 -38789
rect -4726 -38825 -4690 -38789
rect -5021 -38922 -4987 -38848
rect -5022 -38967 -4986 -38922
rect -4923 -38933 -4889 -38841
rect -4825 -38912 -4791 -38825
rect -4727 -38843 -4690 -38825
rect -4826 -38967 -4784 -38912
rect -4727 -38933 -4693 -38843
rect -4629 -38911 -4595 -38825
rect -4532 -38843 -4496 -38789
rect -4632 -38967 -4590 -38911
rect -4531 -38933 -4497 -38843
rect -4433 -38916 -4399 -38825
rect -4338 -38833 -4296 -38789
rect -4436 -38967 -4394 -38916
rect -4335 -38933 -4301 -38833
rect -5022 -39001 -4394 -38967
rect -3775 -38944 -3729 -38691
rect -3769 -38948 -3735 -38944
rect -3579 -38756 -3533 -38691
rect -3573 -38948 -3539 -38756
rect -3383 -38756 -3337 -38691
rect -3377 -38948 -3343 -38756
rect -3301 -38812 -3239 -38683
rect -2938 -38683 -2372 -38645
rect -2938 -38691 -2500 -38683
rect -3153 -38812 -3096 -38762
rect -3301 -38874 -3096 -38812
rect -3153 -38926 -3096 -38874
rect -2938 -38944 -2892 -38691
rect -2932 -38948 -2898 -38944
rect -2742 -38756 -2696 -38691
rect -2736 -38948 -2702 -38756
rect -2546 -38756 -2500 -38691
rect -2445 -38707 -2372 -38683
rect -2327 -38627 -2280 -38492
rect -2223 -38513 -2189 -38410
rect -2130 -38433 -2086 -38364
rect -2227 -38554 -2186 -38513
rect -2125 -38518 -2091 -38433
rect -2027 -38505 -1993 -38410
rect -1934 -38433 -1890 -38364
rect -2029 -38554 -1988 -38505
rect -1929 -38518 -1895 -38433
rect -1831 -38505 -1797 -38410
rect -1737 -38422 -1693 -38364
rect -1835 -38554 -1794 -38505
rect -1733 -38518 -1699 -38422
rect -1635 -38504 -1601 -38410
rect -1638 -38547 -1597 -38504
rect -1638 -38554 -1596 -38547
rect -2227 -38586 -1596 -38554
rect -2227 -38588 -1521 -38586
rect -2327 -38701 -2155 -38627
rect -1771 -38646 -1521 -38588
rect -2540 -38948 -2506 -38756
rect -2445 -38875 -2371 -38707
rect -2327 -38848 -2280 -38701
rect -1771 -38755 -1596 -38646
rect -2224 -38789 -1596 -38755
rect -2224 -38841 -2188 -38789
rect -2026 -38825 -1990 -38789
rect -2321 -38922 -2287 -38848
rect -2322 -38967 -2286 -38922
rect -2223 -38933 -2189 -38841
rect -2125 -38912 -2091 -38825
rect -2027 -38843 -1990 -38825
rect -2126 -38967 -2084 -38912
rect -2027 -38933 -1993 -38843
rect -1929 -38911 -1895 -38825
rect -1832 -38843 -1796 -38789
rect -1932 -38967 -1890 -38911
rect -1831 -38933 -1797 -38843
rect -1733 -38916 -1699 -38825
rect -1638 -38833 -1596 -38789
rect -1736 -38967 -1694 -38916
rect -1635 -38933 -1601 -38833
rect -1357 -38873 -1059 -38293
rect -974 -38295 -842 -38293
rect -312 -38355 -278 -37902
rect 297 -37949 334 -37895
rect 368 -37859 503 -37846
rect 1290 -37859 1324 -37694
rect 1519 -37791 1553 -37683
rect 1617 -37839 1651 -37683
rect 1715 -37791 1749 -37683
rect 1813 -37839 1847 -37683
rect 2026 -37797 2087 -37648
rect 2226 -37797 2260 -37453
rect 2422 -37797 2456 -37453
rect 2026 -37827 2456 -37797
rect 2646 -37804 2682 -37054
rect 2037 -37835 2456 -37827
rect 2504 -37812 2682 -37804
rect 368 -37893 1324 -37859
rect 368 -37900 503 -37893
rect 1372 -37925 1987 -37839
rect 2504 -37848 2691 -37812
rect 2504 -37852 2669 -37848
rect 2504 -37858 2639 -37852
rect 2100 -37908 2174 -37882
rect 2727 -37906 2767 -36970
rect 3026 -37626 3060 -37454
rect 3222 -37562 3256 -37454
rect 3418 -37562 3452 -37454
rect 2585 -37908 2767 -37906
rect 101 -37983 334 -37949
rect 507 -37983 950 -37949
rect -214 -38543 -180 -38147
rect 101 -38355 135 -37983
rect 199 -38453 233 -38047
rect 297 -38355 331 -37983
rect 507 -37984 754 -37983
rect 507 -38047 542 -37984
rect 410 -38344 444 -38047
rect 409 -38450 444 -38344
rect 508 -38355 542 -38047
rect 606 -38346 640 -38047
rect 605 -38450 640 -38346
rect 720 -38354 754 -37984
rect 409 -38453 640 -38450
rect 199 -38487 640 -38453
rect 818 -38543 852 -38046
rect 916 -38354 950 -37983
rect 1682 -38332 1743 -37925
rect 2100 -37946 2767 -37908
rect 2862 -37696 3060 -37626
rect 3497 -37609 3570 -37596
rect 3497 -37637 3670 -37609
rect 3497 -37650 3692 -37637
rect 3497 -37656 3570 -37650
rect 2100 -37947 2586 -37946
rect 2100 -37953 2174 -37947
rect 2515 -37948 2586 -37947
rect 2128 -38298 2162 -37990
rect 2226 -38298 2260 -37990
rect 2324 -38298 2358 -37990
rect 2422 -38298 2456 -37990
rect 2520 -38298 2554 -37990
rect 1682 -38350 2132 -38332
rect 2422 -38350 2457 -38298
rect 1682 -38393 2574 -38350
rect -324 -38608 950 -38543
rect -311 -38873 -181 -38608
rect -5 -38873 125 -38608
rect 312 -38873 442 -38608
rect 758 -38873 888 -38608
rect 1682 -38873 1833 -38393
rect 2059 -38411 2574 -38393
rect 2059 -38873 2183 -38411
rect 2389 -38873 2513 -38411
rect 2862 -38431 2932 -37696
rect 3124 -37793 3158 -37685
rect 3222 -37841 3256 -37685
rect 3320 -37793 3354 -37685
rect 3418 -37841 3452 -37685
rect 3631 -37799 3692 -37650
rect 3831 -37799 3865 -37455
rect 4027 -37799 4061 -37455
rect 3631 -37829 4061 -37799
rect 3642 -37837 4061 -37829
rect 4109 -37812 4244 -37806
rect 4280 -37812 4316 -36485
rect 2977 -37927 3592 -37841
rect 4109 -37850 4316 -37812
rect 4109 -37852 4296 -37850
rect 4109 -37860 4244 -37852
rect 3705 -37910 3779 -37884
rect 4355 -37908 4395 -36415
rect 4190 -37910 4395 -37908
rect 2796 -38477 2932 -38431
rect 3287 -38334 3348 -37927
rect 3705 -37948 4395 -37910
rect 3705 -37949 4191 -37948
rect 3705 -37955 3779 -37949
rect 4120 -37950 4191 -37949
rect 3733 -38300 3767 -37992
rect 3831 -38300 3865 -37992
rect 3929 -38300 3963 -37992
rect 4027 -38300 4061 -37992
rect 4125 -38300 4159 -37992
rect 4650 -38030 4684 -37430
rect 5388 -37674 5422 -37430
rect 5584 -37674 5618 -37430
rect 5780 -37674 5814 -37430
rect 5259 -37711 5814 -37674
rect 5854 -37685 5989 -37677
rect 4719 -37849 4854 -37839
rect 5259 -37849 5296 -37711
rect 5853 -37722 6008 -37685
rect 5853 -37731 5989 -37722
rect 5518 -37768 5653 -37759
rect 6045 -37768 6079 -36399
rect 5518 -37806 6079 -37768
rect 5518 -37813 5653 -37806
rect 4719 -37886 5296 -37849
rect 4719 -37893 4854 -37886
rect 5259 -37940 5296 -37886
rect 5330 -37850 5465 -37837
rect 6115 -37850 6149 -36307
rect 6263 -37337 6991 -37303
rect 6263 -37649 6297 -37337
rect 6361 -37685 6395 -37441
rect 6459 -37649 6493 -37337
rect 6579 -37406 6921 -37372
rect 6579 -37649 6613 -37406
rect 6677 -37685 6711 -37441
rect 6775 -37649 6809 -37406
rect 6212 -37719 6826 -37685
rect 5330 -37884 6149 -37850
rect 6262 -37853 6401 -37799
rect 6792 -37834 6826 -37719
rect 6887 -37758 6921 -37406
rect 6957 -37684 6991 -37337
rect 7137 -37684 7171 -37441
rect 6957 -37718 7171 -37684
rect 7333 -37758 7367 -37441
rect 7643 -37634 7677 -37441
rect 6887 -37792 7367 -37758
rect 7420 -37809 7559 -37755
rect 6792 -37868 6938 -37834
rect 5330 -37891 5465 -37884
rect 4434 -38088 4684 -38030
rect 3287 -38352 3737 -38334
rect 4027 -38352 4062 -38300
rect 3287 -38395 4179 -38352
rect 3287 -38873 3438 -38395
rect 3729 -38413 4179 -38395
rect 3729 -38873 3880 -38413
rect 4022 -38873 4173 -38413
rect 4434 -38543 4499 -38088
rect 4650 -38346 4684 -38088
rect 5063 -37974 5296 -37940
rect 5469 -37974 5912 -37940
rect 4748 -38534 4782 -38138
rect 5063 -38346 5097 -37974
rect 5161 -38444 5195 -38038
rect 5259 -38346 5293 -37974
rect 5469 -37975 5716 -37974
rect 5469 -38038 5504 -37975
rect 5372 -38335 5406 -38038
rect 5371 -38441 5406 -38335
rect 5470 -38346 5504 -38038
rect 5568 -38337 5602 -38038
rect 5567 -38441 5602 -38337
rect 5682 -38345 5716 -37975
rect 5371 -38444 5602 -38441
rect 5161 -38478 5602 -38444
rect 5780 -38534 5814 -38037
rect 5878 -38345 5912 -37974
rect 6261 -37971 6592 -37934
rect 6904 -37930 6938 -37868
rect 7011 -37883 7150 -37829
rect 6904 -37964 7465 -37930
rect 6261 -38054 6298 -37971
rect 6555 -37995 6592 -37971
rect 6555 -38032 6711 -37995
rect 6263 -38243 6297 -38054
rect 6259 -38366 6298 -38243
rect 6361 -38292 6395 -38047
rect 6674 -38053 6711 -38032
rect 6677 -38255 6711 -38053
rect 6773 -38056 7073 -38017
rect 6775 -38255 6809 -38056
rect 7039 -38255 7073 -38056
rect 7137 -38255 7171 -37964
rect 7333 -38238 7367 -38047
rect 7333 -38292 7369 -38238
rect 7431 -38255 7465 -37964
rect 7638 -37973 7681 -37634
rect 7952 -37632 7986 -37441
rect 7948 -37829 7991 -37632
rect 8035 -37815 8174 -37761
rect 7848 -37875 7991 -37829
rect 7542 -38019 7681 -37973
rect 7638 -38064 7681 -38019
rect 7643 -38255 7677 -38064
rect 7741 -38248 7775 -38047
rect 7948 -38066 7991 -37875
rect 6361 -38328 7369 -38292
rect 7736 -38332 7779 -38248
rect 7952 -38255 7986 -38066
rect 8050 -38246 8084 -38047
rect 8045 -38332 8088 -38246
rect 7460 -38366 8092 -38332
rect 6259 -38419 8092 -38366
rect 4364 -38589 4500 -38543
rect 4638 -38599 5912 -38534
rect 4662 -38873 4808 -38599
rect 5107 -38873 5253 -38599
rect 5373 -38873 5519 -38599
rect 5733 -38873 5879 -38599
rect 6297 -38873 6494 -38419
rect 6830 -38873 7027 -38419
rect 7343 -38428 8092 -38419
rect 7343 -38873 7540 -38428
rect 7846 -38873 8043 -38428
rect 8241 -38873 8502 -36190
rect 8938 -36241 16204 -36102
rect 15879 -37121 16146 -37085
rect 10534 -37356 16146 -37121
rect 15879 -37383 16146 -37356
rect 8966 -37715 9184 -37707
rect 16142 -37715 16295 -37676
rect 8966 -37790 16295 -37715
rect 8966 -37796 9184 -37790
rect 16142 -37827 16295 -37790
rect 9948 -37936 9998 -37930
rect 15460 -37936 15558 -37922
rect 9939 -38059 15558 -37936
rect 9948 -38063 9998 -38059
rect 15460 -38086 15558 -38059
rect 16377 -38341 16505 -35429
rect 16630 -38252 16762 -35001
rect 16872 -37676 16961 -34526
rect 18964 -35740 19509 -34202
rect 18381 -36246 84354 -35740
rect 16872 -37827 16969 -37676
rect 18964 -37710 19509 -36246
rect 28710 -36707 28993 -36246
rect 28466 -36735 29131 -36707
rect 34078 -36722 34435 -36655
rect 35256 -36722 35613 -36689
rect 37109 -36718 37392 -36246
rect 28466 -36793 29501 -36735
rect 28466 -36874 28552 -36793
rect 28726 -36830 28761 -36793
rect 29051 -36796 29501 -36793
rect 27614 -36960 28552 -36874
rect 27462 -37250 27592 -37158
rect 27754 -37216 27788 -36960
rect 27852 -37216 27886 -37008
rect 27950 -37216 27984 -36960
rect 28048 -37182 28082 -37008
rect 28629 -37138 28663 -36830
rect 28727 -37138 28761 -36830
rect 28825 -37138 28859 -36830
rect 28923 -37138 28957 -36830
rect 29021 -37138 29055 -36830
rect 28597 -37181 28668 -37180
rect 29009 -37181 29083 -37175
rect 28597 -37182 29083 -37181
rect 28048 -37216 29083 -37182
rect 29440 -37203 29501 -36796
rect 34078 -36911 35613 -36722
rect 36906 -36746 37571 -36718
rect 36906 -36804 37941 -36746
rect 46021 -36757 46304 -36246
rect 55240 -36723 55523 -36246
rect 60589 -36691 60965 -36596
rect 64035 -36657 64342 -36246
rect 62190 -36691 62440 -36664
rect 36906 -36885 36992 -36804
rect 37166 -36841 37201 -36804
rect 37491 -36807 37941 -36804
rect 34078 -36922 34435 -36911
rect 35256 -36956 35613 -36911
rect 36054 -36971 36992 -36885
rect 28049 -37220 29083 -37216
rect 28049 -37222 28598 -37220
rect 27636 -37250 27709 -37244
rect 29009 -37246 29083 -37220
rect 27462 -37291 27709 -37250
rect 27462 -37308 27592 -37291
rect 27636 -37304 27709 -37291
rect 29196 -37289 29981 -37203
rect 35902 -37261 36032 -37169
rect 36194 -37227 36228 -36971
rect 36292 -37227 36326 -37019
rect 36390 -37227 36424 -36971
rect 36488 -37193 36522 -37019
rect 37069 -37149 37103 -36841
rect 37167 -37149 37201 -36841
rect 37265 -37149 37299 -36841
rect 37363 -37149 37397 -36841
rect 37461 -37149 37495 -36841
rect 37037 -37192 37108 -37191
rect 37449 -37192 37523 -37186
rect 37037 -37193 37523 -37192
rect 36488 -37227 37523 -37193
rect 37880 -37214 37941 -36807
rect 42634 -36811 42899 -36780
rect 44160 -36811 44457 -36778
rect 42634 -36978 44457 -36811
rect 45769 -36785 46434 -36757
rect 45769 -36843 46804 -36785
rect 45769 -36924 45855 -36843
rect 46029 -36880 46064 -36843
rect 46354 -36846 46804 -36843
rect 42634 -37045 42899 -36978
rect 44160 -37000 44457 -36978
rect 44917 -37010 45855 -36924
rect 36489 -37231 37523 -37227
rect 36489 -37233 37038 -37231
rect 36076 -37261 36149 -37255
rect 37449 -37257 37523 -37231
rect 28727 -37301 29146 -37293
rect 28727 -37331 29157 -37301
rect 27754 -37546 27788 -37338
rect 27950 -37546 27984 -37338
rect 28146 -37546 28180 -37338
rect 20374 -37672 21002 -37638
rect 16872 -38160 16961 -37827
rect 18066 -37816 19836 -37710
rect 20281 -37806 20315 -37706
rect 20374 -37723 20416 -37672
rect 18170 -37962 18218 -37816
rect 18175 -38133 18209 -37962
rect 18273 -38116 18307 -37925
rect 18364 -37965 18412 -37816
rect 17989 -38160 18134 -38153
rect 16872 -38201 18134 -38160
rect 17989 -38209 18134 -38201
rect 18269 -38167 18311 -38116
rect 18371 -38133 18405 -37965
rect 18469 -38116 18503 -37925
rect 18465 -38167 18507 -38116
rect 18269 -38209 19055 -38167
rect 18916 -38227 19055 -38209
rect 18318 -38252 18463 -38248
rect 16630 -38293 18463 -38252
rect 18318 -38304 18463 -38293
rect 18638 -38336 18783 -38280
rect 18638 -38341 18698 -38336
rect 16377 -38382 18698 -38341
rect 18916 -38409 18958 -38227
rect 18171 -38455 18620 -38418
rect -2322 -39001 -1694 -38967
rect -12522 -39128 -12367 -39126
rect -12502 -39136 -12367 -39128
rect -12997 -39186 -12448 -39184
rect -12037 -39186 -11963 -39160
rect -12997 -39190 -11963 -39186
rect -13292 -39446 -13258 -39190
rect -13194 -39398 -13160 -39190
rect -13096 -39446 -13062 -39190
rect -12998 -39224 -11963 -39190
rect -11850 -39203 -11065 -39117
rect -12998 -39398 -12964 -39224
rect -12449 -39225 -11963 -39224
rect -12449 -39226 -12378 -39225
rect -12037 -39231 -11963 -39225
rect -13432 -39532 -12494 -39446
rect -12580 -39613 -12494 -39532
rect -12417 -39576 -12383 -39268
rect -12319 -39576 -12285 -39268
rect -12221 -39576 -12187 -39268
rect -12123 -39576 -12089 -39268
rect -12025 -39576 -11991 -39268
rect -12320 -39613 -12285 -39576
rect -11606 -39610 -11545 -39203
rect -11995 -39613 -11545 -39610
rect -12580 -39671 -11545 -39613
rect -12580 -39699 -11915 -39671
rect -25977 -42987 -24335 -42872
rect -25977 -43127 -25639 -42987
rect -23728 -44174 -23542 -39776
rect -16396 -39808 -16128 -39776
rect -14343 -39915 -14309 -39911
rect -14349 -40168 -14303 -39915
rect -14147 -40103 -14113 -39911
rect -14153 -40168 -14107 -40103
rect -13951 -40103 -13917 -39911
rect -13727 -39997 -13670 -39933
rect -13870 -40046 -13670 -39997
rect -13957 -40168 -13911 -40103
rect -14349 -40176 -13911 -40168
rect -13870 -40176 -13824 -40046
rect -13727 -40097 -13670 -40046
rect -13506 -39915 -13472 -39911
rect -14553 -40213 -14385 -40183
rect -14560 -40257 -14385 -40213
rect -14349 -40214 -13824 -40176
rect -13512 -40168 -13466 -39915
rect -13310 -40103 -13276 -39911
rect -13316 -40168 -13270 -40103
rect -12896 -39892 -12268 -39858
rect -13114 -40103 -13080 -39911
rect -12896 -39937 -12860 -39892
rect -13120 -40168 -13074 -40103
rect -13512 -40176 -13074 -40168
rect -13019 -40152 -12945 -39984
rect -12895 -40011 -12861 -39937
rect -13019 -40176 -12946 -40152
rect -13716 -40194 -13548 -40183
rect -13751 -40195 -13548 -40194
rect -21820 -41587 -21786 -40996
rect -21520 -40960 -21057 -40926
rect -21824 -41638 -21783 -41587
rect -21608 -41594 -21574 -40996
rect -21520 -41002 -21467 -40960
rect -21613 -41638 -21571 -41594
rect -21510 -41604 -21476 -41002
rect -21412 -41593 -21378 -40996
rect -21311 -41002 -21255 -40960
rect -21417 -41638 -21375 -41593
rect -21299 -41604 -21265 -41002
rect -21201 -41586 -21167 -40996
rect -21113 -41002 -21057 -40960
rect -21824 -41675 -21375 -41638
rect -21205 -41642 -21163 -41586
rect -21103 -41604 -21069 -41002
rect -20614 -41328 -20580 -40925
rect -20410 -40889 -20166 -40851
rect -20615 -41367 -20579 -41328
rect -20410 -40953 -20364 -40889
rect -20403 -41333 -20369 -40953
rect -20305 -41323 -20271 -40925
rect -20212 -40953 -20166 -40889
rect -20207 -41287 -20173 -40953
rect -20312 -41367 -20267 -41323
rect -20615 -41403 -20267 -41367
rect -20210 -41519 -20160 -41287
rect -19709 -41329 -19675 -40926
rect -19505 -40890 -19261 -40852
rect -19976 -41450 -19918 -41355
rect -19710 -41368 -19674 -41329
rect -19505 -40954 -19459 -40890
rect -19498 -41334 -19464 -40954
rect -19400 -41324 -19366 -40926
rect -19307 -40954 -19261 -40890
rect -17594 -40928 -16117 -40815
rect -19302 -41288 -19268 -40954
rect -18425 -41223 -17976 -41205
rect -17594 -41223 -17533 -40928
rect -16867 -41046 -16820 -40928
rect -18937 -41284 -17533 -41223
rect -19407 -41368 -19362 -41324
rect -19710 -41404 -19362 -41368
rect -19580 -41450 -19437 -41443
rect -19976 -41486 -19437 -41450
rect -19976 -41492 -19918 -41486
rect -19580 -41503 -19437 -41486
rect -20817 -41538 -20759 -41525
rect -20708 -41538 -20562 -41522
rect -20210 -41532 -20064 -41519
rect -19305 -41520 -19255 -41288
rect -20817 -41574 -20562 -41538
rect -20266 -41541 -20064 -41532
rect -21205 -41684 -21037 -41642
rect -20817 -41662 -20759 -41574
rect -20708 -41582 -20562 -41574
rect -20521 -41577 -20064 -41541
rect -19899 -41539 -19841 -41527
rect -19803 -41539 -19657 -41523
rect -19305 -41533 -19133 -41520
rect -19899 -41575 -19657 -41539
rect -19361 -41542 -19133 -41533
rect -21079 -41868 -21037 -41684
rect -20614 -41776 -20580 -41617
rect -20521 -41626 -20476 -41577
rect -21088 -41884 -20951 -41868
rect -21726 -41926 -20951 -41884
rect -21820 -42131 -21786 -41960
rect -21726 -41977 -21684 -41926
rect -21825 -42260 -21777 -42131
rect -21722 -42168 -21688 -41977
rect -21624 -42128 -21590 -41960
rect -21530 -41977 -21488 -41926
rect -20618 -41928 -20574 -41776
rect -20516 -41825 -20482 -41626
rect -20418 -41777 -20384 -41617
rect -19899 -41664 -19841 -41575
rect -19803 -41583 -19657 -41575
rect -19616 -41578 -19133 -41542
rect -19709 -41777 -19675 -41618
rect -19616 -41627 -19571 -41578
rect -20424 -41928 -20380 -41777
rect -20747 -41963 -20150 -41928
rect -19713 -41929 -19669 -41777
rect -19611 -41826 -19577 -41627
rect -19513 -41778 -19479 -41618
rect -18937 -41642 -18876 -41284
rect -18308 -41318 -18273 -41284
rect -18405 -41626 -18371 -41318
rect -18307 -41626 -18273 -41318
rect -18209 -41626 -18175 -41318
rect -18111 -41626 -18077 -41318
rect -18013 -41626 -17979 -41318
rect -19324 -41703 -18876 -41642
rect -18437 -41669 -18366 -41668
rect -18025 -41669 -17951 -41663
rect -18437 -41670 -17951 -41669
rect -19519 -41929 -19475 -41778
rect -19324 -41929 -19263 -41703
rect -18663 -41708 -17951 -41670
rect -17594 -41691 -17533 -41284
rect -16860 -41340 -16826 -41046
rect -16762 -41324 -16728 -41032
rect -16671 -41047 -16624 -40928
rect -16969 -41386 -16814 -41374
rect -17006 -41420 -16814 -41386
rect -16969 -41429 -16814 -41420
rect -16768 -41394 -16723 -41324
rect -16664 -41340 -16630 -41047
rect -16429 -41057 -16382 -40928
rect -16422 -41340 -16388 -41057
rect -16324 -41331 -16290 -41032
rect -16328 -41371 -16284 -41331
rect -15436 -41371 -15299 -41301
rect -16328 -41374 -15299 -41371
rect -16768 -41434 -16414 -41394
rect -16376 -41414 -15299 -41374
rect -17104 -41491 -17034 -41489
rect -16699 -41491 -16544 -41482
rect -17104 -41527 -16544 -41491
rect -18663 -41710 -18436 -41708
rect -18025 -41734 -17951 -41708
rect -19009 -41768 -18892 -41753
rect -18490 -41766 -18355 -41758
rect -18510 -41768 -18355 -41766
rect -19009 -41804 -18355 -41768
rect -17838 -41777 -17223 -41691
rect -19009 -41876 -18892 -41804
rect -18510 -41806 -18355 -41804
rect -18490 -41812 -18355 -41806
rect -18307 -41789 -17888 -41781
rect -18307 -41819 -17877 -41789
rect -19842 -41963 -19245 -41929
rect -21631 -42260 -21583 -42128
rect -21526 -42168 -21492 -41977
rect -21302 -42018 -19245 -41963
rect -21302 -42079 -19461 -42018
rect -21302 -42260 -21186 -42079
rect -21960 -42277 -21156 -42260
rect -18307 -42163 -18273 -41819
rect -18111 -42163 -18077 -41819
rect -17938 -41968 -17877 -41819
rect -17698 -41933 -17664 -41777
rect -17600 -41933 -17566 -41825
rect -17502 -41933 -17468 -41777
rect -17404 -41933 -17370 -41825
rect -17104 -41922 -17034 -41527
rect -16699 -41537 -16544 -41527
rect -16457 -41504 -16414 -41434
rect -16457 -41559 -16276 -41504
rect -16457 -41571 -16414 -41559
rect -16864 -41609 -16610 -41573
rect -17816 -41968 -17743 -41962
rect -17938 -41981 -17743 -41968
rect -17916 -42009 -17743 -41981
rect -17816 -42022 -17743 -42009
rect -17306 -41992 -17028 -41922
rect -17698 -42164 -17664 -42056
rect -17502 -42164 -17468 -42056
rect -17306 -42164 -17272 -41992
rect -16864 -41668 -16822 -41609
rect -21960 -42383 -21072 -42277
rect -16860 -42252 -16826 -41668
rect -16652 -41662 -16610 -41609
rect -16555 -41610 -16414 -41571
rect -16649 -42244 -16615 -41662
rect -16555 -41664 -16513 -41610
rect -16653 -42286 -16611 -42244
rect -16551 -42252 -16517 -41664
rect -16453 -42242 -16419 -41644
rect -16242 -41658 -16199 -41414
rect -15436 -41467 -15299 -41414
rect -16016 -41589 -15911 -41517
rect -14560 -40629 -14512 -40257
rect -14441 -40450 -14407 -40291
rect -14349 -40307 -14303 -40214
rect -14343 -40399 -14309 -40307
rect -14245 -40450 -14211 -40291
rect -14153 -40307 -14107 -40214
rect -13957 -40246 -13824 -40214
rect -14147 -40399 -14113 -40307
rect -14049 -40450 -14015 -40291
rect -13957 -40307 -13911 -40246
rect -13788 -40257 -13548 -40195
rect -13512 -40214 -12946 -40176
rect -13951 -40399 -13917 -40307
rect -13788 -40401 -13728 -40257
rect -13604 -40450 -13570 -40291
rect -13512 -40307 -13466 -40214
rect -13506 -40399 -13472 -40307
rect -13408 -40450 -13374 -40291
rect -13316 -40307 -13270 -40214
rect -13120 -40246 -12946 -40214
rect -12901 -40158 -12854 -40011
rect -12797 -40018 -12763 -39926
rect -12700 -39947 -12658 -39892
rect -12798 -40070 -12762 -40018
rect -12699 -40034 -12665 -39947
rect -12601 -40016 -12567 -39926
rect -12506 -39948 -12464 -39892
rect -12601 -40034 -12564 -40016
rect -12503 -40034 -12469 -39948
rect -12405 -40016 -12371 -39926
rect -12310 -39943 -12268 -39892
rect -12600 -40070 -12564 -40034
rect -12406 -40070 -12370 -40016
rect -12307 -40034 -12273 -39943
rect -12209 -40026 -12175 -39926
rect -12212 -40070 -12170 -40026
rect -12798 -40104 -12170 -40070
rect -12901 -40232 -12729 -40158
rect -12345 -40211 -12170 -40104
rect -11643 -39915 -11609 -39911
rect -11649 -40168 -11603 -39915
rect -11447 -40103 -11413 -39911
rect -11453 -40168 -11407 -40103
rect -11251 -40103 -11217 -39911
rect -11027 -39985 -10970 -39933
rect -11175 -40047 -10970 -39985
rect -11257 -40168 -11211 -40103
rect -11649 -40176 -11211 -40168
rect -11175 -40176 -11113 -40047
rect -11027 -40097 -10970 -40047
rect -10806 -39915 -10772 -39911
rect -11853 -40190 -11685 -40183
rect -13310 -40399 -13276 -40307
rect -13212 -40450 -13178 -40291
rect -13120 -40307 -13074 -40246
rect -13114 -40399 -13080 -40307
rect -12901 -40367 -12854 -40232
rect -12345 -40271 -12079 -40211
rect -11875 -40250 -11685 -40190
rect -11853 -40257 -11685 -40250
rect -11649 -40214 -11113 -40176
rect -10812 -40168 -10766 -39915
rect -10610 -40103 -10576 -39911
rect -10616 -40168 -10570 -40103
rect -10196 -39892 -9568 -39858
rect -10414 -40103 -10380 -39911
rect -10196 -39937 -10160 -39892
rect -10420 -40168 -10374 -40103
rect -10812 -40176 -10374 -40168
rect -10319 -40152 -10245 -39984
rect -10195 -40011 -10161 -39937
rect -10319 -40176 -10246 -40152
rect -11016 -40194 -10848 -40183
rect -12801 -40305 -12170 -40271
rect -12801 -40346 -12760 -40305
rect -12895 -40437 -12861 -40367
rect -14450 -40518 -13079 -40450
rect -12900 -40495 -12856 -40437
rect -12797 -40449 -12763 -40346
rect -12699 -40426 -12665 -40341
rect -12603 -40354 -12562 -40305
rect -12704 -40495 -12660 -40426
rect -12601 -40449 -12567 -40354
rect -12503 -40426 -12469 -40341
rect -12409 -40354 -12368 -40305
rect -12212 -40312 -12170 -40305
rect -12508 -40495 -12464 -40426
rect -12405 -40449 -12371 -40354
rect -12307 -40437 -12273 -40341
rect -12212 -40355 -12171 -40312
rect -12311 -40495 -12267 -40437
rect -12209 -40449 -12175 -40355
rect -11741 -40450 -11707 -40291
rect -11649 -40307 -11603 -40214
rect -11643 -40399 -11609 -40307
rect -11545 -40450 -11511 -40291
rect -11453 -40307 -11407 -40214
rect -11257 -40246 -11113 -40214
rect -11447 -40399 -11413 -40307
rect -11349 -40450 -11315 -40291
rect -11257 -40307 -11211 -40246
rect -11076 -40257 -10848 -40194
rect -10812 -40214 -10246 -40176
rect -11251 -40399 -11217 -40307
rect -11076 -40416 -11016 -40257
rect -10904 -40450 -10870 -40291
rect -10812 -40307 -10766 -40214
rect -10806 -40399 -10772 -40307
rect -10708 -40450 -10674 -40291
rect -10616 -40307 -10570 -40214
rect -10420 -40246 -10246 -40214
rect -10201 -40158 -10154 -40011
rect -10097 -40018 -10063 -39926
rect -10000 -39947 -9958 -39892
rect -10098 -40070 -10062 -40018
rect -9999 -40034 -9965 -39947
rect -9901 -40016 -9867 -39926
rect -9806 -39948 -9764 -39892
rect -9901 -40034 -9864 -40016
rect -9803 -40034 -9769 -39948
rect -9705 -40016 -9671 -39926
rect -9610 -39943 -9568 -39892
rect -9900 -40070 -9864 -40034
rect -9706 -40070 -9670 -40016
rect -9607 -40034 -9573 -39943
rect -9509 -40026 -9475 -39926
rect -9512 -40070 -9470 -40026
rect -10098 -40104 -9470 -40070
rect -10201 -40232 -10029 -40158
rect -9645 -40213 -9470 -40104
rect -10610 -40399 -10576 -40307
rect -10512 -40450 -10478 -40291
rect -10420 -40307 -10374 -40246
rect -10414 -40399 -10380 -40307
rect -10201 -40367 -10154 -40232
rect -9645 -40271 -9395 -40213
rect -10101 -40273 -9395 -40271
rect -10101 -40305 -9470 -40273
rect -10101 -40346 -10060 -40305
rect -10195 -40437 -10161 -40367
rect -14202 -40558 -14091 -40518
rect -14213 -40566 -14076 -40558
rect -13391 -40566 -13280 -40518
rect -12900 -40529 -12267 -40495
rect -11750 -40452 -11216 -40450
rect -10913 -40452 -10379 -40450
rect -11750 -40518 -10379 -40452
rect -10200 -40495 -10156 -40437
rect -10097 -40449 -10063 -40346
rect -9999 -40426 -9965 -40341
rect -9903 -40354 -9862 -40305
rect -10004 -40495 -9960 -40426
rect -9901 -40449 -9867 -40354
rect -9803 -40426 -9769 -40341
rect -9709 -40354 -9668 -40305
rect -9512 -40312 -9470 -40305
rect -9808 -40495 -9764 -40426
rect -9705 -40449 -9671 -40354
rect -9607 -40437 -9573 -40341
rect -9512 -40355 -9471 -40312
rect -9611 -40495 -9567 -40437
rect -9509 -40449 -9475 -40355
rect -11593 -40564 -11482 -40518
rect -11410 -40520 -10890 -40518
rect -11616 -40566 -11479 -40564
rect -10715 -40566 -10604 -40518
rect -10200 -40529 -9567 -40495
rect -8150 -40522 -8116 -39928
rect -7944 -39894 -7704 -39860
rect -7944 -39938 -7902 -39894
rect -8978 -40566 -8846 -40564
rect -14230 -40605 -8845 -40566
rect -14213 -40618 -14076 -40605
rect -11616 -40624 -11479 -40605
rect -8978 -40624 -8846 -40605
rect -14561 -40766 -14501 -40629
rect -12051 -40658 -11914 -40647
rect -11105 -40658 -10973 -40648
rect -14230 -40697 -8500 -40658
rect -12051 -40707 -11914 -40697
rect -11105 -40708 -10973 -40697
rect -13824 -40744 -13692 -40736
rect -9301 -40744 -9169 -40734
rect -14560 -41124 -14512 -40766
rect -14230 -40783 -9169 -40744
rect -13824 -40796 -13692 -40783
rect -9301 -40794 -9169 -40783
rect -8539 -40766 -8500 -40697
rect -8158 -40766 -8115 -40522
rect -7938 -40536 -7904 -39938
rect -7840 -40516 -7806 -39928
rect -7746 -39936 -7704 -39894
rect -7844 -40570 -7802 -40516
rect -7742 -40518 -7708 -39936
rect -7943 -40609 -7802 -40570
rect -7747 -40571 -7705 -40518
rect -7531 -40512 -7497 -39928
rect -7535 -40571 -7493 -40512
rect -1357 -39134 8502 -38873
rect 18171 -38506 18212 -38455
rect -1357 -39992 -1059 -39134
rect 252 -39992 513 -39134
rect 1089 -39992 1350 -39134
rect 2129 -39992 2390 -39134
rect 3587 -39992 3848 -39134
rect 4801 -39992 5062 -39134
rect 6747 -39992 7008 -39134
rect 8241 -39992 8502 -39134
rect 18175 -39097 18209 -38506
rect 18382 -38499 18424 -38455
rect 18387 -39097 18421 -38499
rect 18485 -39091 18519 -38489
rect 18578 -38500 18620 -38455
rect 18790 -38451 18958 -38409
rect 18475 -39133 18528 -39091
rect 18583 -39097 18617 -38500
rect 18696 -39091 18730 -38489
rect 18790 -38507 18832 -38451
rect 18684 -39133 18740 -39091
rect 18794 -39097 18828 -38507
rect 18892 -39091 18926 -38489
rect 18882 -39133 18938 -39091
rect 18475 -39167 18938 -39133
rect -7747 -40607 -7493 -40571
rect -7943 -40621 -7900 -40609
rect -8081 -40676 -7900 -40621
rect -7943 -40746 -7900 -40676
rect -7813 -40653 -7658 -40643
rect -7300 -40653 -7168 -40601
rect -7813 -40689 -7168 -40653
rect -7813 -40698 -7658 -40689
rect -8539 -40806 -7981 -40766
rect -7943 -40786 -7589 -40746
rect -8539 -40809 -8029 -40806
rect -14442 -40898 -13908 -40830
rect -13511 -40853 -12878 -40819
rect -14441 -41041 -14407 -40949
rect -14447 -41102 -14401 -41041
rect -14343 -41057 -14309 -40898
rect -14245 -41041 -14211 -40949
rect -14477 -41124 -14401 -41102
rect -14560 -41134 -14401 -41124
rect -14251 -41134 -14205 -41041
rect -14147 -41057 -14113 -40898
rect -14049 -41041 -14015 -40949
rect -14055 -41134 -14009 -41041
rect -13951 -41057 -13917 -40898
rect -13603 -40993 -13569 -40899
rect -13511 -40911 -13467 -40853
rect -13607 -41036 -13566 -40993
rect -13505 -41007 -13471 -40911
rect -13407 -40994 -13373 -40899
rect -13314 -40922 -13270 -40853
rect -13608 -41043 -13566 -41036
rect -13410 -41043 -13369 -40994
rect -13309 -41007 -13275 -40922
rect -13211 -40994 -13177 -40899
rect -13118 -40922 -13074 -40853
rect -13216 -41043 -13175 -40994
rect -13113 -41007 -13079 -40922
rect -13015 -41002 -12981 -40899
rect -12922 -40911 -12878 -40853
rect -12699 -40898 -11208 -40830
rect -10811 -40853 -10178 -40819
rect -12917 -40981 -12883 -40911
rect -13018 -41043 -12977 -41002
rect -13608 -41077 -12977 -41043
rect -14560 -41161 -14009 -41134
rect -14559 -41163 -14009 -41161
rect -14477 -41172 -14009 -41163
rect -13973 -41106 -13805 -41091
rect -13608 -41106 -13433 -41077
rect -13973 -41159 -13433 -41106
rect -12924 -41116 -12877 -40981
rect -12698 -41041 -12664 -40949
rect -12704 -41102 -12658 -41041
rect -12600 -41057 -12566 -40898
rect -12502 -41041 -12468 -40949
rect -13973 -41165 -13805 -41159
rect -14447 -41180 -14009 -41172
rect -14447 -41245 -14401 -41180
rect -14441 -41437 -14407 -41245
rect -14251 -41245 -14205 -41180
rect -14245 -41437 -14211 -41245
rect -14055 -41433 -14009 -41180
rect -14049 -41437 -14015 -41433
rect -13608 -41244 -13433 -41159
rect -13049 -41190 -12877 -41116
rect -13608 -41278 -12980 -41244
rect -13608 -41322 -13566 -41278
rect -13603 -41422 -13569 -41322
rect -13505 -41405 -13471 -41314
rect -13408 -41332 -13372 -41278
rect -13214 -41314 -13178 -41278
rect -13510 -41456 -13468 -41405
rect -13407 -41422 -13373 -41332
rect -13309 -41400 -13275 -41314
rect -13214 -41332 -13177 -41314
rect -13314 -41456 -13272 -41400
rect -13211 -41422 -13177 -41332
rect -13113 -41401 -13079 -41314
rect -13016 -41330 -12980 -41278
rect -13120 -41456 -13078 -41401
rect -13015 -41422 -12981 -41330
rect -12924 -41337 -12877 -41190
rect -12832 -41134 -12658 -41102
rect -12508 -41134 -12462 -41041
rect -12404 -41057 -12370 -40898
rect -12306 -41041 -12272 -40949
rect -12312 -41134 -12266 -41041
rect -12208 -41057 -12174 -40898
rect -12832 -41172 -12266 -41134
rect -12230 -41096 -12062 -41091
rect -12002 -41096 -11942 -41023
rect -12230 -41154 -11942 -41096
rect -11887 -41113 -11827 -40998
rect -11741 -41041 -11707 -40949
rect -11747 -41102 -11701 -41041
rect -11643 -41057 -11609 -40898
rect -11545 -41041 -11511 -40949
rect -11777 -41113 -11701 -41102
rect -12230 -41165 -12062 -41154
rect -12002 -41155 -11942 -41154
rect -11892 -41134 -11701 -41113
rect -11551 -41134 -11505 -41041
rect -11447 -41057 -11413 -40898
rect -11349 -41041 -11315 -40949
rect -11355 -41134 -11309 -41041
rect -11251 -41057 -11217 -40898
rect -10906 -40993 -10860 -40871
rect -10811 -40911 -10767 -40853
rect -10907 -41003 -10860 -40993
rect -10907 -41036 -10866 -41003
rect -10805 -41007 -10771 -40911
rect -10707 -40994 -10673 -40899
rect -10614 -40922 -10570 -40853
rect -10908 -41043 -10866 -41036
rect -10710 -41043 -10669 -40994
rect -10609 -41007 -10575 -40922
rect -10511 -40994 -10477 -40899
rect -10418 -40922 -10374 -40853
rect -10516 -41043 -10475 -40994
rect -10413 -41007 -10379 -40922
rect -10315 -41002 -10281 -40899
rect -10222 -40911 -10178 -40853
rect -9999 -40898 -8583 -40830
rect -10217 -40981 -10183 -40911
rect -10318 -41043 -10277 -41002
rect -10908 -41077 -10277 -41043
rect -11892 -41158 -11309 -41134
rect -12832 -41196 -12759 -41172
rect -12917 -41411 -12883 -41337
rect -12833 -41364 -12759 -41196
rect -12704 -41180 -12266 -41172
rect -12704 -41245 -12658 -41180
rect -12918 -41456 -12882 -41411
rect -12698 -41437 -12664 -41245
rect -13510 -41490 -12882 -41456
rect -12508 -41245 -12462 -41180
rect -12502 -41437 -12468 -41245
rect -12312 -41433 -12266 -41180
rect -12306 -41437 -12272 -41433
rect -12108 -41292 -12051 -41251
rect -11892 -41292 -11847 -41158
rect -11777 -41172 -11309 -41158
rect -11273 -41099 -11105 -41091
rect -10908 -41099 -10733 -41077
rect -11273 -41156 -10733 -41099
rect -10224 -41116 -10177 -40981
rect -9998 -41041 -9964 -40949
rect -10004 -41102 -9958 -41041
rect -9900 -41057 -9866 -40898
rect -9802 -41041 -9768 -40949
rect -11273 -41165 -11105 -41156
rect -11747 -41180 -11309 -41172
rect -11747 -41245 -11701 -41180
rect -12108 -41337 -11847 -41292
rect -12108 -41415 -12051 -41337
rect -11741 -41437 -11707 -41245
rect -11551 -41245 -11505 -41180
rect -11545 -41437 -11511 -41245
rect -11355 -41433 -11309 -41180
rect -11349 -41437 -11315 -41433
rect -10908 -41244 -10733 -41156
rect -10349 -41190 -10177 -41116
rect -10908 -41278 -10280 -41244
rect -10908 -41322 -10866 -41278
rect -10903 -41422 -10869 -41322
rect -10805 -41405 -10771 -41314
rect -10708 -41332 -10672 -41278
rect -10514 -41314 -10478 -41278
rect -10810 -41456 -10768 -41405
rect -10707 -41422 -10673 -41332
rect -10609 -41400 -10575 -41314
rect -10514 -41332 -10477 -41314
rect -10614 -41456 -10572 -41400
rect -10511 -41422 -10477 -41332
rect -10413 -41401 -10379 -41314
rect -10316 -41330 -10280 -41278
rect -10420 -41456 -10378 -41401
rect -10315 -41422 -10281 -41330
rect -10224 -41337 -10177 -41190
rect -10132 -41134 -9958 -41102
rect -9808 -41134 -9762 -41041
rect -9704 -41057 -9670 -40898
rect -9606 -41041 -9572 -40949
rect -9612 -41134 -9566 -41041
rect -9508 -41057 -9474 -40898
rect -10132 -41172 -9566 -41134
rect -9530 -41096 -9362 -41091
rect -9530 -41108 -9327 -41096
rect -9270 -41108 -9210 -41022
rect -9116 -41041 -9082 -40949
rect -9122 -41102 -9076 -41041
rect -9018 -41057 -8984 -40898
rect -8920 -41041 -8886 -40949
rect -9152 -41108 -9076 -41102
rect -9530 -41134 -9076 -41108
rect -8926 -41134 -8880 -41041
rect -8822 -41057 -8788 -40898
rect -8724 -41041 -8690 -40949
rect -8730 -41134 -8684 -41041
rect -8626 -41057 -8592 -40898
rect -8539 -41091 -8500 -40809
rect -8073 -40849 -8029 -40809
rect -9530 -41150 -8684 -41134
rect -9530 -41154 -9327 -41150
rect -9270 -41154 -9210 -41150
rect -9530 -41165 -9362 -41154
rect -9152 -41172 -8684 -41150
rect -8648 -41165 -8480 -41091
rect -8067 -41148 -8033 -40849
rect -7969 -41123 -7935 -40840
rect -10132 -41196 -10059 -41172
rect -10217 -41411 -10183 -41337
rect -10133 -41364 -10059 -41196
rect -10004 -41180 -9566 -41172
rect -10004 -41245 -9958 -41180
rect -10218 -41456 -10182 -41411
rect -9998 -41437 -9964 -41245
rect -10810 -41490 -10182 -41456
rect -9808 -41245 -9762 -41180
rect -9802 -41437 -9768 -41245
rect -9612 -41433 -9566 -41180
rect -9122 -41180 -8684 -41172
rect -9606 -41437 -9572 -41433
rect -9122 -41245 -9076 -41180
rect -9408 -41415 -9351 -41251
rect -9116 -41437 -9082 -41245
rect -8926 -41245 -8880 -41180
rect -8920 -41437 -8886 -41245
rect -8730 -41433 -8684 -41180
rect -8724 -41437 -8690 -41433
rect -7975 -41253 -7928 -41123
rect -7727 -41133 -7693 -40840
rect -7634 -40856 -7589 -40786
rect -7543 -40760 -7388 -40751
rect -7025 -40760 -6883 -40743
rect -7543 -40794 -6883 -40760
rect -7543 -40806 -7388 -40794
rect -7025 -40807 -6883 -40794
rect -7733 -41253 -7686 -41133
rect -7629 -41148 -7595 -40856
rect -7531 -41134 -7497 -40840
rect -7537 -41253 -7490 -41134
rect -7026 -41253 -6921 -41247
rect -8155 -41335 -6921 -41253
rect -7026 -41342 -6921 -41335
rect -16455 -42286 -16413 -42242
rect -16653 -42320 -16413 -42286
rect -16241 -42252 -16207 -41658
rect -21960 -42410 -21156 -42383
rect -22674 -42575 -22616 -42572
rect -20819 -42575 -20761 -42479
rect -22674 -42616 -20761 -42575
rect -22674 -42709 -22616 -42616
rect -22560 -42654 -22502 -42653
rect -19998 -42654 -19940 -42558
rect -22560 -42695 -19940 -42654
rect -22560 -42790 -22502 -42695
rect -19905 -42731 -19847 -42635
rect -22415 -42772 -19847 -42731
rect -22415 -42868 -22357 -42772
rect -22173 -42853 -21190 -42822
rect -22173 -42918 -20895 -42853
rect -22173 -42937 -21190 -42918
rect -22157 -44022 -22123 -43106
rect -22059 -43314 -22025 -42937
rect -21646 -43008 -21205 -42974
rect -21744 -43478 -21710 -43106
rect -21646 -43414 -21612 -43008
rect -21436 -43011 -21205 -43008
rect -21548 -43478 -21514 -43106
rect -21436 -43117 -21401 -43011
rect -21435 -43414 -21401 -43117
rect -21337 -43414 -21303 -43106
rect -21240 -43115 -21205 -43011
rect -21239 -43414 -21205 -43115
rect -21338 -43477 -21303 -43414
rect -21125 -43477 -21091 -43107
rect -21027 -43415 -20993 -42918
rect -21338 -43478 -21091 -43477
rect -20929 -43478 -20895 -43107
rect -21744 -43512 -21511 -43478
rect -21338 -43512 -20895 -43478
rect -22088 -43566 -21953 -43559
rect -21548 -43566 -21511 -43512
rect -22088 -43603 -21511 -43566
rect -22088 -43613 -21953 -43603
rect -21548 -43741 -21511 -43603
rect -21477 -43568 -21342 -43561
rect -20848 -43568 -20790 -43465
rect -21477 -43602 -20790 -43568
rect -21477 -43615 -21342 -43602
rect -21289 -43646 -21154 -43639
rect -20118 -43646 -20060 -43547
rect -18281 -43092 -18247 -42884
rect -18085 -43092 -18051 -42884
rect -17889 -43092 -17855 -42884
rect -17308 -43099 -17274 -42755
rect -17112 -43099 -17078 -42755
rect -16699 -42862 -16665 -42754
rect -16503 -42862 -16469 -42754
rect -16817 -42909 -16744 -42896
rect -16917 -42937 -16744 -42909
rect -16939 -42950 -16744 -42937
rect -16939 -43099 -16878 -42950
rect -16817 -42956 -16744 -42950
rect -16307 -42926 -16273 -42754
rect -16005 -42926 -15935 -41589
rect -6469 -40182 -6435 -40178
rect -6475 -40435 -6429 -40182
rect -6273 -40370 -6239 -40178
rect -6279 -40435 -6233 -40370
rect -6077 -40370 -6043 -40178
rect -5853 -40264 -5796 -40200
rect -5996 -40313 -5796 -40264
rect -6083 -40435 -6037 -40370
rect -6475 -40443 -6037 -40435
rect -5996 -40443 -5950 -40313
rect -5853 -40364 -5796 -40313
rect -5632 -40182 -5598 -40178
rect -6679 -40480 -6511 -40450
rect -6686 -40524 -6511 -40480
rect -6475 -40481 -5950 -40443
rect -5638 -40435 -5592 -40182
rect -5436 -40370 -5402 -40178
rect -5442 -40435 -5396 -40370
rect -5022 -40159 -4394 -40125
rect -5240 -40370 -5206 -40178
rect -5022 -40204 -4986 -40159
rect -5246 -40435 -5200 -40370
rect -5638 -40443 -5200 -40435
rect -5145 -40419 -5071 -40251
rect -5021 -40278 -4987 -40204
rect -5145 -40443 -5072 -40419
rect -5842 -40461 -5674 -40450
rect -5877 -40462 -5674 -40461
rect -6686 -40896 -6638 -40524
rect -6567 -40717 -6533 -40558
rect -6475 -40574 -6429 -40481
rect -6469 -40666 -6435 -40574
rect -6371 -40717 -6337 -40558
rect -6279 -40574 -6233 -40481
rect -6083 -40513 -5950 -40481
rect -6273 -40666 -6239 -40574
rect -6175 -40717 -6141 -40558
rect -6083 -40574 -6037 -40513
rect -5914 -40524 -5674 -40462
rect -5638 -40481 -5072 -40443
rect -6077 -40666 -6043 -40574
rect -5914 -40668 -5854 -40524
rect -5730 -40717 -5696 -40558
rect -5638 -40574 -5592 -40481
rect -5632 -40666 -5598 -40574
rect -5534 -40717 -5500 -40558
rect -5442 -40574 -5396 -40481
rect -5246 -40513 -5072 -40481
rect -5027 -40425 -4980 -40278
rect -4923 -40285 -4889 -40193
rect -4826 -40214 -4784 -40159
rect -4924 -40337 -4888 -40285
rect -4825 -40301 -4791 -40214
rect -4727 -40283 -4693 -40193
rect -4632 -40215 -4590 -40159
rect -4727 -40301 -4690 -40283
rect -4629 -40301 -4595 -40215
rect -4531 -40283 -4497 -40193
rect -4436 -40210 -4394 -40159
rect -4726 -40337 -4690 -40301
rect -4532 -40337 -4496 -40283
rect -4433 -40301 -4399 -40210
rect -4335 -40293 -4301 -40193
rect -4338 -40337 -4296 -40293
rect -4924 -40371 -4296 -40337
rect -5027 -40499 -4855 -40425
rect -4471 -40478 -4296 -40371
rect -3769 -40182 -3735 -40178
rect -3775 -40435 -3729 -40182
rect -3573 -40370 -3539 -40178
rect -3579 -40435 -3533 -40370
rect -3377 -40370 -3343 -40178
rect -3153 -40252 -3096 -40200
rect -3301 -40314 -3096 -40252
rect -3383 -40435 -3337 -40370
rect -3775 -40443 -3337 -40435
rect -3301 -40443 -3239 -40314
rect -3153 -40364 -3096 -40314
rect -2932 -40182 -2898 -40178
rect -3979 -40457 -3811 -40450
rect -5436 -40666 -5402 -40574
rect -5338 -40717 -5304 -40558
rect -5246 -40574 -5200 -40513
rect -5240 -40666 -5206 -40574
rect -5027 -40634 -4980 -40499
rect -4471 -40538 -4205 -40478
rect -4001 -40517 -3811 -40457
rect -3979 -40524 -3811 -40517
rect -3775 -40481 -3239 -40443
rect -2938 -40435 -2892 -40182
rect -2736 -40370 -2702 -40178
rect -2742 -40435 -2696 -40370
rect -2322 -40159 -1694 -40125
rect -2540 -40370 -2506 -40178
rect -2322 -40204 -2286 -40159
rect -2546 -40435 -2500 -40370
rect -2938 -40443 -2500 -40435
rect -2445 -40419 -2371 -40251
rect -2321 -40278 -2287 -40204
rect -2445 -40443 -2372 -40419
rect -4927 -40572 -4296 -40538
rect -4927 -40613 -4886 -40572
rect -5021 -40704 -4987 -40634
rect -6576 -40785 -5205 -40717
rect -5026 -40762 -4982 -40704
rect -4923 -40716 -4889 -40613
rect -4825 -40693 -4791 -40608
rect -4729 -40621 -4688 -40572
rect -4830 -40762 -4786 -40693
rect -4727 -40716 -4693 -40621
rect -4629 -40693 -4595 -40608
rect -4535 -40621 -4494 -40572
rect -4338 -40579 -4296 -40572
rect -4634 -40762 -4590 -40693
rect -4531 -40716 -4497 -40621
rect -4433 -40704 -4399 -40608
rect -4338 -40622 -4297 -40579
rect -4437 -40762 -4393 -40704
rect -4335 -40716 -4301 -40622
rect -3867 -40717 -3833 -40558
rect -3775 -40574 -3729 -40481
rect -3769 -40666 -3735 -40574
rect -3671 -40717 -3637 -40558
rect -3579 -40574 -3533 -40481
rect -3383 -40513 -3239 -40481
rect -3573 -40666 -3539 -40574
rect -3475 -40717 -3441 -40558
rect -3383 -40574 -3337 -40513
rect -2938 -40481 -2372 -40443
rect -3377 -40666 -3343 -40574
rect -3030 -40717 -2996 -40558
rect -2938 -40574 -2892 -40481
rect -2932 -40666 -2898 -40574
rect -2834 -40717 -2800 -40558
rect -2742 -40574 -2696 -40481
rect -2546 -40513 -2372 -40481
rect -2327 -40425 -2280 -40278
rect -2223 -40285 -2189 -40193
rect -2126 -40214 -2084 -40159
rect -2224 -40337 -2188 -40285
rect -2125 -40301 -2091 -40214
rect -2027 -40283 -1993 -40193
rect -1932 -40215 -1890 -40159
rect -2027 -40301 -1990 -40283
rect -1929 -40301 -1895 -40215
rect -1831 -40283 -1797 -40193
rect -1736 -40210 -1694 -40159
rect -2026 -40337 -1990 -40301
rect -1832 -40337 -1796 -40283
rect -1733 -40301 -1699 -40210
rect -1635 -40293 -1601 -40193
rect -1357 -40253 8502 -39992
rect 14248 -39865 14762 -39702
rect 16008 -39865 16229 -39837
rect 14248 -39995 16229 -39865
rect 14248 -40127 14762 -39995
rect -1638 -40337 -1596 -40293
rect -2224 -40371 -1596 -40337
rect -2327 -40499 -2155 -40425
rect -1771 -40480 -1596 -40371
rect -2736 -40666 -2702 -40574
rect -2638 -40717 -2604 -40558
rect -2546 -40574 -2500 -40513
rect -2540 -40666 -2506 -40574
rect -2327 -40634 -2280 -40499
rect -1771 -40538 -1521 -40480
rect -2227 -40540 -1521 -40538
rect -2227 -40572 -1596 -40540
rect -2227 -40613 -2186 -40572
rect -2321 -40704 -2287 -40634
rect -6328 -40825 -6217 -40785
rect -6339 -40833 -6202 -40825
rect -5517 -40833 -5406 -40785
rect -5026 -40796 -4393 -40762
rect -3876 -40719 -3342 -40717
rect -3039 -40719 -2505 -40717
rect -3876 -40785 -2505 -40719
rect -2326 -40762 -2282 -40704
rect -2223 -40716 -2189 -40613
rect -2125 -40693 -2091 -40608
rect -2029 -40621 -1988 -40572
rect -2130 -40762 -2086 -40693
rect -2027 -40716 -1993 -40621
rect -1929 -40693 -1895 -40608
rect -1835 -40621 -1794 -40572
rect -1638 -40579 -1596 -40572
rect -1934 -40762 -1890 -40693
rect -1831 -40716 -1797 -40621
rect -1733 -40704 -1699 -40608
rect -1638 -40622 -1597 -40579
rect -1737 -40762 -1693 -40704
rect -1635 -40716 -1601 -40622
rect -3719 -40831 -3608 -40785
rect -3536 -40787 -3016 -40785
rect -3742 -40833 -3605 -40831
rect -2841 -40833 -2730 -40785
rect -2326 -40796 -1693 -40762
rect -1357 -40831 -1059 -40253
rect -311 -40518 -181 -40253
rect -5 -40518 125 -40253
rect 312 -40518 442 -40253
rect 758 -40518 888 -40253
rect -324 -40583 950 -40518
rect -1357 -40833 -972 -40831
rect -6356 -40872 -971 -40833
rect -6339 -40885 -6202 -40872
rect -3742 -40891 -3605 -40872
rect -1104 -40891 -972 -40872
rect -6687 -41033 -6627 -40896
rect -5950 -41011 -5818 -41003
rect -1427 -41011 -1295 -41001
rect -6686 -41391 -6638 -41033
rect -6356 -41050 -1295 -41011
rect -5950 -41063 -5818 -41050
rect -1427 -41061 -1295 -41050
rect -6568 -41165 -6034 -41097
rect -5637 -41120 -5004 -41086
rect -6567 -41308 -6533 -41216
rect -6573 -41369 -6527 -41308
rect -6469 -41324 -6435 -41165
rect -6371 -41308 -6337 -41216
rect -6603 -41391 -6527 -41369
rect -6686 -41401 -6527 -41391
rect -6377 -41401 -6331 -41308
rect -6273 -41324 -6239 -41165
rect -6175 -41308 -6141 -41216
rect -6181 -41401 -6135 -41308
rect -6077 -41324 -6043 -41165
rect -5729 -41260 -5695 -41166
rect -5637 -41178 -5593 -41120
rect -5733 -41303 -5692 -41260
rect -5631 -41274 -5597 -41178
rect -5533 -41261 -5499 -41166
rect -5440 -41189 -5396 -41120
rect -5734 -41310 -5692 -41303
rect -5536 -41310 -5495 -41261
rect -5435 -41274 -5401 -41189
rect -5337 -41261 -5303 -41166
rect -5244 -41189 -5200 -41120
rect -5342 -41310 -5301 -41261
rect -5239 -41274 -5205 -41189
rect -5141 -41269 -5107 -41166
rect -5048 -41178 -5004 -41120
rect -4825 -41165 -3334 -41097
rect -2937 -41120 -2304 -41086
rect -5043 -41248 -5009 -41178
rect -5144 -41310 -5103 -41269
rect -5734 -41344 -5103 -41310
rect -6686 -41428 -6135 -41401
rect -6685 -41430 -6135 -41428
rect -6603 -41439 -6135 -41430
rect -6099 -41373 -5931 -41358
rect -5734 -41373 -5559 -41344
rect -6099 -41426 -5559 -41373
rect -5050 -41383 -5003 -41248
rect -4824 -41308 -4790 -41216
rect -4830 -41369 -4784 -41308
rect -4726 -41324 -4692 -41165
rect -4628 -41308 -4594 -41216
rect -6099 -41432 -5931 -41426
rect -6573 -41447 -6135 -41439
rect -6573 -41512 -6527 -41447
rect -6567 -41704 -6533 -41512
rect -6377 -41512 -6331 -41447
rect -6371 -41704 -6337 -41512
rect -6181 -41700 -6135 -41447
rect -6175 -41704 -6141 -41700
rect -5734 -41511 -5559 -41426
rect -5175 -41457 -5003 -41383
rect -5734 -41545 -5106 -41511
rect -5734 -41589 -5692 -41545
rect -5729 -41689 -5695 -41589
rect -5631 -41672 -5597 -41581
rect -5534 -41599 -5498 -41545
rect -5340 -41581 -5304 -41545
rect -5636 -41723 -5594 -41672
rect -5533 -41689 -5499 -41599
rect -5435 -41667 -5401 -41581
rect -5340 -41599 -5303 -41581
rect -5440 -41723 -5398 -41667
rect -5337 -41689 -5303 -41599
rect -5239 -41668 -5205 -41581
rect -5142 -41597 -5106 -41545
rect -5246 -41723 -5204 -41668
rect -5141 -41689 -5107 -41597
rect -5050 -41604 -5003 -41457
rect -4958 -41401 -4784 -41369
rect -4634 -41401 -4588 -41308
rect -4530 -41324 -4496 -41165
rect -4432 -41308 -4398 -41216
rect -4438 -41401 -4392 -41308
rect -4334 -41324 -4300 -41165
rect -4958 -41439 -4392 -41401
rect -4013 -41380 -3953 -41265
rect -3867 -41308 -3833 -41216
rect -3873 -41369 -3827 -41308
rect -3769 -41324 -3735 -41165
rect -3671 -41308 -3637 -41216
rect -3903 -41380 -3827 -41369
rect -4018 -41401 -3827 -41380
rect -3677 -41401 -3631 -41308
rect -3573 -41324 -3539 -41165
rect -3475 -41308 -3441 -41216
rect -3481 -41401 -3435 -41308
rect -3377 -41324 -3343 -41165
rect -3032 -41260 -2986 -41138
rect -2937 -41178 -2893 -41120
rect -3033 -41270 -2986 -41260
rect -3033 -41303 -2992 -41270
rect -2931 -41274 -2897 -41178
rect -2833 -41261 -2799 -41166
rect -2740 -41189 -2696 -41120
rect -3034 -41310 -2992 -41303
rect -2836 -41310 -2795 -41261
rect -2735 -41274 -2701 -41189
rect -2637 -41261 -2603 -41166
rect -2544 -41189 -2500 -41120
rect -2642 -41310 -2601 -41261
rect -2539 -41274 -2505 -41189
rect -2441 -41269 -2407 -41166
rect -2348 -41178 -2304 -41120
rect -2125 -41165 -709 -41097
rect -2343 -41248 -2309 -41178
rect -2444 -41310 -2403 -41269
rect -3034 -41344 -2403 -41310
rect -4018 -41425 -3435 -41401
rect -4958 -41463 -4885 -41439
rect -5043 -41678 -5009 -41604
rect -4959 -41631 -4885 -41463
rect -4830 -41447 -4392 -41439
rect -4830 -41512 -4784 -41447
rect -5044 -41723 -5008 -41678
rect -4824 -41704 -4790 -41512
rect -5636 -41757 -5008 -41723
rect -4634 -41512 -4588 -41447
rect -4628 -41704 -4594 -41512
rect -4438 -41700 -4392 -41447
rect -4432 -41704 -4398 -41700
rect -4234 -41559 -4177 -41518
rect -4018 -41559 -3973 -41425
rect -3903 -41439 -3435 -41425
rect -3399 -41366 -3231 -41358
rect -3034 -41366 -2859 -41344
rect -3399 -41423 -2859 -41366
rect -2350 -41383 -2303 -41248
rect -2124 -41308 -2090 -41216
rect -2130 -41369 -2084 -41308
rect -2026 -41324 -1992 -41165
rect -1928 -41308 -1894 -41216
rect -3399 -41432 -3231 -41423
rect -3873 -41447 -3435 -41439
rect -3873 -41512 -3827 -41447
rect -4234 -41604 -3973 -41559
rect -4234 -41682 -4177 -41604
rect -3867 -41704 -3833 -41512
rect -3677 -41512 -3631 -41447
rect -3671 -41704 -3637 -41512
rect -3481 -41700 -3435 -41447
rect -3475 -41704 -3441 -41700
rect -3034 -41511 -2859 -41423
rect -2475 -41457 -2303 -41383
rect -3034 -41545 -2406 -41511
rect -3034 -41589 -2992 -41545
rect -3029 -41689 -2995 -41589
rect -2931 -41672 -2897 -41581
rect -2834 -41599 -2798 -41545
rect -2640 -41581 -2604 -41545
rect -2936 -41723 -2894 -41672
rect -2833 -41689 -2799 -41599
rect -2735 -41667 -2701 -41581
rect -2640 -41599 -2603 -41581
rect -2740 -41723 -2698 -41667
rect -2637 -41689 -2603 -41599
rect -2539 -41668 -2505 -41581
rect -2442 -41597 -2406 -41545
rect -2546 -41723 -2504 -41668
rect -2441 -41689 -2407 -41597
rect -2350 -41604 -2303 -41457
rect -2258 -41401 -2084 -41369
rect -1934 -41401 -1888 -41308
rect -1830 -41324 -1796 -41165
rect -1732 -41308 -1698 -41216
rect -1738 -41401 -1692 -41308
rect -1634 -41324 -1600 -41165
rect -2258 -41439 -1692 -41401
rect -1656 -41363 -1488 -41358
rect -1656 -41375 -1453 -41363
rect -1396 -41375 -1336 -41289
rect -1242 -41308 -1208 -41216
rect -1248 -41369 -1202 -41308
rect -1144 -41324 -1110 -41165
rect -1046 -41308 -1012 -41216
rect -1278 -41375 -1202 -41369
rect -1656 -41401 -1202 -41375
rect -1052 -41401 -1006 -41308
rect -948 -41324 -914 -41165
rect -850 -41308 -816 -41216
rect -856 -41401 -810 -41308
rect -752 -41324 -718 -41165
rect -312 -41224 -278 -40771
rect -214 -40979 -180 -40583
rect 199 -40673 640 -40639
rect 101 -41143 135 -40771
rect 199 -41079 233 -40673
rect 409 -40676 640 -40673
rect 297 -41143 331 -40771
rect 409 -40782 444 -40676
rect 410 -41079 444 -40782
rect 508 -41079 542 -40771
rect 605 -40780 640 -40676
rect 606 -41079 640 -40780
rect 507 -41142 542 -41079
rect 720 -41142 754 -40772
rect 818 -41080 852 -40583
rect 1682 -40733 1833 -40253
rect 2059 -40715 2183 -40253
rect 2389 -40715 2513 -40253
rect 2796 -40695 2932 -40649
rect 2059 -40733 2574 -40715
rect 507 -41143 754 -41142
rect 916 -41143 950 -40772
rect 101 -41177 334 -41143
rect 507 -41177 950 -41143
rect 1682 -40776 2574 -40733
rect 1682 -40794 2132 -40776
rect -463 -41277 -278 -41224
rect -1656 -41417 -810 -41401
rect -1656 -41421 -1453 -41417
rect -1396 -41421 -1336 -41417
rect -1656 -41432 -1488 -41421
rect -1278 -41439 -810 -41417
rect -2258 -41463 -2185 -41439
rect -2343 -41678 -2309 -41604
rect -2259 -41631 -2185 -41463
rect -2130 -41447 -1692 -41439
rect -2130 -41512 -2084 -41447
rect -2344 -41723 -2308 -41678
rect -2124 -41704 -2090 -41512
rect -2936 -41757 -2308 -41723
rect -1934 -41512 -1888 -41447
rect -1928 -41704 -1894 -41512
rect -1738 -41700 -1692 -41447
rect -1248 -41447 -810 -41439
rect -1732 -41704 -1698 -41700
rect -1248 -41512 -1202 -41447
rect -1534 -41682 -1477 -41518
rect -1242 -41704 -1208 -41512
rect -1052 -41512 -1006 -41447
rect -1046 -41704 -1012 -41512
rect -856 -41700 -810 -41447
rect -850 -41704 -816 -41700
rect -6898 -42127 -6762 -42081
rect -17491 -43112 -17356 -43106
rect -17511 -43114 -17356 -43112
rect -18573 -43139 -18443 -43122
rect -18399 -43139 -18326 -43126
rect -19108 -43145 -19050 -43144
rect -18573 -43145 -18326 -43139
rect -19108 -43180 -18326 -43145
rect -17718 -43150 -17356 -43114
rect -17308 -43129 -16878 -43099
rect -17308 -43137 -16889 -43129
rect -16699 -43141 -16665 -42985
rect -16601 -43093 -16567 -42985
rect -16503 -43141 -16469 -42985
rect -16405 -43093 -16371 -42985
rect -16307 -42996 -15935 -42926
rect -17511 -43152 -17356 -43150
rect -17491 -43160 -17356 -43152
rect -19108 -43213 -18443 -43180
rect -18399 -43186 -18326 -43180
rect -19108 -43281 -19050 -43213
rect -18573 -43272 -18443 -43213
rect -17986 -43210 -17437 -43208
rect -17026 -43210 -16952 -43184
rect -17986 -43214 -16952 -43210
rect -18281 -43470 -18247 -43214
rect -18183 -43422 -18149 -43214
rect -18085 -43470 -18051 -43214
rect -17987 -43248 -16952 -43214
rect -16839 -43227 -16054 -43141
rect -17987 -43422 -17953 -43248
rect -17438 -43249 -16952 -43248
rect -17438 -43250 -17367 -43249
rect -17026 -43255 -16952 -43249
rect -18421 -43556 -17483 -43470
rect -21289 -43684 -20060 -43646
rect -21289 -43693 -21154 -43684
rect -20953 -43730 -20818 -43721
rect -19193 -43730 -19135 -43633
rect -17569 -43637 -17483 -43556
rect -17406 -43600 -17372 -43292
rect -17308 -43600 -17274 -43292
rect -17210 -43600 -17176 -43292
rect -17112 -43600 -17078 -43292
rect -17014 -43600 -16980 -43292
rect -17309 -43637 -17274 -43600
rect -16595 -43634 -16534 -43227
rect -16984 -43637 -16534 -43634
rect -17569 -43695 -16534 -43637
rect -6858 -43658 -6824 -42127
rect -4418 -42200 -4282 -42154
rect -4418 -42453 -4378 -42200
rect -4421 -42589 -4375 -42453
rect -312 -41687 -278 -41277
rect -243 -41231 -108 -41224
rect 297 -41231 334 -41177
rect 1682 -41201 1743 -40794
rect 2422 -40828 2457 -40776
rect 2128 -41136 2162 -40828
rect 2226 -41136 2260 -40828
rect 2324 -41136 2358 -40828
rect 2422 -41136 2456 -40828
rect 2520 -41136 2554 -40828
rect 2100 -41179 2174 -41173
rect 2515 -41179 2586 -41178
rect 2100 -41180 2586 -41179
rect -243 -41268 334 -41231
rect -243 -41278 -108 -41268
rect 297 -41406 334 -41268
rect 368 -41233 503 -41226
rect 368 -41267 1324 -41233
rect 368 -41280 503 -41267
rect 556 -41311 691 -41304
rect 1119 -41311 1255 -41304
rect 556 -41349 1255 -41311
rect 556 -41358 691 -41349
rect 1119 -41350 1255 -41349
rect 297 -41443 852 -41406
rect 892 -41440 1084 -41386
rect 1290 -41432 1324 -41267
rect 1372 -41287 1987 -41201
rect 2100 -41218 2767 -41180
rect 2100 -41244 2174 -41218
rect 2585 -41220 2767 -41218
rect 2504 -41274 2639 -41268
rect 2504 -41278 2669 -41274
rect 426 -41687 460 -41443
rect 622 -41687 656 -41443
rect 818 -41687 852 -41443
rect 1038 -41524 1084 -41440
rect 1284 -41502 1455 -41432
rect 1519 -41443 1553 -41335
rect 1617 -41443 1651 -41287
rect 1715 -41443 1749 -41335
rect 1813 -41443 1847 -41287
rect 2037 -41299 2456 -41291
rect 2026 -41329 2456 -41299
rect 2504 -41314 2691 -41278
rect 2504 -41322 2682 -41314
rect 1421 -41674 1455 -41502
rect 1892 -41478 1965 -41472
rect 2026 -41478 2087 -41329
rect 1892 -41491 2087 -41478
rect 1892 -41519 2065 -41491
rect 1892 -41532 1965 -41519
rect 1617 -41674 1651 -41566
rect 1813 -41674 1847 -41566
rect 2226 -41673 2260 -41329
rect 2422 -41673 2456 -41329
rect 2646 -42072 2682 -41322
rect 2527 -42118 2682 -42072
rect 2727 -42156 2767 -41220
rect 2862 -41430 2932 -40695
rect 3287 -40731 3438 -40253
rect 3729 -40713 3880 -40253
rect 4022 -40713 4173 -40253
rect 4662 -40527 4808 -40253
rect 5107 -40527 5253 -40253
rect 5373 -40527 5519 -40253
rect 5733 -40527 5879 -40253
rect 4364 -40583 4500 -40537
rect 3729 -40731 4179 -40713
rect 3287 -40774 4179 -40731
rect 3287 -40792 3737 -40774
rect 3287 -41199 3348 -40792
rect 4027 -40826 4062 -40774
rect 3733 -41134 3767 -40826
rect 3831 -41134 3865 -40826
rect 3929 -41134 3963 -40826
rect 4027 -41134 4061 -40826
rect 4125 -41134 4159 -40826
rect 4434 -41038 4499 -40583
rect 4638 -40592 5912 -40527
rect 4650 -41038 4684 -40780
rect 4748 -40988 4782 -40592
rect 5161 -40682 5602 -40648
rect 4434 -41096 4684 -41038
rect 3705 -41177 3779 -41171
rect 4120 -41177 4191 -41176
rect 3705 -41178 4191 -41177
rect 2977 -41285 3592 -41199
rect 3705 -41216 4395 -41178
rect 3705 -41242 3779 -41216
rect 4190 -41218 4395 -41216
rect 4109 -41274 4244 -41266
rect 4109 -41276 4296 -41274
rect 2862 -41500 3060 -41430
rect 3124 -41441 3158 -41333
rect 3222 -41441 3256 -41285
rect 3320 -41441 3354 -41333
rect 3418 -41441 3452 -41285
rect 3642 -41297 4061 -41289
rect 3631 -41327 4061 -41297
rect 4109 -41314 4316 -41276
rect 4109 -41320 4244 -41314
rect 3026 -41672 3060 -41500
rect 3497 -41476 3570 -41470
rect 3631 -41476 3692 -41327
rect 3497 -41489 3692 -41476
rect 3497 -41517 3670 -41489
rect 3497 -41530 3570 -41517
rect 3222 -41672 3256 -41564
rect 3418 -41672 3452 -41564
rect 3831 -41671 3865 -41327
rect 4027 -41671 4061 -41327
rect 2631 -42202 2767 -42156
rect 4280 -42641 4316 -41314
rect 2795 -42677 4316 -42641
rect 2795 -42789 2831 -42677
rect 4355 -42711 4395 -41218
rect 4650 -41696 4684 -41096
rect 5063 -41152 5097 -40780
rect 5161 -41088 5195 -40682
rect 5371 -40685 5602 -40682
rect 5259 -41152 5293 -40780
rect 5371 -40791 5406 -40685
rect 5372 -41088 5406 -40791
rect 5470 -41088 5504 -40780
rect 5567 -40789 5602 -40685
rect 5568 -41088 5602 -40789
rect 5469 -41151 5504 -41088
rect 5682 -41151 5716 -40781
rect 5780 -41089 5814 -40592
rect 6297 -40707 6494 -40253
rect 6830 -40707 7027 -40253
rect 7343 -40698 7540 -40253
rect 7846 -40698 8043 -40253
rect 8241 -40680 8502 -40253
rect 9786 -40190 9850 -40167
rect 15151 -40190 15234 -39995
rect 16008 -40017 16229 -39995
rect 9786 -40273 15234 -40190
rect 9786 -40285 9850 -40273
rect 19091 -40351 19240 -37816
rect 19652 -38346 19836 -37816
rect 20276 -37850 20318 -37806
rect 20379 -37814 20413 -37723
rect 20477 -37796 20511 -37706
rect 20570 -37728 20612 -37672
rect 20476 -37850 20512 -37796
rect 20575 -37814 20609 -37728
rect 20673 -37796 20707 -37706
rect 20764 -37727 20806 -37672
rect 20670 -37814 20707 -37796
rect 20771 -37814 20805 -37727
rect 20869 -37798 20903 -37706
rect 20966 -37717 21002 -37672
rect 20967 -37791 21001 -37717
rect 20670 -37850 20706 -37814
rect 20868 -37850 20904 -37798
rect 20276 -37884 20904 -37850
rect 20276 -37993 20451 -37884
rect 20960 -37938 21007 -37791
rect 21051 -37932 21125 -37764
rect 21186 -37883 21220 -37691
rect 20201 -38051 20451 -37993
rect 20835 -38012 21007 -37938
rect 20201 -38053 20907 -38051
rect 20276 -38085 20907 -38053
rect 20276 -38092 20318 -38085
rect 20277 -38135 20318 -38092
rect 20281 -38229 20315 -38135
rect 20379 -38217 20413 -38121
rect 20474 -38134 20515 -38085
rect 20373 -38275 20417 -38217
rect 20477 -38229 20511 -38134
rect 20575 -38206 20609 -38121
rect 20668 -38134 20709 -38085
rect 20570 -38275 20614 -38206
rect 20673 -38229 20707 -38134
rect 20771 -38206 20805 -38121
rect 20866 -38126 20907 -38085
rect 20766 -38275 20810 -38206
rect 20869 -38229 20903 -38126
rect 20960 -38147 21007 -38012
rect 21052 -37956 21125 -37932
rect 21180 -37948 21226 -37883
rect 21382 -37883 21416 -37691
rect 21376 -37948 21422 -37883
rect 21578 -37695 21612 -37691
rect 21572 -37948 21618 -37695
rect 21776 -37765 21833 -37713
rect 21776 -37827 21981 -37765
rect 21776 -37877 21833 -37827
rect 21180 -37956 21618 -37948
rect 21052 -37994 21618 -37956
rect 21919 -37956 21981 -37827
rect 22023 -37883 22057 -37691
rect 22017 -37948 22063 -37883
rect 22219 -37883 22253 -37691
rect 22213 -37948 22259 -37883
rect 22415 -37695 22449 -37691
rect 22409 -37948 22455 -37695
rect 23074 -37672 23702 -37638
rect 22981 -37806 23015 -37706
rect 23074 -37723 23116 -37672
rect 22976 -37850 23018 -37806
rect 23079 -37814 23113 -37723
rect 23177 -37796 23211 -37706
rect 23270 -37728 23312 -37672
rect 23176 -37850 23212 -37796
rect 23275 -37814 23309 -37728
rect 23373 -37796 23407 -37706
rect 23464 -37727 23506 -37672
rect 23370 -37814 23407 -37796
rect 23471 -37814 23505 -37727
rect 23569 -37798 23603 -37706
rect 23666 -37717 23702 -37672
rect 23667 -37791 23701 -37717
rect 23370 -37850 23406 -37814
rect 23568 -37850 23604 -37798
rect 22976 -37884 23604 -37850
rect 22017 -37956 22455 -37948
rect 21052 -38026 21226 -37994
rect 21180 -38087 21226 -38026
rect 20967 -38217 21001 -38147
rect 21186 -38179 21220 -38087
rect 20962 -38275 21006 -38217
rect 21284 -38230 21318 -38071
rect 21376 -38087 21422 -37994
rect 21382 -38179 21416 -38087
rect 21480 -38230 21514 -38071
rect 21572 -38087 21618 -37994
rect 21919 -37994 22455 -37956
rect 21919 -38026 22063 -37994
rect 21578 -38179 21612 -38087
rect 21676 -38230 21710 -38071
rect 22017 -38087 22063 -38026
rect 22023 -38179 22057 -38087
rect 22121 -38230 22155 -38071
rect 22213 -38087 22259 -37994
rect 22219 -38179 22253 -38087
rect 22317 -38230 22351 -38071
rect 22409 -38087 22455 -37994
rect 22491 -37970 22659 -37963
rect 22491 -38030 22681 -37970
rect 22976 -37991 23151 -37884
rect 23660 -37938 23707 -37791
rect 23751 -37932 23825 -37764
rect 23886 -37883 23920 -37691
rect 22491 -38037 22659 -38030
rect 22885 -38051 23151 -37991
rect 23535 -38012 23707 -37938
rect 22415 -38179 22449 -38087
rect 22513 -38230 22547 -38071
rect 22976 -38085 23607 -38051
rect 22976 -38092 23018 -38085
rect 22977 -38135 23018 -38092
rect 22981 -38229 23015 -38135
rect 23079 -38217 23113 -38121
rect 23174 -38134 23215 -38085
rect 20373 -38309 21006 -38275
rect 21185 -38232 21719 -38230
rect 22022 -38232 22556 -38230
rect 21185 -38298 22556 -38232
rect 23073 -38275 23117 -38217
rect 23177 -38229 23211 -38134
rect 23275 -38206 23309 -38121
rect 23368 -38134 23409 -38085
rect 23270 -38275 23314 -38206
rect 23373 -38229 23407 -38134
rect 23471 -38206 23505 -38121
rect 23566 -38126 23607 -38085
rect 23466 -38275 23510 -38206
rect 23569 -38229 23603 -38126
rect 23660 -38147 23707 -38012
rect 23752 -37956 23825 -37932
rect 23880 -37948 23926 -37883
rect 24082 -37883 24116 -37691
rect 24076 -37948 24122 -37883
rect 24278 -37695 24312 -37691
rect 24272 -37948 24318 -37695
rect 24476 -37777 24533 -37713
rect 24476 -37826 24676 -37777
rect 24476 -37877 24533 -37826
rect 23880 -37956 24318 -37948
rect 23752 -37994 24318 -37956
rect 24630 -37956 24676 -37826
rect 24723 -37883 24757 -37691
rect 24717 -37948 24763 -37883
rect 24919 -37883 24953 -37691
rect 24913 -37948 24959 -37883
rect 25115 -37695 25149 -37691
rect 25109 -37948 25155 -37695
rect 28727 -37675 28761 -37331
rect 28923 -37675 28957 -37331
rect 29096 -37480 29157 -37331
rect 29336 -37445 29370 -37289
rect 29434 -37445 29468 -37337
rect 29532 -37445 29566 -37289
rect 35902 -37302 36149 -37261
rect 36984 -37289 37119 -37281
rect 36964 -37291 37119 -37289
rect 35902 -37319 36032 -37302
rect 36076 -37315 36149 -37302
rect 36757 -37327 37119 -37291
rect 37636 -37300 38421 -37214
rect 44765 -37300 44895 -37208
rect 45057 -37266 45091 -37010
rect 45155 -37266 45189 -37058
rect 45253 -37266 45287 -37010
rect 45351 -37232 45385 -37058
rect 45932 -37188 45966 -36880
rect 46030 -37188 46064 -36880
rect 46128 -37188 46162 -36880
rect 46226 -37188 46260 -36880
rect 46324 -37188 46358 -36880
rect 45900 -37231 45971 -37230
rect 46312 -37231 46386 -37225
rect 45900 -37232 46386 -37231
rect 45351 -37266 46386 -37232
rect 46743 -37253 46804 -36846
rect 51498 -36814 51724 -36805
rect 53151 -36814 53397 -36734
rect 51498 -36947 53397 -36814
rect 54967 -36751 55632 -36723
rect 54967 -36809 56002 -36751
rect 54967 -36890 55053 -36809
rect 55227 -36846 55262 -36809
rect 55552 -36812 56002 -36809
rect 51498 -37039 51724 -36947
rect 53151 -36954 53397 -36947
rect 54115 -36976 55053 -36890
rect 45352 -37270 46386 -37266
rect 45352 -37272 45901 -37270
rect 44939 -37300 45012 -37294
rect 46312 -37296 46386 -37270
rect 36964 -37329 37119 -37327
rect 36984 -37335 37119 -37329
rect 37167 -37312 37586 -37304
rect 29630 -37445 29664 -37337
rect 37167 -37342 37597 -37312
rect 29218 -37480 29291 -37474
rect 29096 -37493 29291 -37480
rect 29118 -37521 29291 -37493
rect 29218 -37534 29291 -37521
rect 29728 -37504 30100 -37434
rect 29336 -37676 29370 -37568
rect 29532 -37676 29566 -37568
rect 29728 -37676 29762 -37504
rect 24717 -37956 25155 -37948
rect 23752 -38026 23926 -37994
rect 23880 -38087 23926 -38026
rect 23667 -38217 23701 -38147
rect 23886 -38179 23920 -38087
rect 23662 -38275 23706 -38217
rect 23984 -38230 24018 -38071
rect 24076 -38087 24122 -37994
rect 24082 -38179 24116 -38087
rect 24180 -38230 24214 -38071
rect 24272 -38087 24318 -37994
rect 24354 -37974 24522 -37963
rect 24354 -37975 24557 -37974
rect 24354 -38037 24594 -37975
rect 24630 -37994 25155 -37956
rect 24630 -38026 24763 -37994
rect 24278 -38179 24312 -38087
rect 24376 -38230 24410 -38071
rect 24534 -38181 24594 -38037
rect 24717 -38087 24763 -38026
rect 24723 -38179 24757 -38087
rect 24821 -38230 24855 -38071
rect 24913 -38087 24959 -37994
rect 24919 -38179 24953 -38087
rect 25017 -38230 25051 -38071
rect 25109 -38087 25155 -37994
rect 25191 -37993 25359 -37963
rect 25191 -38037 25366 -37993
rect 25115 -38179 25149 -38087
rect 25213 -38230 25247 -38071
rect 21410 -38346 21521 -38298
rect 21696 -38300 22216 -38298
rect 22288 -38344 22399 -38298
rect 23073 -38309 23706 -38275
rect 23885 -38298 25256 -38230
rect 22285 -38346 22422 -38344
rect 24086 -38346 24197 -38298
rect 24897 -38338 25008 -38298
rect 24882 -38346 25019 -38338
rect 19651 -38385 25036 -38346
rect 19652 -38404 19784 -38385
rect 22285 -38404 22422 -38385
rect 24882 -38398 25019 -38385
rect 25318 -38409 25366 -38037
rect 19975 -38524 20107 -38514
rect 24498 -38524 24630 -38516
rect 19975 -38563 25036 -38524
rect 25307 -38546 25367 -38409
rect 19975 -38574 20107 -38563
rect 24498 -38576 24630 -38563
rect 19389 -38678 20805 -38610
rect 20984 -38633 21617 -38599
rect 19398 -38837 19432 -38678
rect 19496 -38821 19530 -38729
rect 19490 -38914 19536 -38821
rect 19594 -38837 19628 -38678
rect 19692 -38821 19726 -38729
rect 19686 -38914 19732 -38821
rect 19790 -38837 19824 -38678
rect 19888 -38821 19922 -38729
rect 19882 -38882 19928 -38821
rect 19882 -38888 19958 -38882
rect 20016 -38888 20076 -38802
rect 20280 -38837 20314 -38678
rect 20378 -38821 20412 -38729
rect 20168 -38876 20336 -38871
rect 20133 -38888 20336 -38876
rect 19882 -38914 20336 -38888
rect 19490 -38930 20336 -38914
rect 19490 -38952 19958 -38930
rect 20016 -38934 20076 -38930
rect 20133 -38934 20336 -38930
rect 20168 -38945 20336 -38934
rect 20372 -38914 20418 -38821
rect 20476 -38837 20510 -38678
rect 20574 -38821 20608 -38729
rect 20568 -38914 20614 -38821
rect 20672 -38837 20706 -38678
rect 20984 -38691 21028 -38633
rect 20770 -38821 20804 -38729
rect 20989 -38761 21023 -38691
rect 20764 -38882 20810 -38821
rect 20764 -38914 20938 -38882
rect 20372 -38952 20938 -38914
rect 19490 -38960 19928 -38952
rect 19490 -39213 19536 -38960
rect 19496 -39217 19530 -39213
rect 19686 -39025 19732 -38960
rect 19692 -39217 19726 -39025
rect 19882 -39025 19928 -38960
rect 20372 -38960 20810 -38952
rect 19888 -39217 19922 -39025
rect 20157 -39195 20214 -39031
rect 20372 -39213 20418 -38960
rect 20378 -39217 20412 -39213
rect 20568 -39025 20614 -38960
rect 20574 -39217 20608 -39025
rect 20764 -39025 20810 -38960
rect 20865 -38976 20938 -38952
rect 20983 -38896 21030 -38761
rect 21087 -38782 21121 -38679
rect 21180 -38702 21224 -38633
rect 21083 -38823 21124 -38782
rect 21185 -38787 21219 -38702
rect 21283 -38774 21317 -38679
rect 21376 -38702 21420 -38633
rect 21281 -38823 21322 -38774
rect 21381 -38787 21415 -38702
rect 21479 -38774 21513 -38679
rect 21573 -38691 21617 -38633
rect 21475 -38823 21516 -38774
rect 21577 -38787 21611 -38691
rect 21666 -38773 21712 -38651
rect 22014 -38678 23505 -38610
rect 23684 -38633 24317 -38599
rect 21666 -38783 21713 -38773
rect 21672 -38816 21713 -38783
rect 21672 -38823 21714 -38816
rect 21083 -38857 21714 -38823
rect 22023 -38837 22057 -38678
rect 22121 -38821 22155 -38729
rect 21539 -38879 21714 -38857
rect 21911 -38879 22079 -38871
rect 20983 -38970 21155 -38896
rect 21539 -38936 22079 -38879
rect 20770 -39217 20804 -39025
rect 20865 -39144 20939 -38976
rect 20983 -39117 21030 -38970
rect 21539 -39024 21714 -38936
rect 21911 -38945 22079 -38936
rect 22115 -38914 22161 -38821
rect 22219 -38837 22253 -38678
rect 22317 -38821 22351 -38729
rect 22311 -38914 22357 -38821
rect 22415 -38837 22449 -38678
rect 22513 -38821 22547 -38729
rect 22507 -38882 22553 -38821
rect 22507 -38893 22583 -38882
rect 22633 -38893 22693 -38778
rect 22980 -38837 23014 -38678
rect 23078 -38821 23112 -38729
rect 22507 -38914 22698 -38893
rect 22115 -38938 22698 -38914
rect 22115 -38952 22583 -38938
rect 22115 -38960 22553 -38952
rect 21086 -39058 21714 -39024
rect 21086 -39110 21122 -39058
rect 21284 -39094 21320 -39058
rect 20989 -39191 21023 -39117
rect 20988 -39236 21024 -39191
rect 21087 -39202 21121 -39110
rect 21185 -39181 21219 -39094
rect 21283 -39112 21320 -39094
rect 21184 -39236 21226 -39181
rect 21283 -39202 21317 -39112
rect 21381 -39180 21415 -39094
rect 21478 -39112 21514 -39058
rect 21378 -39236 21420 -39180
rect 21479 -39202 21513 -39112
rect 21577 -39185 21611 -39094
rect 21672 -39102 21714 -39058
rect 21574 -39236 21616 -39185
rect 21675 -39202 21709 -39102
rect 20988 -39270 21616 -39236
rect 22115 -39213 22161 -38960
rect 22121 -39217 22155 -39213
rect 22311 -39025 22357 -38960
rect 22317 -39217 22351 -39025
rect 22507 -39025 22553 -38960
rect 22513 -39217 22547 -39025
rect 22653 -39072 22698 -38938
rect 23072 -38914 23118 -38821
rect 23176 -38837 23210 -38678
rect 23274 -38821 23308 -38729
rect 23268 -38914 23314 -38821
rect 23372 -38837 23406 -38678
rect 23684 -38691 23728 -38633
rect 23470 -38821 23504 -38729
rect 23689 -38761 23723 -38691
rect 23464 -38882 23510 -38821
rect 23464 -38914 23638 -38882
rect 23072 -38952 23638 -38914
rect 23072 -38960 23510 -38952
rect 22857 -39072 22914 -39031
rect 22653 -39117 22914 -39072
rect 22857 -39195 22914 -39117
rect 23072 -39213 23118 -38960
rect 23078 -39217 23112 -39213
rect 23268 -39025 23314 -38960
rect 23274 -39217 23308 -39025
rect 23464 -39025 23510 -38960
rect 23565 -38976 23638 -38952
rect 23683 -38896 23730 -38761
rect 23787 -38782 23821 -38679
rect 23880 -38702 23924 -38633
rect 23783 -38823 23824 -38782
rect 23885 -38787 23919 -38702
rect 23983 -38774 24017 -38679
rect 24076 -38702 24120 -38633
rect 23981 -38823 24022 -38774
rect 24081 -38787 24115 -38702
rect 24179 -38774 24213 -38679
rect 24273 -38691 24317 -38633
rect 24714 -38678 25248 -38610
rect 24175 -38823 24216 -38774
rect 24277 -38787 24311 -38691
rect 24375 -38773 24409 -38679
rect 24372 -38816 24413 -38773
rect 24372 -38823 24414 -38816
rect 23783 -38857 24414 -38823
rect 24723 -38837 24757 -38678
rect 24821 -38821 24855 -38729
rect 24239 -38886 24414 -38857
rect 24611 -38886 24779 -38871
rect 23683 -38970 23855 -38896
rect 24239 -38939 24779 -38886
rect 23470 -39217 23504 -39025
rect 23565 -39144 23639 -38976
rect 23683 -39117 23730 -38970
rect 24239 -39024 24414 -38939
rect 24611 -38945 24779 -38939
rect 24815 -38914 24861 -38821
rect 24919 -38837 24953 -38678
rect 25017 -38821 25051 -38729
rect 25011 -38914 25057 -38821
rect 25115 -38837 25149 -38678
rect 25213 -38821 25247 -38729
rect 25207 -38882 25253 -38821
rect 25207 -38904 25283 -38882
rect 25318 -38904 25366 -38546
rect 25207 -38914 25366 -38904
rect 24815 -38941 25366 -38914
rect 24815 -38943 25365 -38941
rect 24815 -38952 25283 -38943
rect 24815 -38960 25253 -38952
rect 23786 -39058 24414 -39024
rect 23786 -39110 23822 -39058
rect 23984 -39094 24020 -39058
rect 23689 -39191 23723 -39117
rect 23688 -39236 23724 -39191
rect 23787 -39202 23821 -39110
rect 23885 -39181 23919 -39094
rect 23983 -39112 24020 -39094
rect 23884 -39236 23926 -39181
rect 23983 -39202 24017 -39112
rect 24081 -39180 24115 -39094
rect 24178 -39112 24214 -39058
rect 24078 -39236 24120 -39180
rect 24179 -39202 24213 -39112
rect 24277 -39185 24311 -39094
rect 24372 -39102 24414 -39058
rect 24274 -39236 24316 -39185
rect 24375 -39202 24409 -39102
rect 23688 -39270 24316 -39236
rect 24815 -39213 24861 -38960
rect 24821 -39217 24855 -39213
rect 25011 -39025 25057 -38960
rect 25017 -39217 25051 -39025
rect 25207 -39025 25253 -38960
rect 25213 -39217 25247 -39025
rect 27728 -38611 27762 -38267
rect 27924 -38611 27958 -38267
rect 28337 -38374 28371 -38266
rect 28533 -38374 28567 -38266
rect 28219 -38421 28292 -38408
rect 28119 -38449 28292 -38421
rect 28097 -38462 28292 -38449
rect 28097 -38611 28158 -38462
rect 28219 -38468 28292 -38462
rect 28729 -38438 28763 -38266
rect 27728 -38641 28158 -38611
rect 27728 -38649 28147 -38641
rect 28337 -38653 28371 -38497
rect 28435 -38605 28469 -38497
rect 28533 -38653 28567 -38497
rect 28631 -38605 28665 -38497
rect 28729 -38508 29007 -38438
rect 27372 -38722 27599 -38720
rect 28010 -38722 28084 -38696
rect 27372 -38760 28084 -38722
rect 28197 -38739 28812 -38653
rect 21421 -39571 21581 -39439
rect 21428 -39754 21563 -39571
rect 21418 -39886 21578 -39754
rect 21941 -40205 21975 -39761
rect 22137 -40205 22171 -39761
rect 22379 -39693 25303 -39596
rect 21941 -40206 22171 -40205
rect 21315 -40219 21447 -40209
rect 21758 -40218 21893 -40212
rect 21738 -40219 21893 -40218
rect 21315 -40255 21893 -40219
rect 21941 -40243 22185 -40206
rect 21315 -40269 21447 -40255
rect 21738 -40258 21893 -40255
rect 21758 -40266 21893 -40258
rect 22151 -40278 22185 -40243
rect 22281 -40278 22341 -40218
rect 19886 -40351 21482 -40308
rect 18037 -40373 21482 -40351
rect 21668 -40311 21827 -40310
rect 21668 -40316 21828 -40311
rect 21976 -40316 22111 -40310
rect 21668 -40355 22111 -40316
rect 21668 -40356 21882 -40355
rect 21668 -40369 21828 -40356
rect 21976 -40364 22111 -40355
rect 22151 -40339 22341 -40278
rect 21668 -40370 21827 -40369
rect 18037 -40440 20066 -40373
rect 9465 -40494 9524 -40487
rect 9465 -40577 13441 -40494
rect 9465 -40582 9524 -40577
rect 7343 -40707 8092 -40698
rect 6259 -40760 8092 -40707
rect 5469 -41152 5716 -41151
rect 5878 -41152 5912 -40781
rect 6259 -40883 6298 -40760
rect 7460 -40794 8092 -40760
rect 6361 -40834 7369 -40798
rect 6263 -41072 6297 -40883
rect 5063 -41186 5296 -41152
rect 5469 -41186 5912 -41152
rect 6261 -41155 6298 -41072
rect 6361 -41079 6395 -40834
rect 6677 -41073 6711 -40871
rect 6775 -41070 6809 -40871
rect 7039 -41070 7073 -40871
rect 6674 -41094 6711 -41073
rect 6555 -41131 6711 -41094
rect 6773 -41109 7073 -41070
rect 6555 -41155 6592 -41131
rect 4719 -41240 4854 -41233
rect 5259 -41240 5296 -41186
rect 6261 -41192 6592 -41155
rect 7137 -41162 7171 -40871
rect 7333 -40888 7369 -40834
rect 7333 -41079 7367 -40888
rect 7431 -41162 7465 -40871
rect 7643 -41062 7677 -40871
rect 7736 -40878 7779 -40794
rect 7638 -41107 7681 -41062
rect 7741 -41079 7775 -40878
rect 7952 -41060 7986 -40871
rect 8045 -40880 8088 -40794
rect 7542 -41153 7681 -41107
rect 6904 -41196 7465 -41162
rect 4719 -41277 5296 -41240
rect 4719 -41287 4854 -41277
rect 5259 -41415 5296 -41277
rect 5330 -41242 5465 -41235
rect 5330 -41276 6149 -41242
rect 6904 -41258 6938 -41196
rect 5330 -41289 5465 -41276
rect 5518 -41320 5653 -41313
rect 5518 -41358 6079 -41320
rect 5518 -41367 5653 -41358
rect 5853 -41404 5989 -41395
rect 5259 -41452 5814 -41415
rect 5853 -41441 6008 -41404
rect 5854 -41449 5989 -41441
rect 5388 -41696 5422 -41452
rect 5584 -41696 5618 -41452
rect 5780 -41696 5814 -41452
rect -1621 -42825 2831 -42789
rect 2893 -42745 4395 -42711
rect 6045 -42727 6079 -41358
rect -1621 -42873 -1572 -42825
rect 789 -42869 925 -42860
rect 2893 -42869 2927 -42745
rect 5739 -42761 6079 -42727
rect 2972 -42800 3108 -42797
rect 5739 -42800 5773 -42761
rect 2972 -42834 5773 -42800
rect 5877 -42819 6013 -42813
rect 6115 -42819 6149 -41276
rect 6262 -41327 6401 -41273
rect 6792 -41292 6938 -41258
rect 6792 -41407 6826 -41292
rect 7011 -41297 7150 -41243
rect 6212 -41441 6826 -41407
rect 6887 -41368 7367 -41334
rect 6263 -41789 6297 -41477
rect 6361 -41685 6395 -41441
rect 6459 -41789 6493 -41477
rect 6579 -41720 6613 -41477
rect 6677 -41685 6711 -41441
rect 6775 -41720 6809 -41477
rect 6887 -41720 6921 -41368
rect 6579 -41754 6921 -41720
rect 6957 -41442 7171 -41408
rect 6957 -41789 6991 -41442
rect 7137 -41685 7171 -41442
rect 6263 -41823 6991 -41789
rect 7333 -41685 7367 -41368
rect 7420 -41371 7559 -41317
rect 7638 -41492 7681 -41153
rect 7948 -41251 7991 -41060
rect 8050 -41079 8084 -40880
rect 8241 -40941 9396 -40680
rect 12778 -40766 13063 -40708
rect 13358 -40766 13441 -40577
rect 18166 -40592 18210 -40440
rect 18170 -40751 18204 -40592
rect 18268 -40742 18302 -40543
rect 18360 -40591 18404 -40440
rect 12778 -40794 17738 -40766
rect 18076 -40794 18222 -40786
rect 12778 -40830 18222 -40794
rect 18263 -40791 18308 -40742
rect 18366 -40751 18400 -40591
rect 19112 -40592 19156 -40440
rect 19116 -40751 19150 -40592
rect 19214 -40742 19248 -40543
rect 19306 -40591 19350 -40440
rect 18263 -40792 18657 -40791
rect 18263 -40827 18706 -40792
rect 19022 -40794 19168 -40786
rect 12778 -40860 17738 -40830
rect 18076 -40846 18222 -40830
rect 18518 -40836 18706 -40827
rect 18963 -40830 19168 -40794
rect 19209 -40791 19254 -40742
rect 19312 -40751 19346 -40591
rect 19209 -40827 19879 -40791
rect 18574 -40852 18706 -40836
rect 19022 -40846 19168 -40830
rect 19464 -40836 19879 -40827
rect 12778 -40927 13063 -40860
rect 18299 -40883 18442 -40866
rect 17841 -40919 18442 -40883
rect 7848 -41297 7991 -41251
rect 7643 -41685 7677 -41492
rect 7948 -41494 7991 -41297
rect 8035 -41365 8174 -41311
rect 7952 -41685 7986 -41494
rect 2972 -42843 3108 -42834
rect 5877 -42853 6149 -42819
rect 5877 -42859 6013 -42853
rect -1708 -42919 -1572 -42873
rect 756 -42903 2927 -42869
rect 789 -42906 925 -42903
rect 8241 -42936 8502 -40941
rect -5550 -42958 -4918 -42949
rect -3050 -42958 -2418 -42949
rect -550 -42958 82 -42949
rect 1950 -42958 2582 -42949
rect 4450 -42958 5082 -42949
rect 7434 -42958 8502 -42936
rect -6751 -42959 -4918 -42958
rect -4251 -42959 8502 -42958
rect -6751 -43011 8502 -42959
rect -6751 -43134 -6712 -43011
rect -5550 -43045 -4212 -43011
rect -3050 -43045 -2418 -43011
rect -6649 -43085 -5641 -43049
rect -6747 -43323 -6713 -43134
rect -6749 -43406 -6712 -43323
rect -6649 -43330 -6615 -43085
rect -6333 -43324 -6299 -43122
rect -6235 -43321 -6201 -43122
rect -5971 -43321 -5937 -43122
rect -6336 -43345 -6299 -43324
rect -6455 -43382 -6299 -43345
rect -6237 -43360 -5937 -43321
rect -6455 -43406 -6418 -43382
rect -6749 -43443 -6418 -43406
rect -5873 -43413 -5839 -43122
rect -5677 -43139 -5641 -43085
rect -5677 -43330 -5643 -43139
rect -5579 -43413 -5545 -43122
rect -5367 -43313 -5333 -43122
rect -5274 -43129 -5231 -43045
rect -5039 -43046 -4212 -43045
rect -5372 -43358 -5329 -43313
rect -5269 -43330 -5235 -43129
rect -5058 -43311 -5024 -43122
rect -4965 -43131 -4922 -43046
rect -5468 -43404 -5329 -43358
rect -6106 -43447 -5545 -43413
rect -6106 -43509 -6072 -43447
rect -6748 -43578 -6609 -43524
rect -6218 -43543 -6072 -43509
rect -6218 -43658 -6184 -43543
rect -5999 -43548 -5860 -43494
rect -6858 -43692 -6184 -43658
rect -6123 -43619 -5643 -43585
rect -17569 -43723 -16904 -43695
rect -21548 -43778 -20993 -43741
rect -20953 -43765 -19135 -43730
rect -20953 -43767 -20799 -43765
rect -20953 -43775 -20818 -43767
rect -19193 -43770 -19135 -43765
rect -21419 -44022 -21385 -43778
rect -21223 -44022 -21189 -43778
rect -21027 -44022 -20993 -43778
rect -8448 -43886 -8248 -43862
rect -18829 -44022 -8248 -43886
rect -8448 -44033 -8248 -44022
rect -6747 -44040 -6713 -43728
rect -6649 -43936 -6615 -43692
rect -6551 -44040 -6517 -43728
rect -6431 -43971 -6397 -43728
rect -6333 -43936 -6299 -43692
rect -6235 -43971 -6201 -43728
rect -6123 -43971 -6089 -43619
rect -6431 -44005 -6089 -43971
rect -6053 -43693 -5839 -43659
rect -6053 -44040 -6019 -43693
rect -6747 -44074 -6019 -44040
rect -5873 -43936 -5839 -43693
rect -5677 -43936 -5643 -43619
rect -5590 -43622 -5451 -43568
rect -5372 -43743 -5329 -43404
rect -5062 -43502 -5019 -43311
rect -4960 -43330 -4926 -43131
rect -4251 -43134 -4212 -43046
rect -4149 -43085 -3141 -43049
rect -4421 -43295 -4375 -43159
rect -5162 -43548 -5019 -43502
rect -5367 -43936 -5333 -43743
rect -5062 -43745 -5019 -43548
rect -4975 -43616 -4836 -43562
rect -5058 -43936 -5024 -43745
rect -7311 -44140 -7148 -44120
rect -26388 -44360 -23542 -44174
rect -19006 -44276 -7148 -44140
rect -4415 -43658 -4381 -43295
rect -4247 -43323 -4213 -43134
rect -4249 -43406 -4212 -43323
rect -4149 -43330 -4115 -43085
rect -3833 -43324 -3799 -43122
rect -3735 -43321 -3701 -43122
rect -3471 -43321 -3437 -43122
rect -3836 -43345 -3799 -43324
rect -3955 -43382 -3799 -43345
rect -3737 -43360 -3437 -43321
rect -3955 -43406 -3918 -43382
rect -4249 -43443 -3918 -43406
rect -3373 -43413 -3339 -43122
rect -3177 -43139 -3141 -43085
rect -3177 -43330 -3143 -43139
rect -3079 -43413 -3045 -43122
rect -2867 -43313 -2833 -43122
rect -2774 -43129 -2731 -43045
rect -2872 -43358 -2829 -43313
rect -2769 -43330 -2735 -43129
rect -2558 -43311 -2524 -43122
rect -2465 -43131 -2422 -43045
rect -2968 -43404 -2829 -43358
rect -3866 -43474 -3727 -43420
rect -3606 -43447 -3045 -43413
rect -3606 -43509 -3572 -43447
rect -4248 -43578 -4109 -43524
rect -3718 -43543 -3572 -43509
rect -3718 -43658 -3684 -43543
rect -3499 -43548 -3360 -43494
rect -4415 -43692 -3684 -43658
rect -3623 -43619 -3143 -43585
rect -4247 -44040 -4213 -43728
rect -4149 -43936 -4115 -43692
rect -4051 -44040 -4017 -43728
rect -3931 -43971 -3897 -43728
rect -3833 -43936 -3799 -43692
rect -3735 -43971 -3701 -43728
rect -3623 -43971 -3589 -43619
rect -3931 -44005 -3589 -43971
rect -3553 -43693 -3339 -43659
rect -3553 -44040 -3519 -43693
rect -4247 -44074 -3519 -44040
rect -3373 -43936 -3339 -43693
rect -3177 -43936 -3143 -43619
rect -3090 -43622 -2951 -43568
rect -2872 -43743 -2829 -43404
rect -2788 -43468 -2649 -43414
rect -2562 -43502 -2519 -43311
rect -2460 -43330 -2426 -43131
rect -1751 -43134 -1712 -43011
rect -550 -43045 82 -43011
rect -1649 -43085 -641 -43049
rect -2662 -43548 -2519 -43502
rect -2867 -43936 -2833 -43743
rect -2562 -43745 -2519 -43548
rect -2475 -43616 -2336 -43562
rect -2558 -43936 -2524 -43745
rect -1873 -43291 -1827 -43155
rect -1867 -43658 -1833 -43291
rect -1747 -43323 -1713 -43134
rect -1749 -43406 -1712 -43323
rect -1649 -43330 -1615 -43085
rect -1333 -43324 -1299 -43122
rect -1235 -43321 -1201 -43122
rect -971 -43321 -937 -43122
rect -1336 -43345 -1299 -43324
rect -1455 -43382 -1299 -43345
rect -1237 -43360 -937 -43321
rect -1455 -43406 -1418 -43382
rect -1749 -43443 -1418 -43406
rect -873 -43413 -839 -43122
rect -677 -43139 -641 -43085
rect -677 -43330 -643 -43139
rect -579 -43413 -545 -43122
rect -367 -43313 -333 -43122
rect -274 -43129 -231 -43045
rect -372 -43358 -329 -43313
rect -269 -43330 -235 -43129
rect -58 -43311 -24 -43122
rect 35 -43131 78 -43045
rect -468 -43404 -329 -43358
rect -1366 -43474 -1227 -43420
rect -1106 -43447 -545 -43413
rect -1106 -43509 -1072 -43447
rect -1748 -43578 -1609 -43524
rect -1218 -43543 -1072 -43509
rect -1218 -43658 -1184 -43543
rect -999 -43548 -860 -43494
rect -1867 -43692 -1184 -43658
rect -1123 -43619 -643 -43585
rect -1747 -44040 -1713 -43728
rect -1649 -43936 -1615 -43692
rect -1551 -44040 -1517 -43728
rect -1431 -43971 -1397 -43728
rect -1333 -43936 -1299 -43692
rect -1235 -43971 -1201 -43728
rect -1123 -43971 -1089 -43619
rect -1431 -44005 -1089 -43971
rect -1053 -43693 -839 -43659
rect -1053 -44040 -1019 -43693
rect -1747 -44074 -1019 -44040
rect -873 -43936 -839 -43693
rect -677 -43936 -643 -43619
rect -590 -43622 -451 -43568
rect -372 -43743 -329 -43404
rect -288 -43468 -149 -43414
rect -62 -43502 -19 -43311
rect 40 -43330 74 -43131
rect 749 -43134 788 -43011
rect 1950 -43045 2582 -43011
rect 851 -43085 1859 -43049
rect -162 -43548 -19 -43502
rect -367 -43936 -333 -43743
rect -62 -43745 -19 -43548
rect 25 -43616 164 -43562
rect -58 -43936 -24 -43745
rect 607 -43291 653 -43155
rect 613 -43658 647 -43291
rect 753 -43323 787 -43134
rect 751 -43406 788 -43323
rect 851 -43330 885 -43085
rect 1167 -43324 1201 -43122
rect 1265 -43321 1299 -43122
rect 1529 -43321 1563 -43122
rect 1164 -43345 1201 -43324
rect 1045 -43382 1201 -43345
rect 1263 -43360 1563 -43321
rect 1045 -43406 1082 -43382
rect 751 -43443 1082 -43406
rect 1627 -43413 1661 -43122
rect 1823 -43139 1859 -43085
rect 1823 -43330 1857 -43139
rect 1921 -43413 1955 -43122
rect 2133 -43313 2167 -43122
rect 2226 -43129 2269 -43045
rect 2128 -43358 2171 -43313
rect 2231 -43330 2265 -43129
rect 2442 -43311 2476 -43122
rect 2535 -43131 2578 -43045
rect 2032 -43404 2171 -43358
rect 1134 -43474 1273 -43420
rect 1394 -43447 1955 -43413
rect 1394 -43509 1428 -43447
rect 752 -43578 891 -43524
rect 1282 -43543 1428 -43509
rect 1282 -43658 1316 -43543
rect 1501 -43548 1640 -43494
rect 613 -43692 1316 -43658
rect 1377 -43619 1857 -43585
rect 613 -43693 647 -43692
rect 753 -44040 787 -43728
rect 851 -43936 885 -43692
rect 949 -44040 983 -43728
rect 1069 -43971 1103 -43728
rect 1167 -43936 1201 -43692
rect 1265 -43971 1299 -43728
rect 1377 -43971 1411 -43619
rect 1069 -44005 1411 -43971
rect 1447 -43693 1661 -43659
rect 1447 -44040 1481 -43693
rect 753 -44074 1481 -44040
rect 1627 -43936 1661 -43693
rect 1823 -43936 1857 -43619
rect 1910 -43622 2049 -43568
rect 2128 -43743 2171 -43404
rect 2212 -43468 2351 -43414
rect 2438 -43502 2481 -43311
rect 2540 -43330 2574 -43131
rect 3249 -43134 3288 -43011
rect 4450 -43045 5082 -43011
rect 3351 -43085 4359 -43049
rect 3024 -43291 3070 -43155
rect 3029 -43292 3064 -43291
rect 2338 -43548 2481 -43502
rect 2133 -43936 2167 -43743
rect 2438 -43745 2481 -43548
rect 2525 -43616 2664 -43562
rect 3029 -43658 3063 -43292
rect 3253 -43323 3287 -43134
rect 3251 -43406 3288 -43323
rect 3351 -43330 3385 -43085
rect 3667 -43324 3701 -43122
rect 3765 -43321 3799 -43122
rect 4029 -43321 4063 -43122
rect 3664 -43345 3701 -43324
rect 3545 -43382 3701 -43345
rect 3763 -43360 4063 -43321
rect 3545 -43406 3582 -43382
rect 3251 -43443 3582 -43406
rect 4127 -43413 4161 -43122
rect 4323 -43139 4359 -43085
rect 4323 -43330 4357 -43139
rect 4421 -43413 4455 -43122
rect 4633 -43313 4667 -43122
rect 4726 -43129 4769 -43045
rect 4628 -43358 4671 -43313
rect 4731 -43330 4765 -43129
rect 4942 -43311 4976 -43122
rect 5035 -43131 5078 -43045
rect 4532 -43404 4671 -43358
rect 3894 -43447 4455 -43413
rect 3894 -43509 3928 -43447
rect 3252 -43578 3391 -43524
rect 3782 -43543 3928 -43509
rect 3782 -43658 3816 -43543
rect 4001 -43548 4140 -43494
rect 3029 -43692 3816 -43658
rect 3877 -43619 4357 -43585
rect 2442 -43936 2476 -43745
rect 3253 -44040 3287 -43728
rect 3351 -43936 3385 -43692
rect 3449 -44040 3483 -43728
rect 3569 -43971 3603 -43728
rect 3667 -43936 3701 -43692
rect 3765 -43971 3799 -43728
rect 3877 -43971 3911 -43619
rect 3569 -44005 3911 -43971
rect 3947 -43693 4161 -43659
rect 3947 -44040 3981 -43693
rect 3253 -44074 3981 -44040
rect 4127 -43936 4161 -43693
rect 4323 -43936 4357 -43619
rect 4410 -43622 4549 -43568
rect 4628 -43743 4671 -43404
rect 4938 -43502 4981 -43311
rect 5040 -43330 5074 -43131
rect 6249 -43134 6288 -43011
rect 6351 -43085 7359 -43049
rect 7434 -43063 8502 -43011
rect 5929 -43291 5975 -43155
rect 4838 -43548 4981 -43502
rect 4633 -43936 4667 -43743
rect 4938 -43745 4981 -43548
rect 5025 -43616 5164 -43562
rect 5935 -43658 5969 -43291
rect 6253 -43323 6287 -43134
rect 6251 -43406 6288 -43323
rect 6351 -43330 6385 -43085
rect 6667 -43324 6701 -43122
rect 6765 -43321 6799 -43122
rect 7029 -43321 7063 -43122
rect 6664 -43345 6701 -43324
rect 6545 -43382 6701 -43345
rect 6763 -43360 7063 -43321
rect 6545 -43406 6582 -43382
rect 6251 -43443 6582 -43406
rect 7127 -43413 7161 -43122
rect 7323 -43139 7359 -43085
rect 7323 -43330 7357 -43139
rect 7421 -43413 7455 -43122
rect 7633 -43313 7667 -43122
rect 7726 -43129 7769 -43063
rect 7628 -43358 7671 -43313
rect 7731 -43330 7765 -43129
rect 7942 -43311 7976 -43122
rect 8035 -43131 8078 -43063
rect 7532 -43404 7671 -43358
rect 6894 -43447 7455 -43413
rect 6894 -43509 6928 -43447
rect 6252 -43578 6391 -43524
rect 6782 -43543 6928 -43509
rect 6782 -43658 6816 -43543
rect 7001 -43548 7140 -43494
rect 5935 -43692 6816 -43658
rect 6877 -43619 7357 -43585
rect 4942 -43936 4976 -43745
rect 6253 -44040 6287 -43728
rect 6351 -43936 6385 -43692
rect 6449 -44040 6483 -43728
rect 6569 -43971 6603 -43728
rect 6667 -43936 6701 -43692
rect 6765 -43971 6799 -43728
rect 6877 -43971 6911 -43619
rect 6569 -44005 6911 -43971
rect 6947 -43693 7161 -43659
rect 6947 -44040 6981 -43693
rect 6253 -44074 6981 -44040
rect 7127 -43936 7161 -43693
rect 7323 -43936 7357 -43619
rect 7410 -43622 7549 -43568
rect 7628 -43743 7671 -43404
rect 7938 -43502 7981 -43311
rect 8040 -43330 8074 -43131
rect 7838 -43548 7981 -43502
rect 7633 -43936 7667 -43743
rect 7938 -43745 7981 -43548
rect 8025 -43616 8164 -43562
rect 7942 -43936 7976 -43745
rect -19006 -44277 -18868 -44276
rect -22212 -44322 -22054 -44289
rect -7311 -44295 -7148 -44276
rect -19144 -44322 -19007 -44317
rect -22212 -44374 -19007 -44322
rect -22212 -44405 -22054 -44374
rect -19144 -44375 -19007 -44374
rect 9135 -41735 9396 -40941
rect 17841 -40972 17877 -40919
rect 18299 -40926 18442 -40919
rect 13760 -41134 17877 -40972
rect 18169 -41001 18517 -40965
rect 9618 -41297 9687 -41279
rect 14831 -41297 14942 -41134
rect 9618 -41408 14942 -41297
rect 9618 -41418 9687 -41408
rect 18169 -41040 18205 -41001
rect 18170 -41443 18204 -41040
rect 18381 -41415 18415 -41035
rect 18472 -41045 18517 -41001
rect 18374 -41479 18420 -41415
rect 18479 -41443 18513 -41045
rect 18574 -41081 18624 -40852
rect 19245 -40883 19388 -40866
rect 18962 -40919 19388 -40883
rect 19245 -40926 19388 -40919
rect 19115 -41001 19463 -40965
rect 18577 -41415 18611 -41081
rect 18572 -41479 18618 -41415
rect 19115 -41040 19151 -41001
rect 18374 -41517 18618 -41479
rect 19116 -41443 19150 -41040
rect 19327 -41415 19361 -41035
rect 19418 -41045 19463 -41001
rect 19320 -41479 19366 -41415
rect 19425 -41443 19459 -41045
rect 19520 -41081 19570 -40836
rect 19523 -41415 19557 -41081
rect 19610 -41101 19670 -40935
rect 19845 -41023 19879 -40836
rect 19934 -40933 19968 -40562
rect 20032 -40870 20066 -40440
rect 20244 -40463 20685 -40429
rect 20244 -40466 20475 -40463
rect 20130 -40932 20164 -40562
rect 20244 -40570 20279 -40466
rect 20244 -40869 20278 -40570
rect 20342 -40869 20376 -40561
rect 20440 -40572 20475 -40466
rect 20440 -40869 20474 -40572
rect 20342 -40932 20377 -40869
rect 20130 -40933 20377 -40932
rect 20553 -40933 20587 -40561
rect 20651 -40869 20685 -40463
rect 20749 -40933 20783 -40561
rect 21064 -40769 21098 -40373
rect 21166 -40389 21482 -40373
rect 21166 -40424 21481 -40389
rect 19934 -40967 20377 -40933
rect 20550 -40967 20783 -40933
rect 21162 -40954 21196 -40561
rect 21400 -40730 21481 -40424
rect 21843 -40727 21877 -40415
rect 21941 -40643 21975 -40415
rect 22053 -40643 22087 -40415
rect 22151 -40623 22185 -40339
rect 22281 -40352 22341 -40339
rect 21941 -40678 22087 -40643
rect 21810 -40730 22289 -40727
rect 22379 -40730 22449 -39693
rect 21400 -40888 22449 -40730
rect 21784 -40931 22449 -40888
rect 22506 -40572 22576 -39838
rect 22673 -40514 22707 -39693
rect 22771 -40570 22805 -39806
rect 23073 -40514 23107 -39693
rect 23003 -40570 23137 -40557
rect 22506 -40626 22735 -40572
rect 22771 -40604 23137 -40570
rect 20381 -41023 20516 -41016
rect 19840 -41057 20516 -41023
rect 20381 -41070 20516 -41057
rect 20550 -41021 20587 -40967
rect 21162 -40990 21439 -40954
rect 20992 -41021 21127 -41014
rect 20550 -41058 21127 -41021
rect 20193 -41101 20328 -41094
rect 19610 -41139 20328 -41101
rect 20193 -41148 20328 -41139
rect 19857 -41185 19992 -41176
rect 19725 -41220 19992 -41185
rect 20550 -41196 20587 -41058
rect 20992 -41068 21127 -41058
rect 19725 -41317 19785 -41220
rect 19838 -41222 19992 -41220
rect 19857 -41230 19992 -41222
rect 20032 -41233 20587 -41196
rect 19518 -41479 19564 -41415
rect 19320 -41517 19564 -41479
rect 20032 -41477 20066 -41233
rect 20228 -41477 20262 -41233
rect 20424 -41477 20458 -41233
rect 21162 -41477 21196 -40990
rect 21308 -41014 21439 -40990
rect 21793 -41090 21827 -40931
rect 21891 -41074 21925 -40982
rect 21681 -41198 21849 -41124
rect 21885 -41167 21931 -41074
rect 21989 -41090 22023 -40931
rect 22087 -41074 22121 -40982
rect 22081 -41167 22127 -41074
rect 22185 -41090 22219 -40931
rect 22283 -41074 22317 -40982
rect 22277 -41135 22323 -41074
rect 22506 -41135 22576 -40626
rect 22277 -41167 22576 -41135
rect 21885 -41205 22576 -41167
rect 21885 -41213 22323 -41205
rect 21885 -41466 21931 -41213
rect 21891 -41470 21925 -41466
rect 22081 -41278 22127 -41213
rect 22087 -41470 22121 -41278
rect 22277 -41278 22323 -41213
rect 22283 -41470 22317 -41278
rect 22771 -41399 22805 -40604
rect 23003 -40611 23137 -40604
rect 23171 -40560 23205 -39806
rect 23279 -40560 23397 -40548
rect 23171 -40594 23397 -40560
rect 23171 -41399 23205 -40594
rect 23279 -40606 23397 -40594
rect 23550 -40570 23620 -40389
rect 23673 -40514 23707 -39693
rect 23550 -40624 23724 -40570
rect 23771 -40580 23805 -39806
rect 24073 -40514 24107 -39693
rect 24003 -40580 24137 -40572
rect 23771 -40619 24137 -40580
rect 23771 -41399 23805 -40619
rect 24003 -40626 24137 -40619
rect 24171 -40587 24205 -39806
rect 24356 -40587 24474 -40575
rect 24171 -40621 24474 -40587
rect 24171 -41399 24205 -40621
rect 24356 -40633 24474 -40621
rect 24541 -40577 24611 -40390
rect 24673 -40514 24707 -39693
rect 24541 -40631 24724 -40577
rect 24771 -40581 24805 -39806
rect 25073 -40514 25107 -39693
rect 25171 -40571 25205 -39806
rect 25252 -40571 25370 -40563
rect 24996 -40581 25130 -40574
rect 24771 -40620 25130 -40581
rect 24771 -41399 24805 -40620
rect 24996 -40628 25130 -40620
rect 25171 -40605 25373 -40571
rect 25171 -41399 25205 -40605
rect 25252 -40621 25370 -40605
rect 27383 -39832 27459 -38760
rect 27598 -38761 28084 -38760
rect 27598 -38762 27669 -38761
rect 28010 -38767 28084 -38761
rect 27630 -39112 27664 -38804
rect 27728 -39112 27762 -38804
rect 27826 -39112 27860 -38804
rect 27924 -39112 27958 -38804
rect 28022 -39112 28056 -38804
rect 27727 -39164 27762 -39112
rect 28441 -39146 28502 -38739
rect 28931 -38903 29001 -38508
rect 29175 -38762 29209 -38178
rect 29382 -38144 29622 -38110
rect 29382 -38186 29424 -38144
rect 29171 -38821 29213 -38762
rect 29386 -38768 29420 -38186
rect 29484 -38766 29518 -38178
rect 29580 -38188 29622 -38144
rect 29383 -38821 29425 -38768
rect 29171 -38857 29425 -38821
rect 29480 -38820 29522 -38766
rect 29582 -38786 29616 -38188
rect 29794 -38772 29828 -38178
rect 29480 -38859 29621 -38820
rect 29578 -38871 29621 -38859
rect 29336 -38903 29491 -38893
rect 28931 -38939 29491 -38903
rect 28931 -38941 29001 -38939
rect 29336 -38948 29491 -38939
rect 29578 -38926 29759 -38871
rect 29578 -38996 29621 -38926
rect 29066 -39010 29221 -39001
rect 29029 -39044 29221 -39010
rect 29066 -39056 29221 -39044
rect 29267 -39036 29621 -38996
rect 29793 -39016 29836 -38772
rect 30030 -38841 30100 -37504
rect 36194 -37557 36228 -37349
rect 36390 -37557 36424 -37349
rect 36586 -37557 36620 -37349
rect 31167 -38536 31201 -38036
rect 31346 -38000 31667 -37966
rect 31166 -38582 31201 -38536
rect 31346 -38582 31386 -38000
rect 31435 -38040 31470 -38000
rect 31436 -38544 31470 -38040
rect 31534 -38537 31568 -38036
rect 31632 -38039 31667 -38000
rect 31166 -38622 31386 -38582
rect 31531 -38657 31569 -38537
rect 31632 -38544 31666 -38039
rect 31762 -38620 31796 -38036
rect 32088 -38550 32122 -38036
rect 32316 -38326 32350 -38036
rect 37167 -37686 37201 -37342
rect 37363 -37686 37397 -37342
rect 37536 -37491 37597 -37342
rect 37776 -37456 37810 -37300
rect 37874 -37456 37908 -37348
rect 37972 -37456 38006 -37300
rect 44765 -37341 45012 -37300
rect 45847 -37328 45982 -37320
rect 45827 -37330 45982 -37328
rect 38070 -37456 38104 -37348
rect 44765 -37358 44895 -37341
rect 44939 -37354 45012 -37341
rect 45620 -37366 45982 -37330
rect 46499 -37339 47284 -37253
rect 53963 -37266 54093 -37174
rect 54255 -37232 54289 -36976
rect 54353 -37232 54387 -37024
rect 54451 -37232 54485 -36976
rect 54549 -37198 54583 -37024
rect 55130 -37154 55164 -36846
rect 55228 -37154 55262 -36846
rect 55326 -37154 55360 -36846
rect 55424 -37154 55458 -36846
rect 55522 -37154 55556 -36846
rect 55098 -37197 55169 -37196
rect 55510 -37197 55584 -37191
rect 55098 -37198 55584 -37197
rect 54549 -37232 55584 -37198
rect 55941 -37219 56002 -36812
rect 60589 -36842 62440 -36691
rect 63721 -36685 64386 -36657
rect 63721 -36743 64756 -36685
rect 63721 -36824 63807 -36743
rect 63981 -36780 64016 -36743
rect 64306 -36746 64756 -36743
rect 60589 -36910 60965 -36842
rect 62190 -36893 62440 -36842
rect 62869 -36910 63807 -36824
rect 62717 -37200 62847 -37108
rect 63009 -37166 63043 -36910
rect 63107 -37166 63141 -36958
rect 63205 -37166 63239 -36910
rect 63303 -37132 63337 -36958
rect 63884 -37088 63918 -36780
rect 63982 -37088 64016 -36780
rect 64080 -37088 64114 -36780
rect 64178 -37088 64212 -36780
rect 64276 -37088 64310 -36780
rect 63852 -37131 63923 -37130
rect 64264 -37131 64338 -37125
rect 63852 -37132 64338 -37131
rect 63303 -37166 64338 -37132
rect 64695 -37153 64756 -36746
rect 69365 -36697 69703 -36601
rect 73141 -36640 73481 -36246
rect 78595 -36636 78865 -36515
rect 80608 -36636 80903 -36594
rect 82477 -36602 82688 -36246
rect 71353 -36697 71621 -36656
rect 69365 -36828 71621 -36697
rect 72874 -36668 73539 -36640
rect 72874 -36726 73909 -36668
rect 72874 -36807 72960 -36726
rect 73134 -36763 73169 -36726
rect 73459 -36729 73909 -36726
rect 69365 -36892 69703 -36828
rect 71353 -36896 71621 -36828
rect 72022 -36893 72960 -36807
rect 63304 -37170 64338 -37166
rect 63304 -37172 63853 -37170
rect 62891 -37200 62964 -37194
rect 64264 -37196 64338 -37170
rect 54550 -37236 55584 -37232
rect 54550 -37238 55099 -37236
rect 54137 -37266 54210 -37260
rect 55510 -37262 55584 -37236
rect 53963 -37307 54210 -37266
rect 55045 -37294 55180 -37286
rect 55025 -37296 55180 -37294
rect 53963 -37324 54093 -37307
rect 54137 -37320 54210 -37307
rect 54818 -37332 55180 -37296
rect 55697 -37305 56482 -37219
rect 62717 -37241 62964 -37200
rect 63799 -37228 63934 -37220
rect 63779 -37230 63934 -37228
rect 62717 -37258 62847 -37241
rect 62891 -37254 62964 -37241
rect 63572 -37266 63934 -37230
rect 64451 -37239 65236 -37153
rect 71870 -37183 72000 -37091
rect 72162 -37149 72196 -36893
rect 72260 -37149 72294 -36941
rect 72358 -37149 72392 -36893
rect 72456 -37115 72490 -36941
rect 73037 -37071 73071 -36763
rect 73135 -37071 73169 -36763
rect 73233 -37071 73267 -36763
rect 73331 -37071 73365 -36763
rect 73429 -37071 73463 -36763
rect 73005 -37114 73076 -37113
rect 73417 -37114 73491 -37108
rect 73005 -37115 73491 -37114
rect 72456 -37149 73491 -37115
rect 73848 -37136 73909 -36729
rect 78595 -36775 80903 -36636
rect 82238 -36630 82903 -36602
rect 82238 -36688 83273 -36630
rect 82238 -36769 82324 -36688
rect 82498 -36725 82533 -36688
rect 82823 -36691 83273 -36688
rect 78595 -36800 78865 -36775
rect 80608 -36867 80903 -36775
rect 81386 -36855 82324 -36769
rect 72457 -37153 73491 -37149
rect 72457 -37155 73006 -37153
rect 72044 -37183 72117 -37177
rect 73417 -37179 73491 -37153
rect 71870 -37224 72117 -37183
rect 72952 -37211 73087 -37203
rect 72932 -37213 73087 -37211
rect 63779 -37268 63934 -37266
rect 63799 -37274 63934 -37268
rect 63982 -37251 64401 -37243
rect 63982 -37281 64412 -37251
rect 55025 -37334 55180 -37332
rect 45827 -37368 45982 -37366
rect 45847 -37374 45982 -37368
rect 46030 -37351 46449 -37343
rect 46030 -37381 46460 -37351
rect 37658 -37491 37731 -37485
rect 37536 -37504 37731 -37491
rect 37558 -37532 37731 -37504
rect 37658 -37545 37731 -37532
rect 38168 -37515 38540 -37445
rect 37776 -37687 37810 -37579
rect 37972 -37687 38006 -37579
rect 38168 -37687 38202 -37515
rect 32315 -38419 32352 -38326
rect 32315 -38456 32452 -38419
rect 32088 -38584 32247 -38550
rect 31911 -38620 32049 -38609
rect 31167 -38695 31569 -38657
rect 31636 -38654 32049 -38620
rect 30930 -38706 31068 -38696
rect 30540 -38740 31068 -38706
rect 30019 -38913 30124 -38841
rect 30540 -39016 30583 -38740
rect 30930 -38750 31068 -38740
rect 30986 -38841 31124 -38832
rect 30776 -38875 31124 -38841
rect 30776 -39002 30848 -38875
rect 30986 -38886 31124 -38875
rect 30776 -39011 30860 -39002
rect 28052 -39164 28502 -39146
rect 27610 -39207 28502 -39164
rect 27610 -39225 28059 -39207
rect 28441 -39502 28502 -39207
rect 29175 -39384 29209 -39090
rect 29267 -39106 29312 -39036
rect 29659 -39056 30583 -39016
rect 29707 -39059 30583 -39056
rect 29168 -39502 29215 -39384
rect 29273 -39398 29307 -39106
rect 29371 -39383 29405 -39090
rect 29613 -39373 29647 -39090
rect 29707 -39099 29751 -39059
rect 30781 -39081 30860 -39011
rect 29364 -39502 29411 -39383
rect 29606 -39502 29653 -39373
rect 29711 -39398 29745 -39099
rect 31069 -39323 31103 -39032
rect 31067 -39434 31104 -39323
rect 31167 -39340 31201 -38695
rect 31396 -38765 31434 -38695
rect 31636 -38733 31670 -38654
rect 31911 -38663 32049 -38654
rect 31386 -38903 31440 -38765
rect 31539 -38767 31670 -38733
rect 31736 -38750 31874 -38696
rect 32121 -38765 32175 -38627
rect 32213 -38628 32247 -38584
rect 32213 -38682 32379 -38628
rect 31539 -39340 31573 -38767
rect 32213 -38797 32247 -38682
rect 32299 -38797 32353 -38780
rect 31637 -38836 31796 -38801
rect 32213 -38802 32353 -38797
rect 32185 -38831 32353 -38802
rect 31637 -39340 31671 -38836
rect 31762 -39340 31796 -38836
rect 31860 -39323 31894 -38832
rect 31990 -39322 32024 -38832
rect 30530 -39438 31141 -39434
rect 31859 -39438 31896 -39323
rect 31987 -39438 32024 -39322
rect 32088 -39340 32122 -38832
rect 32185 -38836 32247 -38831
rect 32186 -39340 32220 -38836
rect 32299 -38839 32353 -38831
rect 32414 -38949 32452 -38456
rect 32414 -38987 32706 -38949
rect 32316 -39321 32350 -39032
rect 32414 -39037 32452 -38987
rect 32314 -39438 32351 -39321
rect 32414 -39340 32448 -39037
rect 30530 -39502 32464 -39438
rect 28441 -39547 32464 -39502
rect 28441 -39615 30643 -39547
rect 30991 -39599 32464 -39547
rect 9135 -41996 10105 -41735
rect 9283 -42439 9431 -42391
rect 9127 -42574 9250 -42530
rect 8968 -42701 9125 -42661
rect 8968 -44232 9022 -42701
rect 9182 -43005 9236 -42574
rect 9083 -43059 9236 -43005
rect 9083 -44232 9137 -43059
rect 9227 -44137 9281 -44107
rect 9325 -44137 9379 -42439
rect 9844 -43776 10105 -41996
rect 26587 -39888 27459 -39832
rect 32668 -39882 32706 -38987
rect 26587 -39964 30693 -39888
rect 26587 -39978 27459 -39964
rect 11368 -42251 11402 -42247
rect 11362 -42504 11408 -42251
rect 11564 -42439 11598 -42247
rect 11558 -42504 11604 -42439
rect 11760 -42439 11794 -42247
rect 12029 -42433 12086 -42269
rect 11754 -42504 11800 -42439
rect 12250 -42251 12284 -42247
rect 11362 -42512 11800 -42504
rect 12244 -42504 12290 -42251
rect 12446 -42439 12480 -42247
rect 12440 -42504 12486 -42439
rect 12860 -42228 13488 -42194
rect 12642 -42439 12676 -42247
rect 12860 -42273 12896 -42228
rect 12636 -42504 12682 -42439
rect 12244 -42512 12682 -42504
rect 12737 -42488 12811 -42320
rect 12861 -42347 12895 -42273
rect 12737 -42512 12810 -42488
rect 11362 -42534 11830 -42512
rect 12040 -42530 12208 -42519
rect 11888 -42534 11948 -42530
rect 12005 -42534 12208 -42530
rect 11362 -42550 12208 -42534
rect 11270 -42786 11304 -42627
rect 11362 -42643 11408 -42550
rect 11368 -42735 11402 -42643
rect 11466 -42786 11500 -42627
rect 11558 -42643 11604 -42550
rect 11754 -42576 12208 -42550
rect 11754 -42582 11830 -42576
rect 11564 -42735 11598 -42643
rect 11662 -42786 11696 -42627
rect 11754 -42643 11800 -42582
rect 11760 -42735 11794 -42643
rect 11888 -42662 11948 -42576
rect 12005 -42588 12208 -42576
rect 12040 -42593 12208 -42588
rect 12244 -42550 12810 -42512
rect 12152 -42786 12186 -42627
rect 12244 -42643 12290 -42550
rect 12250 -42735 12284 -42643
rect 12348 -42786 12382 -42627
rect 12440 -42643 12486 -42550
rect 12636 -42582 12810 -42550
rect 12855 -42494 12902 -42347
rect 12959 -42354 12993 -42262
rect 13056 -42283 13098 -42228
rect 12958 -42406 12994 -42354
rect 13057 -42370 13091 -42283
rect 13155 -42352 13189 -42262
rect 13250 -42284 13292 -42228
rect 13155 -42370 13192 -42352
rect 13253 -42370 13287 -42284
rect 13351 -42352 13385 -42262
rect 13446 -42279 13488 -42228
rect 13156 -42406 13192 -42370
rect 13350 -42406 13386 -42352
rect 13449 -42370 13483 -42279
rect 13547 -42362 13581 -42262
rect 13544 -42406 13586 -42362
rect 12958 -42440 13586 -42406
rect 12855 -42568 13027 -42494
rect 13411 -42528 13586 -42440
rect 13993 -42251 14027 -42247
rect 13987 -42504 14033 -42251
rect 14189 -42439 14223 -42247
rect 14183 -42504 14229 -42439
rect 14385 -42439 14419 -42247
rect 14729 -42347 14786 -42269
rect 14525 -42392 14786 -42347
rect 14379 -42504 14425 -42439
rect 13987 -42512 14425 -42504
rect 13783 -42528 13951 -42519
rect 12446 -42735 12480 -42643
rect 12544 -42786 12578 -42627
rect 12636 -42643 12682 -42582
rect 12642 -42735 12676 -42643
rect 12855 -42703 12902 -42568
rect 13411 -42585 13951 -42528
rect 13411 -42607 13586 -42585
rect 13783 -42593 13951 -42585
rect 13987 -42526 14455 -42512
rect 14525 -42526 14570 -42392
rect 14729 -42433 14786 -42392
rect 14950 -42251 14984 -42247
rect 14944 -42504 14990 -42251
rect 15146 -42439 15180 -42247
rect 15140 -42504 15186 -42439
rect 15560 -42228 16188 -42194
rect 15342 -42439 15376 -42247
rect 15560 -42273 15596 -42228
rect 15336 -42504 15382 -42439
rect 14944 -42512 15382 -42504
rect 15437 -42488 15511 -42320
rect 15561 -42347 15595 -42273
rect 15437 -42512 15510 -42488
rect 13987 -42550 14570 -42526
rect 12955 -42641 13586 -42607
rect 12955 -42682 12996 -42641
rect 12861 -42773 12895 -42703
rect 11261 -42854 12677 -42786
rect 12856 -42831 12900 -42773
rect 12959 -42785 12993 -42682
rect 13057 -42762 13091 -42677
rect 13153 -42690 13194 -42641
rect 13052 -42831 13096 -42762
rect 13155 -42785 13189 -42690
rect 13253 -42762 13287 -42677
rect 13347 -42690 13388 -42641
rect 13544 -42648 13586 -42641
rect 13248 -42831 13292 -42762
rect 13351 -42785 13385 -42690
rect 13449 -42773 13483 -42677
rect 13544 -42681 13585 -42648
rect 13538 -42691 13585 -42681
rect 13445 -42831 13489 -42773
rect 13538 -42813 13584 -42691
rect 13895 -42786 13929 -42627
rect 13987 -42643 14033 -42550
rect 13993 -42735 14027 -42643
rect 14091 -42786 14125 -42627
rect 14183 -42643 14229 -42550
rect 14379 -42571 14570 -42550
rect 14379 -42582 14455 -42571
rect 14189 -42735 14223 -42643
rect 14287 -42786 14321 -42627
rect 14379 -42643 14425 -42582
rect 14385 -42735 14419 -42643
rect 14505 -42686 14565 -42571
rect 14944 -42550 15510 -42512
rect 14852 -42786 14886 -42627
rect 14944 -42643 14990 -42550
rect 14950 -42735 14984 -42643
rect 15048 -42786 15082 -42627
rect 15140 -42643 15186 -42550
rect 15336 -42582 15510 -42550
rect 15555 -42494 15602 -42347
rect 15659 -42354 15693 -42262
rect 15756 -42283 15798 -42228
rect 15658 -42406 15694 -42354
rect 15757 -42370 15791 -42283
rect 15855 -42352 15889 -42262
rect 15950 -42284 15992 -42228
rect 15855 -42370 15892 -42352
rect 15953 -42370 15987 -42284
rect 16051 -42352 16085 -42262
rect 16146 -42279 16188 -42228
rect 15856 -42406 15892 -42370
rect 16050 -42406 16086 -42352
rect 16149 -42370 16183 -42279
rect 16247 -42362 16281 -42262
rect 16244 -42406 16286 -42362
rect 15658 -42440 16286 -42406
rect 15555 -42568 15727 -42494
rect 16111 -42525 16286 -42440
rect 16693 -42251 16727 -42247
rect 16687 -42504 16733 -42251
rect 16889 -42439 16923 -42247
rect 16883 -42504 16929 -42439
rect 17085 -42439 17119 -42247
rect 17079 -42504 17125 -42439
rect 16687 -42512 17125 -42504
rect 16483 -42525 16651 -42519
rect 15146 -42735 15180 -42643
rect 15244 -42786 15278 -42627
rect 15336 -42643 15382 -42582
rect 15342 -42735 15376 -42643
rect 15555 -42703 15602 -42568
rect 16111 -42578 16651 -42525
rect 16111 -42607 16286 -42578
rect 16483 -42593 16651 -42578
rect 16687 -42521 17155 -42512
rect 16687 -42523 17237 -42521
rect 16687 -42550 17238 -42523
rect 15655 -42641 16286 -42607
rect 15655 -42682 15696 -42641
rect 15561 -42773 15595 -42703
rect 12856 -42865 13489 -42831
rect 13886 -42854 15377 -42786
rect 15556 -42831 15600 -42773
rect 15659 -42785 15693 -42682
rect 15757 -42762 15791 -42677
rect 15853 -42690 15894 -42641
rect 15752 -42831 15796 -42762
rect 15855 -42785 15889 -42690
rect 15953 -42762 15987 -42677
rect 16047 -42690 16088 -42641
rect 16244 -42648 16286 -42641
rect 15948 -42831 15992 -42762
rect 16051 -42785 16085 -42690
rect 16149 -42773 16183 -42677
rect 16244 -42691 16285 -42648
rect 16145 -42831 16189 -42773
rect 16247 -42785 16281 -42691
rect 16595 -42786 16629 -42627
rect 16687 -42643 16733 -42550
rect 16693 -42735 16727 -42643
rect 16791 -42786 16825 -42627
rect 16883 -42643 16929 -42550
rect 17079 -42560 17238 -42550
rect 17079 -42582 17155 -42560
rect 16889 -42735 16923 -42643
rect 16987 -42786 17021 -42627
rect 17079 -42643 17125 -42582
rect 17085 -42735 17119 -42643
rect 15556 -42865 16189 -42831
rect 16586 -42854 17120 -42786
rect 11847 -42901 11979 -42890
rect 16370 -42901 16502 -42888
rect 11847 -42940 16908 -42901
rect 17190 -42918 17238 -42560
rect 11847 -42950 11979 -42940
rect 16370 -42948 16502 -42940
rect 17179 -43055 17239 -42918
rect 11524 -43079 11656 -43060
rect 14157 -43079 14294 -43060
rect 16754 -43079 16891 -43066
rect 11523 -43118 16908 -43079
rect 11524 -43120 11889 -43118
rect 11628 -43776 11889 -43120
rect 12245 -43189 12878 -43155
rect 13282 -43166 13393 -43118
rect 14157 -43120 14294 -43118
rect 13568 -43166 14088 -43164
rect 14160 -43166 14271 -43120
rect 12153 -43329 12187 -43235
rect 12245 -43247 12289 -43189
rect 12149 -43372 12190 -43329
rect 12251 -43343 12285 -43247
rect 12349 -43330 12383 -43235
rect 12442 -43258 12486 -43189
rect 12148 -43379 12190 -43372
rect 12346 -43379 12387 -43330
rect 12447 -43343 12481 -43258
rect 12545 -43330 12579 -43235
rect 12638 -43258 12682 -43189
rect 12540 -43379 12581 -43330
rect 12643 -43343 12677 -43258
rect 12741 -43338 12775 -43235
rect 12834 -43247 12878 -43189
rect 13057 -43232 14428 -43166
rect 13057 -43234 13591 -43232
rect 13894 -43234 14428 -43232
rect 14945 -43189 15578 -43155
rect 15958 -43166 16069 -43118
rect 16754 -43126 16891 -43118
rect 16769 -43166 16880 -43126
rect 12839 -43317 12873 -43247
rect 12738 -43379 12779 -43338
rect 12148 -43411 12779 -43379
rect 12073 -43413 12779 -43411
rect 12073 -43471 12323 -43413
rect 12832 -43452 12879 -43317
rect 13058 -43377 13092 -43285
rect 13052 -43438 13098 -43377
rect 13156 -43393 13190 -43234
rect 13254 -43377 13288 -43285
rect 12148 -43580 12323 -43471
rect 12707 -43526 12879 -43452
rect 12148 -43614 12776 -43580
rect 12148 -43658 12190 -43614
rect 12153 -43758 12187 -43658
rect 12251 -43741 12285 -43650
rect 12348 -43668 12384 -43614
rect 12542 -43650 12578 -43614
rect 9844 -44037 11889 -43776
rect 12246 -43792 12288 -43741
rect 12349 -43758 12383 -43668
rect 12447 -43736 12481 -43650
rect 12542 -43668 12579 -43650
rect 12442 -43792 12484 -43736
rect 12545 -43758 12579 -43668
rect 12643 -43737 12677 -43650
rect 12740 -43666 12776 -43614
rect 12636 -43792 12678 -43737
rect 12741 -43758 12775 -43666
rect 12832 -43673 12879 -43526
rect 12924 -43470 13098 -43438
rect 13248 -43470 13294 -43377
rect 13352 -43393 13386 -43234
rect 13450 -43377 13484 -43285
rect 13444 -43470 13490 -43377
rect 13548 -43393 13582 -43234
rect 13895 -43377 13929 -43285
rect 12924 -43508 13490 -43470
rect 13889 -43438 13935 -43377
rect 13993 -43393 14027 -43234
rect 14091 -43377 14125 -43285
rect 13791 -43470 13935 -43438
rect 14085 -43470 14131 -43377
rect 14189 -43393 14223 -43234
rect 14287 -43377 14321 -43285
rect 14281 -43470 14327 -43377
rect 14385 -43393 14419 -43234
rect 14853 -43329 14887 -43235
rect 14945 -43247 14989 -43189
rect 14849 -43372 14890 -43329
rect 14951 -43343 14985 -43247
rect 15049 -43330 15083 -43235
rect 15142 -43258 15186 -43189
rect 14848 -43379 14890 -43372
rect 15046 -43379 15087 -43330
rect 15147 -43343 15181 -43258
rect 15245 -43330 15279 -43235
rect 15338 -43258 15382 -43189
rect 15240 -43379 15281 -43330
rect 15343 -43343 15377 -43258
rect 15441 -43338 15475 -43235
rect 15534 -43247 15578 -43189
rect 15757 -43234 17128 -43166
rect 15539 -43317 15573 -43247
rect 15438 -43379 15479 -43338
rect 14848 -43413 15479 -43379
rect 12924 -43532 12997 -43508
rect 12839 -43747 12873 -43673
rect 12923 -43700 12997 -43532
rect 13052 -43516 13490 -43508
rect 13052 -43581 13098 -43516
rect 12838 -43792 12874 -43747
rect 13058 -43773 13092 -43581
rect 12246 -43826 12874 -43792
rect 13248 -43581 13294 -43516
rect 13254 -43773 13288 -43581
rect 13444 -43769 13490 -43516
rect 13791 -43508 14327 -43470
rect 14363 -43434 14531 -43427
rect 14363 -43494 14553 -43434
rect 14757 -43473 15023 -43413
rect 15532 -43452 15579 -43317
rect 15758 -43377 15792 -43285
rect 15752 -43438 15798 -43377
rect 15856 -43393 15890 -43234
rect 15954 -43377 15988 -43285
rect 14363 -43501 14531 -43494
rect 13450 -43773 13484 -43769
rect 13648 -43637 13705 -43587
rect 13791 -43637 13853 -43508
rect 13889 -43516 14327 -43508
rect 13889 -43581 13935 -43516
rect 13648 -43699 13853 -43637
rect 13648 -43751 13705 -43699
rect 13895 -43773 13929 -43581
rect 14085 -43581 14131 -43516
rect 14091 -43773 14125 -43581
rect 14281 -43769 14327 -43516
rect 14287 -43773 14321 -43769
rect 14848 -43580 15023 -43473
rect 15407 -43526 15579 -43452
rect 14848 -43614 15476 -43580
rect 14848 -43658 14890 -43614
rect 14853 -43758 14887 -43658
rect 14951 -43741 14985 -43650
rect 15048 -43668 15084 -43614
rect 15242 -43650 15278 -43614
rect 14946 -43792 14988 -43741
rect 15049 -43758 15083 -43668
rect 15147 -43736 15181 -43650
rect 15242 -43668 15279 -43650
rect 15142 -43792 15184 -43736
rect 15245 -43758 15279 -43668
rect 15343 -43737 15377 -43650
rect 15440 -43666 15476 -43614
rect 15336 -43792 15378 -43737
rect 15441 -43758 15475 -43666
rect 15532 -43673 15579 -43526
rect 15624 -43470 15798 -43438
rect 15948 -43470 15994 -43377
rect 16052 -43393 16086 -43234
rect 16150 -43377 16184 -43285
rect 16144 -43470 16190 -43377
rect 16248 -43393 16282 -43234
rect 16406 -43427 16466 -43283
rect 16595 -43377 16629 -43285
rect 15624 -43508 16190 -43470
rect 16226 -43489 16466 -43427
rect 16589 -43438 16635 -43377
rect 16693 -43393 16727 -43234
rect 16791 -43377 16825 -43285
rect 16502 -43470 16635 -43438
rect 16785 -43470 16831 -43377
rect 16889 -43393 16923 -43234
rect 16987 -43377 17021 -43285
rect 16981 -43470 17027 -43377
rect 17085 -43393 17119 -43234
rect 17190 -43427 17238 -43055
rect 16226 -43490 16429 -43489
rect 16226 -43501 16394 -43490
rect 15624 -43532 15697 -43508
rect 15539 -43747 15573 -43673
rect 15623 -43700 15697 -43532
rect 15752 -43516 16190 -43508
rect 15752 -43581 15798 -43516
rect 15538 -43792 15574 -43747
rect 15758 -43773 15792 -43581
rect 14946 -43826 15574 -43792
rect 15948 -43581 15994 -43516
rect 15954 -43773 15988 -43581
rect 16144 -43769 16190 -43516
rect 16502 -43508 17027 -43470
rect 17063 -43471 17238 -43427
rect 17063 -43501 17231 -43471
rect 16150 -43773 16184 -43769
rect 16348 -43638 16405 -43587
rect 16502 -43638 16548 -43508
rect 16589 -43516 17027 -43508
rect 16589 -43581 16635 -43516
rect 16348 -43687 16548 -43638
rect 16348 -43751 16405 -43687
rect 16595 -43773 16629 -43581
rect 16785 -43581 16831 -43516
rect 16791 -43773 16825 -43581
rect 16981 -43769 17027 -43516
rect 16987 -43773 17021 -43769
rect 26587 -43728 26733 -39978
rect 27383 -40146 27459 -39978
rect 27383 -40222 27525 -40146
rect 27449 -40611 27525 -40222
rect 28458 -40188 29123 -40160
rect 28458 -40246 29493 -40188
rect 28458 -40327 28544 -40246
rect 28718 -40283 28753 -40246
rect 29043 -40249 29493 -40246
rect 27606 -40413 28544 -40327
rect 27449 -40703 27584 -40611
rect 27746 -40669 27780 -40413
rect 27844 -40669 27878 -40461
rect 27942 -40669 27976 -40413
rect 28040 -40635 28074 -40461
rect 28621 -40591 28655 -40283
rect 28719 -40591 28753 -40283
rect 28817 -40591 28851 -40283
rect 28915 -40591 28949 -40283
rect 29013 -40591 29047 -40283
rect 28589 -40634 28660 -40633
rect 29001 -40634 29075 -40628
rect 28589 -40635 29075 -40634
rect 28040 -40669 29075 -40635
rect 29432 -40656 29493 -40249
rect 28041 -40673 29075 -40669
rect 28041 -40675 28590 -40673
rect 27628 -40703 27701 -40697
rect 29001 -40699 29075 -40673
rect 27449 -40720 27701 -40703
rect 27454 -40744 27701 -40720
rect 28536 -40731 28671 -40723
rect 28516 -40733 28671 -40731
rect 27454 -40761 27584 -40744
rect 27628 -40757 27701 -40744
rect 28309 -40769 28671 -40733
rect 29188 -40742 29973 -40656
rect 28516 -40771 28671 -40769
rect 28536 -40777 28671 -40771
rect 28719 -40754 29138 -40746
rect 28719 -40784 29149 -40754
rect 27746 -40999 27780 -40791
rect 27942 -40999 27976 -40791
rect 28138 -40999 28172 -40791
rect 28719 -41128 28753 -40784
rect 28915 -41128 28949 -40784
rect 29088 -40933 29149 -40784
rect 29328 -40898 29362 -40742
rect 29426 -40898 29460 -40790
rect 29524 -40898 29558 -40742
rect 29622 -40898 29656 -40790
rect 29210 -40933 29283 -40927
rect 29088 -40946 29283 -40933
rect 29110 -40974 29283 -40946
rect 29210 -40987 29283 -40974
rect 29720 -40957 30092 -40887
rect 29328 -41129 29362 -41021
rect 29524 -41129 29558 -41021
rect 29720 -41129 29754 -40957
rect 27720 -42064 27754 -41720
rect 27916 -42064 27950 -41720
rect 28329 -41827 28363 -41719
rect 28525 -41827 28559 -41719
rect 28211 -41874 28284 -41861
rect 28111 -41902 28284 -41874
rect 28089 -41915 28284 -41902
rect 28089 -42064 28150 -41915
rect 28211 -41921 28284 -41915
rect 28721 -41891 28755 -41719
rect 27720 -42094 28150 -42064
rect 27720 -42102 28139 -42094
rect 28329 -42106 28363 -41950
rect 28427 -42058 28461 -41950
rect 28525 -42106 28559 -41950
rect 28623 -42058 28657 -41950
rect 28721 -41961 28999 -41891
rect 24721 -43730 26733 -43728
rect 27364 -42175 27591 -42173
rect 28002 -42175 28076 -42149
rect 27364 -42213 28076 -42175
rect 28189 -42192 28804 -42106
rect 27590 -42214 28076 -42213
rect 27590 -42215 27661 -42214
rect 28002 -42220 28076 -42214
rect 27622 -42565 27656 -42257
rect 27720 -42565 27754 -42257
rect 27818 -42565 27852 -42257
rect 27916 -42565 27950 -42257
rect 28014 -42565 28048 -42257
rect 27719 -42617 27754 -42565
rect 28433 -42599 28494 -42192
rect 28923 -42356 28993 -41961
rect 29167 -42215 29201 -41631
rect 29374 -41597 29614 -41563
rect 29374 -41639 29416 -41597
rect 29163 -42274 29205 -42215
rect 29378 -42221 29412 -41639
rect 29476 -42219 29510 -41631
rect 29572 -41641 29614 -41597
rect 29375 -42274 29417 -42221
rect 29163 -42310 29417 -42274
rect 29472 -42273 29514 -42219
rect 29574 -42239 29608 -41641
rect 29786 -42225 29820 -41631
rect 29472 -42312 29613 -42273
rect 29570 -42324 29613 -42312
rect 29328 -42356 29483 -42346
rect 28923 -42392 29483 -42356
rect 28923 -42394 28993 -42392
rect 29328 -42401 29483 -42392
rect 29570 -42379 29751 -42324
rect 29570 -42449 29613 -42379
rect 29058 -42463 29213 -42454
rect 29021 -42497 29213 -42463
rect 29058 -42509 29213 -42497
rect 29259 -42489 29613 -42449
rect 29785 -42469 29828 -42225
rect 30022 -42294 30092 -40957
rect 30267 -40245 30359 -40160
rect 30290 -42220 30333 -40245
rect 30617 -40668 30693 -39964
rect 30919 -39920 32706 -39882
rect 30919 -40298 30957 -39920
rect 32126 -40219 32791 -40191
rect 32126 -40277 33161 -40219
rect 30896 -40352 30969 -40298
rect 32126 -40358 32212 -40277
rect 32386 -40314 32421 -40277
rect 32711 -40280 33161 -40277
rect 31274 -40444 32212 -40358
rect 31122 -40668 31252 -40642
rect 30617 -40734 31252 -40668
rect 31414 -40700 31448 -40444
rect 31512 -40700 31546 -40492
rect 31610 -40700 31644 -40444
rect 31708 -40666 31742 -40492
rect 32289 -40622 32323 -40314
rect 32387 -40622 32421 -40314
rect 32485 -40622 32519 -40314
rect 32583 -40622 32617 -40314
rect 32681 -40622 32715 -40314
rect 32257 -40665 32328 -40664
rect 32669 -40665 32743 -40659
rect 32257 -40666 32743 -40665
rect 31708 -40700 32743 -40666
rect 33100 -40687 33161 -40280
rect 36168 -38622 36202 -38278
rect 36364 -38622 36398 -38278
rect 36777 -38385 36811 -38277
rect 36973 -38385 37007 -38277
rect 36659 -38432 36732 -38419
rect 36559 -38460 36732 -38432
rect 36537 -38473 36732 -38460
rect 36537 -38622 36598 -38473
rect 36659 -38479 36732 -38473
rect 37169 -38449 37203 -38277
rect 36168 -38652 36598 -38622
rect 36168 -38660 36587 -38652
rect 36777 -38664 36811 -38508
rect 36875 -38616 36909 -38508
rect 36973 -38664 37007 -38508
rect 37071 -38616 37105 -38508
rect 37169 -38519 37447 -38449
rect 31709 -40704 32743 -40700
rect 31709 -40706 32258 -40704
rect 31296 -40734 31369 -40728
rect 32669 -40730 32743 -40704
rect 30617 -40744 31369 -40734
rect 31122 -40775 31369 -40744
rect 32204 -40762 32339 -40754
rect 32184 -40764 32339 -40762
rect 31122 -40792 31252 -40775
rect 31296 -40788 31369 -40775
rect 31149 -40842 31225 -40792
rect 31977 -40800 32339 -40764
rect 32856 -40773 33641 -40687
rect 32184 -40802 32339 -40800
rect 32204 -40808 32339 -40802
rect 32387 -40785 32806 -40777
rect 32387 -40815 32817 -40785
rect 31414 -41030 31448 -40822
rect 31610 -41030 31644 -40822
rect 31806 -41030 31840 -40822
rect 32387 -41159 32421 -40815
rect 32583 -41159 32617 -40815
rect 32756 -40964 32817 -40815
rect 32996 -40929 33030 -40773
rect 33094 -40929 33128 -40821
rect 33192 -40929 33226 -40773
rect 33290 -40929 33324 -40821
rect 32878 -40964 32951 -40958
rect 32756 -40977 32951 -40964
rect 32778 -41005 32951 -40977
rect 32878 -41018 32951 -41005
rect 33388 -40988 33760 -40918
rect 32996 -41160 33030 -41052
rect 33192 -41160 33226 -41052
rect 33388 -41160 33422 -40988
rect 31388 -42095 31422 -41751
rect 31584 -42095 31618 -41751
rect 31997 -41858 32031 -41750
rect 32193 -41858 32227 -41750
rect 31879 -41905 31952 -41892
rect 31779 -41933 31952 -41905
rect 31757 -41946 31952 -41933
rect 31757 -42095 31818 -41946
rect 31879 -41952 31952 -41946
rect 32389 -41922 32423 -41750
rect 31388 -42125 31818 -42095
rect 31388 -42133 31807 -42125
rect 31997 -42137 32031 -41981
rect 32095 -42089 32129 -41981
rect 32193 -42137 32227 -41981
rect 32291 -42089 32325 -41981
rect 32389 -41992 32667 -41922
rect 30290 -42263 30575 -42220
rect 30011 -42366 30116 -42294
rect 30532 -42469 30575 -42263
rect 28044 -42617 28494 -42599
rect 27602 -42660 28494 -42617
rect 27602 -42678 28051 -42660
rect 28433 -42955 28494 -42660
rect 29167 -42837 29201 -42543
rect 29259 -42559 29304 -42489
rect 29651 -42509 30575 -42469
rect 29699 -42512 30575 -42509
rect 29160 -42955 29207 -42837
rect 29265 -42851 29299 -42559
rect 29363 -42836 29397 -42543
rect 29605 -42826 29639 -42543
rect 29699 -42552 29743 -42512
rect 29356 -42955 29403 -42836
rect 29598 -42955 29645 -42826
rect 29703 -42851 29737 -42552
rect 28433 -43068 29910 -42955
rect 31032 -42206 31259 -42204
rect 31670 -42206 31744 -42180
rect 31032 -42244 31744 -42206
rect 31857 -42223 32472 -42137
rect 31258 -42245 31744 -42244
rect 31258 -42246 31329 -42245
rect 31670 -42251 31744 -42245
rect 31290 -42596 31324 -42288
rect 31388 -42596 31422 -42288
rect 31486 -42596 31520 -42288
rect 31584 -42596 31618 -42288
rect 31682 -42596 31716 -42288
rect 31387 -42648 31422 -42596
rect 32101 -42630 32162 -42223
rect 32591 -42387 32661 -41992
rect 32835 -42246 32869 -41662
rect 33042 -41628 33282 -41594
rect 33042 -41670 33084 -41628
rect 32831 -42305 32873 -42246
rect 33046 -42252 33080 -41670
rect 33144 -42250 33178 -41662
rect 33240 -41672 33282 -41628
rect 33043 -42305 33085 -42252
rect 32831 -42341 33085 -42305
rect 33140 -42304 33182 -42250
rect 33242 -42270 33276 -41672
rect 33454 -42256 33488 -41662
rect 33140 -42343 33281 -42304
rect 33238 -42355 33281 -42343
rect 32996 -42387 33151 -42377
rect 32591 -42423 33151 -42387
rect 32591 -42425 32661 -42423
rect 32996 -42432 33151 -42423
rect 33238 -42410 33419 -42355
rect 33238 -42480 33281 -42410
rect 32726 -42494 32881 -42485
rect 32689 -42528 32881 -42494
rect 32726 -42540 32881 -42528
rect 32927 -42520 33281 -42480
rect 33453 -42500 33496 -42256
rect 33690 -42325 33760 -40988
rect 33679 -42397 33784 -42325
rect 34185 -42500 34408 -42410
rect 31712 -42648 32162 -42630
rect 31270 -42691 32162 -42648
rect 31270 -42709 31719 -42691
rect 32101 -42986 32162 -42691
rect 32835 -42868 32869 -42574
rect 32927 -42590 32972 -42520
rect 33319 -42540 34521 -42500
rect 33367 -42543 34521 -42540
rect 32828 -42986 32875 -42868
rect 32933 -42882 32967 -42590
rect 33031 -42867 33065 -42574
rect 33273 -42857 33307 -42574
rect 33367 -42583 33411 -42543
rect 34185 -42580 34408 -42543
rect 33024 -42986 33071 -42867
rect 33266 -42986 33313 -42857
rect 33371 -42882 33405 -42583
rect 32101 -43099 33578 -42986
rect 24721 -43898 26752 -43730
rect 24721 -43899 26676 -43898
rect 9227 -44191 9379 -44137
rect 9227 -44232 9281 -44191
rect 35812 -38733 36039 -38731
rect 36450 -38733 36524 -38707
rect 35812 -38771 36524 -38733
rect 36637 -38750 37252 -38664
rect 35823 -39621 35899 -38771
rect 36038 -38772 36524 -38771
rect 36038 -38773 36109 -38772
rect 36450 -38778 36524 -38772
rect 36070 -39123 36104 -38815
rect 36168 -39123 36202 -38815
rect 36266 -39123 36300 -38815
rect 36364 -39123 36398 -38815
rect 36462 -39123 36496 -38815
rect 36167 -39175 36202 -39123
rect 36881 -39157 36942 -38750
rect 37371 -38914 37441 -38519
rect 37615 -38773 37649 -38189
rect 37822 -38155 38062 -38121
rect 37822 -38197 37864 -38155
rect 37611 -38832 37653 -38773
rect 37826 -38779 37860 -38197
rect 37924 -38777 37958 -38189
rect 38020 -38199 38062 -38155
rect 37823 -38832 37865 -38779
rect 37611 -38868 37865 -38832
rect 37920 -38831 37962 -38777
rect 38022 -38797 38056 -38199
rect 38234 -38783 38268 -38189
rect 37920 -38870 38061 -38831
rect 38018 -38882 38061 -38870
rect 37776 -38914 37931 -38904
rect 37371 -38950 37931 -38914
rect 37371 -38952 37441 -38950
rect 37776 -38959 37931 -38950
rect 38018 -38937 38199 -38882
rect 38018 -39007 38061 -38937
rect 37506 -39021 37661 -39012
rect 37469 -39055 37661 -39021
rect 37506 -39067 37661 -39055
rect 37707 -39047 38061 -39007
rect 38233 -39027 38276 -38783
rect 38470 -38852 38540 -37515
rect 45057 -37596 45091 -37388
rect 45253 -37596 45287 -37388
rect 45449 -37596 45483 -37388
rect 46030 -37725 46064 -37381
rect 46226 -37725 46260 -37381
rect 46399 -37530 46460 -37381
rect 46639 -37495 46673 -37339
rect 46737 -37495 46771 -37387
rect 46835 -37495 46869 -37339
rect 55045 -37340 55180 -37334
rect 55228 -37317 55647 -37309
rect 55228 -37347 55658 -37317
rect 46933 -37495 46967 -37387
rect 46521 -37530 46594 -37524
rect 46399 -37543 46594 -37530
rect 46421 -37571 46594 -37543
rect 46521 -37584 46594 -37571
rect 47031 -37554 47403 -37484
rect 46639 -37726 46673 -37618
rect 46835 -37726 46869 -37618
rect 47031 -37726 47065 -37554
rect 39607 -38547 39641 -38047
rect 39786 -38011 40107 -37977
rect 39606 -38593 39641 -38547
rect 39786 -38593 39826 -38011
rect 39875 -38051 39910 -38011
rect 39876 -38555 39910 -38051
rect 39974 -38548 40008 -38047
rect 40072 -38050 40107 -38011
rect 39606 -38633 39826 -38593
rect 39971 -38668 40009 -38548
rect 40072 -38555 40106 -38050
rect 40202 -38631 40236 -38047
rect 40528 -38561 40562 -38047
rect 40756 -38337 40790 -38047
rect 40755 -38430 40792 -38337
rect 40755 -38467 40892 -38430
rect 40528 -38595 40687 -38561
rect 40351 -38631 40489 -38620
rect 39607 -38706 40009 -38668
rect 40076 -38665 40489 -38631
rect 39370 -38717 39508 -38707
rect 38980 -38751 39508 -38717
rect 38459 -38924 38564 -38852
rect 38980 -39027 39023 -38751
rect 39370 -38761 39508 -38751
rect 39426 -38852 39564 -38843
rect 39216 -38886 39564 -38852
rect 39216 -39013 39288 -38886
rect 39426 -38897 39564 -38886
rect 39216 -39022 39300 -39013
rect 36492 -39175 36942 -39157
rect 36050 -39218 36942 -39175
rect 36050 -39236 36499 -39218
rect 35167 -39767 35899 -39621
rect 36881 -39513 36942 -39218
rect 37615 -39395 37649 -39101
rect 37707 -39117 37752 -39047
rect 38099 -39067 39023 -39027
rect 38147 -39070 39023 -39067
rect 37608 -39513 37655 -39395
rect 37713 -39409 37747 -39117
rect 37811 -39394 37845 -39101
rect 38053 -39384 38087 -39101
rect 38147 -39110 38191 -39070
rect 39221 -39092 39300 -39022
rect 37804 -39513 37851 -39394
rect 38046 -39513 38093 -39384
rect 38151 -39409 38185 -39110
rect 39509 -39334 39543 -39043
rect 39507 -39445 39544 -39334
rect 39607 -39351 39641 -38706
rect 39836 -38776 39874 -38706
rect 40076 -38744 40110 -38665
rect 40351 -38674 40489 -38665
rect 39826 -38914 39880 -38776
rect 39979 -38778 40110 -38744
rect 40176 -38761 40314 -38707
rect 40561 -38776 40615 -38638
rect 40653 -38639 40687 -38595
rect 40653 -38693 40819 -38639
rect 39979 -39351 40013 -38778
rect 40653 -38808 40687 -38693
rect 40739 -38808 40793 -38791
rect 40077 -38847 40236 -38812
rect 40653 -38813 40793 -38808
rect 40625 -38842 40793 -38813
rect 40077 -39351 40111 -38847
rect 40202 -39351 40236 -38847
rect 40300 -39334 40334 -38843
rect 40430 -39333 40464 -38843
rect 38970 -39449 39581 -39445
rect 40299 -39449 40336 -39334
rect 40427 -39449 40464 -39333
rect 40528 -39351 40562 -38843
rect 40625 -38847 40687 -38842
rect 40626 -39351 40660 -38847
rect 40739 -38850 40793 -38842
rect 40854 -38960 40892 -38467
rect 40854 -38998 41146 -38960
rect 40756 -39332 40790 -39043
rect 40854 -39048 40892 -38998
rect 40754 -39449 40791 -39332
rect 40854 -39351 40888 -39048
rect 38970 -39513 40904 -39449
rect 36881 -39558 40904 -39513
rect 36881 -39626 39083 -39558
rect 39431 -39610 40904 -39558
rect 35167 -43750 35313 -39767
rect 35823 -39899 35899 -39767
rect 41108 -39893 41146 -38998
rect 35823 -39975 39133 -39899
rect 35823 -40157 35899 -39975
rect 35823 -40233 35965 -40157
rect 35889 -40622 35965 -40233
rect 36898 -40199 37563 -40171
rect 36898 -40257 37933 -40199
rect 36898 -40338 36984 -40257
rect 37158 -40294 37193 -40257
rect 37483 -40260 37933 -40257
rect 36046 -40424 36984 -40338
rect 35889 -40714 36024 -40622
rect 36186 -40680 36220 -40424
rect 36284 -40680 36318 -40472
rect 36382 -40680 36416 -40424
rect 36480 -40646 36514 -40472
rect 37061 -40602 37095 -40294
rect 37159 -40602 37193 -40294
rect 37257 -40602 37291 -40294
rect 37355 -40602 37389 -40294
rect 37453 -40602 37487 -40294
rect 37029 -40645 37100 -40644
rect 37441 -40645 37515 -40639
rect 37029 -40646 37515 -40645
rect 36480 -40680 37515 -40646
rect 37872 -40667 37933 -40260
rect 36481 -40684 37515 -40680
rect 36481 -40686 37030 -40684
rect 36068 -40714 36141 -40708
rect 37441 -40710 37515 -40684
rect 35889 -40731 36141 -40714
rect 35894 -40755 36141 -40731
rect 36976 -40742 37111 -40734
rect 36956 -40744 37111 -40742
rect 35894 -40772 36024 -40755
rect 36068 -40768 36141 -40755
rect 36749 -40780 37111 -40744
rect 37628 -40753 38413 -40667
rect 36956 -40782 37111 -40780
rect 36976 -40788 37111 -40782
rect 37159 -40765 37578 -40757
rect 37159 -40795 37589 -40765
rect 36186 -41010 36220 -40802
rect 36382 -41010 36416 -40802
rect 36578 -41010 36612 -40802
rect 37159 -41139 37193 -40795
rect 37355 -41139 37389 -40795
rect 37528 -40944 37589 -40795
rect 37768 -40909 37802 -40753
rect 37866 -40909 37900 -40801
rect 37964 -40909 37998 -40753
rect 38062 -40909 38096 -40801
rect 37650 -40944 37723 -40938
rect 37528 -40957 37723 -40944
rect 37550 -40985 37723 -40957
rect 37650 -40998 37723 -40985
rect 38160 -40968 38532 -40898
rect 37768 -41140 37802 -41032
rect 37964 -41140 37998 -41032
rect 38160 -41140 38194 -40968
rect 36160 -42075 36194 -41731
rect 36356 -42075 36390 -41731
rect 36769 -41838 36803 -41730
rect 36965 -41838 36999 -41730
rect 36651 -41885 36724 -41872
rect 36551 -41913 36724 -41885
rect 36529 -41926 36724 -41913
rect 36529 -42075 36590 -41926
rect 36651 -41932 36724 -41926
rect 37161 -41902 37195 -41730
rect 36160 -42105 36590 -42075
rect 36160 -42113 36579 -42105
rect 36769 -42117 36803 -41961
rect 36867 -42069 36901 -41961
rect 36965 -42117 36999 -41961
rect 37063 -42069 37097 -41961
rect 37161 -41972 37439 -41902
rect 35804 -42186 36031 -42184
rect 36442 -42186 36516 -42160
rect 35804 -42224 36516 -42186
rect 36629 -42203 37244 -42117
rect 36030 -42225 36516 -42224
rect 36030 -42226 36101 -42225
rect 36442 -42231 36516 -42225
rect 36062 -42576 36096 -42268
rect 36160 -42576 36194 -42268
rect 36258 -42576 36292 -42268
rect 36356 -42576 36390 -42268
rect 36454 -42576 36488 -42268
rect 36159 -42628 36194 -42576
rect 36873 -42610 36934 -42203
rect 37363 -42367 37433 -41972
rect 37607 -42226 37641 -41642
rect 37814 -41608 38054 -41574
rect 37814 -41650 37856 -41608
rect 37603 -42285 37645 -42226
rect 37818 -42232 37852 -41650
rect 37916 -42230 37950 -41642
rect 38012 -41652 38054 -41608
rect 37815 -42285 37857 -42232
rect 37603 -42321 37857 -42285
rect 37912 -42284 37954 -42230
rect 38014 -42250 38048 -41652
rect 38226 -42236 38260 -41642
rect 37912 -42323 38053 -42284
rect 38010 -42335 38053 -42323
rect 37768 -42367 37923 -42357
rect 37363 -42403 37923 -42367
rect 37363 -42405 37433 -42403
rect 37768 -42412 37923 -42403
rect 38010 -42390 38191 -42335
rect 38010 -42460 38053 -42390
rect 37498 -42474 37653 -42465
rect 37461 -42508 37653 -42474
rect 37498 -42520 37653 -42508
rect 37699 -42500 38053 -42460
rect 38225 -42480 38268 -42236
rect 38462 -42305 38532 -40968
rect 38707 -40256 38799 -40171
rect 38730 -42231 38773 -40256
rect 39057 -40679 39133 -39975
rect 39359 -39931 41146 -39893
rect 39359 -40309 39397 -39931
rect 40566 -40230 41231 -40202
rect 40566 -40288 41601 -40230
rect 39336 -40363 39409 -40309
rect 40566 -40369 40652 -40288
rect 40826 -40325 40861 -40288
rect 41151 -40291 41601 -40288
rect 39714 -40455 40652 -40369
rect 39562 -40679 39692 -40653
rect 39057 -40745 39692 -40679
rect 39854 -40711 39888 -40455
rect 39952 -40711 39986 -40503
rect 40050 -40711 40084 -40455
rect 40148 -40677 40182 -40503
rect 40729 -40633 40763 -40325
rect 40827 -40633 40861 -40325
rect 40925 -40633 40959 -40325
rect 41023 -40633 41057 -40325
rect 41121 -40633 41155 -40325
rect 40697 -40676 40768 -40675
rect 41109 -40676 41183 -40670
rect 40697 -40677 41183 -40676
rect 40148 -40711 41183 -40677
rect 41540 -40698 41601 -40291
rect 45031 -38661 45065 -38317
rect 45227 -38661 45261 -38317
rect 45640 -38424 45674 -38316
rect 45836 -38424 45870 -38316
rect 45522 -38471 45595 -38458
rect 45422 -38499 45595 -38471
rect 45400 -38512 45595 -38499
rect 45400 -38661 45461 -38512
rect 45522 -38518 45595 -38512
rect 46032 -38488 46066 -38316
rect 45031 -38691 45461 -38661
rect 45031 -38699 45450 -38691
rect 45640 -38703 45674 -38547
rect 45738 -38655 45772 -38547
rect 45836 -38703 45870 -38547
rect 45934 -38655 45968 -38547
rect 46032 -38558 46310 -38488
rect 44675 -38772 44902 -38770
rect 45313 -38772 45387 -38746
rect 44675 -38810 45387 -38772
rect 45500 -38789 46115 -38703
rect 40149 -40715 41183 -40711
rect 40149 -40717 40698 -40715
rect 39736 -40745 39809 -40739
rect 41109 -40741 41183 -40715
rect 39057 -40755 39809 -40745
rect 39562 -40786 39809 -40755
rect 40644 -40773 40779 -40765
rect 40624 -40775 40779 -40773
rect 39562 -40803 39692 -40786
rect 39736 -40799 39809 -40786
rect 39589 -40853 39665 -40803
rect 40417 -40811 40779 -40775
rect 41296 -40784 42081 -40698
rect 40624 -40813 40779 -40811
rect 40644 -40819 40779 -40813
rect 40827 -40796 41246 -40788
rect 40827 -40826 41257 -40796
rect 39854 -41041 39888 -40833
rect 40050 -41041 40084 -40833
rect 40246 -41041 40280 -40833
rect 40827 -41170 40861 -40826
rect 41023 -41170 41057 -40826
rect 41196 -40975 41257 -40826
rect 41436 -40940 41470 -40784
rect 41534 -40940 41568 -40832
rect 41632 -40940 41666 -40784
rect 41730 -40940 41764 -40832
rect 41318 -40975 41391 -40969
rect 41196 -40988 41391 -40975
rect 41218 -41016 41391 -40988
rect 41318 -41029 41391 -41016
rect 41828 -40999 42200 -40929
rect 41436 -41171 41470 -41063
rect 41632 -41171 41666 -41063
rect 41828 -41171 41862 -40999
rect 39828 -42106 39862 -41762
rect 40024 -42106 40058 -41762
rect 40437 -41869 40471 -41761
rect 40633 -41869 40667 -41761
rect 40319 -41916 40392 -41903
rect 40219 -41944 40392 -41916
rect 40197 -41957 40392 -41944
rect 40197 -42106 40258 -41957
rect 40319 -41963 40392 -41957
rect 40829 -41933 40863 -41761
rect 39828 -42136 40258 -42106
rect 39828 -42144 40247 -42136
rect 40437 -42148 40471 -41992
rect 40535 -42100 40569 -41992
rect 40633 -42148 40667 -41992
rect 40731 -42100 40765 -41992
rect 40829 -42003 41107 -41933
rect 38730 -42274 39015 -42231
rect 38451 -42377 38556 -42305
rect 38972 -42480 39015 -42274
rect 36484 -42628 36934 -42610
rect 36042 -42671 36934 -42628
rect 36042 -42689 36491 -42671
rect 36873 -42966 36934 -42671
rect 37607 -42848 37641 -42554
rect 37699 -42570 37744 -42500
rect 38091 -42520 39015 -42480
rect 38139 -42523 39015 -42520
rect 37600 -42966 37647 -42848
rect 37705 -42862 37739 -42570
rect 37803 -42847 37837 -42554
rect 38045 -42837 38079 -42554
rect 38139 -42563 38183 -42523
rect 37796 -42966 37843 -42847
rect 38038 -42966 38085 -42837
rect 38143 -42862 38177 -42563
rect 36873 -43079 38350 -42966
rect 39472 -42217 39699 -42215
rect 40110 -42217 40184 -42191
rect 39472 -42255 40184 -42217
rect 40297 -42234 40912 -42148
rect 39698 -42256 40184 -42255
rect 39698 -42257 39769 -42256
rect 40110 -42262 40184 -42256
rect 39730 -42607 39764 -42299
rect 39828 -42607 39862 -42299
rect 39926 -42607 39960 -42299
rect 40024 -42607 40058 -42299
rect 40122 -42607 40156 -42299
rect 39827 -42659 39862 -42607
rect 40541 -42641 40602 -42234
rect 41031 -42398 41101 -42003
rect 41275 -42257 41309 -41673
rect 41482 -41639 41722 -41605
rect 41482 -41681 41524 -41639
rect 41271 -42316 41313 -42257
rect 41486 -42263 41520 -41681
rect 41584 -42261 41618 -41673
rect 41680 -41683 41722 -41639
rect 41483 -42316 41525 -42263
rect 41271 -42352 41525 -42316
rect 41580 -42315 41622 -42261
rect 41682 -42281 41716 -41683
rect 41894 -42267 41928 -41673
rect 41580 -42354 41721 -42315
rect 41678 -42366 41721 -42354
rect 41436 -42398 41591 -42388
rect 41031 -42434 41591 -42398
rect 41031 -42436 41101 -42434
rect 41436 -42443 41591 -42434
rect 41678 -42421 41859 -42366
rect 41678 -42491 41721 -42421
rect 41166 -42505 41321 -42496
rect 41129 -42539 41321 -42505
rect 41166 -42551 41321 -42539
rect 41367 -42531 41721 -42491
rect 41893 -42511 41936 -42267
rect 42130 -42336 42200 -40999
rect 42119 -42408 42224 -42336
rect 42634 -42511 42971 -42348
rect 40152 -42659 40602 -42641
rect 39710 -42702 40602 -42659
rect 39710 -42720 40159 -42702
rect 40541 -42997 40602 -42702
rect 41275 -42879 41309 -42585
rect 41367 -42601 41412 -42531
rect 41759 -42551 42971 -42511
rect 41807 -42554 42971 -42551
rect 41268 -42997 41315 -42879
rect 41373 -42893 41407 -42601
rect 41471 -42878 41505 -42585
rect 41713 -42868 41747 -42585
rect 41807 -42594 41851 -42554
rect 41464 -42997 41511 -42878
rect 41706 -42997 41753 -42868
rect 41811 -42893 41845 -42594
rect 42634 -42679 42971 -42554
rect 40541 -43110 42018 -42997
rect 35144 -43897 35347 -43750
rect 42275 -43931 42592 -43640
rect 42292 -44711 42558 -43931
rect 44686 -39748 44762 -38810
rect 44901 -38811 45387 -38810
rect 44901 -38812 44972 -38811
rect 45313 -38817 45387 -38811
rect 44933 -39162 44967 -38854
rect 45031 -39162 45065 -38854
rect 45129 -39162 45163 -38854
rect 45227 -39162 45261 -38854
rect 45325 -39162 45359 -38854
rect 45030 -39214 45065 -39162
rect 45744 -39196 45805 -38789
rect 46234 -38953 46304 -38558
rect 46478 -38812 46512 -38228
rect 46685 -38194 46925 -38160
rect 46685 -38236 46727 -38194
rect 46474 -38871 46516 -38812
rect 46689 -38818 46723 -38236
rect 46787 -38816 46821 -38228
rect 46883 -38238 46925 -38194
rect 46686 -38871 46728 -38818
rect 46474 -38907 46728 -38871
rect 46783 -38870 46825 -38816
rect 46885 -38836 46919 -38238
rect 47097 -38822 47131 -38228
rect 46783 -38909 46924 -38870
rect 46881 -38921 46924 -38909
rect 46639 -38953 46794 -38943
rect 46234 -38989 46794 -38953
rect 46234 -38991 46304 -38989
rect 46639 -38998 46794 -38989
rect 46881 -38976 47062 -38921
rect 46881 -39046 46924 -38976
rect 46369 -39060 46524 -39051
rect 46332 -39094 46524 -39060
rect 46369 -39106 46524 -39094
rect 46570 -39086 46924 -39046
rect 47096 -39066 47139 -38822
rect 47333 -38891 47403 -37554
rect 54255 -37562 54289 -37354
rect 54451 -37562 54485 -37354
rect 54647 -37562 54681 -37354
rect 55228 -37691 55262 -37347
rect 55424 -37691 55458 -37347
rect 55597 -37496 55658 -37347
rect 55837 -37461 55871 -37305
rect 55935 -37461 55969 -37353
rect 56033 -37461 56067 -37305
rect 56131 -37461 56165 -37353
rect 55719 -37496 55792 -37490
rect 55597 -37509 55792 -37496
rect 55619 -37537 55792 -37509
rect 55719 -37550 55792 -37537
rect 56229 -37520 56601 -37450
rect 55837 -37692 55871 -37584
rect 56033 -37692 56067 -37584
rect 56229 -37692 56263 -37520
rect 48470 -38586 48504 -38086
rect 48649 -38050 48970 -38016
rect 48469 -38632 48504 -38586
rect 48649 -38632 48689 -38050
rect 48738 -38090 48773 -38050
rect 48739 -38594 48773 -38090
rect 48837 -38587 48871 -38086
rect 48935 -38089 48970 -38050
rect 48469 -38672 48689 -38632
rect 48834 -38707 48872 -38587
rect 48935 -38594 48969 -38089
rect 49065 -38670 49099 -38086
rect 49391 -38600 49425 -38086
rect 49619 -38376 49653 -38086
rect 49618 -38469 49655 -38376
rect 49618 -38506 49755 -38469
rect 49391 -38634 49550 -38600
rect 49214 -38670 49352 -38659
rect 48470 -38745 48872 -38707
rect 48939 -38704 49352 -38670
rect 48233 -38756 48371 -38746
rect 47843 -38790 48371 -38756
rect 47322 -38963 47427 -38891
rect 47843 -39066 47886 -38790
rect 48233 -38800 48371 -38790
rect 48289 -38891 48427 -38882
rect 48079 -38925 48427 -38891
rect 48079 -39052 48151 -38925
rect 48289 -38936 48427 -38925
rect 48079 -39061 48163 -39052
rect 45355 -39214 45805 -39196
rect 44913 -39257 45805 -39214
rect 44913 -39275 45362 -39257
rect 45744 -39552 45805 -39257
rect 46478 -39434 46512 -39140
rect 46570 -39156 46615 -39086
rect 46962 -39106 47886 -39066
rect 47010 -39109 47886 -39106
rect 46471 -39552 46518 -39434
rect 46576 -39448 46610 -39156
rect 46674 -39433 46708 -39140
rect 46916 -39423 46950 -39140
rect 47010 -39149 47054 -39109
rect 48084 -39131 48163 -39061
rect 46667 -39552 46714 -39433
rect 46909 -39552 46956 -39423
rect 47014 -39448 47048 -39149
rect 48372 -39373 48406 -39082
rect 48370 -39484 48407 -39373
rect 48470 -39390 48504 -38745
rect 48699 -38815 48737 -38745
rect 48939 -38783 48973 -38704
rect 49214 -38713 49352 -38704
rect 48689 -38953 48743 -38815
rect 48842 -38817 48973 -38783
rect 49039 -38800 49177 -38746
rect 49424 -38815 49478 -38677
rect 49516 -38678 49550 -38634
rect 49516 -38732 49682 -38678
rect 48842 -39390 48876 -38817
rect 49516 -38847 49550 -38732
rect 49602 -38847 49656 -38830
rect 48940 -38886 49099 -38851
rect 49516 -38852 49656 -38847
rect 49488 -38881 49656 -38852
rect 48940 -39390 48974 -38886
rect 49065 -39390 49099 -38886
rect 49163 -39373 49197 -38882
rect 49293 -39372 49327 -38882
rect 47833 -39488 48444 -39484
rect 49162 -39488 49199 -39373
rect 49290 -39488 49327 -39372
rect 49391 -39390 49425 -38882
rect 49488 -38886 49550 -38881
rect 49489 -39390 49523 -38886
rect 49602 -38889 49656 -38881
rect 49717 -38999 49755 -38506
rect 49717 -39037 50009 -38999
rect 49619 -39371 49653 -39082
rect 49717 -39087 49755 -39037
rect 49617 -39488 49654 -39371
rect 49717 -39390 49751 -39087
rect 47833 -39552 49767 -39488
rect 45744 -39597 49767 -39552
rect 45744 -39665 47946 -39597
rect 48294 -39649 49767 -39597
rect 44036 -39894 44762 -39748
rect 44036 -43895 44182 -39894
rect 44686 -39938 44762 -39894
rect 49971 -39932 50009 -39037
rect 44686 -40014 47996 -39938
rect 44686 -40196 44762 -40014
rect 44686 -40272 44828 -40196
rect 44752 -40661 44828 -40272
rect 45761 -40238 46426 -40210
rect 45761 -40296 46796 -40238
rect 45761 -40377 45847 -40296
rect 46021 -40333 46056 -40296
rect 46346 -40299 46796 -40296
rect 44909 -40463 45847 -40377
rect 44752 -40753 44887 -40661
rect 45049 -40719 45083 -40463
rect 45147 -40719 45181 -40511
rect 45245 -40719 45279 -40463
rect 45343 -40685 45377 -40511
rect 45924 -40641 45958 -40333
rect 46022 -40641 46056 -40333
rect 46120 -40641 46154 -40333
rect 46218 -40641 46252 -40333
rect 46316 -40641 46350 -40333
rect 45892 -40684 45963 -40683
rect 46304 -40684 46378 -40678
rect 45892 -40685 46378 -40684
rect 45343 -40719 46378 -40685
rect 46735 -40706 46796 -40299
rect 45344 -40723 46378 -40719
rect 45344 -40725 45893 -40723
rect 44931 -40753 45004 -40747
rect 46304 -40749 46378 -40723
rect 44752 -40770 45004 -40753
rect 44757 -40794 45004 -40770
rect 45839 -40781 45974 -40773
rect 45819 -40783 45974 -40781
rect 44757 -40811 44887 -40794
rect 44931 -40807 45004 -40794
rect 45612 -40819 45974 -40783
rect 46491 -40792 47276 -40706
rect 45819 -40821 45974 -40819
rect 45839 -40827 45974 -40821
rect 46022 -40804 46441 -40796
rect 46022 -40834 46452 -40804
rect 45049 -41049 45083 -40841
rect 45245 -41049 45279 -40841
rect 45441 -41049 45475 -40841
rect 46022 -41178 46056 -40834
rect 46218 -41178 46252 -40834
rect 46391 -40983 46452 -40834
rect 46631 -40948 46665 -40792
rect 46729 -40948 46763 -40840
rect 46827 -40948 46861 -40792
rect 46925 -40948 46959 -40840
rect 46513 -40983 46586 -40977
rect 46391 -40996 46586 -40983
rect 46413 -41024 46586 -40996
rect 46513 -41037 46586 -41024
rect 47023 -41007 47395 -40937
rect 46631 -41179 46665 -41071
rect 46827 -41179 46861 -41071
rect 47023 -41179 47057 -41007
rect 45023 -42114 45057 -41770
rect 45219 -42114 45253 -41770
rect 45632 -41877 45666 -41769
rect 45828 -41877 45862 -41769
rect 45514 -41924 45587 -41911
rect 45414 -41952 45587 -41924
rect 45392 -41965 45587 -41952
rect 45392 -42114 45453 -41965
rect 45514 -41971 45587 -41965
rect 46024 -41941 46058 -41769
rect 45023 -42144 45453 -42114
rect 45023 -42152 45442 -42144
rect 45632 -42156 45666 -42000
rect 45730 -42108 45764 -42000
rect 45828 -42156 45862 -42000
rect 45926 -42108 45960 -42000
rect 46024 -42011 46302 -41941
rect 44667 -42225 44894 -42223
rect 45305 -42225 45379 -42199
rect 44667 -42263 45379 -42225
rect 45492 -42242 46107 -42156
rect 44893 -42264 45379 -42263
rect 44893 -42265 44964 -42264
rect 45305 -42270 45379 -42264
rect 44925 -42615 44959 -42307
rect 45023 -42615 45057 -42307
rect 45121 -42615 45155 -42307
rect 45219 -42615 45253 -42307
rect 45317 -42615 45351 -42307
rect 45022 -42667 45057 -42615
rect 45736 -42649 45797 -42242
rect 46226 -42406 46296 -42011
rect 46470 -42265 46504 -41681
rect 46677 -41647 46917 -41613
rect 46677 -41689 46719 -41647
rect 46466 -42324 46508 -42265
rect 46681 -42271 46715 -41689
rect 46779 -42269 46813 -41681
rect 46875 -41691 46917 -41647
rect 46678 -42324 46720 -42271
rect 46466 -42360 46720 -42324
rect 46775 -42323 46817 -42269
rect 46877 -42289 46911 -41691
rect 47089 -42275 47123 -41681
rect 46775 -42362 46916 -42323
rect 46873 -42374 46916 -42362
rect 46631 -42406 46786 -42396
rect 46226 -42442 46786 -42406
rect 46226 -42444 46296 -42442
rect 46631 -42451 46786 -42442
rect 46873 -42429 47054 -42374
rect 46873 -42499 46916 -42429
rect 46361 -42513 46516 -42504
rect 46324 -42547 46516 -42513
rect 46361 -42559 46516 -42547
rect 46562 -42539 46916 -42499
rect 47088 -42519 47131 -42275
rect 47325 -42344 47395 -41007
rect 47570 -40295 47662 -40210
rect 47593 -42270 47636 -40295
rect 47920 -40718 47996 -40014
rect 48222 -39970 50009 -39932
rect 48222 -40348 48260 -39970
rect 49429 -40269 50094 -40241
rect 49429 -40327 50464 -40269
rect 48199 -40402 48272 -40348
rect 49429 -40408 49515 -40327
rect 49689 -40364 49724 -40327
rect 50014 -40330 50464 -40327
rect 48577 -40494 49515 -40408
rect 48425 -40718 48555 -40692
rect 47920 -40784 48555 -40718
rect 48717 -40750 48751 -40494
rect 48815 -40750 48849 -40542
rect 48913 -40750 48947 -40494
rect 49011 -40716 49045 -40542
rect 49592 -40672 49626 -40364
rect 49690 -40672 49724 -40364
rect 49788 -40672 49822 -40364
rect 49886 -40672 49920 -40364
rect 49984 -40672 50018 -40364
rect 49560 -40715 49631 -40714
rect 49972 -40715 50046 -40709
rect 49560 -40716 50046 -40715
rect 49011 -40750 50046 -40716
rect 50403 -40737 50464 -40330
rect 54229 -38627 54263 -38283
rect 54425 -38627 54459 -38283
rect 54838 -38390 54872 -38282
rect 55034 -38390 55068 -38282
rect 54720 -38437 54793 -38424
rect 54620 -38465 54793 -38437
rect 54598 -38478 54793 -38465
rect 54598 -38627 54659 -38478
rect 54720 -38484 54793 -38478
rect 55230 -38454 55264 -38282
rect 54229 -38657 54659 -38627
rect 54229 -38665 54648 -38657
rect 54838 -38669 54872 -38513
rect 54936 -38621 54970 -38513
rect 55034 -38669 55068 -38513
rect 55132 -38621 55166 -38513
rect 55230 -38524 55508 -38454
rect 49012 -40754 50046 -40750
rect 49012 -40756 49561 -40754
rect 48599 -40784 48672 -40778
rect 49972 -40780 50046 -40754
rect 47920 -40794 48672 -40784
rect 48425 -40825 48672 -40794
rect 49507 -40812 49642 -40804
rect 49487 -40814 49642 -40812
rect 48425 -40842 48555 -40825
rect 48599 -40838 48672 -40825
rect 48452 -40892 48528 -40842
rect 49280 -40850 49642 -40814
rect 50159 -40823 50944 -40737
rect 49487 -40852 49642 -40850
rect 49507 -40858 49642 -40852
rect 49690 -40835 50109 -40827
rect 49690 -40865 50120 -40835
rect 48717 -41080 48751 -40872
rect 48913 -41080 48947 -40872
rect 49109 -41080 49143 -40872
rect 49690 -41209 49724 -40865
rect 49886 -41209 49920 -40865
rect 50059 -41014 50120 -40865
rect 50299 -40979 50333 -40823
rect 50397 -40979 50431 -40871
rect 50495 -40979 50529 -40823
rect 50593 -40979 50627 -40871
rect 50181 -41014 50254 -41008
rect 50059 -41027 50254 -41014
rect 50081 -41055 50254 -41027
rect 50181 -41068 50254 -41055
rect 50691 -41038 51063 -40968
rect 50299 -41210 50333 -41102
rect 50495 -41210 50529 -41102
rect 50691 -41210 50725 -41038
rect 48691 -42145 48725 -41801
rect 48887 -42145 48921 -41801
rect 49300 -41908 49334 -41800
rect 49496 -41908 49530 -41800
rect 49182 -41955 49255 -41942
rect 49082 -41983 49255 -41955
rect 49060 -41996 49255 -41983
rect 49060 -42145 49121 -41996
rect 49182 -42002 49255 -41996
rect 49692 -41972 49726 -41800
rect 48691 -42175 49121 -42145
rect 48691 -42183 49110 -42175
rect 49300 -42187 49334 -42031
rect 49398 -42139 49432 -42031
rect 49496 -42187 49530 -42031
rect 49594 -42139 49628 -42031
rect 49692 -42042 49970 -41972
rect 47593 -42313 47878 -42270
rect 47314 -42416 47419 -42344
rect 47835 -42519 47878 -42313
rect 45347 -42667 45797 -42649
rect 44905 -42710 45797 -42667
rect 44905 -42728 45354 -42710
rect 45736 -43005 45797 -42710
rect 46470 -42887 46504 -42593
rect 46562 -42609 46607 -42539
rect 46954 -42559 47878 -42519
rect 47002 -42562 47878 -42559
rect 46463 -43005 46510 -42887
rect 46568 -42901 46602 -42609
rect 46666 -42886 46700 -42593
rect 46908 -42876 46942 -42593
rect 47002 -42602 47046 -42562
rect 46659 -43005 46706 -42886
rect 46901 -43005 46948 -42876
rect 47006 -42901 47040 -42602
rect 45736 -43118 47213 -43005
rect 48335 -42256 48562 -42254
rect 48973 -42256 49047 -42230
rect 48335 -42294 49047 -42256
rect 49160 -42273 49775 -42187
rect 48561 -42295 49047 -42294
rect 48561 -42296 48632 -42295
rect 48973 -42301 49047 -42295
rect 48593 -42646 48627 -42338
rect 48691 -42646 48725 -42338
rect 48789 -42646 48823 -42338
rect 48887 -42646 48921 -42338
rect 48985 -42646 49019 -42338
rect 48690 -42698 48725 -42646
rect 49404 -42680 49465 -42273
rect 49894 -42437 49964 -42042
rect 50138 -42296 50172 -41712
rect 50345 -41678 50585 -41644
rect 50345 -41720 50387 -41678
rect 50134 -42355 50176 -42296
rect 50349 -42302 50383 -41720
rect 50447 -42300 50481 -41712
rect 50543 -41722 50585 -41678
rect 50346 -42355 50388 -42302
rect 50134 -42391 50388 -42355
rect 50443 -42354 50485 -42300
rect 50545 -42320 50579 -41722
rect 50757 -42306 50791 -41712
rect 50443 -42393 50584 -42354
rect 50541 -42405 50584 -42393
rect 50299 -42437 50454 -42427
rect 49894 -42473 50454 -42437
rect 49894 -42475 49964 -42473
rect 50299 -42482 50454 -42473
rect 50541 -42460 50722 -42405
rect 50541 -42530 50584 -42460
rect 50029 -42544 50184 -42535
rect 49992 -42578 50184 -42544
rect 50029 -42590 50184 -42578
rect 50230 -42570 50584 -42530
rect 50756 -42550 50799 -42306
rect 50993 -42375 51063 -41038
rect 50982 -42447 51087 -42375
rect 51512 -42550 51726 -42435
rect 49015 -42698 49465 -42680
rect 48573 -42741 49465 -42698
rect 48573 -42759 49022 -42741
rect 49404 -43036 49465 -42741
rect 50138 -42918 50172 -42624
rect 50230 -42640 50275 -42570
rect 50622 -42590 51824 -42550
rect 50670 -42593 51824 -42590
rect 50131 -43036 50178 -42918
rect 50236 -42932 50270 -42640
rect 50334 -42917 50368 -42624
rect 50576 -42907 50610 -42624
rect 50670 -42633 50714 -42593
rect 50327 -43036 50374 -42917
rect 50569 -43036 50616 -42907
rect 50674 -42932 50708 -42633
rect 51512 -42655 51726 -42593
rect 49404 -43149 50881 -43036
rect 42309 -44720 42549 -44711
rect 53873 -38738 54100 -38736
rect 54511 -38738 54585 -38712
rect 53873 -38776 54585 -38738
rect 54698 -38755 55313 -38669
rect 53884 -39647 53960 -38776
rect 54099 -38777 54585 -38776
rect 54099 -38778 54170 -38777
rect 54511 -38783 54585 -38777
rect 54131 -39128 54165 -38820
rect 54229 -39128 54263 -38820
rect 54327 -39128 54361 -38820
rect 54425 -39128 54459 -38820
rect 54523 -39128 54557 -38820
rect 54228 -39180 54263 -39128
rect 54942 -39162 55003 -38755
rect 55432 -38919 55502 -38524
rect 55676 -38778 55710 -38194
rect 55883 -38160 56123 -38126
rect 55883 -38202 55925 -38160
rect 55672 -38837 55714 -38778
rect 55887 -38784 55921 -38202
rect 55985 -38782 56019 -38194
rect 56081 -38204 56123 -38160
rect 55884 -38837 55926 -38784
rect 55672 -38873 55926 -38837
rect 55981 -38836 56023 -38782
rect 56083 -38802 56117 -38204
rect 56295 -38788 56329 -38194
rect 55981 -38875 56122 -38836
rect 56079 -38887 56122 -38875
rect 55837 -38919 55992 -38909
rect 55432 -38955 55992 -38919
rect 55432 -38957 55502 -38955
rect 55837 -38964 55992 -38955
rect 56079 -38942 56260 -38887
rect 56079 -39012 56122 -38942
rect 55567 -39026 55722 -39017
rect 55530 -39060 55722 -39026
rect 55567 -39072 55722 -39060
rect 55768 -39052 56122 -39012
rect 56294 -39032 56337 -38788
rect 56531 -38857 56601 -37520
rect 63009 -37496 63043 -37288
rect 63205 -37496 63239 -37288
rect 63401 -37496 63435 -37288
rect 63982 -37625 64016 -37281
rect 64178 -37625 64212 -37281
rect 64351 -37430 64412 -37281
rect 64591 -37395 64625 -37239
rect 64689 -37395 64723 -37287
rect 64787 -37395 64821 -37239
rect 71870 -37241 72000 -37224
rect 72044 -37237 72117 -37224
rect 72725 -37249 73087 -37213
rect 73604 -37222 74389 -37136
rect 81234 -37145 81364 -37053
rect 81526 -37111 81560 -36855
rect 81624 -37111 81658 -36903
rect 81722 -37111 81756 -36855
rect 81820 -37077 81854 -36903
rect 82401 -37033 82435 -36725
rect 82499 -37033 82533 -36725
rect 82597 -37033 82631 -36725
rect 82695 -37033 82729 -36725
rect 82793 -37033 82827 -36725
rect 82369 -37076 82440 -37075
rect 82781 -37076 82855 -37070
rect 82369 -37077 82855 -37076
rect 81820 -37111 82855 -37077
rect 83212 -37098 83273 -36691
rect 81821 -37115 82855 -37111
rect 81821 -37117 82370 -37115
rect 81408 -37145 81481 -37139
rect 82781 -37141 82855 -37115
rect 81234 -37186 81481 -37145
rect 82316 -37173 82451 -37165
rect 82296 -37175 82451 -37173
rect 81234 -37203 81364 -37186
rect 81408 -37199 81481 -37186
rect 82089 -37211 82451 -37175
rect 82968 -37184 83753 -37098
rect 82296 -37213 82451 -37211
rect 82316 -37219 82451 -37213
rect 82499 -37196 82918 -37188
rect 72932 -37251 73087 -37249
rect 72952 -37257 73087 -37251
rect 73135 -37234 73554 -37226
rect 73135 -37264 73565 -37234
rect 64885 -37395 64919 -37287
rect 64473 -37430 64546 -37424
rect 64351 -37443 64546 -37430
rect 64373 -37471 64546 -37443
rect 64473 -37484 64546 -37471
rect 64983 -37454 65355 -37384
rect 64591 -37626 64625 -37518
rect 64787 -37626 64821 -37518
rect 64983 -37626 65017 -37454
rect 57668 -38552 57702 -38052
rect 57847 -38016 58168 -37982
rect 57667 -38598 57702 -38552
rect 57847 -38598 57887 -38016
rect 57936 -38056 57971 -38016
rect 57937 -38560 57971 -38056
rect 58035 -38553 58069 -38052
rect 58133 -38055 58168 -38016
rect 57667 -38638 57887 -38598
rect 58032 -38673 58070 -38553
rect 58133 -38560 58167 -38055
rect 58263 -38636 58297 -38052
rect 58589 -38566 58623 -38052
rect 58817 -38342 58851 -38052
rect 58816 -38435 58853 -38342
rect 58816 -38472 58953 -38435
rect 58589 -38600 58748 -38566
rect 58412 -38636 58550 -38625
rect 57668 -38711 58070 -38673
rect 58137 -38670 58550 -38636
rect 57431 -38722 57569 -38712
rect 57041 -38756 57569 -38722
rect 56520 -38929 56625 -38857
rect 57041 -39032 57084 -38756
rect 57431 -38766 57569 -38756
rect 57487 -38857 57625 -38848
rect 57277 -38891 57625 -38857
rect 57277 -39018 57349 -38891
rect 57487 -38902 57625 -38891
rect 57277 -39027 57361 -39018
rect 54553 -39180 55003 -39162
rect 54111 -39223 55003 -39180
rect 54111 -39241 54560 -39223
rect 54942 -39518 55003 -39223
rect 55676 -39400 55710 -39106
rect 55768 -39122 55813 -39052
rect 56160 -39072 57084 -39032
rect 56208 -39075 57084 -39072
rect 55669 -39518 55716 -39400
rect 55774 -39414 55808 -39122
rect 55872 -39399 55906 -39106
rect 56114 -39389 56148 -39106
rect 56208 -39115 56252 -39075
rect 57282 -39097 57361 -39027
rect 55865 -39518 55912 -39399
rect 56107 -39518 56154 -39389
rect 56212 -39414 56246 -39115
rect 57570 -39339 57604 -39048
rect 57568 -39450 57605 -39339
rect 57668 -39356 57702 -38711
rect 57897 -38781 57935 -38711
rect 58137 -38749 58171 -38670
rect 58412 -38679 58550 -38670
rect 57887 -38919 57941 -38781
rect 58040 -38783 58171 -38749
rect 58237 -38766 58375 -38712
rect 58622 -38781 58676 -38643
rect 58714 -38644 58748 -38600
rect 58714 -38698 58880 -38644
rect 58040 -39356 58074 -38783
rect 58714 -38813 58748 -38698
rect 58800 -38813 58854 -38796
rect 58138 -38852 58297 -38817
rect 58714 -38818 58854 -38813
rect 58686 -38847 58854 -38818
rect 58138 -39356 58172 -38852
rect 58263 -39356 58297 -38852
rect 58361 -39339 58395 -38848
rect 58491 -39338 58525 -38848
rect 57031 -39454 57642 -39450
rect 58360 -39454 58397 -39339
rect 58488 -39454 58525 -39338
rect 58589 -39356 58623 -38848
rect 58686 -38852 58748 -38847
rect 58687 -39356 58721 -38852
rect 58800 -38855 58854 -38847
rect 58915 -38965 58953 -38472
rect 58915 -39003 59207 -38965
rect 58817 -39337 58851 -39048
rect 58915 -39053 58953 -39003
rect 58815 -39454 58852 -39337
rect 58915 -39356 58949 -39053
rect 57031 -39518 58965 -39454
rect 54942 -39563 58965 -39518
rect 54942 -39631 57144 -39563
rect 57492 -39615 58965 -39563
rect 53173 -39808 53960 -39647
rect 53173 -43729 53334 -39808
rect 53884 -39904 53960 -39808
rect 59169 -39898 59207 -39003
rect 53884 -39980 57194 -39904
rect 53884 -40162 53960 -39980
rect 53884 -40238 54026 -40162
rect 53950 -40627 54026 -40238
rect 54959 -40204 55624 -40176
rect 54959 -40262 55994 -40204
rect 54959 -40343 55045 -40262
rect 55219 -40299 55254 -40262
rect 55544 -40265 55994 -40262
rect 54107 -40429 55045 -40343
rect 53950 -40719 54085 -40627
rect 54247 -40685 54281 -40429
rect 54345 -40685 54379 -40477
rect 54443 -40685 54477 -40429
rect 54541 -40651 54575 -40477
rect 55122 -40607 55156 -40299
rect 55220 -40607 55254 -40299
rect 55318 -40607 55352 -40299
rect 55416 -40607 55450 -40299
rect 55514 -40607 55548 -40299
rect 55090 -40650 55161 -40649
rect 55502 -40650 55576 -40644
rect 55090 -40651 55576 -40650
rect 54541 -40685 55576 -40651
rect 55933 -40672 55994 -40265
rect 54542 -40689 55576 -40685
rect 54542 -40691 55091 -40689
rect 54129 -40719 54202 -40713
rect 55502 -40715 55576 -40689
rect 53950 -40736 54202 -40719
rect 53955 -40760 54202 -40736
rect 55037 -40747 55172 -40739
rect 55017 -40749 55172 -40747
rect 53955 -40777 54085 -40760
rect 54129 -40773 54202 -40760
rect 54810 -40785 55172 -40749
rect 55689 -40758 56474 -40672
rect 55017 -40787 55172 -40785
rect 55037 -40793 55172 -40787
rect 55220 -40770 55639 -40762
rect 55220 -40800 55650 -40770
rect 54247 -41015 54281 -40807
rect 54443 -41015 54477 -40807
rect 54639 -41015 54673 -40807
rect 55220 -41144 55254 -40800
rect 55416 -41144 55450 -40800
rect 55589 -40949 55650 -40800
rect 55829 -40914 55863 -40758
rect 55927 -40914 55961 -40806
rect 56025 -40914 56059 -40758
rect 56123 -40914 56157 -40806
rect 55711 -40949 55784 -40943
rect 55589 -40962 55784 -40949
rect 55611 -40990 55784 -40962
rect 55711 -41003 55784 -40990
rect 56221 -40973 56593 -40903
rect 55829 -41145 55863 -41037
rect 56025 -41145 56059 -41037
rect 56221 -41145 56255 -40973
rect 54221 -42080 54255 -41736
rect 54417 -42080 54451 -41736
rect 54830 -41843 54864 -41735
rect 55026 -41843 55060 -41735
rect 54712 -41890 54785 -41877
rect 54612 -41918 54785 -41890
rect 54590 -41931 54785 -41918
rect 54590 -42080 54651 -41931
rect 54712 -41937 54785 -41931
rect 55222 -41907 55256 -41735
rect 54221 -42110 54651 -42080
rect 54221 -42118 54640 -42110
rect 54830 -42122 54864 -41966
rect 54928 -42074 54962 -41966
rect 55026 -42122 55060 -41966
rect 55124 -42074 55158 -41966
rect 55222 -41977 55500 -41907
rect 53865 -42191 54092 -42189
rect 54503 -42191 54577 -42165
rect 53865 -42229 54577 -42191
rect 54690 -42208 55305 -42122
rect 54091 -42230 54577 -42229
rect 54091 -42231 54162 -42230
rect 54503 -42236 54577 -42230
rect 54123 -42581 54157 -42273
rect 54221 -42581 54255 -42273
rect 54319 -42581 54353 -42273
rect 54417 -42581 54451 -42273
rect 54515 -42581 54549 -42273
rect 54220 -42633 54255 -42581
rect 54934 -42615 54995 -42208
rect 55424 -42372 55494 -41977
rect 55668 -42231 55702 -41647
rect 55875 -41613 56115 -41579
rect 55875 -41655 55917 -41613
rect 55664 -42290 55706 -42231
rect 55879 -42237 55913 -41655
rect 55977 -42235 56011 -41647
rect 56073 -41657 56115 -41613
rect 55876 -42290 55918 -42237
rect 55664 -42326 55918 -42290
rect 55973 -42289 56015 -42235
rect 56075 -42255 56109 -41657
rect 56287 -42241 56321 -41647
rect 55973 -42328 56114 -42289
rect 56071 -42340 56114 -42328
rect 55829 -42372 55984 -42362
rect 55424 -42408 55984 -42372
rect 55424 -42410 55494 -42408
rect 55829 -42417 55984 -42408
rect 56071 -42395 56252 -42340
rect 56071 -42465 56114 -42395
rect 55559 -42479 55714 -42470
rect 55522 -42513 55714 -42479
rect 55559 -42525 55714 -42513
rect 55760 -42505 56114 -42465
rect 56286 -42485 56329 -42241
rect 56523 -42310 56593 -40973
rect 56768 -40261 56860 -40176
rect 56791 -42236 56834 -40261
rect 57118 -40684 57194 -39980
rect 57420 -39936 59207 -39898
rect 57420 -40314 57458 -39936
rect 58627 -40235 59292 -40207
rect 58627 -40293 59662 -40235
rect 57397 -40368 57470 -40314
rect 58627 -40374 58713 -40293
rect 58887 -40330 58922 -40293
rect 59212 -40296 59662 -40293
rect 57775 -40460 58713 -40374
rect 57623 -40684 57753 -40658
rect 57118 -40750 57753 -40684
rect 57915 -40716 57949 -40460
rect 58013 -40716 58047 -40508
rect 58111 -40716 58145 -40460
rect 58209 -40682 58243 -40508
rect 58790 -40638 58824 -40330
rect 58888 -40638 58922 -40330
rect 58986 -40638 59020 -40330
rect 59084 -40638 59118 -40330
rect 59182 -40638 59216 -40330
rect 58758 -40681 58829 -40680
rect 59170 -40681 59244 -40675
rect 58758 -40682 59244 -40681
rect 58209 -40716 59244 -40682
rect 59601 -40703 59662 -40296
rect 62983 -38561 63017 -38217
rect 63179 -38561 63213 -38217
rect 63592 -38324 63626 -38216
rect 63788 -38324 63822 -38216
rect 63474 -38371 63547 -38358
rect 63374 -38399 63547 -38371
rect 63352 -38412 63547 -38399
rect 63352 -38561 63413 -38412
rect 63474 -38418 63547 -38412
rect 63984 -38388 64018 -38216
rect 62983 -38591 63413 -38561
rect 62983 -38599 63402 -38591
rect 63592 -38603 63626 -38447
rect 63690 -38555 63724 -38447
rect 63788 -38603 63822 -38447
rect 63886 -38555 63920 -38447
rect 63984 -38458 64262 -38388
rect 62627 -38672 62854 -38670
rect 63265 -38672 63339 -38646
rect 58210 -40720 59244 -40716
rect 58210 -40722 58759 -40720
rect 57797 -40750 57870 -40744
rect 59170 -40746 59244 -40720
rect 57118 -40760 57870 -40750
rect 57623 -40791 57870 -40760
rect 58705 -40778 58840 -40770
rect 58685 -40780 58840 -40778
rect 57623 -40808 57753 -40791
rect 57797 -40804 57870 -40791
rect 57650 -40858 57726 -40808
rect 58478 -40816 58840 -40780
rect 59357 -40789 60142 -40703
rect 58685 -40818 58840 -40816
rect 58705 -40824 58840 -40818
rect 58888 -40801 59307 -40793
rect 58888 -40831 59318 -40801
rect 57915 -41046 57949 -40838
rect 58111 -41046 58145 -40838
rect 58307 -41046 58341 -40838
rect 58888 -41175 58922 -40831
rect 59084 -41175 59118 -40831
rect 59257 -40980 59318 -40831
rect 59497 -40945 59531 -40789
rect 59595 -40945 59629 -40837
rect 59693 -40945 59727 -40789
rect 59791 -40945 59825 -40837
rect 59379 -40980 59452 -40974
rect 59257 -40993 59452 -40980
rect 59279 -41021 59452 -40993
rect 59379 -41034 59452 -41021
rect 59889 -41004 60261 -40934
rect 59497 -41176 59531 -41068
rect 59693 -41176 59727 -41068
rect 59889 -41176 59923 -41004
rect 57889 -42111 57923 -41767
rect 58085 -42111 58119 -41767
rect 58498 -41874 58532 -41766
rect 58694 -41874 58728 -41766
rect 58380 -41921 58453 -41908
rect 58280 -41949 58453 -41921
rect 58258 -41962 58453 -41949
rect 58258 -42111 58319 -41962
rect 58380 -41968 58453 -41962
rect 58890 -41938 58924 -41766
rect 57889 -42141 58319 -42111
rect 57889 -42149 58308 -42141
rect 58498 -42153 58532 -41997
rect 58596 -42105 58630 -41997
rect 58694 -42153 58728 -41997
rect 58792 -42105 58826 -41997
rect 58890 -42008 59168 -41938
rect 56791 -42279 57076 -42236
rect 56512 -42382 56617 -42310
rect 57033 -42485 57076 -42279
rect 54545 -42633 54995 -42615
rect 54103 -42676 54995 -42633
rect 54103 -42694 54552 -42676
rect 54934 -42971 54995 -42676
rect 55668 -42853 55702 -42559
rect 55760 -42575 55805 -42505
rect 56152 -42525 57076 -42485
rect 56200 -42528 57076 -42525
rect 55661 -42971 55708 -42853
rect 55766 -42867 55800 -42575
rect 55864 -42852 55898 -42559
rect 56106 -42842 56140 -42559
rect 56200 -42568 56244 -42528
rect 55857 -42971 55904 -42852
rect 56099 -42971 56146 -42842
rect 56204 -42867 56238 -42568
rect 54934 -43084 56411 -42971
rect 57533 -42222 57760 -42220
rect 58171 -42222 58245 -42196
rect 57533 -42260 58245 -42222
rect 58358 -42239 58973 -42153
rect 57759 -42261 58245 -42260
rect 57759 -42262 57830 -42261
rect 58171 -42267 58245 -42261
rect 57791 -42612 57825 -42304
rect 57889 -42612 57923 -42304
rect 57987 -42612 58021 -42304
rect 58085 -42612 58119 -42304
rect 58183 -42612 58217 -42304
rect 57888 -42664 57923 -42612
rect 58602 -42646 58663 -42239
rect 59092 -42403 59162 -42008
rect 59336 -42262 59370 -41678
rect 59543 -41644 59783 -41610
rect 59543 -41686 59585 -41644
rect 59332 -42321 59374 -42262
rect 59547 -42268 59581 -41686
rect 59645 -42266 59679 -41678
rect 59741 -41688 59783 -41644
rect 59544 -42321 59586 -42268
rect 59332 -42357 59586 -42321
rect 59641 -42320 59683 -42266
rect 59743 -42286 59777 -41688
rect 59955 -42272 59989 -41678
rect 59641 -42359 59782 -42320
rect 59739 -42371 59782 -42359
rect 59497 -42403 59652 -42393
rect 59092 -42439 59652 -42403
rect 59092 -42441 59162 -42439
rect 59497 -42448 59652 -42439
rect 59739 -42426 59920 -42371
rect 59739 -42496 59782 -42426
rect 59227 -42510 59382 -42501
rect 59190 -42544 59382 -42510
rect 59227 -42556 59382 -42544
rect 59428 -42536 59782 -42496
rect 59954 -42516 59997 -42272
rect 60191 -42341 60261 -41004
rect 60180 -42413 60285 -42341
rect 60638 -42516 60930 -42347
rect 58213 -42664 58663 -42646
rect 57771 -42707 58663 -42664
rect 57771 -42725 58220 -42707
rect 58602 -43002 58663 -42707
rect 59336 -42884 59370 -42590
rect 59428 -42606 59473 -42536
rect 59820 -42556 61022 -42516
rect 59868 -42559 61022 -42556
rect 59329 -43002 59376 -42884
rect 59434 -42898 59468 -42606
rect 59532 -42883 59566 -42590
rect 59774 -42873 59808 -42590
rect 59868 -42599 59912 -42559
rect 59525 -43002 59572 -42883
rect 59767 -43002 59814 -42873
rect 59872 -42898 59906 -42599
rect 60638 -42646 60930 -42559
rect 58602 -43115 60079 -43002
rect 53155 -43896 53349 -43729
rect 62627 -38710 63339 -38672
rect 63452 -38689 64067 -38603
rect 62638 -39674 62714 -38710
rect 62853 -38711 63339 -38710
rect 62853 -38712 62924 -38711
rect 63265 -38717 63339 -38711
rect 62885 -39062 62919 -38754
rect 62983 -39062 63017 -38754
rect 63081 -39062 63115 -38754
rect 63179 -39062 63213 -38754
rect 63277 -39062 63311 -38754
rect 62982 -39114 63017 -39062
rect 63696 -39096 63757 -38689
rect 64186 -38853 64256 -38458
rect 64430 -38712 64464 -38128
rect 64637 -38094 64877 -38060
rect 64637 -38136 64679 -38094
rect 64426 -38771 64468 -38712
rect 64641 -38718 64675 -38136
rect 64739 -38716 64773 -38128
rect 64835 -38138 64877 -38094
rect 64638 -38771 64680 -38718
rect 64426 -38807 64680 -38771
rect 64735 -38770 64777 -38716
rect 64837 -38736 64871 -38138
rect 65049 -38722 65083 -38128
rect 64735 -38809 64876 -38770
rect 64833 -38821 64876 -38809
rect 64591 -38853 64746 -38843
rect 64186 -38889 64746 -38853
rect 64186 -38891 64256 -38889
rect 64591 -38898 64746 -38889
rect 64833 -38876 65014 -38821
rect 64833 -38946 64876 -38876
rect 64321 -38960 64476 -38951
rect 64284 -38994 64476 -38960
rect 64321 -39006 64476 -38994
rect 64522 -38986 64876 -38946
rect 65048 -38966 65091 -38722
rect 65285 -38791 65355 -37454
rect 72162 -37479 72196 -37271
rect 72358 -37479 72392 -37271
rect 72554 -37479 72588 -37271
rect 73135 -37608 73169 -37264
rect 73331 -37608 73365 -37264
rect 73504 -37413 73565 -37264
rect 73744 -37378 73778 -37222
rect 73842 -37378 73876 -37270
rect 73940 -37378 73974 -37222
rect 82499 -37226 82929 -37196
rect 74038 -37378 74072 -37270
rect 73626 -37413 73699 -37407
rect 73504 -37426 73699 -37413
rect 73526 -37454 73699 -37426
rect 73626 -37467 73699 -37454
rect 74136 -37437 74508 -37367
rect 73744 -37609 73778 -37501
rect 73940 -37609 73974 -37501
rect 74136 -37609 74170 -37437
rect 66422 -38486 66456 -37986
rect 66601 -37950 66922 -37916
rect 66421 -38532 66456 -38486
rect 66601 -38532 66641 -37950
rect 66690 -37990 66725 -37950
rect 66691 -38494 66725 -37990
rect 66789 -38487 66823 -37986
rect 66887 -37989 66922 -37950
rect 66421 -38572 66641 -38532
rect 66786 -38607 66824 -38487
rect 66887 -38494 66921 -37989
rect 67017 -38570 67051 -37986
rect 67343 -38500 67377 -37986
rect 67571 -38276 67605 -37986
rect 67570 -38369 67607 -38276
rect 67570 -38406 67707 -38369
rect 67343 -38534 67502 -38500
rect 67166 -38570 67304 -38559
rect 66422 -38645 66824 -38607
rect 66891 -38604 67304 -38570
rect 66185 -38656 66323 -38646
rect 65795 -38690 66323 -38656
rect 65274 -38863 65379 -38791
rect 65795 -38966 65838 -38690
rect 66185 -38700 66323 -38690
rect 66241 -38791 66379 -38782
rect 66031 -38825 66379 -38791
rect 66031 -38952 66103 -38825
rect 66241 -38836 66379 -38825
rect 66031 -38961 66115 -38952
rect 63307 -39114 63757 -39096
rect 62865 -39157 63757 -39114
rect 62865 -39175 63314 -39157
rect 63696 -39452 63757 -39157
rect 64430 -39334 64464 -39040
rect 64522 -39056 64567 -38986
rect 64914 -39006 65838 -38966
rect 64962 -39009 65838 -39006
rect 64423 -39452 64470 -39334
rect 64528 -39348 64562 -39056
rect 64626 -39333 64660 -39040
rect 64868 -39323 64902 -39040
rect 64962 -39049 65006 -39009
rect 66036 -39031 66115 -38961
rect 64619 -39452 64666 -39333
rect 64861 -39452 64908 -39323
rect 64966 -39348 65000 -39049
rect 66324 -39273 66358 -38982
rect 66322 -39384 66359 -39273
rect 66422 -39290 66456 -38645
rect 66651 -38715 66689 -38645
rect 66891 -38683 66925 -38604
rect 67166 -38613 67304 -38604
rect 66641 -38853 66695 -38715
rect 66794 -38717 66925 -38683
rect 66991 -38700 67129 -38646
rect 67376 -38715 67430 -38577
rect 67468 -38578 67502 -38534
rect 67468 -38632 67634 -38578
rect 66794 -39290 66828 -38717
rect 67468 -38747 67502 -38632
rect 67554 -38747 67608 -38730
rect 66892 -38786 67051 -38751
rect 67468 -38752 67608 -38747
rect 67440 -38781 67608 -38752
rect 66892 -39290 66926 -38786
rect 67017 -39290 67051 -38786
rect 67115 -39273 67149 -38782
rect 67245 -39272 67279 -38782
rect 65785 -39388 66396 -39384
rect 67114 -39388 67151 -39273
rect 67242 -39388 67279 -39272
rect 67343 -39290 67377 -38782
rect 67440 -38786 67502 -38781
rect 67441 -39290 67475 -38786
rect 67554 -38789 67608 -38781
rect 67669 -38899 67707 -38406
rect 67669 -38937 67961 -38899
rect 67571 -39271 67605 -38982
rect 67669 -38987 67707 -38937
rect 67569 -39388 67606 -39271
rect 67669 -39290 67703 -38987
rect 65785 -39452 67719 -39388
rect 63696 -39497 67719 -39452
rect 63696 -39565 65898 -39497
rect 66246 -39549 67719 -39497
rect 61925 -39838 62714 -39674
rect 67923 -39832 67961 -38937
rect 61925 -39891 65948 -39838
rect 61925 -44461 62142 -39891
rect 62638 -39914 65948 -39891
rect 62638 -40096 62714 -39914
rect 62638 -40172 62780 -40096
rect 62704 -40561 62780 -40172
rect 63713 -40138 64378 -40110
rect 63713 -40196 64748 -40138
rect 63713 -40277 63799 -40196
rect 63973 -40233 64008 -40196
rect 64298 -40199 64748 -40196
rect 62861 -40363 63799 -40277
rect 62704 -40653 62839 -40561
rect 63001 -40619 63035 -40363
rect 63099 -40619 63133 -40411
rect 63197 -40619 63231 -40363
rect 63295 -40585 63329 -40411
rect 63876 -40541 63910 -40233
rect 63974 -40541 64008 -40233
rect 64072 -40541 64106 -40233
rect 64170 -40541 64204 -40233
rect 64268 -40541 64302 -40233
rect 63844 -40584 63915 -40583
rect 64256 -40584 64330 -40578
rect 63844 -40585 64330 -40584
rect 63295 -40619 64330 -40585
rect 64687 -40606 64748 -40199
rect 63296 -40623 64330 -40619
rect 63296 -40625 63845 -40623
rect 62883 -40653 62956 -40647
rect 64256 -40649 64330 -40623
rect 62704 -40670 62956 -40653
rect 62709 -40694 62956 -40670
rect 63791 -40681 63926 -40673
rect 63771 -40683 63926 -40681
rect 62709 -40711 62839 -40694
rect 62883 -40707 62956 -40694
rect 63564 -40719 63926 -40683
rect 64443 -40692 65228 -40606
rect 63771 -40721 63926 -40719
rect 63791 -40727 63926 -40721
rect 63974 -40704 64393 -40696
rect 63974 -40734 64404 -40704
rect 63001 -40949 63035 -40741
rect 63197 -40949 63231 -40741
rect 63393 -40949 63427 -40741
rect 63974 -41078 64008 -40734
rect 64170 -41078 64204 -40734
rect 64343 -40883 64404 -40734
rect 64583 -40848 64617 -40692
rect 64681 -40848 64715 -40740
rect 64779 -40848 64813 -40692
rect 64877 -40848 64911 -40740
rect 64465 -40883 64538 -40877
rect 64343 -40896 64538 -40883
rect 64365 -40924 64538 -40896
rect 64465 -40937 64538 -40924
rect 64975 -40907 65347 -40837
rect 64583 -41079 64617 -40971
rect 64779 -41079 64813 -40971
rect 64975 -41079 65009 -40907
rect 62975 -42014 63009 -41670
rect 63171 -42014 63205 -41670
rect 63584 -41777 63618 -41669
rect 63780 -41777 63814 -41669
rect 63466 -41824 63539 -41811
rect 63366 -41852 63539 -41824
rect 63344 -41865 63539 -41852
rect 63344 -42014 63405 -41865
rect 63466 -41871 63539 -41865
rect 63976 -41841 64010 -41669
rect 62792 -42027 62927 -42021
rect 62772 -42029 62927 -42027
rect 62244 -42065 62927 -42029
rect 62975 -42044 63405 -42014
rect 62975 -42052 63394 -42044
rect 63584 -42056 63618 -41900
rect 63682 -42008 63716 -41900
rect 63780 -42056 63814 -41900
rect 63878 -42008 63912 -41900
rect 63976 -41911 64254 -41841
rect 62427 -43092 62563 -42065
rect 62772 -42067 62927 -42065
rect 62792 -42075 62927 -42067
rect 62619 -42125 62846 -42123
rect 63257 -42125 63331 -42099
rect 62619 -42163 63331 -42125
rect 63444 -42142 64059 -42056
rect 62845 -42164 63331 -42163
rect 62845 -42165 62916 -42164
rect 63257 -42170 63331 -42164
rect 62877 -42515 62911 -42207
rect 62975 -42515 63009 -42207
rect 63073 -42515 63107 -42207
rect 63171 -42515 63205 -42207
rect 63269 -42515 63303 -42207
rect 62974 -42567 63009 -42515
rect 63688 -42549 63749 -42142
rect 64178 -42306 64248 -41911
rect 64422 -42165 64456 -41581
rect 64629 -41547 64869 -41513
rect 64629 -41589 64671 -41547
rect 64418 -42224 64460 -42165
rect 64633 -42171 64667 -41589
rect 64731 -42169 64765 -41581
rect 64827 -41591 64869 -41547
rect 64630 -42224 64672 -42171
rect 64418 -42260 64672 -42224
rect 64727 -42223 64769 -42169
rect 64829 -42189 64863 -41591
rect 65041 -42175 65075 -41581
rect 64727 -42262 64868 -42223
rect 64825 -42274 64868 -42262
rect 64583 -42306 64738 -42296
rect 64178 -42342 64738 -42306
rect 64178 -42344 64248 -42342
rect 64583 -42351 64738 -42342
rect 64825 -42329 65006 -42274
rect 64825 -42399 64868 -42329
rect 64313 -42413 64468 -42404
rect 64276 -42447 64468 -42413
rect 64313 -42459 64468 -42447
rect 64514 -42439 64868 -42399
rect 65040 -42419 65083 -42175
rect 65277 -42244 65347 -40907
rect 65522 -40195 65614 -40110
rect 65545 -42170 65588 -40195
rect 65872 -40618 65948 -39914
rect 66174 -39870 67961 -39832
rect 66174 -40248 66212 -39870
rect 67381 -40169 68046 -40141
rect 67381 -40227 68416 -40169
rect 66151 -40302 66224 -40248
rect 67381 -40308 67467 -40227
rect 67641 -40264 67676 -40227
rect 67966 -40230 68416 -40227
rect 66529 -40394 67467 -40308
rect 66377 -40618 66507 -40592
rect 65872 -40684 66507 -40618
rect 66669 -40650 66703 -40394
rect 66767 -40650 66801 -40442
rect 66865 -40650 66899 -40394
rect 66963 -40616 66997 -40442
rect 67544 -40572 67578 -40264
rect 67642 -40572 67676 -40264
rect 67740 -40572 67774 -40264
rect 67838 -40572 67872 -40264
rect 67936 -40572 67970 -40264
rect 67512 -40615 67583 -40614
rect 67924 -40615 67998 -40609
rect 67512 -40616 67998 -40615
rect 66963 -40650 67998 -40616
rect 68355 -40637 68416 -40230
rect 72136 -38544 72170 -38200
rect 72332 -38544 72366 -38200
rect 72745 -38307 72779 -38199
rect 72941 -38307 72975 -38199
rect 72627 -38354 72700 -38341
rect 72527 -38382 72700 -38354
rect 72505 -38395 72700 -38382
rect 72505 -38544 72566 -38395
rect 72627 -38401 72700 -38395
rect 73137 -38371 73171 -38199
rect 72136 -38574 72566 -38544
rect 72136 -38582 72555 -38574
rect 72745 -38586 72779 -38430
rect 72843 -38538 72877 -38430
rect 72941 -38586 72975 -38430
rect 73039 -38538 73073 -38430
rect 73137 -38441 73415 -38371
rect 71780 -38655 72007 -38653
rect 72418 -38655 72492 -38629
rect 66964 -40654 67998 -40650
rect 66964 -40656 67513 -40654
rect 66551 -40684 66624 -40678
rect 67924 -40680 67998 -40654
rect 65872 -40694 66624 -40684
rect 66377 -40725 66624 -40694
rect 67459 -40712 67594 -40704
rect 67439 -40714 67594 -40712
rect 66377 -40742 66507 -40725
rect 66551 -40738 66624 -40725
rect 66404 -40792 66480 -40742
rect 67232 -40750 67594 -40714
rect 68111 -40723 68896 -40637
rect 67439 -40752 67594 -40750
rect 67459 -40758 67594 -40752
rect 67642 -40735 68061 -40727
rect 67642 -40765 68072 -40735
rect 66669 -40980 66703 -40772
rect 66865 -40980 66899 -40772
rect 67061 -40980 67095 -40772
rect 67642 -41109 67676 -40765
rect 67838 -41109 67872 -40765
rect 68011 -40914 68072 -40765
rect 68251 -40879 68285 -40723
rect 68349 -40879 68383 -40771
rect 68447 -40879 68481 -40723
rect 68545 -40879 68579 -40771
rect 68133 -40914 68206 -40908
rect 68011 -40927 68206 -40914
rect 68033 -40955 68206 -40927
rect 68133 -40968 68206 -40955
rect 68643 -40938 69015 -40868
rect 68251 -41110 68285 -41002
rect 68447 -41110 68481 -41002
rect 68643 -41110 68677 -40938
rect 66643 -42045 66677 -41701
rect 66839 -42045 66873 -41701
rect 67252 -41808 67286 -41700
rect 67448 -41808 67482 -41700
rect 67134 -41855 67207 -41842
rect 67034 -41883 67207 -41855
rect 67012 -41896 67207 -41883
rect 67012 -42045 67073 -41896
rect 67134 -41902 67207 -41896
rect 67644 -41872 67678 -41700
rect 66460 -42058 66595 -42052
rect 66440 -42060 66595 -42058
rect 66026 -42096 66595 -42060
rect 66643 -42075 67073 -42045
rect 66643 -42083 67062 -42075
rect 67252 -42087 67286 -41931
rect 67350 -42039 67384 -41931
rect 67448 -42087 67482 -41931
rect 67546 -42039 67580 -41931
rect 67644 -41942 67922 -41872
rect 65545 -42213 65830 -42170
rect 65266 -42316 65371 -42244
rect 65787 -42419 65830 -42213
rect 63299 -42567 63749 -42549
rect 62857 -42610 63749 -42567
rect 62857 -42628 63306 -42610
rect 63688 -42905 63749 -42610
rect 64422 -42787 64456 -42493
rect 64514 -42509 64559 -42439
rect 64906 -42459 65830 -42419
rect 64954 -42462 65830 -42459
rect 64415 -42905 64462 -42787
rect 64520 -42801 64554 -42509
rect 64618 -42786 64652 -42493
rect 64860 -42776 64894 -42493
rect 64954 -42502 64998 -42462
rect 64611 -42905 64658 -42786
rect 64853 -42905 64900 -42776
rect 64958 -42801 64992 -42502
rect 63688 -43018 65165 -42905
rect 66026 -43092 66162 -42096
rect 66440 -42098 66595 -42096
rect 66460 -42106 66595 -42098
rect 66287 -42156 66514 -42154
rect 66925 -42156 66999 -42130
rect 66287 -42194 66999 -42156
rect 67112 -42173 67727 -42087
rect 66513 -42195 66999 -42194
rect 66513 -42196 66584 -42195
rect 66925 -42201 66999 -42195
rect 66545 -42546 66579 -42238
rect 66643 -42546 66677 -42238
rect 66741 -42546 66775 -42238
rect 66839 -42546 66873 -42238
rect 66937 -42546 66971 -42238
rect 66642 -42598 66677 -42546
rect 67356 -42580 67417 -42173
rect 67846 -42337 67916 -41942
rect 68090 -42196 68124 -41612
rect 68297 -41578 68537 -41544
rect 68297 -41620 68339 -41578
rect 68086 -42255 68128 -42196
rect 68301 -42202 68335 -41620
rect 68399 -42200 68433 -41612
rect 68495 -41622 68537 -41578
rect 68298 -42255 68340 -42202
rect 68086 -42291 68340 -42255
rect 68395 -42254 68437 -42200
rect 68497 -42220 68531 -41622
rect 68709 -42206 68743 -41612
rect 68395 -42293 68536 -42254
rect 68493 -42305 68536 -42293
rect 68251 -42337 68406 -42327
rect 67846 -42373 68406 -42337
rect 67846 -42375 67916 -42373
rect 68251 -42382 68406 -42373
rect 68493 -42360 68674 -42305
rect 68493 -42430 68536 -42360
rect 67981 -42444 68136 -42435
rect 67944 -42478 68136 -42444
rect 67981 -42490 68136 -42478
rect 68182 -42470 68536 -42430
rect 68708 -42450 68751 -42206
rect 68945 -42275 69015 -40938
rect 68934 -42347 69039 -42275
rect 69403 -42450 69664 -42289
rect 66967 -42598 67417 -42580
rect 66525 -42641 67417 -42598
rect 66525 -42659 66974 -42641
rect 67356 -42936 67417 -42641
rect 68090 -42818 68124 -42524
rect 68182 -42540 68227 -42470
rect 68574 -42490 69776 -42450
rect 68622 -42493 69776 -42490
rect 68083 -42936 68130 -42818
rect 68188 -42832 68222 -42540
rect 68286 -42817 68320 -42524
rect 68528 -42807 68562 -42524
rect 68622 -42533 68666 -42493
rect 68279 -42936 68326 -42817
rect 68521 -42936 68568 -42807
rect 68626 -42832 68660 -42533
rect 69403 -42593 69664 -42493
rect 67356 -43049 68833 -42936
rect 62427 -43228 66162 -43092
rect 61868 -44744 62212 -44461
rect 8987 -45477 9123 -45475
rect 62427 -45477 62563 -43228
rect 71780 -38693 72492 -38655
rect 72605 -38672 73220 -38586
rect 71791 -39715 71867 -38693
rect 72006 -38694 72492 -38693
rect 72006 -38695 72077 -38694
rect 72418 -38700 72492 -38694
rect 72038 -39045 72072 -38737
rect 72136 -39045 72170 -38737
rect 72234 -39045 72268 -38737
rect 72332 -39045 72366 -38737
rect 72430 -39045 72464 -38737
rect 72135 -39097 72170 -39045
rect 72849 -39079 72910 -38672
rect 73339 -38836 73409 -38441
rect 73583 -38695 73617 -38111
rect 73790 -38077 74030 -38043
rect 73790 -38119 73832 -38077
rect 73579 -38754 73621 -38695
rect 73794 -38701 73828 -38119
rect 73892 -38699 73926 -38111
rect 73988 -38121 74030 -38077
rect 73791 -38754 73833 -38701
rect 73579 -38790 73833 -38754
rect 73888 -38753 73930 -38699
rect 73990 -38719 74024 -38121
rect 74202 -38705 74236 -38111
rect 73888 -38792 74029 -38753
rect 73986 -38804 74029 -38792
rect 73744 -38836 73899 -38826
rect 73339 -38872 73899 -38836
rect 73339 -38874 73409 -38872
rect 73744 -38881 73899 -38872
rect 73986 -38859 74167 -38804
rect 73986 -38929 74029 -38859
rect 73474 -38943 73629 -38934
rect 73437 -38977 73629 -38943
rect 73474 -38989 73629 -38977
rect 73675 -38969 74029 -38929
rect 74201 -38949 74244 -38705
rect 74438 -38774 74508 -37437
rect 81526 -37441 81560 -37233
rect 81722 -37441 81756 -37233
rect 81918 -37441 81952 -37233
rect 82499 -37570 82533 -37226
rect 82695 -37570 82729 -37226
rect 82868 -37375 82929 -37226
rect 83108 -37340 83142 -37184
rect 83206 -37340 83240 -37232
rect 83304 -37340 83338 -37184
rect 83402 -37340 83436 -37232
rect 82990 -37375 83063 -37369
rect 82868 -37388 83063 -37375
rect 82890 -37416 83063 -37388
rect 82990 -37429 83063 -37416
rect 83500 -37399 83872 -37329
rect 83108 -37571 83142 -37463
rect 83304 -37571 83338 -37463
rect 83500 -37571 83534 -37399
rect 75575 -38469 75609 -37969
rect 75754 -37933 76075 -37899
rect 75574 -38515 75609 -38469
rect 75754 -38515 75794 -37933
rect 75843 -37973 75878 -37933
rect 75844 -38477 75878 -37973
rect 75942 -38470 75976 -37969
rect 76040 -37972 76075 -37933
rect 75574 -38555 75794 -38515
rect 75939 -38590 75977 -38470
rect 76040 -38477 76074 -37972
rect 76170 -38553 76204 -37969
rect 76496 -38483 76530 -37969
rect 76724 -38259 76758 -37969
rect 76723 -38352 76760 -38259
rect 76723 -38389 76860 -38352
rect 76496 -38517 76655 -38483
rect 76319 -38553 76457 -38542
rect 75575 -38628 75977 -38590
rect 76044 -38587 76457 -38553
rect 75338 -38639 75476 -38629
rect 74948 -38673 75476 -38639
rect 74427 -38846 74532 -38774
rect 74948 -38949 74991 -38673
rect 75338 -38683 75476 -38673
rect 75394 -38774 75532 -38765
rect 75184 -38808 75532 -38774
rect 75184 -38935 75256 -38808
rect 75394 -38819 75532 -38808
rect 75184 -38944 75268 -38935
rect 72460 -39097 72910 -39079
rect 72018 -39140 72910 -39097
rect 72018 -39158 72467 -39140
rect 72849 -39435 72910 -39140
rect 73583 -39317 73617 -39023
rect 73675 -39039 73720 -38969
rect 74067 -38989 74991 -38949
rect 74115 -38992 74991 -38989
rect 73576 -39435 73623 -39317
rect 73681 -39331 73715 -39039
rect 73779 -39316 73813 -39023
rect 74021 -39306 74055 -39023
rect 74115 -39032 74159 -38992
rect 75189 -39014 75268 -38944
rect 73772 -39435 73819 -39316
rect 74014 -39435 74061 -39306
rect 74119 -39331 74153 -39032
rect 75477 -39256 75511 -38965
rect 75475 -39367 75512 -39256
rect 75575 -39273 75609 -38628
rect 75804 -38698 75842 -38628
rect 76044 -38666 76078 -38587
rect 76319 -38596 76457 -38587
rect 75794 -38836 75848 -38698
rect 75947 -38700 76078 -38666
rect 76144 -38683 76282 -38629
rect 76529 -38698 76583 -38560
rect 76621 -38561 76655 -38517
rect 76621 -38615 76787 -38561
rect 75947 -39273 75981 -38700
rect 76621 -38730 76655 -38615
rect 76707 -38730 76761 -38713
rect 76045 -38769 76204 -38734
rect 76621 -38735 76761 -38730
rect 76593 -38764 76761 -38735
rect 76045 -39273 76079 -38769
rect 76170 -39273 76204 -38769
rect 76268 -39256 76302 -38765
rect 76398 -39255 76432 -38765
rect 74938 -39371 75549 -39367
rect 76267 -39371 76304 -39256
rect 76395 -39371 76432 -39255
rect 76496 -39273 76530 -38765
rect 76593 -38769 76655 -38764
rect 76594 -39273 76628 -38769
rect 76707 -38772 76761 -38764
rect 76822 -38882 76860 -38389
rect 76822 -38920 77114 -38882
rect 76724 -39254 76758 -38965
rect 76822 -38970 76860 -38920
rect 76722 -39371 76759 -39254
rect 76822 -39273 76856 -38970
rect 74938 -39435 76872 -39371
rect 72849 -39480 76872 -39435
rect 72849 -39548 75051 -39480
rect 75399 -39532 76872 -39480
rect 71116 -39821 71867 -39715
rect 77076 -39815 77114 -38920
rect 71116 -39885 75101 -39821
rect 71116 -43721 71286 -39885
rect 71791 -39897 75101 -39885
rect 71791 -40079 71867 -39897
rect 71791 -40155 71933 -40079
rect 71857 -40544 71933 -40155
rect 72866 -40121 73531 -40093
rect 72866 -40179 73901 -40121
rect 72866 -40260 72952 -40179
rect 73126 -40216 73161 -40179
rect 73451 -40182 73901 -40179
rect 72014 -40346 72952 -40260
rect 71857 -40636 71992 -40544
rect 72154 -40602 72188 -40346
rect 72252 -40602 72286 -40394
rect 72350 -40602 72384 -40346
rect 72448 -40568 72482 -40394
rect 73029 -40524 73063 -40216
rect 73127 -40524 73161 -40216
rect 73225 -40524 73259 -40216
rect 73323 -40524 73357 -40216
rect 73421 -40524 73455 -40216
rect 72997 -40567 73068 -40566
rect 73409 -40567 73483 -40561
rect 72997 -40568 73483 -40567
rect 72448 -40602 73483 -40568
rect 73840 -40589 73901 -40182
rect 72449 -40606 73483 -40602
rect 72449 -40608 72998 -40606
rect 72036 -40636 72109 -40630
rect 73409 -40632 73483 -40606
rect 71857 -40653 72109 -40636
rect 71862 -40677 72109 -40653
rect 72944 -40664 73079 -40656
rect 72924 -40666 73079 -40664
rect 71862 -40694 71992 -40677
rect 72036 -40690 72109 -40677
rect 72717 -40702 73079 -40666
rect 73596 -40675 74381 -40589
rect 72924 -40704 73079 -40702
rect 72944 -40710 73079 -40704
rect 73127 -40687 73546 -40679
rect 73127 -40717 73557 -40687
rect 72154 -40932 72188 -40724
rect 72350 -40932 72384 -40724
rect 72546 -40932 72580 -40724
rect 73127 -41061 73161 -40717
rect 73323 -41061 73357 -40717
rect 73496 -40866 73557 -40717
rect 73736 -40831 73770 -40675
rect 73834 -40831 73868 -40723
rect 73932 -40831 73966 -40675
rect 74030 -40831 74064 -40723
rect 73618 -40866 73691 -40860
rect 73496 -40879 73691 -40866
rect 73518 -40907 73691 -40879
rect 73618 -40920 73691 -40907
rect 74128 -40890 74500 -40820
rect 73736 -41062 73770 -40954
rect 73932 -41062 73966 -40954
rect 74128 -41062 74162 -40890
rect 72128 -41997 72162 -41653
rect 72324 -41997 72358 -41653
rect 72737 -41760 72771 -41652
rect 72933 -41760 72967 -41652
rect 72619 -41807 72692 -41794
rect 72519 -41835 72692 -41807
rect 72497 -41848 72692 -41835
rect 72497 -41997 72558 -41848
rect 72619 -41854 72692 -41848
rect 73129 -41824 73163 -41652
rect 71945 -42010 72080 -42004
rect 71925 -42012 72080 -42010
rect 71397 -42048 72080 -42012
rect 72128 -42027 72558 -41997
rect 72128 -42035 72547 -42027
rect 72737 -42039 72771 -41883
rect 72835 -41991 72869 -41883
rect 72933 -42039 72967 -41883
rect 73031 -41991 73065 -41883
rect 73129 -41894 73407 -41824
rect 71580 -43075 71716 -42048
rect 71925 -42050 72080 -42048
rect 71945 -42058 72080 -42050
rect 71772 -42108 71999 -42106
rect 72410 -42108 72484 -42082
rect 71772 -42146 72484 -42108
rect 72597 -42125 73212 -42039
rect 71998 -42147 72484 -42146
rect 71998 -42148 72069 -42147
rect 72410 -42153 72484 -42147
rect 72030 -42498 72064 -42190
rect 72128 -42498 72162 -42190
rect 72226 -42498 72260 -42190
rect 72324 -42498 72358 -42190
rect 72422 -42498 72456 -42190
rect 72127 -42550 72162 -42498
rect 72841 -42532 72902 -42125
rect 73331 -42289 73401 -41894
rect 73575 -42148 73609 -41564
rect 73782 -41530 74022 -41496
rect 73782 -41572 73824 -41530
rect 73571 -42207 73613 -42148
rect 73786 -42154 73820 -41572
rect 73884 -42152 73918 -41564
rect 73980 -41574 74022 -41530
rect 73783 -42207 73825 -42154
rect 73571 -42243 73825 -42207
rect 73880 -42206 73922 -42152
rect 73982 -42172 74016 -41574
rect 74194 -42158 74228 -41564
rect 73880 -42245 74021 -42206
rect 73978 -42257 74021 -42245
rect 73736 -42289 73891 -42279
rect 73331 -42325 73891 -42289
rect 73331 -42327 73401 -42325
rect 73736 -42334 73891 -42325
rect 73978 -42312 74159 -42257
rect 73978 -42382 74021 -42312
rect 73466 -42396 73621 -42387
rect 73429 -42430 73621 -42396
rect 73466 -42442 73621 -42430
rect 73667 -42422 74021 -42382
rect 74193 -42402 74236 -42158
rect 74430 -42227 74500 -40890
rect 74675 -40178 74767 -40093
rect 74698 -42153 74741 -40178
rect 75025 -40601 75101 -39897
rect 75327 -39853 77114 -39815
rect 75327 -40231 75365 -39853
rect 76534 -40152 77199 -40124
rect 76534 -40210 77569 -40152
rect 75304 -40285 75377 -40231
rect 76534 -40291 76620 -40210
rect 76794 -40247 76829 -40210
rect 77119 -40213 77569 -40210
rect 75682 -40377 76620 -40291
rect 75530 -40601 75660 -40575
rect 75025 -40667 75660 -40601
rect 75822 -40633 75856 -40377
rect 75920 -40633 75954 -40425
rect 76018 -40633 76052 -40377
rect 76116 -40599 76150 -40425
rect 76697 -40555 76731 -40247
rect 76795 -40555 76829 -40247
rect 76893 -40555 76927 -40247
rect 76991 -40555 77025 -40247
rect 77089 -40555 77123 -40247
rect 76665 -40598 76736 -40597
rect 77077 -40598 77151 -40592
rect 76665 -40599 77151 -40598
rect 76116 -40633 77151 -40599
rect 77508 -40620 77569 -40213
rect 81500 -38506 81534 -38162
rect 81696 -38506 81730 -38162
rect 82109 -38269 82143 -38161
rect 82305 -38269 82339 -38161
rect 81991 -38316 82064 -38303
rect 81891 -38344 82064 -38316
rect 81869 -38357 82064 -38344
rect 81869 -38506 81930 -38357
rect 81991 -38363 82064 -38357
rect 82501 -38333 82535 -38161
rect 81500 -38536 81930 -38506
rect 81500 -38544 81919 -38536
rect 82109 -38548 82143 -38392
rect 82207 -38500 82241 -38392
rect 82305 -38548 82339 -38392
rect 82403 -38500 82437 -38392
rect 82501 -38403 82779 -38333
rect 81144 -38617 81371 -38615
rect 81782 -38617 81856 -38591
rect 76117 -40637 77151 -40633
rect 76117 -40639 76666 -40637
rect 75704 -40667 75777 -40661
rect 77077 -40663 77151 -40637
rect 75025 -40677 75777 -40667
rect 75530 -40708 75777 -40677
rect 76612 -40695 76747 -40687
rect 76592 -40697 76747 -40695
rect 75530 -40725 75660 -40708
rect 75704 -40721 75777 -40708
rect 75557 -40775 75633 -40725
rect 76385 -40733 76747 -40697
rect 77264 -40706 78049 -40620
rect 76592 -40735 76747 -40733
rect 76612 -40741 76747 -40735
rect 76795 -40718 77214 -40710
rect 76795 -40748 77225 -40718
rect 75822 -40963 75856 -40755
rect 76018 -40963 76052 -40755
rect 76214 -40963 76248 -40755
rect 76795 -41092 76829 -40748
rect 76991 -41092 77025 -40748
rect 77164 -40897 77225 -40748
rect 77404 -40862 77438 -40706
rect 77502 -40862 77536 -40754
rect 77600 -40862 77634 -40706
rect 77698 -40862 77732 -40754
rect 77286 -40897 77359 -40891
rect 77164 -40910 77359 -40897
rect 77186 -40938 77359 -40910
rect 77286 -40951 77359 -40938
rect 77796 -40921 78168 -40851
rect 77404 -41093 77438 -40985
rect 77600 -41093 77634 -40985
rect 77796 -41093 77830 -40921
rect 75796 -42028 75830 -41684
rect 75992 -42028 76026 -41684
rect 76405 -41791 76439 -41683
rect 76601 -41791 76635 -41683
rect 76287 -41838 76360 -41825
rect 76187 -41866 76360 -41838
rect 76165 -41879 76360 -41866
rect 76165 -42028 76226 -41879
rect 76287 -41885 76360 -41879
rect 76797 -41855 76831 -41683
rect 75613 -42041 75748 -42035
rect 75593 -42043 75748 -42041
rect 75179 -42079 75748 -42043
rect 75796 -42058 76226 -42028
rect 75796 -42066 76215 -42058
rect 76405 -42070 76439 -41914
rect 76503 -42022 76537 -41914
rect 76601 -42070 76635 -41914
rect 76699 -42022 76733 -41914
rect 76797 -41925 77075 -41855
rect 74698 -42196 74983 -42153
rect 74419 -42299 74524 -42227
rect 74940 -42402 74983 -42196
rect 72452 -42550 72902 -42532
rect 72010 -42593 72902 -42550
rect 72010 -42611 72459 -42593
rect 72841 -42888 72902 -42593
rect 73575 -42770 73609 -42476
rect 73667 -42492 73712 -42422
rect 74059 -42442 74983 -42402
rect 74107 -42445 74983 -42442
rect 73568 -42888 73615 -42770
rect 73673 -42784 73707 -42492
rect 73771 -42769 73805 -42476
rect 74013 -42759 74047 -42476
rect 74107 -42485 74151 -42445
rect 73764 -42888 73811 -42769
rect 74006 -42888 74053 -42759
rect 74111 -42784 74145 -42485
rect 72841 -43001 74318 -42888
rect 75179 -43075 75315 -42079
rect 75593 -42081 75748 -42079
rect 75613 -42089 75748 -42081
rect 75440 -42139 75667 -42137
rect 76078 -42139 76152 -42113
rect 75440 -42177 76152 -42139
rect 76265 -42156 76880 -42070
rect 75666 -42178 76152 -42177
rect 75666 -42179 75737 -42178
rect 76078 -42184 76152 -42178
rect 75698 -42529 75732 -42221
rect 75796 -42529 75830 -42221
rect 75894 -42529 75928 -42221
rect 75992 -42529 76026 -42221
rect 76090 -42529 76124 -42221
rect 75795 -42581 75830 -42529
rect 76509 -42563 76570 -42156
rect 76999 -42320 77069 -41925
rect 77243 -42179 77277 -41595
rect 77450 -41561 77690 -41527
rect 77450 -41603 77492 -41561
rect 77239 -42238 77281 -42179
rect 77454 -42185 77488 -41603
rect 77552 -42183 77586 -41595
rect 77648 -41605 77690 -41561
rect 77451 -42238 77493 -42185
rect 77239 -42274 77493 -42238
rect 77548 -42237 77590 -42183
rect 77650 -42203 77684 -41605
rect 77862 -42189 77896 -41595
rect 77548 -42276 77689 -42237
rect 77646 -42288 77689 -42276
rect 77404 -42320 77559 -42310
rect 76999 -42356 77559 -42320
rect 76999 -42358 77069 -42356
rect 77404 -42365 77559 -42356
rect 77646 -42343 77827 -42288
rect 77646 -42413 77689 -42343
rect 77134 -42427 77289 -42418
rect 77097 -42461 77289 -42427
rect 77134 -42473 77289 -42461
rect 77335 -42453 77689 -42413
rect 77861 -42433 77904 -42189
rect 78098 -42258 78168 -40921
rect 78087 -42330 78192 -42258
rect 78689 -42433 78791 -42395
rect 76120 -42581 76570 -42563
rect 75678 -42624 76570 -42581
rect 75678 -42642 76127 -42624
rect 76509 -42919 76570 -42624
rect 77243 -42801 77277 -42507
rect 77335 -42523 77380 -42453
rect 77727 -42473 78929 -42433
rect 77775 -42476 78929 -42473
rect 77236 -42919 77283 -42801
rect 77341 -42815 77375 -42523
rect 77439 -42800 77473 -42507
rect 77681 -42790 77715 -42507
rect 77775 -42516 77819 -42476
rect 78689 -42506 78791 -42476
rect 77432 -42919 77479 -42800
rect 77674 -42919 77721 -42790
rect 77779 -42815 77813 -42516
rect 76509 -43032 77986 -42919
rect 71580 -43211 75315 -43075
rect 71077 -43901 71323 -43721
rect -24214 -45613 62563 -45477
rect -24214 -45618 -22243 -45613
rect -24214 -45776 -24078 -45618
rect 71580 -45776 71716 -43211
rect 81144 -38655 81856 -38617
rect 81969 -38634 82584 -38548
rect 81155 -39636 81231 -38655
rect 81370 -38656 81856 -38655
rect 81370 -38657 81441 -38656
rect 81782 -38662 81856 -38656
rect 81402 -39007 81436 -38699
rect 81500 -39007 81534 -38699
rect 81598 -39007 81632 -38699
rect 81696 -39007 81730 -38699
rect 81794 -39007 81828 -38699
rect 81499 -39059 81534 -39007
rect 82213 -39041 82274 -38634
rect 82703 -38798 82773 -38403
rect 82947 -38657 82981 -38073
rect 83154 -38039 83394 -38005
rect 83154 -38081 83196 -38039
rect 82943 -38716 82985 -38657
rect 83158 -38663 83192 -38081
rect 83256 -38661 83290 -38073
rect 83352 -38083 83394 -38039
rect 83155 -38716 83197 -38663
rect 82943 -38752 83197 -38716
rect 83252 -38715 83294 -38661
rect 83354 -38681 83388 -38083
rect 83566 -38667 83600 -38073
rect 83252 -38754 83393 -38715
rect 83350 -38766 83393 -38754
rect 83108 -38798 83263 -38788
rect 82703 -38834 83263 -38798
rect 82703 -38836 82773 -38834
rect 83108 -38843 83263 -38834
rect 83350 -38821 83531 -38766
rect 83350 -38891 83393 -38821
rect 82838 -38905 82993 -38896
rect 82801 -38939 82993 -38905
rect 82838 -38951 82993 -38939
rect 83039 -38931 83393 -38891
rect 83565 -38911 83608 -38667
rect 83802 -38736 83872 -37399
rect 84939 -38431 84973 -37931
rect 85118 -37895 85439 -37861
rect 84938 -38477 84973 -38431
rect 85118 -38477 85158 -37895
rect 85207 -37935 85242 -37895
rect 85208 -38439 85242 -37935
rect 85306 -38432 85340 -37931
rect 85404 -37934 85439 -37895
rect 84938 -38517 85158 -38477
rect 85303 -38552 85341 -38432
rect 85404 -38439 85438 -37934
rect 85534 -38515 85568 -37931
rect 85860 -38445 85894 -37931
rect 86088 -38221 86122 -37931
rect 86087 -38314 86124 -38221
rect 86087 -38351 86224 -38314
rect 85860 -38479 86019 -38445
rect 85683 -38515 85821 -38504
rect 84939 -38590 85341 -38552
rect 85408 -38549 85821 -38515
rect 84702 -38601 84840 -38591
rect 84312 -38635 84840 -38601
rect 83791 -38808 83896 -38736
rect 84312 -38911 84355 -38635
rect 84702 -38645 84840 -38635
rect 84758 -38736 84896 -38727
rect 84548 -38770 84896 -38736
rect 84548 -38897 84620 -38770
rect 84758 -38781 84896 -38770
rect 84548 -38906 84632 -38897
rect 81824 -39059 82274 -39041
rect 81382 -39102 82274 -39059
rect 81382 -39120 81831 -39102
rect 82213 -39397 82274 -39102
rect 82947 -39279 82981 -38985
rect 83039 -39001 83084 -38931
rect 83431 -38951 84355 -38911
rect 83479 -38954 84355 -38951
rect 82940 -39397 82987 -39279
rect 83045 -39293 83079 -39001
rect 83143 -39278 83177 -38985
rect 83385 -39268 83419 -38985
rect 83479 -38994 83523 -38954
rect 84553 -38976 84632 -38906
rect 83136 -39397 83183 -39278
rect 83378 -39397 83425 -39268
rect 83483 -39293 83517 -38994
rect 84841 -39218 84875 -38927
rect 84839 -39329 84876 -39218
rect 84939 -39235 84973 -38590
rect 85168 -38660 85206 -38590
rect 85408 -38628 85442 -38549
rect 85683 -38558 85821 -38549
rect 85158 -38798 85212 -38660
rect 85311 -38662 85442 -38628
rect 85508 -38645 85646 -38591
rect 85893 -38660 85947 -38522
rect 85985 -38523 86019 -38479
rect 85985 -38577 86151 -38523
rect 85311 -39235 85345 -38662
rect 85985 -38692 86019 -38577
rect 86071 -38692 86125 -38675
rect 85409 -38731 85568 -38696
rect 85985 -38697 86125 -38692
rect 85957 -38726 86125 -38697
rect 85409 -39235 85443 -38731
rect 85534 -39235 85568 -38731
rect 85632 -39218 85666 -38727
rect 85762 -39217 85796 -38727
rect 84302 -39333 84913 -39329
rect 85631 -39333 85668 -39218
rect 85759 -39333 85796 -39217
rect 85860 -39235 85894 -38727
rect 85957 -38731 86019 -38726
rect 85958 -39235 85992 -38731
rect 86071 -38734 86125 -38726
rect 86186 -38844 86224 -38351
rect 86186 -38882 86478 -38844
rect 86088 -39216 86122 -38927
rect 86186 -38932 86224 -38882
rect 86086 -39333 86123 -39216
rect 86186 -39235 86220 -38932
rect 84302 -39397 86236 -39333
rect 82213 -39442 86236 -39397
rect 82213 -39510 84415 -39442
rect 84763 -39494 86236 -39442
rect 80392 -39783 81273 -39636
rect 86440 -39777 86478 -38882
rect 80392 -39859 84465 -39783
rect 80392 -39862 81273 -39859
rect 80392 -44464 80618 -39862
rect 81155 -40041 81231 -39862
rect 81155 -40117 81297 -40041
rect 81221 -40506 81297 -40117
rect 82230 -40083 82895 -40055
rect 82230 -40141 83265 -40083
rect 82230 -40222 82316 -40141
rect 82490 -40178 82525 -40141
rect 82815 -40144 83265 -40141
rect 81378 -40308 82316 -40222
rect 81221 -40598 81356 -40506
rect 81518 -40564 81552 -40308
rect 81616 -40564 81650 -40356
rect 81714 -40564 81748 -40308
rect 81812 -40530 81846 -40356
rect 82393 -40486 82427 -40178
rect 82491 -40486 82525 -40178
rect 82589 -40486 82623 -40178
rect 82687 -40486 82721 -40178
rect 82785 -40486 82819 -40178
rect 82361 -40529 82432 -40528
rect 82773 -40529 82847 -40523
rect 82361 -40530 82847 -40529
rect 81812 -40564 82847 -40530
rect 83204 -40551 83265 -40144
rect 81813 -40568 82847 -40564
rect 81813 -40570 82362 -40568
rect 81400 -40598 81473 -40592
rect 82773 -40594 82847 -40568
rect 81221 -40615 81473 -40598
rect 81226 -40639 81473 -40615
rect 82308 -40626 82443 -40618
rect 82288 -40628 82443 -40626
rect 81226 -40656 81356 -40639
rect 81400 -40652 81473 -40639
rect 82081 -40664 82443 -40628
rect 82960 -40637 83745 -40551
rect 82288 -40666 82443 -40664
rect 82308 -40672 82443 -40666
rect 82491 -40649 82910 -40641
rect 82491 -40679 82921 -40649
rect 81518 -40894 81552 -40686
rect 81714 -40894 81748 -40686
rect 81910 -40894 81944 -40686
rect 82491 -41023 82525 -40679
rect 82687 -41023 82721 -40679
rect 82860 -40828 82921 -40679
rect 83100 -40793 83134 -40637
rect 83198 -40793 83232 -40685
rect 83296 -40793 83330 -40637
rect 83394 -40793 83428 -40685
rect 82982 -40828 83055 -40822
rect 82860 -40841 83055 -40828
rect 82882 -40869 83055 -40841
rect 82982 -40882 83055 -40869
rect 83492 -40852 83864 -40782
rect 83100 -41024 83134 -40916
rect 83296 -41024 83330 -40916
rect 83492 -41024 83526 -40852
rect 81492 -41959 81526 -41615
rect 81688 -41959 81722 -41615
rect 82101 -41722 82135 -41614
rect 82297 -41722 82331 -41614
rect 81983 -41769 82056 -41756
rect 81883 -41797 82056 -41769
rect 81861 -41810 82056 -41797
rect 81861 -41959 81922 -41810
rect 81983 -41816 82056 -41810
rect 82493 -41786 82527 -41614
rect 81309 -41972 81444 -41966
rect 81289 -41974 81444 -41972
rect 80761 -42010 81444 -41974
rect 81492 -41989 81922 -41959
rect 81492 -41997 81911 -41989
rect 82101 -42001 82135 -41845
rect 82199 -41953 82233 -41845
rect 82297 -42001 82331 -41845
rect 82395 -41953 82429 -41845
rect 82493 -41856 82771 -41786
rect 80944 -43037 81080 -42010
rect 81289 -42012 81444 -42010
rect 81309 -42020 81444 -42012
rect 81136 -42070 81363 -42068
rect 81774 -42070 81848 -42044
rect 81136 -42108 81848 -42070
rect 81961 -42087 82576 -42001
rect 81362 -42109 81848 -42108
rect 81362 -42110 81433 -42109
rect 81774 -42115 81848 -42109
rect 81394 -42460 81428 -42152
rect 81492 -42460 81526 -42152
rect 81590 -42460 81624 -42152
rect 81688 -42460 81722 -42152
rect 81786 -42460 81820 -42152
rect 81491 -42512 81526 -42460
rect 82205 -42494 82266 -42087
rect 82695 -42251 82765 -41856
rect 82939 -42110 82973 -41526
rect 83146 -41492 83386 -41458
rect 83146 -41534 83188 -41492
rect 82935 -42169 82977 -42110
rect 83150 -42116 83184 -41534
rect 83248 -42114 83282 -41526
rect 83344 -41536 83386 -41492
rect 83147 -42169 83189 -42116
rect 82935 -42205 83189 -42169
rect 83244 -42168 83286 -42114
rect 83346 -42134 83380 -41536
rect 83558 -42120 83592 -41526
rect 83244 -42207 83385 -42168
rect 83342 -42219 83385 -42207
rect 83100 -42251 83255 -42241
rect 82695 -42287 83255 -42251
rect 82695 -42289 82765 -42287
rect 83100 -42296 83255 -42287
rect 83342 -42274 83523 -42219
rect 83342 -42344 83385 -42274
rect 82830 -42358 82985 -42349
rect 82793 -42392 82985 -42358
rect 82830 -42404 82985 -42392
rect 83031 -42384 83385 -42344
rect 83557 -42364 83600 -42120
rect 83794 -42189 83864 -40852
rect 84039 -40140 84131 -40055
rect 84062 -42115 84105 -40140
rect 84389 -40563 84465 -39859
rect 84691 -39815 86478 -39777
rect 84691 -40193 84729 -39815
rect 85898 -40114 86563 -40086
rect 85898 -40172 86933 -40114
rect 84668 -40247 84741 -40193
rect 85898 -40253 85984 -40172
rect 86158 -40209 86193 -40172
rect 86483 -40175 86933 -40172
rect 85046 -40339 85984 -40253
rect 84894 -40563 85024 -40537
rect 84389 -40629 85024 -40563
rect 85186 -40595 85220 -40339
rect 85284 -40595 85318 -40387
rect 85382 -40595 85416 -40339
rect 85480 -40561 85514 -40387
rect 86061 -40517 86095 -40209
rect 86159 -40517 86193 -40209
rect 86257 -40517 86291 -40209
rect 86355 -40517 86389 -40209
rect 86453 -40517 86487 -40209
rect 86029 -40560 86100 -40559
rect 86441 -40560 86515 -40554
rect 86029 -40561 86515 -40560
rect 85480 -40595 86515 -40561
rect 86872 -40582 86933 -40175
rect 85481 -40599 86515 -40595
rect 85481 -40601 86030 -40599
rect 85068 -40629 85141 -40623
rect 86441 -40625 86515 -40599
rect 84389 -40639 85141 -40629
rect 84894 -40670 85141 -40639
rect 85976 -40657 86111 -40649
rect 85956 -40659 86111 -40657
rect 84894 -40687 85024 -40670
rect 85068 -40683 85141 -40670
rect 84921 -40737 84997 -40687
rect 85749 -40695 86111 -40659
rect 86628 -40668 87413 -40582
rect 85956 -40697 86111 -40695
rect 85976 -40703 86111 -40697
rect 86159 -40680 86578 -40672
rect 86159 -40710 86589 -40680
rect 85186 -40925 85220 -40717
rect 85382 -40925 85416 -40717
rect 85578 -40925 85612 -40717
rect 86159 -41054 86193 -40710
rect 86355 -41054 86389 -40710
rect 86528 -40859 86589 -40710
rect 86768 -40824 86802 -40668
rect 86866 -40824 86900 -40716
rect 86964 -40824 86998 -40668
rect 87062 -40824 87096 -40716
rect 86650 -40859 86723 -40853
rect 86528 -40872 86723 -40859
rect 86550 -40900 86723 -40872
rect 86650 -40913 86723 -40900
rect 87160 -40883 87532 -40813
rect 86768 -41055 86802 -40947
rect 86964 -41055 86998 -40947
rect 87160 -41055 87194 -40883
rect 85160 -41990 85194 -41646
rect 85356 -41990 85390 -41646
rect 85769 -41753 85803 -41645
rect 85965 -41753 85999 -41645
rect 85651 -41800 85724 -41787
rect 85551 -41828 85724 -41800
rect 85529 -41841 85724 -41828
rect 85529 -41990 85590 -41841
rect 85651 -41847 85724 -41841
rect 86161 -41817 86195 -41645
rect 84977 -42003 85112 -41997
rect 84957 -42005 85112 -42003
rect 84543 -42041 85112 -42005
rect 85160 -42020 85590 -41990
rect 85160 -42028 85579 -42020
rect 85769 -42032 85803 -41876
rect 85867 -41984 85901 -41876
rect 85965 -42032 85999 -41876
rect 86063 -41984 86097 -41876
rect 86161 -41887 86439 -41817
rect 84062 -42158 84347 -42115
rect 83783 -42261 83888 -42189
rect 84304 -42364 84347 -42158
rect 81816 -42512 82266 -42494
rect 81374 -42555 82266 -42512
rect 81374 -42573 81823 -42555
rect 82205 -42850 82266 -42555
rect 82939 -42732 82973 -42438
rect 83031 -42454 83076 -42384
rect 83423 -42404 84347 -42364
rect 83471 -42407 84347 -42404
rect 82932 -42850 82979 -42732
rect 83037 -42746 83071 -42454
rect 83135 -42731 83169 -42438
rect 83377 -42721 83411 -42438
rect 83471 -42447 83515 -42407
rect 83128 -42850 83175 -42731
rect 83370 -42850 83417 -42721
rect 83475 -42746 83509 -42447
rect 82205 -42963 83682 -42850
rect 84543 -43037 84679 -42041
rect 84957 -42043 85112 -42041
rect 84977 -42051 85112 -42043
rect 84804 -42101 85031 -42099
rect 85442 -42101 85516 -42075
rect 84804 -42139 85516 -42101
rect 85629 -42118 86244 -42032
rect 85030 -42140 85516 -42139
rect 85030 -42141 85101 -42140
rect 85442 -42146 85516 -42140
rect 85062 -42491 85096 -42183
rect 85160 -42491 85194 -42183
rect 85258 -42491 85292 -42183
rect 85356 -42491 85390 -42183
rect 85454 -42491 85488 -42183
rect 85159 -42543 85194 -42491
rect 85873 -42525 85934 -42118
rect 86363 -42282 86433 -41887
rect 86607 -42141 86641 -41557
rect 86814 -41523 87054 -41489
rect 86814 -41565 86856 -41523
rect 86603 -42200 86645 -42141
rect 86818 -42147 86852 -41565
rect 86916 -42145 86950 -41557
rect 87012 -41567 87054 -41523
rect 86815 -42200 86857 -42147
rect 86603 -42236 86857 -42200
rect 86912 -42199 86954 -42145
rect 87014 -42165 87048 -41567
rect 87226 -42151 87260 -41557
rect 86912 -42238 87053 -42199
rect 87010 -42250 87053 -42238
rect 86768 -42282 86923 -42272
rect 86363 -42318 86923 -42282
rect 86363 -42320 86433 -42318
rect 86768 -42327 86923 -42318
rect 87010 -42305 87191 -42250
rect 87010 -42375 87053 -42305
rect 86498 -42389 86653 -42380
rect 86461 -42423 86653 -42389
rect 86498 -42435 86653 -42423
rect 86699 -42415 87053 -42375
rect 87225 -42395 87268 -42151
rect 87462 -42220 87532 -40883
rect 87451 -42292 87556 -42220
rect 88080 -42395 88439 -42245
rect 85484 -42543 85934 -42525
rect 85042 -42586 85934 -42543
rect 85042 -42604 85491 -42586
rect 85873 -42881 85934 -42586
rect 86607 -42763 86641 -42469
rect 86699 -42485 86744 -42415
rect 87091 -42435 88439 -42395
rect 87139 -42438 88439 -42435
rect 86600 -42881 86647 -42763
rect 86705 -42777 86739 -42485
rect 86803 -42762 86837 -42469
rect 87045 -42752 87079 -42469
rect 87139 -42478 87183 -42438
rect 86796 -42881 86843 -42762
rect 87038 -42881 87085 -42752
rect 87143 -42777 87177 -42478
rect 88080 -42588 88439 -42438
rect 85873 -42994 87350 -42881
rect 80944 -43173 84679 -43037
rect 80303 -44740 80690 -44464
rect -24214 -45912 71716 -45776
rect -24214 -46146 -24078 -45912
rect 80968 -46146 81104 -43173
rect -24214 -46282 81104 -46146
rect -7309 -46786 17635 -46650
rect -24059 -47023 11109 -46888
rect -29448 -54911 -29178 -54761
rect -28849 -54911 -28729 -52231
rect -28236 -52262 -28144 -52236
rect -28644 -52296 -28144 -52262
rect -28236 -52380 -28144 -52296
rect -28644 -52414 -28144 -52380
rect -28236 -52498 -28144 -52414
rect -28644 -52532 -28144 -52498
rect -28236 -52616 -28144 -52532
rect -28644 -52650 -28144 -52616
rect -28236 -52734 -28144 -52650
rect -28644 -52768 -28144 -52734
rect -28236 -52852 -28144 -52768
rect -28644 -52886 -28144 -52852
rect -28236 -52970 -28144 -52886
rect -28644 -53004 -28144 -52970
rect -28236 -53088 -28144 -53004
rect -28644 -53122 -28144 -53088
rect -28236 -53206 -28144 -53122
rect -28644 -53240 -28144 -53206
rect 8944 -52313 20212 -51980
rect -28236 -53324 -28144 -53240
rect -28644 -53358 -28144 -53324
rect -28236 -53442 -28144 -53358
rect -28644 -53476 -28144 -53442
rect -28236 -53560 -28144 -53476
rect -28644 -53594 -28144 -53560
rect -28236 -53678 -28144 -53594
rect -28644 -53712 -28144 -53678
rect -13640 -53099 -13606 -53095
rect -13646 -53352 -13600 -53099
rect -13444 -53287 -13410 -53095
rect -13450 -53352 -13404 -53287
rect -13248 -53287 -13214 -53095
rect -13024 -53181 -12967 -53117
rect -13167 -53230 -12967 -53181
rect -13254 -53352 -13208 -53287
rect -13646 -53360 -13208 -53352
rect -13167 -53360 -13121 -53230
rect -13024 -53281 -12967 -53230
rect -12803 -53099 -12769 -53095
rect -13850 -53397 -13682 -53367
rect -28236 -53796 -28144 -53712
rect -28644 -53830 -28144 -53796
rect -28236 -53914 -28144 -53830
rect -28644 -53948 -28144 -53914
rect -28236 -54032 -28144 -53948
rect -28644 -54066 -28144 -54032
rect -28236 -54150 -28144 -54066
rect -28644 -54184 -28144 -54150
rect -28236 -54268 -28144 -54184
rect -28644 -54302 -28144 -54268
rect -28236 -54386 -28144 -54302
rect -28644 -54420 -28144 -54386
rect -28236 -54504 -28144 -54420
rect -28644 -54538 -28144 -54504
rect -28236 -54622 -28144 -54538
rect -28644 -54656 -28144 -54622
rect -21239 -54126 -21205 -53882
rect -21043 -54126 -21009 -53882
rect -20847 -54126 -20813 -53882
rect -21239 -54163 -20684 -54126
rect -20721 -54301 -20684 -54163
rect -20279 -54301 -20144 -54291
rect -20721 -54338 -20144 -54301
rect -20721 -54392 -20684 -54338
rect -20279 -54345 -20144 -54338
rect -28236 -54740 -28144 -54656
rect -28644 -54774 -28144 -54740
rect -28236 -54858 -28144 -54774
rect -28644 -54892 -28144 -54858
rect -21337 -54426 -20894 -54392
rect -20721 -54426 -20488 -54392
rect -21337 -54797 -21303 -54426
rect -21141 -54427 -20894 -54426
rect -29448 -55189 -28729 -54911
rect -28236 -54976 -28144 -54892
rect -28644 -55010 -28144 -54976
rect -28236 -55094 -28144 -55010
rect -28644 -55128 -28144 -55094
rect -29448 -56093 -29178 -55189
rect -28849 -55802 -28729 -55189
rect -28236 -55212 -28144 -55128
rect -28644 -55246 -28144 -55212
rect -28236 -55330 -28144 -55246
rect -28644 -55364 -28144 -55330
rect -21239 -54986 -21205 -54489
rect -21141 -54797 -21107 -54427
rect -20929 -54490 -20894 -54427
rect -21027 -54789 -20993 -54490
rect -21027 -54893 -20992 -54789
rect -20929 -54798 -20895 -54490
rect -20831 -54787 -20797 -54490
rect -20831 -54893 -20796 -54787
rect -20718 -54798 -20684 -54426
rect -21027 -54896 -20796 -54893
rect -20620 -54896 -20586 -54490
rect -20522 -54798 -20488 -54426
rect -21027 -54930 -20586 -54896
rect -20207 -54897 -20173 -54590
rect -20109 -54798 -20075 -53882
rect -19653 -54363 -19516 -54346
rect -19240 -54348 -19206 -54004
rect -19044 -54348 -19010 -54004
rect -18631 -54111 -18597 -54003
rect -18435 -54111 -18401 -54003
rect -18749 -54158 -18676 -54145
rect -18849 -54186 -18676 -54158
rect -18871 -54199 -18676 -54186
rect -18871 -54348 -18810 -54199
rect -18749 -54205 -18676 -54199
rect -18239 -54175 -18205 -54003
rect -16891 -54039 -15414 -53926
rect -18239 -54176 -17835 -54175
rect -18239 -54234 -17771 -54176
rect -19423 -54361 -19288 -54355
rect -19443 -54363 -19288 -54361
rect -19653 -54399 -19288 -54363
rect -19240 -54378 -18810 -54348
rect -19240 -54386 -18821 -54378
rect -18631 -54390 -18597 -54234
rect -18533 -54342 -18499 -54234
rect -18435 -54390 -18401 -54234
rect -18337 -54342 -18303 -54234
rect -18239 -54245 -17835 -54234
rect -17722 -54334 -17273 -54316
rect -16891 -54334 -16830 -54039
rect -16164 -54157 -16117 -54039
rect -18198 -54390 -16830 -54334
rect -19653 -54404 -19516 -54399
rect -19443 -54401 -19288 -54399
rect -19423 -54409 -19288 -54401
rect -18771 -54395 -16830 -54390
rect -18771 -54476 -18137 -54395
rect -17605 -54429 -17570 -54395
rect -19338 -54849 -19304 -54541
rect -19240 -54849 -19206 -54541
rect -19142 -54849 -19108 -54541
rect -19044 -54849 -19010 -54541
rect -18946 -54849 -18912 -54541
rect -19241 -54897 -19206 -54849
rect -18527 -54883 -18466 -54476
rect -18198 -54478 -18137 -54476
rect -17702 -54737 -17668 -54429
rect -17604 -54737 -17570 -54429
rect -17506 -54737 -17472 -54429
rect -17408 -54737 -17374 -54429
rect -17310 -54737 -17276 -54429
rect -17734 -54780 -17663 -54779
rect -17322 -54780 -17248 -54774
rect -17734 -54781 -17248 -54780
rect -17960 -54819 -17248 -54781
rect -16891 -54802 -16830 -54395
rect -16157 -54451 -16123 -54157
rect -16059 -54435 -16025 -54143
rect -15968 -54158 -15921 -54039
rect -16266 -54497 -16111 -54485
rect -16303 -54531 -16111 -54497
rect -16266 -54540 -16111 -54531
rect -16065 -54505 -16020 -54435
rect -15961 -54451 -15927 -54158
rect -15726 -54168 -15679 -54039
rect -15719 -54451 -15685 -54168
rect -15621 -54442 -15587 -54143
rect -15625 -54482 -15581 -54442
rect -15625 -54485 -14485 -54482
rect -16065 -54545 -15711 -54505
rect -15673 -54525 -14485 -54485
rect -16401 -54602 -16331 -54600
rect -15996 -54602 -15841 -54593
rect -16401 -54638 -15841 -54602
rect -17960 -54821 -17733 -54819
rect -17322 -54845 -17248 -54819
rect -18916 -54897 -18466 -54883
rect -20392 -54986 -18436 -54897
rect -17135 -54888 -16520 -54802
rect -21971 -55210 -21910 -55032
rect -21337 -55049 -18436 -54986
rect -21337 -55051 -20063 -55049
rect -19683 -55210 -19630 -55114
rect -28236 -55448 -28144 -55364
rect -28644 -55482 -28144 -55448
rect -28236 -55566 -28144 -55482
rect -28644 -55600 -28144 -55566
rect -21971 -55246 -19630 -55210
rect -21971 -55248 -21910 -55246
rect -17604 -54900 -17185 -54892
rect -17604 -54930 -17174 -54900
rect -17604 -55274 -17570 -54930
rect -17408 -55274 -17374 -54930
rect -17235 -55079 -17174 -54930
rect -16995 -55044 -16961 -54888
rect -16897 -55044 -16863 -54936
rect -16799 -55044 -16765 -54888
rect -16701 -55044 -16667 -54936
rect -16401 -55033 -16331 -54638
rect -15996 -54648 -15841 -54638
rect -15754 -54615 -15711 -54545
rect -15754 -54670 -15573 -54615
rect -15754 -54682 -15711 -54670
rect -16161 -54720 -15907 -54684
rect -17113 -55079 -17040 -55073
rect -17235 -55092 -17040 -55079
rect -17213 -55120 -17040 -55092
rect -17113 -55133 -17040 -55120
rect -16603 -55103 -16325 -55033
rect -16995 -55275 -16961 -55167
rect -16799 -55275 -16765 -55167
rect -16603 -55275 -16569 -55103
rect -16161 -54779 -16119 -54720
rect -16157 -55363 -16123 -54779
rect -15949 -54773 -15907 -54720
rect -15852 -54721 -15711 -54682
rect -15946 -55355 -15912 -54773
rect -15852 -54775 -15810 -54721
rect -15950 -55397 -15908 -55355
rect -15848 -55363 -15814 -54775
rect -15750 -55353 -15716 -54755
rect -15539 -54769 -15496 -54525
rect -15313 -54700 -15208 -54628
rect -15752 -55397 -15710 -55353
rect -15950 -55431 -15710 -55397
rect -15538 -55363 -15504 -54769
rect -28236 -55684 -28144 -55600
rect -28644 -55718 -28144 -55684
rect -28236 -55802 -28172 -55718
rect -28849 -55836 -28172 -55802
rect -28849 -56038 -28729 -55836
rect -28236 -55866 -28172 -55836
rect -28138 -55914 -27982 -55842
rect -28849 -56072 -28236 -56038
rect -28849 -56093 -28729 -56072
rect -29448 -56274 -28729 -56093
rect -28070 -56188 -28036 -55914
rect -28070 -56222 -27428 -56188
rect -29448 -56308 -28236 -56274
rect -29448 -56371 -28729 -56308
rect -21712 -56272 -21652 -56073
rect -21182 -56257 -21148 -55913
rect -20986 -56257 -20952 -55913
rect -20573 -56020 -20539 -55912
rect -20377 -56020 -20343 -55912
rect -20691 -56067 -20618 -56054
rect -20791 -56095 -20618 -56067
rect -20813 -56108 -20618 -56095
rect -20813 -56257 -20752 -56108
rect -20691 -56114 -20618 -56108
rect -20181 -56084 -20147 -55912
rect -19409 -56062 -19375 -55818
rect -19213 -56062 -19179 -55818
rect -19017 -56062 -18983 -55818
rect -19584 -56073 -19449 -56065
rect -19944 -56084 -19449 -56073
rect -20181 -56108 -19449 -56084
rect -19409 -56099 -18854 -56062
rect -21365 -56270 -21230 -56264
rect -21385 -56272 -21230 -56270
rect -21712 -56308 -21230 -56272
rect -21182 -56287 -20752 -56257
rect -21182 -56295 -20763 -56287
rect -20573 -56299 -20539 -56143
rect -20475 -56251 -20441 -56143
rect -20377 -56299 -20343 -56143
rect -20279 -56251 -20245 -56143
rect -20181 -56154 -19903 -56108
rect -19603 -56110 -19449 -56108
rect -19584 -56119 -19449 -56110
rect -19699 -56156 -19641 -56148
rect -19248 -56156 -19113 -56147
rect -19725 -56194 -19113 -56156
rect -21712 -56310 -21652 -56308
rect -21385 -56310 -21230 -56308
rect -21365 -56318 -21230 -56310
rect -29448 -57168 -29178 -56371
rect -28849 -56510 -28729 -56371
rect -27836 -56458 -27428 -56424
rect -28849 -56544 -28236 -56510
rect -21838 -56368 -21311 -56366
rect -20900 -56368 -20826 -56342
rect -21838 -56406 -20826 -56368
rect -20713 -56385 -20098 -56299
rect -21838 -56511 -21798 -56406
rect -21312 -56407 -20826 -56406
rect -21312 -56408 -21241 -56407
rect -20900 -56413 -20826 -56407
rect -28849 -56746 -28729 -56544
rect -27836 -56694 -27428 -56660
rect -28849 -56780 -28236 -56746
rect -21855 -56748 -21795 -56511
rect -21280 -56758 -21246 -56450
rect -21182 -56758 -21148 -56450
rect -21084 -56758 -21050 -56450
rect -20986 -56758 -20952 -56450
rect -20888 -56758 -20854 -56450
rect -28849 -56982 -28729 -56780
rect -21183 -56810 -21148 -56758
rect -20469 -56792 -20408 -56385
rect -20010 -56513 -19952 -56376
rect -19796 -56379 -19738 -56279
rect -19699 -56285 -19641 -56194
rect -19248 -56201 -19113 -56194
rect -19060 -56238 -18925 -56225
rect -19601 -56272 -18925 -56238
rect -19601 -56379 -19567 -56272
rect -19060 -56279 -18925 -56272
rect -18891 -56237 -18854 -56099
rect -18449 -56237 -18314 -56227
rect -18891 -56274 -18314 -56237
rect -18891 -56328 -18854 -56274
rect -18449 -56281 -18314 -56274
rect -18279 -56299 -18245 -55818
rect -17578 -56203 -17544 -55995
rect -17382 -56203 -17348 -55995
rect -17186 -56203 -17152 -55995
rect -16605 -56210 -16571 -55866
rect -16409 -56210 -16375 -55866
rect -15996 -55973 -15962 -55865
rect -15800 -55973 -15766 -55865
rect -16114 -56020 -16041 -56007
rect -16214 -56048 -16041 -56020
rect -16236 -56061 -16041 -56048
rect -16236 -56210 -16175 -56061
rect -16114 -56067 -16041 -56061
rect -15604 -56037 -15570 -55865
rect -15302 -56037 -15232 -54700
rect -16788 -56223 -16653 -56217
rect -16808 -56225 -16653 -56223
rect -17870 -56250 -17740 -56233
rect -17696 -56250 -17623 -56237
rect -17870 -56291 -17623 -56250
rect -17015 -56261 -16653 -56225
rect -16605 -56240 -16175 -56210
rect -16605 -56248 -16186 -56240
rect -15996 -56252 -15962 -56096
rect -15898 -56204 -15864 -56096
rect -15800 -56252 -15766 -56096
rect -15702 -56204 -15668 -56096
rect -15604 -56107 -15232 -56037
rect -16808 -56263 -16653 -56261
rect -16788 -56271 -16653 -56263
rect -17870 -56299 -17740 -56291
rect -17696 -56297 -17623 -56291
rect -19796 -56413 -19567 -56379
rect -19507 -56362 -19064 -56328
rect -18891 -56362 -18658 -56328
rect -19796 -56416 -19738 -56413
rect -19507 -56733 -19473 -56362
rect -19311 -56363 -19064 -56362
rect -20858 -56810 -19689 -56792
rect -27836 -56930 -27428 -56896
rect -28849 -57016 -28236 -56982
rect -21300 -56871 -19689 -56810
rect -20859 -56907 -19689 -56871
rect -28849 -57168 -28729 -57016
rect -19804 -56925 -19689 -56907
rect -19409 -56922 -19375 -56425
rect -19311 -56733 -19277 -56363
rect -19099 -56426 -19064 -56363
rect -19197 -56725 -19163 -56426
rect -19197 -56829 -19162 -56725
rect -19099 -56734 -19065 -56426
rect -19001 -56723 -18967 -56426
rect -19001 -56829 -18966 -56723
rect -18888 -56734 -18854 -56362
rect -19197 -56832 -18966 -56829
rect -18790 -56832 -18756 -56426
rect -18692 -56734 -18658 -56362
rect -18279 -56333 -17740 -56299
rect -17283 -56321 -16734 -56319
rect -16323 -56321 -16249 -56295
rect -17283 -56325 -16249 -56321
rect -19197 -56866 -18756 -56832
rect -18377 -56895 -18343 -56526
rect -18279 -56734 -18245 -56333
rect -17870 -56383 -17740 -56333
rect -17578 -56581 -17544 -56325
rect -17480 -56533 -17446 -56325
rect -17382 -56581 -17348 -56325
rect -17284 -56359 -16249 -56325
rect -16136 -56338 -15351 -56252
rect -17284 -56533 -17250 -56359
rect -16735 -56360 -16249 -56359
rect -16735 -56361 -16664 -56360
rect -16323 -56366 -16249 -56360
rect -17718 -56667 -16780 -56581
rect -16866 -56748 -16780 -56667
rect -16703 -56711 -16669 -56403
rect -16605 -56711 -16571 -56403
rect -16507 -56711 -16473 -56403
rect -16409 -56711 -16375 -56403
rect -16311 -56711 -16277 -56403
rect -16606 -56748 -16571 -56711
rect -15892 -56745 -15831 -56338
rect -16281 -56748 -15831 -56745
rect -16866 -56806 -15831 -56748
rect -16866 -56834 -16201 -56806
rect -16830 -56895 -16620 -56834
rect -18578 -56922 -16620 -56895
rect -19507 -56925 -16620 -56922
rect -19804 -57050 -16620 -56925
rect -15698 -56884 -15430 -56834
rect -14668 -56884 -14485 -54525
rect -13857 -53441 -13682 -53397
rect -13646 -53398 -13121 -53360
rect -12809 -53352 -12763 -53099
rect -12607 -53287 -12573 -53095
rect -12613 -53352 -12567 -53287
rect -12193 -53076 -11565 -53042
rect -12411 -53287 -12377 -53095
rect -12193 -53121 -12157 -53076
rect -12417 -53352 -12371 -53287
rect -12809 -53360 -12371 -53352
rect -12316 -53336 -12242 -53168
rect -12192 -53195 -12158 -53121
rect -12316 -53360 -12243 -53336
rect -13013 -53378 -12845 -53367
rect -13048 -53379 -12845 -53378
rect -13857 -53813 -13809 -53441
rect -13738 -53634 -13704 -53475
rect -13646 -53491 -13600 -53398
rect -13640 -53583 -13606 -53491
rect -13542 -53634 -13508 -53475
rect -13450 -53491 -13404 -53398
rect -13254 -53430 -13121 -53398
rect -13444 -53583 -13410 -53491
rect -13346 -53634 -13312 -53475
rect -13254 -53491 -13208 -53430
rect -13085 -53441 -12845 -53379
rect -12809 -53398 -12243 -53360
rect -13248 -53583 -13214 -53491
rect -13085 -53585 -13025 -53441
rect -12901 -53634 -12867 -53475
rect -12809 -53491 -12763 -53398
rect -12803 -53583 -12769 -53491
rect -12705 -53634 -12671 -53475
rect -12613 -53491 -12567 -53398
rect -12417 -53430 -12243 -53398
rect -12198 -53342 -12151 -53195
rect -12094 -53202 -12060 -53110
rect -11997 -53131 -11955 -53076
rect -12095 -53254 -12059 -53202
rect -11996 -53218 -11962 -53131
rect -11898 -53200 -11864 -53110
rect -11803 -53132 -11761 -53076
rect -11898 -53218 -11861 -53200
rect -11800 -53218 -11766 -53132
rect -11702 -53200 -11668 -53110
rect -11607 -53127 -11565 -53076
rect -11897 -53254 -11861 -53218
rect -11703 -53254 -11667 -53200
rect -11604 -53218 -11570 -53127
rect -11506 -53210 -11472 -53110
rect -11509 -53254 -11467 -53210
rect -12095 -53288 -11467 -53254
rect -12198 -53416 -12026 -53342
rect -11642 -53395 -11467 -53288
rect -10940 -53099 -10906 -53095
rect -10946 -53352 -10900 -53099
rect -10744 -53287 -10710 -53095
rect -10750 -53352 -10704 -53287
rect -10548 -53287 -10514 -53095
rect -10324 -53169 -10267 -53117
rect -10472 -53231 -10267 -53169
rect -10554 -53352 -10508 -53287
rect -10946 -53360 -10508 -53352
rect -10472 -53360 -10410 -53231
rect -10324 -53281 -10267 -53231
rect -10103 -53099 -10069 -53095
rect -11150 -53374 -10982 -53367
rect -12607 -53583 -12573 -53491
rect -12509 -53634 -12475 -53475
rect -12417 -53491 -12371 -53430
rect -12411 -53583 -12377 -53491
rect -12198 -53551 -12151 -53416
rect -11642 -53455 -11376 -53395
rect -11172 -53434 -10982 -53374
rect -11150 -53441 -10982 -53434
rect -10946 -53398 -10410 -53360
rect -10109 -53352 -10063 -53099
rect -9907 -53287 -9873 -53095
rect -9913 -53352 -9867 -53287
rect -9493 -53076 -8865 -53042
rect -9711 -53287 -9677 -53095
rect -9493 -53121 -9457 -53076
rect -9717 -53352 -9671 -53287
rect -10109 -53360 -9671 -53352
rect -9616 -53336 -9542 -53168
rect -9492 -53195 -9458 -53121
rect -9616 -53360 -9543 -53336
rect -10313 -53378 -10145 -53367
rect -12098 -53489 -11467 -53455
rect -12098 -53530 -12057 -53489
rect -12192 -53621 -12158 -53551
rect -13747 -53702 -12376 -53634
rect -12197 -53679 -12153 -53621
rect -12094 -53633 -12060 -53530
rect -11996 -53610 -11962 -53525
rect -11900 -53538 -11859 -53489
rect -12001 -53679 -11957 -53610
rect -11898 -53633 -11864 -53538
rect -11800 -53610 -11766 -53525
rect -11706 -53538 -11665 -53489
rect -11509 -53496 -11467 -53489
rect -11805 -53679 -11761 -53610
rect -11702 -53633 -11668 -53538
rect -11604 -53621 -11570 -53525
rect -11509 -53539 -11468 -53496
rect -11608 -53679 -11564 -53621
rect -11506 -53633 -11472 -53539
rect -11038 -53634 -11004 -53475
rect -10946 -53491 -10900 -53398
rect -10940 -53583 -10906 -53491
rect -10842 -53634 -10808 -53475
rect -10750 -53491 -10704 -53398
rect -10554 -53430 -10410 -53398
rect -10744 -53583 -10710 -53491
rect -10646 -53634 -10612 -53475
rect -10554 -53491 -10508 -53430
rect -10373 -53441 -10145 -53378
rect -10109 -53398 -9543 -53360
rect -10548 -53583 -10514 -53491
rect -10373 -53600 -10313 -53441
rect -10201 -53634 -10167 -53475
rect -10109 -53491 -10063 -53398
rect -10103 -53583 -10069 -53491
rect -10005 -53634 -9971 -53475
rect -9913 -53491 -9867 -53398
rect -9717 -53430 -9543 -53398
rect -9498 -53342 -9451 -53195
rect -9394 -53202 -9360 -53110
rect -9297 -53131 -9255 -53076
rect -9395 -53254 -9359 -53202
rect -9296 -53218 -9262 -53131
rect -9198 -53200 -9164 -53110
rect -9103 -53132 -9061 -53076
rect -9198 -53218 -9161 -53200
rect -9100 -53218 -9066 -53132
rect -9002 -53200 -8968 -53110
rect -8907 -53127 -8865 -53076
rect -9197 -53254 -9161 -53218
rect -9003 -53254 -8967 -53200
rect -8904 -53218 -8870 -53127
rect -8806 -53210 -8772 -53110
rect -8809 -53254 -8767 -53210
rect -9395 -53288 -8767 -53254
rect -9498 -53416 -9326 -53342
rect -8942 -53397 -8767 -53288
rect -9907 -53583 -9873 -53491
rect -9809 -53634 -9775 -53475
rect -9717 -53491 -9671 -53430
rect -9711 -53583 -9677 -53491
rect -9498 -53551 -9451 -53416
rect -8942 -53455 -8692 -53397
rect -9398 -53457 -8692 -53455
rect -9398 -53489 -8767 -53457
rect -9398 -53530 -9357 -53489
rect -9492 -53621 -9458 -53551
rect -13499 -53742 -13388 -53702
rect -13510 -53750 -13373 -53742
rect -12688 -53750 -12577 -53702
rect -12197 -53713 -11564 -53679
rect -11047 -53636 -10513 -53634
rect -10210 -53636 -9676 -53634
rect -11047 -53702 -9676 -53636
rect -9497 -53679 -9453 -53621
rect -9394 -53633 -9360 -53530
rect -9296 -53610 -9262 -53525
rect -9200 -53538 -9159 -53489
rect -9301 -53679 -9257 -53610
rect -9198 -53633 -9164 -53538
rect -9100 -53610 -9066 -53525
rect -9006 -53538 -8965 -53489
rect -8809 -53496 -8767 -53489
rect -9105 -53679 -9061 -53610
rect -9002 -53633 -8968 -53538
rect -8904 -53621 -8870 -53525
rect -8809 -53539 -8768 -53496
rect -8908 -53679 -8864 -53621
rect -8806 -53633 -8772 -53539
rect -10890 -53748 -10779 -53702
rect -10707 -53704 -10187 -53702
rect -10913 -53750 -10776 -53748
rect -10012 -53750 -9901 -53702
rect -9497 -53713 -8864 -53679
rect -7474 -53699 -7440 -53105
rect -7268 -53071 -7028 -53037
rect -7268 -53115 -7226 -53071
rect -8275 -53750 -8143 -53748
rect -13527 -53789 -8142 -53750
rect -13510 -53802 -13373 -53789
rect -10913 -53808 -10776 -53789
rect -8275 -53808 -8143 -53789
rect -13858 -53950 -13798 -53813
rect -11348 -53842 -11211 -53831
rect -10402 -53842 -10270 -53832
rect -13527 -53881 -7797 -53842
rect -11348 -53891 -11211 -53881
rect -10402 -53892 -10270 -53881
rect -13121 -53928 -12989 -53920
rect -8598 -53928 -8466 -53918
rect -13857 -54308 -13809 -53950
rect -13527 -53967 -8466 -53928
rect -7836 -53943 -7797 -53881
rect -7482 -53943 -7439 -53699
rect -7262 -53713 -7228 -53115
rect -7164 -53693 -7130 -53105
rect -7070 -53113 -7028 -53071
rect -7168 -53747 -7126 -53693
rect -7066 -53695 -7032 -53113
rect -7267 -53786 -7126 -53747
rect -7071 -53748 -7029 -53695
rect -6855 -53689 -6821 -53105
rect -6859 -53748 -6817 -53689
rect -6044 -53197 -5316 -53163
rect -6044 -53509 -6010 -53197
rect -5946 -53545 -5912 -53301
rect -5848 -53509 -5814 -53197
rect -5728 -53266 -5386 -53232
rect -5728 -53509 -5694 -53266
rect -5630 -53545 -5596 -53301
rect -5532 -53509 -5498 -53266
rect -6155 -53579 -5481 -53545
rect -7071 -53784 -6817 -53748
rect -7267 -53798 -7224 -53786
rect -7405 -53853 -7224 -53798
rect -7267 -53923 -7224 -53853
rect -7137 -53830 -6982 -53820
rect -6597 -53830 -6465 -53759
rect -7137 -53866 -6465 -53830
rect -7137 -53875 -6982 -53866
rect -13121 -53980 -12989 -53967
rect -8598 -53978 -8466 -53967
rect -7840 -53983 -7305 -53943
rect -7267 -53963 -6913 -53923
rect -7840 -53986 -7353 -53983
rect -13739 -54082 -13205 -54014
rect -12808 -54037 -12175 -54003
rect -13738 -54225 -13704 -54133
rect -13744 -54286 -13698 -54225
rect -13640 -54241 -13606 -54082
rect -13542 -54225 -13508 -54133
rect -13774 -54308 -13698 -54286
rect -13857 -54318 -13698 -54308
rect -13548 -54318 -13502 -54225
rect -13444 -54241 -13410 -54082
rect -13346 -54225 -13312 -54133
rect -13352 -54318 -13306 -54225
rect -13248 -54241 -13214 -54082
rect -12900 -54177 -12866 -54083
rect -12808 -54095 -12764 -54037
rect -12904 -54220 -12863 -54177
rect -12802 -54191 -12768 -54095
rect -12704 -54178 -12670 -54083
rect -12611 -54106 -12567 -54037
rect -12905 -54227 -12863 -54220
rect -12707 -54227 -12666 -54178
rect -12606 -54191 -12572 -54106
rect -12508 -54178 -12474 -54083
rect -12415 -54106 -12371 -54037
rect -12513 -54227 -12472 -54178
rect -12410 -54191 -12376 -54106
rect -12312 -54186 -12278 -54083
rect -12219 -54095 -12175 -54037
rect -11996 -54082 -10505 -54014
rect -10108 -54037 -9475 -54003
rect -12214 -54165 -12180 -54095
rect -12315 -54227 -12274 -54186
rect -12905 -54261 -12274 -54227
rect -13857 -54345 -13306 -54318
rect -13856 -54347 -13306 -54345
rect -13774 -54356 -13306 -54347
rect -13270 -54290 -13102 -54275
rect -12905 -54290 -12730 -54261
rect -13270 -54343 -12730 -54290
rect -12221 -54300 -12174 -54165
rect -11995 -54225 -11961 -54133
rect -12001 -54286 -11955 -54225
rect -11897 -54241 -11863 -54082
rect -11799 -54225 -11765 -54133
rect -13270 -54349 -13102 -54343
rect -13744 -54364 -13306 -54356
rect -13744 -54429 -13698 -54364
rect -13738 -54621 -13704 -54429
rect -13548 -54429 -13502 -54364
rect -13542 -54621 -13508 -54429
rect -13352 -54617 -13306 -54364
rect -13346 -54621 -13312 -54617
rect -12905 -54428 -12730 -54343
rect -12346 -54374 -12174 -54300
rect -12905 -54462 -12277 -54428
rect -12905 -54506 -12863 -54462
rect -12900 -54606 -12866 -54506
rect -12802 -54589 -12768 -54498
rect -12705 -54516 -12669 -54462
rect -12511 -54498 -12475 -54462
rect -12807 -54640 -12765 -54589
rect -12704 -54606 -12670 -54516
rect -12606 -54584 -12572 -54498
rect -12511 -54516 -12474 -54498
rect -12611 -54640 -12569 -54584
rect -12508 -54606 -12474 -54516
rect -12410 -54585 -12376 -54498
rect -12313 -54514 -12277 -54462
rect -12417 -54640 -12375 -54585
rect -12312 -54606 -12278 -54514
rect -12221 -54521 -12174 -54374
rect -12129 -54318 -11955 -54286
rect -11805 -54318 -11759 -54225
rect -11701 -54241 -11667 -54082
rect -11603 -54225 -11569 -54133
rect -11609 -54318 -11563 -54225
rect -11505 -54241 -11471 -54082
rect -12129 -54356 -11563 -54318
rect -11527 -54280 -11359 -54275
rect -11299 -54280 -11239 -54207
rect -11527 -54338 -11239 -54280
rect -11184 -54297 -11124 -54182
rect -11038 -54225 -11004 -54133
rect -11044 -54286 -10998 -54225
rect -10940 -54241 -10906 -54082
rect -10842 -54225 -10808 -54133
rect -11074 -54297 -10998 -54286
rect -11527 -54349 -11359 -54338
rect -11299 -54339 -11239 -54338
rect -11189 -54318 -10998 -54297
rect -10848 -54318 -10802 -54225
rect -10744 -54241 -10710 -54082
rect -10646 -54225 -10612 -54133
rect -10652 -54318 -10606 -54225
rect -10548 -54241 -10514 -54082
rect -10203 -54177 -10157 -54055
rect -10108 -54095 -10064 -54037
rect -10204 -54187 -10157 -54177
rect -10204 -54220 -10163 -54187
rect -10102 -54191 -10068 -54095
rect -10004 -54178 -9970 -54083
rect -9911 -54106 -9867 -54037
rect -10205 -54227 -10163 -54220
rect -10007 -54227 -9966 -54178
rect -9906 -54191 -9872 -54106
rect -9808 -54178 -9774 -54083
rect -9715 -54106 -9671 -54037
rect -9813 -54227 -9772 -54178
rect -9710 -54191 -9676 -54106
rect -9612 -54186 -9578 -54083
rect -9519 -54095 -9475 -54037
rect -9296 -54082 -7880 -54014
rect -9514 -54165 -9480 -54095
rect -9615 -54227 -9574 -54186
rect -10205 -54261 -9574 -54227
rect -11189 -54342 -10606 -54318
rect -12129 -54380 -12056 -54356
rect -12214 -54595 -12180 -54521
rect -12130 -54548 -12056 -54380
rect -12001 -54364 -11563 -54356
rect -12001 -54429 -11955 -54364
rect -12215 -54640 -12179 -54595
rect -11995 -54621 -11961 -54429
rect -12807 -54674 -12179 -54640
rect -11805 -54429 -11759 -54364
rect -11799 -54621 -11765 -54429
rect -11609 -54617 -11563 -54364
rect -11603 -54621 -11569 -54617
rect -11405 -54476 -11348 -54435
rect -11189 -54476 -11144 -54342
rect -11074 -54356 -10606 -54342
rect -10570 -54283 -10402 -54275
rect -10205 -54283 -10030 -54261
rect -10570 -54340 -10030 -54283
rect -9521 -54300 -9474 -54165
rect -9295 -54225 -9261 -54133
rect -9301 -54286 -9255 -54225
rect -9197 -54241 -9163 -54082
rect -9099 -54225 -9065 -54133
rect -10570 -54349 -10402 -54340
rect -11044 -54364 -10606 -54356
rect -11044 -54429 -10998 -54364
rect -11405 -54521 -11144 -54476
rect -11405 -54599 -11348 -54521
rect -11038 -54621 -11004 -54429
rect -10848 -54429 -10802 -54364
rect -10842 -54621 -10808 -54429
rect -10652 -54617 -10606 -54364
rect -10646 -54621 -10612 -54617
rect -10205 -54428 -10030 -54340
rect -9646 -54374 -9474 -54300
rect -10205 -54462 -9577 -54428
rect -10205 -54506 -10163 -54462
rect -10200 -54606 -10166 -54506
rect -10102 -54589 -10068 -54498
rect -10005 -54516 -9969 -54462
rect -9811 -54498 -9775 -54462
rect -10107 -54640 -10065 -54589
rect -10004 -54606 -9970 -54516
rect -9906 -54584 -9872 -54498
rect -9811 -54516 -9774 -54498
rect -9911 -54640 -9869 -54584
rect -9808 -54606 -9774 -54516
rect -9710 -54585 -9676 -54498
rect -9613 -54514 -9577 -54462
rect -9717 -54640 -9675 -54585
rect -9612 -54606 -9578 -54514
rect -9521 -54521 -9474 -54374
rect -9429 -54318 -9255 -54286
rect -9105 -54318 -9059 -54225
rect -9001 -54241 -8967 -54082
rect -8903 -54225 -8869 -54133
rect -8909 -54318 -8863 -54225
rect -8805 -54241 -8771 -54082
rect -9429 -54356 -8863 -54318
rect -8827 -54280 -8659 -54275
rect -8827 -54292 -8624 -54280
rect -8567 -54292 -8507 -54206
rect -8413 -54225 -8379 -54133
rect -8419 -54286 -8373 -54225
rect -8315 -54241 -8281 -54082
rect -8217 -54225 -8183 -54133
rect -8449 -54292 -8373 -54286
rect -8827 -54318 -8373 -54292
rect -8223 -54318 -8177 -54225
rect -8119 -54241 -8085 -54082
rect -8021 -54225 -7987 -54133
rect -8027 -54318 -7981 -54225
rect -7923 -54241 -7889 -54082
rect -7836 -54275 -7797 -53986
rect -7397 -54026 -7353 -53986
rect -8827 -54334 -7981 -54318
rect -8827 -54338 -8624 -54334
rect -8567 -54338 -8507 -54334
rect -8827 -54349 -8659 -54338
rect -8449 -54356 -7981 -54334
rect -7945 -54349 -7777 -54275
rect -7391 -54325 -7357 -54026
rect -7293 -54300 -7259 -54017
rect -9429 -54380 -9356 -54356
rect -9514 -54595 -9480 -54521
rect -9430 -54548 -9356 -54380
rect -9301 -54364 -8863 -54356
rect -9301 -54429 -9255 -54364
rect -9515 -54640 -9479 -54595
rect -9295 -54621 -9261 -54429
rect -10107 -54674 -9479 -54640
rect -9105 -54429 -9059 -54364
rect -9099 -54621 -9065 -54429
rect -8909 -54617 -8863 -54364
rect -8419 -54364 -7981 -54356
rect -8903 -54621 -8869 -54617
rect -8419 -54429 -8373 -54364
rect -8705 -54599 -8648 -54435
rect -8413 -54621 -8379 -54429
rect -8223 -54429 -8177 -54364
rect -8217 -54621 -8183 -54429
rect -8027 -54617 -7981 -54364
rect -8021 -54621 -7987 -54617
rect -7723 -54430 -7445 -54429
rect -7299 -54430 -7252 -54300
rect -7051 -54310 -7017 -54017
rect -6958 -54033 -6913 -53963
rect -6867 -53937 -6712 -53928
rect -6867 -53971 -6305 -53937
rect -6867 -53983 -6712 -53971
rect -7057 -54430 -7010 -54310
rect -6953 -54325 -6919 -54033
rect -6855 -54311 -6821 -54017
rect -6861 -54430 -6814 -54311
rect -7723 -54512 -6732 -54430
rect -19804 -57056 -19689 -57050
rect -27836 -57166 -27428 -57132
rect -29448 -57218 -28729 -57168
rect -29448 -57252 -28236 -57218
rect -29448 -57446 -28729 -57252
rect -27836 -57402 -27428 -57368
rect -29448 -58329 -29178 -57446
rect -28849 -57454 -28729 -57446
rect -28849 -57488 -28236 -57454
rect -28849 -57690 -28729 -57488
rect -27836 -57638 -27428 -57604
rect -28849 -57724 -28236 -57690
rect -28849 -57926 -28729 -57724
rect -28104 -57802 -27948 -57730
rect -28644 -57842 -28236 -57808
rect -28849 -57960 -28236 -57926
rect -28849 -58162 -28729 -57960
rect -28644 -58078 -28236 -58044
rect -28849 -58196 -28236 -58162
rect -28849 -58329 -28729 -58196
rect -28056 -58206 -28022 -57802
rect -27836 -57874 -27428 -57840
rect -28056 -58240 -27428 -58206
rect -28644 -58314 -28236 -58280
rect -29448 -58398 -28729 -58329
rect -29448 -58432 -28236 -58398
rect -29448 -58607 -28729 -58432
rect -27836 -58476 -27428 -58442
rect -28644 -58550 -28236 -58516
rect -29448 -59163 -29178 -58607
rect -28849 -58634 -28729 -58607
rect -28849 -58668 -28236 -58634
rect -28849 -58870 -28729 -58668
rect -28644 -58786 -28236 -58752
rect -28117 -58763 -27977 -58661
rect -27836 -58712 -27428 -58678
rect -28849 -58904 -28236 -58870
rect -28849 -59106 -28729 -58904
rect -28644 -59022 -28236 -58988
rect -28059 -59106 -28025 -58763
rect -27836 -58948 -27428 -58914
rect -28849 -59140 -28236 -59106
rect -28059 -59140 -27902 -59106
rect -28849 -59342 -28729 -59140
rect -28644 -59258 -28236 -59224
rect -28172 -59339 -27995 -59263
rect -27936 -59280 -27902 -59140
rect -27936 -59314 -27428 -59280
rect -28849 -59376 -28236 -59342
rect -28849 -59418 -28729 -59376
rect -28116 -59815 -28055 -59339
rect -27836 -59550 -27428 -59516
rect -26527 -57171 -19689 -57056
rect -15698 -57067 -14485 -56884
rect -11902 -55015 -10425 -54902
rect -12733 -55310 -12284 -55292
rect -11902 -55310 -11841 -55015
rect -11175 -55133 -11128 -55015
rect -12733 -55353 -11841 -55310
rect -12616 -55405 -12581 -55353
rect -12291 -55371 -11841 -55353
rect -12713 -55713 -12679 -55405
rect -12615 -55713 -12581 -55405
rect -12517 -55713 -12483 -55405
rect -12419 -55713 -12385 -55405
rect -12321 -55713 -12287 -55405
rect -11902 -55778 -11841 -55371
rect -11168 -55427 -11134 -55133
rect -11070 -55411 -11036 -55119
rect -10979 -55134 -10932 -55015
rect -11277 -55473 -11122 -55461
rect -11314 -55507 -11122 -55473
rect -11277 -55516 -11122 -55507
rect -11076 -55481 -11031 -55411
rect -10972 -55427 -10938 -55134
rect -10737 -55144 -10690 -55015
rect -10730 -55427 -10696 -55144
rect -10632 -55418 -10598 -55119
rect -10636 -55458 -10592 -55418
rect -10636 -55461 -7556 -55458
rect -11076 -55521 -10722 -55481
rect -10684 -55501 -7556 -55461
rect -11412 -55578 -11342 -55576
rect -11007 -55578 -10852 -55569
rect -11412 -55614 -10852 -55578
rect -13258 -55855 -13072 -55798
rect -12798 -55853 -12663 -55845
rect -12818 -55855 -12663 -55853
rect -13258 -55891 -12663 -55855
rect -12146 -55864 -11531 -55778
rect -13258 -55952 -13072 -55891
rect -12818 -55893 -12663 -55891
rect -12798 -55899 -12663 -55893
rect -12615 -55876 -12196 -55868
rect -12615 -55906 -12185 -55876
rect -12615 -56250 -12581 -55906
rect -12419 -56250 -12385 -55906
rect -12246 -56055 -12185 -55906
rect -12006 -56020 -11972 -55864
rect -11908 -56020 -11874 -55912
rect -11810 -56020 -11776 -55864
rect -11712 -56020 -11678 -55912
rect -11412 -56009 -11342 -55614
rect -11007 -55624 -10852 -55614
rect -10765 -55591 -10722 -55521
rect -10765 -55646 -10584 -55591
rect -10765 -55658 -10722 -55646
rect -11172 -55696 -10918 -55660
rect -12124 -56055 -12051 -56049
rect -12246 -56068 -12051 -56055
rect -12224 -56096 -12051 -56068
rect -12124 -56109 -12051 -56096
rect -11614 -56079 -11336 -56009
rect -12006 -56251 -11972 -56143
rect -11810 -56251 -11776 -56143
rect -11614 -56251 -11580 -56079
rect -11172 -55755 -11130 -55696
rect -11168 -56339 -11134 -55755
rect -10960 -55749 -10918 -55696
rect -10863 -55697 -10722 -55658
rect -10957 -56331 -10923 -55749
rect -10863 -55751 -10821 -55697
rect -10961 -56373 -10919 -56331
rect -10859 -56339 -10825 -55751
rect -10761 -56329 -10727 -55731
rect -10550 -55745 -10507 -55501
rect -7732 -55580 -7556 -55501
rect -10324 -55676 -10219 -55604
rect -10763 -56373 -10721 -56329
rect -10961 -56407 -10721 -56373
rect -10549 -56339 -10515 -55745
rect -15698 -57099 -15430 -57067
rect -28147 -62311 -28010 -59815
rect -27236 -60736 -26896 -60567
rect -26527 -60736 -26412 -57171
rect -18084 -57441 -14546 -57235
rect -14754 -57443 -14546 -57441
rect -15693 -57701 -15425 -57654
rect -27236 -60851 -26412 -60736
rect -23096 -57887 -15425 -57701
rect -12589 -57179 -12555 -56971
rect -12393 -57179 -12359 -56971
rect -12197 -57179 -12163 -56971
rect -11616 -57186 -11582 -56842
rect -11420 -57186 -11386 -56842
rect -11007 -56949 -10973 -56841
rect -10811 -56949 -10777 -56841
rect -11125 -56996 -11052 -56983
rect -11225 -57024 -11052 -56996
rect -11247 -57037 -11052 -57024
rect -11247 -57186 -11186 -57037
rect -11125 -57043 -11052 -57037
rect -10615 -57013 -10581 -56841
rect -10313 -57013 -10243 -55676
rect -6339 -56230 -6305 -53971
rect -6155 -55119 -6121 -53579
rect -6045 -53713 -5906 -53659
rect -5515 -53694 -5481 -53579
rect -5420 -53618 -5386 -53266
rect -5350 -53544 -5316 -53197
rect -5170 -53544 -5136 -53301
rect -5350 -53578 -5136 -53544
rect -4974 -53618 -4940 -53301
rect -4664 -53494 -4630 -53301
rect -5420 -53652 -4940 -53618
rect -4887 -53669 -4748 -53615
rect -5515 -53728 -5369 -53694
rect -6046 -53831 -5715 -53794
rect -5663 -53817 -5524 -53763
rect -5403 -53790 -5369 -53728
rect -5296 -53743 -5157 -53689
rect -5403 -53824 -4842 -53790
rect -6046 -53914 -6009 -53831
rect -5752 -53855 -5715 -53831
rect -5752 -53892 -5596 -53855
rect -6044 -54103 -6010 -53914
rect -6048 -54226 -6009 -54103
rect -5946 -54152 -5912 -53907
rect -5633 -53913 -5596 -53892
rect -5630 -54115 -5596 -53913
rect -5534 -53916 -5234 -53877
rect -5532 -54115 -5498 -53916
rect -5268 -54115 -5234 -53916
rect -5170 -54115 -5136 -53824
rect -4974 -54098 -4940 -53907
rect -4974 -54152 -4938 -54098
rect -4876 -54115 -4842 -53824
rect -4669 -53833 -4626 -53494
rect -4355 -53492 -4321 -53301
rect -4359 -53689 -4316 -53492
rect -4272 -53675 -4133 -53621
rect -4459 -53735 -4316 -53689
rect -4585 -53823 -4446 -53769
rect -4765 -53879 -4626 -53833
rect -4669 -53924 -4626 -53879
rect -4664 -54115 -4630 -53924
rect -4566 -54108 -4532 -53907
rect -4359 -53926 -4316 -53735
rect -5946 -54188 -4938 -54152
rect -4571 -54192 -4528 -54108
rect -4355 -54115 -4321 -53926
rect -4257 -54106 -4223 -53907
rect -3544 -53197 -2816 -53163
rect -3544 -53509 -3510 -53197
rect -3446 -53545 -3412 -53301
rect -3348 -53509 -3314 -53197
rect -3228 -53266 -2886 -53232
rect -3228 -53509 -3194 -53266
rect -3130 -53545 -3096 -53301
rect -3032 -53509 -2998 -53266
rect -3712 -53579 -2981 -53545
rect -3712 -53942 -3678 -53579
rect -3545 -53713 -3406 -53659
rect -3015 -53694 -2981 -53579
rect -2920 -53618 -2886 -53266
rect -2850 -53544 -2816 -53197
rect -2670 -53544 -2636 -53301
rect -2850 -53578 -2636 -53544
rect -2474 -53618 -2440 -53301
rect -2164 -53494 -2130 -53301
rect -2920 -53652 -2440 -53618
rect -2387 -53669 -2248 -53615
rect -3015 -53728 -2869 -53694
rect -3546 -53831 -3215 -53794
rect -3163 -53817 -3024 -53763
rect -2903 -53790 -2869 -53728
rect -2796 -53743 -2657 -53689
rect -2903 -53824 -2342 -53790
rect -3546 -53914 -3509 -53831
rect -3252 -53855 -3215 -53831
rect -3252 -53892 -3096 -53855
rect -3718 -54078 -3672 -53942
rect -3544 -54103 -3510 -53914
rect -4262 -54191 -4219 -54106
rect -3548 -54191 -3509 -54103
rect -3446 -54152 -3412 -53907
rect -3133 -53913 -3096 -53892
rect -3130 -54115 -3096 -53913
rect -3034 -53916 -2734 -53877
rect -3032 -54115 -2998 -53916
rect -2768 -54115 -2734 -53916
rect -2670 -54115 -2636 -53824
rect -2474 -54098 -2440 -53907
rect -2474 -54152 -2438 -54098
rect -2376 -54115 -2342 -53824
rect -2169 -53833 -2126 -53494
rect -1855 -53492 -1821 -53301
rect -1859 -53689 -1816 -53492
rect -1772 -53675 -1633 -53621
rect -1959 -53735 -1816 -53689
rect -2085 -53823 -1946 -53769
rect -2265 -53879 -2126 -53833
rect -2169 -53924 -2126 -53879
rect -2164 -54115 -2130 -53924
rect -2066 -54108 -2032 -53907
rect -1859 -53926 -1816 -53735
rect -3446 -54188 -2438 -54152
rect -4336 -54192 -3509 -54191
rect -2071 -54192 -2028 -54108
rect -1855 -54115 -1821 -53926
rect -1757 -54106 -1723 -53907
rect -1044 -53197 -316 -53163
rect -1044 -53509 -1010 -53197
rect -946 -53545 -912 -53301
rect -848 -53509 -814 -53197
rect -728 -53266 -386 -53232
rect -728 -53509 -694 -53266
rect -630 -53545 -596 -53301
rect -532 -53509 -498 -53266
rect -1164 -53579 -481 -53545
rect -1164 -53946 -1130 -53579
rect -1045 -53713 -906 -53659
rect -515 -53694 -481 -53579
rect -420 -53618 -386 -53266
rect -350 -53544 -316 -53197
rect -170 -53544 -136 -53301
rect -350 -53578 -136 -53544
rect 26 -53618 60 -53301
rect 336 -53494 370 -53301
rect -420 -53652 60 -53618
rect 113 -53669 252 -53615
rect -515 -53728 -369 -53694
rect -1046 -53831 -715 -53794
rect -663 -53817 -524 -53763
rect -403 -53790 -369 -53728
rect -296 -53743 -157 -53689
rect -403 -53824 158 -53790
rect -1046 -53914 -1009 -53831
rect -752 -53855 -715 -53831
rect -752 -53892 -596 -53855
rect -1170 -54082 -1124 -53946
rect -1044 -54103 -1010 -53914
rect -1762 -54192 -1719 -54106
rect -4847 -54226 -3509 -54192
rect -2347 -54226 -1715 -54192
rect -1048 -54226 -1009 -54103
rect -946 -54152 -912 -53907
rect -633 -53913 -596 -53892
rect -630 -54115 -596 -53913
rect -534 -53916 -234 -53877
rect -532 -54115 -498 -53916
rect -268 -54115 -234 -53916
rect -170 -54115 -136 -53824
rect 26 -54098 60 -53907
rect 26 -54152 62 -54098
rect 124 -54115 158 -53824
rect 331 -53833 374 -53494
rect 645 -53492 679 -53301
rect 641 -53689 684 -53492
rect 728 -53675 867 -53621
rect 541 -53735 684 -53689
rect 415 -53823 554 -53769
rect 235 -53879 374 -53833
rect 331 -53924 374 -53879
rect 336 -54115 370 -53924
rect 434 -54108 468 -53907
rect 641 -53926 684 -53735
rect -946 -54188 62 -54152
rect 429 -54192 472 -54108
rect 645 -54115 679 -53926
rect 743 -54106 777 -53907
rect 1456 -53197 2184 -53163
rect 1456 -53509 1490 -53197
rect 1316 -53545 1350 -53544
rect 1554 -53545 1588 -53301
rect 1652 -53509 1686 -53197
rect 1772 -53266 2114 -53232
rect 1772 -53509 1806 -53266
rect 1870 -53545 1904 -53301
rect 1968 -53509 2002 -53266
rect 1316 -53579 2019 -53545
rect 1316 -53946 1350 -53579
rect 1455 -53713 1594 -53659
rect 1985 -53694 2019 -53579
rect 2080 -53618 2114 -53266
rect 2150 -53544 2184 -53197
rect 2330 -53544 2364 -53301
rect 2150 -53578 2364 -53544
rect 2526 -53618 2560 -53301
rect 2836 -53494 2870 -53301
rect 2080 -53652 2560 -53618
rect 2613 -53669 2752 -53615
rect 1985 -53728 2131 -53694
rect 1454 -53831 1785 -53794
rect 1837 -53817 1976 -53763
rect 2097 -53790 2131 -53728
rect 2204 -53743 2343 -53689
rect 2097 -53824 2658 -53790
rect 1454 -53914 1491 -53831
rect 1748 -53855 1785 -53831
rect 1748 -53892 1904 -53855
rect 1310 -54082 1356 -53946
rect 1456 -54103 1490 -53914
rect 738 -54192 781 -54106
rect 153 -54226 785 -54192
rect 1452 -54226 1491 -54103
rect 1554 -54152 1588 -53907
rect 1867 -53913 1904 -53892
rect 1870 -54115 1904 -53913
rect 1966 -53916 2266 -53877
rect 1968 -54115 2002 -53916
rect 2232 -54115 2266 -53916
rect 2330 -54115 2364 -53824
rect 2526 -54098 2560 -53907
rect 2526 -54152 2562 -54098
rect 2624 -54115 2658 -53824
rect 2831 -53833 2874 -53494
rect 3145 -53492 3179 -53301
rect 3956 -53197 4684 -53163
rect 3141 -53689 3184 -53492
rect 3956 -53509 3990 -53197
rect 4054 -53545 4088 -53301
rect 4152 -53509 4186 -53197
rect 4272 -53266 4614 -53232
rect 4272 -53509 4306 -53266
rect 4370 -53545 4404 -53301
rect 4468 -53509 4502 -53266
rect 3732 -53579 4519 -53545
rect 3228 -53675 3367 -53621
rect 3041 -53735 3184 -53689
rect 2915 -53823 3054 -53769
rect 2735 -53879 2874 -53833
rect 2831 -53924 2874 -53879
rect 2836 -54115 2870 -53924
rect 2934 -54108 2968 -53907
rect 3141 -53926 3184 -53735
rect 1554 -54188 2562 -54152
rect 2929 -54192 2972 -54108
rect 3145 -54115 3179 -53926
rect 3243 -54106 3277 -53907
rect 3732 -53945 3766 -53579
rect 3955 -53713 4094 -53659
rect 4485 -53694 4519 -53579
rect 4580 -53618 4614 -53266
rect 4650 -53544 4684 -53197
rect 4830 -53544 4864 -53301
rect 4650 -53578 4864 -53544
rect 5026 -53618 5060 -53301
rect 5336 -53494 5370 -53301
rect 4580 -53652 5060 -53618
rect 5113 -53669 5252 -53615
rect 4485 -53728 4631 -53694
rect 3954 -53831 4285 -53794
rect 4597 -53790 4631 -53728
rect 4704 -53743 4843 -53689
rect 4597 -53824 5158 -53790
rect 3954 -53914 3991 -53831
rect 4248 -53855 4285 -53831
rect 4248 -53892 4404 -53855
rect 3732 -53946 3767 -53945
rect 3727 -54082 3773 -53946
rect 3956 -54103 3990 -53914
rect 3238 -54192 3281 -54106
rect 2653 -54226 3285 -54192
rect 3952 -54226 3991 -54103
rect 4054 -54152 4088 -53907
rect 4367 -53913 4404 -53892
rect 4370 -54115 4404 -53913
rect 4466 -53916 4766 -53877
rect 4468 -54115 4502 -53916
rect 4732 -54115 4766 -53916
rect 4830 -54115 4864 -53824
rect 5026 -54098 5060 -53907
rect 5026 -54152 5062 -54098
rect 5124 -54115 5158 -53824
rect 5331 -53833 5374 -53494
rect 5645 -53492 5679 -53301
rect 6956 -53197 7684 -53163
rect 5641 -53689 5684 -53492
rect 6956 -53509 6990 -53197
rect 7054 -53545 7088 -53301
rect 7152 -53509 7186 -53197
rect 7272 -53266 7614 -53232
rect 7272 -53509 7306 -53266
rect 7370 -53545 7404 -53301
rect 7468 -53509 7502 -53266
rect 6638 -53579 7519 -53545
rect 5728 -53675 5867 -53621
rect 5541 -53735 5684 -53689
rect 5235 -53879 5374 -53833
rect 5331 -53924 5374 -53879
rect 5336 -54115 5370 -53924
rect 5434 -54108 5468 -53907
rect 5641 -53926 5684 -53735
rect 4054 -54188 5062 -54152
rect 5429 -54192 5472 -54108
rect 5645 -54115 5679 -53926
rect 5743 -54106 5777 -53907
rect 6638 -53946 6672 -53579
rect 6955 -53713 7094 -53659
rect 7485 -53694 7519 -53579
rect 7580 -53618 7614 -53266
rect 7650 -53544 7684 -53197
rect 7830 -53544 7864 -53301
rect 7650 -53578 7864 -53544
rect 8026 -53618 8060 -53301
rect 8336 -53494 8370 -53301
rect 7580 -53652 8060 -53618
rect 8113 -53669 8252 -53615
rect 7485 -53728 7631 -53694
rect 6954 -53831 7285 -53794
rect 7597 -53790 7631 -53728
rect 7704 -53743 7843 -53689
rect 7597 -53824 8158 -53790
rect 6954 -53914 6991 -53831
rect 7248 -53855 7285 -53831
rect 7248 -53892 7404 -53855
rect 6632 -54082 6678 -53946
rect 6956 -54103 6990 -53914
rect 5738 -54192 5781 -54106
rect 5153 -54226 5785 -54192
rect 6952 -54226 6991 -54103
rect 7054 -54152 7088 -53907
rect 7367 -53913 7404 -53892
rect 7370 -54115 7404 -53913
rect 7466 -53916 7766 -53877
rect 7468 -54115 7502 -53916
rect 7732 -54115 7766 -53916
rect 7830 -54115 7864 -53824
rect 8026 -54098 8060 -53907
rect 8026 -54152 8062 -54098
rect 8124 -54115 8158 -53824
rect 8331 -53833 8374 -53494
rect 8645 -53492 8679 -53301
rect 8641 -53689 8684 -53492
rect 8728 -53675 8867 -53621
rect 8541 -53735 8684 -53689
rect 8235 -53879 8374 -53833
rect 8331 -53924 8374 -53879
rect 8336 -54115 8370 -53924
rect 8434 -54108 8468 -53907
rect 8641 -53926 8684 -53735
rect 7054 -54188 8062 -54152
rect 8429 -54174 8472 -54108
rect 8645 -54115 8679 -53926
rect 8743 -54106 8777 -53907
rect 8738 -54174 8781 -54106
rect 8944 -54174 9205 -52313
rect 17559 -52637 17756 -52456
rect 17215 -53112 17496 -52903
rect 9429 -53315 9629 -53281
rect 16855 -53315 17217 -53269
rect 9429 -53487 17217 -53315
rect 9429 -53652 9629 -53487
rect 16855 -53540 17217 -53487
rect 8137 -54226 9205 -54174
rect 16615 -54213 16907 -54212
rect -6048 -54278 9205 -54226
rect -6048 -54279 -4215 -54278
rect -3548 -54279 9205 -54278
rect -5616 -54299 -5082 -54279
rect -4847 -54288 -4215 -54279
rect -2347 -54288 -1715 -54279
rect 153 -54288 785 -54279
rect 2653 -54288 3285 -54279
rect 5153 -54288 5785 -54279
rect -5607 -54458 -5573 -54299
rect -5509 -54442 -5475 -54350
rect -5515 -54535 -5469 -54442
rect -5411 -54458 -5377 -54299
rect -5313 -54442 -5279 -54350
rect -5319 -54535 -5273 -54442
rect -5215 -54458 -5181 -54299
rect 8137 -54301 9205 -54279
rect -5117 -54442 -5083 -54350
rect -1005 -54364 -869 -54318
rect 1492 -54334 1628 -54331
rect -918 -54412 -869 -54364
rect 1459 -54368 3630 -54334
rect 1492 -54377 1628 -54368
rect -5123 -54503 -5077 -54442
rect -4100 -54503 -4054 -54437
rect -918 -54448 3534 -54412
rect -5123 -54535 -4054 -54503
rect -5515 -54573 -4054 -54535
rect -5515 -54581 -5077 -54573
rect -5515 -54834 -5469 -54581
rect -5509 -54838 -5475 -54834
rect -5319 -54646 -5273 -54581
rect -5313 -54838 -5279 -54646
rect -5123 -54646 -5077 -54581
rect -5117 -54838 -5083 -54646
rect -3718 -54784 -3672 -54648
rect 3498 -54560 3534 -54448
rect 3596 -54492 3630 -54368
rect 6580 -54384 6716 -54378
rect 3675 -54403 3811 -54394
rect 3675 -54437 6476 -54403
rect 6580 -54418 6852 -54384
rect 6580 -54424 6716 -54418
rect 3675 -54440 3811 -54437
rect 6442 -54476 6476 -54437
rect 3596 -54526 5098 -54492
rect 6442 -54510 6782 -54476
rect -6195 -55165 -6059 -55119
rect -3715 -55037 -3675 -54784
rect -3715 -55083 -3579 -55037
rect -6339 -56293 -6155 -56230
rect -6318 -56294 -6155 -56293
rect -11799 -57199 -11664 -57193
rect -11819 -57201 -11664 -57199
rect -12026 -57237 -11664 -57201
rect -11616 -57216 -11186 -57186
rect -11616 -57224 -11197 -57216
rect -11007 -57228 -10973 -57072
rect -10909 -57180 -10875 -57072
rect -10811 -57228 -10777 -57072
rect -10713 -57180 -10679 -57072
rect -10615 -57083 -10243 -57013
rect -5864 -55725 -5830 -55533
rect -5870 -55790 -5824 -55725
rect -5668 -55725 -5634 -55533
rect -5674 -55790 -5628 -55725
rect -5472 -55537 -5438 -55533
rect -5478 -55790 -5432 -55537
rect -4933 -55514 -4305 -55480
rect -5026 -55648 -4992 -55548
rect -4933 -55565 -4891 -55514
rect -5031 -55692 -4989 -55648
rect -4928 -55656 -4894 -55565
rect -4830 -55638 -4796 -55548
rect -4737 -55570 -4695 -55514
rect -4831 -55692 -4795 -55638
rect -4732 -55656 -4698 -55570
rect -4634 -55638 -4600 -55548
rect -4543 -55569 -4501 -55514
rect -4637 -55656 -4600 -55638
rect -4536 -55656 -4502 -55569
rect -4438 -55640 -4404 -55548
rect -4341 -55559 -4305 -55514
rect -4340 -55633 -4306 -55559
rect -4637 -55692 -4601 -55656
rect -4439 -55692 -4403 -55640
rect -5031 -55726 -4403 -55692
rect -5870 -55798 -5432 -55790
rect -5900 -55807 -5432 -55798
rect -5982 -55809 -5432 -55807
rect -5983 -55836 -5432 -55809
rect -5983 -55846 -5824 -55836
rect -5983 -56204 -5935 -55846
rect -5900 -55868 -5824 -55846
rect -5870 -55929 -5824 -55868
rect -5864 -56021 -5830 -55929
rect -5766 -56072 -5732 -55913
rect -5674 -55929 -5628 -55836
rect -5668 -56021 -5634 -55929
rect -5570 -56072 -5536 -55913
rect -5478 -55929 -5432 -55836
rect -5396 -55811 -5228 -55805
rect -5031 -55811 -4856 -55726
rect -4347 -55780 -4300 -55633
rect -4256 -55774 -4182 -55606
rect -4121 -55725 -4087 -55533
rect -5396 -55864 -4856 -55811
rect -4472 -55854 -4300 -55780
rect -5396 -55879 -5228 -55864
rect -5031 -55893 -4856 -55864
rect -5472 -56021 -5438 -55929
rect -5374 -56072 -5340 -55913
rect -5031 -55927 -4400 -55893
rect -5031 -55934 -4989 -55927
rect -5030 -55977 -4989 -55934
rect -5026 -56071 -4992 -55977
rect -4928 -56059 -4894 -55963
rect -4833 -55976 -4792 -55927
rect -5865 -56140 -5331 -56072
rect -4934 -56117 -4890 -56059
rect -4830 -56071 -4796 -55976
rect -4732 -56048 -4698 -55963
rect -4639 -55976 -4598 -55927
rect -4737 -56117 -4693 -56048
rect -4634 -56071 -4600 -55976
rect -4536 -56048 -4502 -55963
rect -4441 -55968 -4400 -55927
rect -4541 -56117 -4497 -56048
rect -4438 -56071 -4404 -55968
rect -4347 -55989 -4300 -55854
rect -4255 -55798 -4182 -55774
rect -4127 -55790 -4081 -55725
rect -3925 -55725 -3891 -55533
rect -3931 -55790 -3885 -55725
rect -3729 -55537 -3695 -55533
rect -3735 -55790 -3689 -55537
rect -3531 -55633 -3474 -55555
rect -3531 -55678 -3270 -55633
rect -3531 -55719 -3474 -55678
rect -4127 -55798 -3689 -55790
rect -4255 -55836 -3689 -55798
rect -4255 -55868 -4081 -55836
rect -4127 -55929 -4081 -55868
rect -4340 -56059 -4306 -55989
rect -4121 -56021 -4087 -55929
rect -4345 -56117 -4301 -56059
rect -4023 -56072 -3989 -55913
rect -3931 -55929 -3885 -55836
rect -3925 -56021 -3891 -55929
rect -3827 -56072 -3793 -55913
rect -3735 -55929 -3689 -55836
rect -3653 -55816 -3485 -55805
rect -3315 -55812 -3270 -55678
rect -3164 -55725 -3130 -55533
rect -3170 -55790 -3124 -55725
rect -2968 -55725 -2934 -55533
rect -2974 -55790 -2928 -55725
rect -2772 -55537 -2738 -55533
rect -2778 -55790 -2732 -55537
rect -2233 -55514 -1605 -55480
rect -2326 -55648 -2292 -55548
rect -2233 -55565 -2191 -55514
rect -2331 -55692 -2289 -55648
rect -2228 -55656 -2194 -55565
rect -2130 -55638 -2096 -55548
rect -2037 -55570 -1995 -55514
rect -2131 -55692 -2095 -55638
rect -2032 -55656 -1998 -55570
rect -1934 -55638 -1900 -55548
rect -1843 -55569 -1801 -55514
rect -1937 -55656 -1900 -55638
rect -1836 -55656 -1802 -55569
rect -1738 -55640 -1704 -55548
rect -1641 -55559 -1605 -55514
rect -1640 -55633 -1606 -55559
rect -1937 -55692 -1901 -55656
rect -1739 -55692 -1703 -55640
rect -2331 -55726 -1703 -55692
rect -3170 -55798 -2732 -55790
rect -3200 -55812 -2732 -55798
rect -3425 -55816 -3365 -55815
rect -3653 -55874 -3365 -55816
rect -3315 -55836 -2732 -55812
rect -3315 -55857 -3124 -55836
rect -3653 -55879 -3485 -55874
rect -3729 -56021 -3695 -55929
rect -3631 -56072 -3597 -55913
rect -3425 -55947 -3365 -55874
rect -3310 -55972 -3250 -55857
rect -3200 -55868 -3124 -55857
rect -3170 -55929 -3124 -55868
rect -3164 -56021 -3130 -55929
rect -3066 -56072 -3032 -55913
rect -2974 -55929 -2928 -55836
rect -2968 -56021 -2934 -55929
rect -2870 -56072 -2836 -55913
rect -2778 -55929 -2732 -55836
rect -2696 -55814 -2528 -55805
rect -2331 -55814 -2156 -55726
rect -1647 -55780 -1600 -55633
rect -1556 -55774 -1482 -55606
rect -1421 -55725 -1387 -55533
rect -2696 -55871 -2156 -55814
rect -1772 -55854 -1600 -55780
rect -2696 -55879 -2528 -55871
rect -2331 -55893 -2156 -55871
rect -2772 -56021 -2738 -55929
rect -2674 -56072 -2640 -55913
rect -2331 -55927 -1700 -55893
rect -2331 -55934 -2289 -55927
rect -2330 -55967 -2289 -55934
rect -2330 -55977 -2283 -55967
rect -4934 -56151 -4301 -56117
rect -4122 -56140 -2631 -56072
rect -2329 -56099 -2283 -55977
rect -2228 -56059 -2194 -55963
rect -2133 -55976 -2092 -55927
rect -2234 -56117 -2190 -56059
rect -2130 -56071 -2096 -55976
rect -2032 -56048 -1998 -55963
rect -1939 -55976 -1898 -55927
rect -2037 -56117 -1993 -56048
rect -1934 -56071 -1900 -55976
rect -1836 -56048 -1802 -55963
rect -1741 -55968 -1700 -55927
rect -1841 -56117 -1797 -56048
rect -1738 -56071 -1704 -55968
rect -1647 -55989 -1600 -55854
rect -1555 -55798 -1482 -55774
rect -1427 -55790 -1381 -55725
rect -1225 -55725 -1191 -55533
rect -1231 -55790 -1185 -55725
rect -1029 -55537 -995 -55533
rect -1035 -55790 -989 -55537
rect -831 -55719 -774 -55555
rect -539 -55725 -505 -55533
rect -1427 -55798 -989 -55790
rect -545 -55790 -499 -55725
rect -343 -55725 -309 -55533
rect -349 -55790 -303 -55725
rect -147 -55537 -113 -55533
rect -153 -55790 -107 -55537
rect -545 -55798 -107 -55790
rect -1555 -55836 -989 -55798
rect -1555 -55868 -1381 -55836
rect -1640 -56059 -1606 -55989
rect -1645 -56117 -1601 -56059
rect -2234 -56151 -1601 -56117
rect -1427 -55929 -1381 -55868
rect -1421 -56021 -1387 -55929
rect -1323 -56072 -1289 -55913
rect -1231 -55929 -1185 -55836
rect -1225 -56021 -1191 -55929
rect -1127 -56072 -1093 -55913
rect -1035 -55929 -989 -55836
rect -693 -55820 -633 -55816
rect -575 -55820 -107 -55798
rect 3498 -54596 5019 -54560
rect 3334 -55081 3470 -55035
rect 3230 -55165 3385 -55119
rect -693 -55836 -107 -55820
rect -693 -55862 -499 -55836
rect -1029 -56021 -995 -55929
rect -931 -56072 -897 -55913
rect -693 -55948 -633 -55862
rect -575 -55868 -499 -55862
rect -545 -55929 -499 -55868
rect -539 -56021 -505 -55929
rect -441 -56072 -407 -55913
rect -349 -55929 -303 -55836
rect -343 -56021 -309 -55929
rect -245 -56072 -211 -55913
rect -153 -55929 -107 -55836
rect -147 -56021 -113 -55929
rect -49 -56072 -15 -55913
rect -1422 -56140 -6 -56072
rect 391 -55960 425 -55550
rect 1129 -55794 1163 -55550
rect 1325 -55794 1359 -55550
rect 1521 -55794 1555 -55550
rect 1000 -55831 1555 -55794
rect 1741 -55797 1787 -55713
rect 2124 -55735 2158 -55563
rect 2320 -55671 2354 -55563
rect 2516 -55671 2550 -55563
rect 240 -56013 425 -55960
rect 460 -55969 595 -55959
rect 1000 -55969 1037 -55831
rect 1595 -55851 1787 -55797
rect 1987 -55805 2158 -55735
rect 2595 -55718 2668 -55705
rect 2595 -55746 2768 -55718
rect 2595 -55759 2790 -55746
rect 2595 -55765 2668 -55759
rect 1259 -55888 1394 -55879
rect 1822 -55888 1958 -55887
rect 1259 -55926 1958 -55888
rect 1259 -55933 1394 -55926
rect 1822 -55933 1958 -55926
rect 460 -56006 1037 -55969
rect 460 -56013 595 -56006
rect -5984 -56341 -5924 -56204
rect -3474 -56273 -3337 -56263
rect -2528 -56273 -2396 -56262
rect -514 -56273 -382 -56263
rect -5653 -56312 -382 -56273
rect -3474 -56323 -3337 -56312
rect -2528 -56322 -2396 -56312
rect -514 -56323 -382 -56312
rect -5983 -56713 -5935 -56341
rect -5636 -56365 -5499 -56352
rect -3039 -56365 -2902 -56346
rect -271 -56365 -139 -56346
rect -5653 -56404 -138 -56365
rect -5636 -56412 -5499 -56404
rect -5625 -56452 -5514 -56412
rect -4814 -56452 -4703 -56404
rect -3039 -56406 -2902 -56404
rect -5873 -56520 -4502 -56452
rect -4323 -56475 -3690 -56441
rect -3016 -56452 -2905 -56406
rect -2833 -56452 -2313 -56450
rect -2138 -56452 -2027 -56404
rect -5864 -56679 -5830 -56520
rect -5766 -56663 -5732 -56571
rect -5983 -56757 -5808 -56713
rect -5976 -56787 -5808 -56757
rect -5772 -56756 -5726 -56663
rect -5668 -56679 -5634 -56520
rect -5570 -56663 -5536 -56571
rect -5576 -56756 -5530 -56663
rect -5472 -56679 -5438 -56520
rect -5374 -56663 -5340 -56571
rect -5380 -56724 -5334 -56663
rect -5027 -56679 -4993 -56520
rect -4929 -56663 -4895 -56571
rect -5380 -56756 -5247 -56724
rect -5772 -56794 -5247 -56756
rect -4935 -56756 -4889 -56663
rect -4831 -56679 -4797 -56520
rect -4733 -56663 -4699 -56571
rect -4739 -56756 -4693 -56663
rect -4635 -56679 -4601 -56520
rect -4323 -56533 -4279 -56475
rect -4537 -56663 -4503 -56571
rect -4318 -56603 -4284 -56533
rect -4543 -56724 -4497 -56663
rect -4543 -56756 -4369 -56724
rect -5772 -56802 -5334 -56794
rect -5772 -57055 -5726 -56802
rect -5766 -57059 -5732 -57055
rect -5576 -56867 -5530 -56802
rect -5570 -57059 -5536 -56867
rect -5380 -56867 -5334 -56802
rect -5374 -57059 -5340 -56867
rect -5293 -56924 -5247 -56794
rect -4935 -56794 -4369 -56756
rect -4935 -56802 -4497 -56794
rect -5150 -56924 -5093 -56873
rect -5293 -56973 -5093 -56924
rect -5150 -57037 -5093 -56973
rect -4935 -57055 -4889 -56802
rect -4929 -57059 -4895 -57055
rect -4739 -56867 -4693 -56802
rect -4733 -57059 -4699 -56867
rect -4543 -56867 -4497 -56802
rect -4442 -56818 -4369 -56794
rect -4324 -56738 -4277 -56603
rect -4220 -56624 -4186 -56521
rect -4127 -56544 -4083 -56475
rect -4224 -56665 -4183 -56624
rect -4122 -56629 -4088 -56544
rect -4024 -56616 -3990 -56521
rect -3931 -56544 -3887 -56475
rect -4026 -56665 -3985 -56616
rect -3926 -56629 -3892 -56544
rect -3828 -56616 -3794 -56521
rect -3734 -56533 -3690 -56475
rect -3173 -56518 -1802 -56452
rect -3173 -56520 -2639 -56518
rect -2336 -56520 -1802 -56518
rect -1623 -56475 -990 -56441
rect -3832 -56665 -3791 -56616
rect -3730 -56629 -3696 -56533
rect -3632 -56615 -3598 -56521
rect -3635 -56658 -3594 -56615
rect -3635 -56665 -3593 -56658
rect -4224 -56699 -3593 -56665
rect -3164 -56679 -3130 -56520
rect -3066 -56663 -3032 -56571
rect -4324 -56812 -4152 -56738
rect -3768 -56759 -3502 -56699
rect -3276 -56720 -3108 -56713
rect -4537 -57059 -4503 -56867
rect -4442 -56986 -4368 -56818
rect -4324 -56959 -4277 -56812
rect -3768 -56866 -3593 -56759
rect -3298 -56780 -3108 -56720
rect -3276 -56787 -3108 -56780
rect -3072 -56756 -3026 -56663
rect -2968 -56679 -2934 -56520
rect -2870 -56663 -2836 -56571
rect -2876 -56756 -2830 -56663
rect -2772 -56679 -2738 -56520
rect -2674 -56663 -2640 -56571
rect -2680 -56724 -2634 -56663
rect -2499 -56713 -2439 -56554
rect -2327 -56679 -2293 -56520
rect -2229 -56663 -2195 -56571
rect -2680 -56756 -2536 -56724
rect -3072 -56794 -2536 -56756
rect -2499 -56776 -2271 -56713
rect -2439 -56787 -2271 -56776
rect -2235 -56756 -2189 -56663
rect -2131 -56679 -2097 -56520
rect -2033 -56663 -1999 -56571
rect -2039 -56756 -1993 -56663
rect -1935 -56679 -1901 -56520
rect -1623 -56533 -1579 -56475
rect -1837 -56663 -1803 -56571
rect -1618 -56603 -1584 -56533
rect -1843 -56724 -1797 -56663
rect -1843 -56756 -1669 -56724
rect -3072 -56802 -2634 -56794
rect -4221 -56900 -3593 -56866
rect -4221 -56952 -4185 -56900
rect -4023 -56936 -3987 -56900
rect -4318 -57033 -4284 -56959
rect -4319 -57078 -4283 -57033
rect -4220 -57044 -4186 -56952
rect -4122 -57023 -4088 -56936
rect -4024 -56954 -3987 -56936
rect -4123 -57078 -4081 -57023
rect -4024 -57044 -3990 -56954
rect -3926 -57022 -3892 -56936
rect -3829 -56954 -3793 -56900
rect -3929 -57078 -3887 -57022
rect -3828 -57044 -3794 -56954
rect -3730 -57027 -3696 -56936
rect -3635 -56944 -3593 -56900
rect -3733 -57078 -3691 -57027
rect -3632 -57044 -3598 -56944
rect -4319 -57112 -3691 -57078
rect -3072 -57055 -3026 -56802
rect -3066 -57059 -3032 -57055
rect -2876 -56867 -2830 -56802
rect -2870 -57059 -2836 -56867
rect -2680 -56867 -2634 -56802
rect -2674 -57059 -2640 -56867
rect -2598 -56923 -2536 -56794
rect -2235 -56794 -1669 -56756
rect -2235 -56802 -1797 -56794
rect -2450 -56923 -2393 -56873
rect -2598 -56985 -2393 -56923
rect -2450 -57037 -2393 -56985
rect -2235 -57055 -2189 -56802
rect -2229 -57059 -2195 -57055
rect -2039 -56867 -1993 -56802
rect -2033 -57059 -1999 -56867
rect -1843 -56867 -1797 -56802
rect -1742 -56818 -1669 -56794
rect -1624 -56738 -1577 -56603
rect -1520 -56624 -1486 -56521
rect -1427 -56544 -1383 -56475
rect -1524 -56665 -1483 -56624
rect -1422 -56629 -1388 -56544
rect -1324 -56616 -1290 -56521
rect -1231 -56544 -1187 -56475
rect -1326 -56665 -1285 -56616
rect -1226 -56629 -1192 -56544
rect -1128 -56616 -1094 -56521
rect -1034 -56533 -990 -56475
rect -1132 -56665 -1091 -56616
rect -1030 -56629 -996 -56533
rect -932 -56615 -898 -56521
rect -935 -56658 -894 -56615
rect -935 -56665 -893 -56658
rect -1524 -56697 -893 -56665
rect -1524 -56699 -818 -56697
rect -1624 -56812 -1452 -56738
rect -1068 -56757 -818 -56699
rect -1837 -57059 -1803 -56867
rect -1742 -56986 -1668 -56818
rect -1624 -56959 -1577 -56812
rect -1068 -56866 -893 -56757
rect -1521 -56900 -893 -56866
rect -1521 -56952 -1485 -56900
rect -1323 -56936 -1287 -56900
rect -1618 -57033 -1584 -56959
rect -1619 -57078 -1583 -57033
rect -1520 -57044 -1486 -56952
rect -1422 -57023 -1388 -56936
rect -1324 -56954 -1287 -56936
rect -1423 -57078 -1381 -57023
rect -1324 -57044 -1290 -56954
rect -1226 -57022 -1192 -56936
rect -1129 -56954 -1093 -56900
rect -1229 -57078 -1187 -57022
rect -1128 -57044 -1094 -56954
rect -1030 -57027 -996 -56936
rect -935 -56944 -893 -56900
rect -1033 -57078 -991 -57027
rect -932 -57044 -898 -56944
rect -654 -56984 -356 -56404
rect -271 -56406 -139 -56404
rect 391 -56466 425 -56013
rect 1000 -56060 1037 -56006
rect 1071 -55970 1206 -55957
rect 1993 -55970 2027 -55805
rect 2222 -55902 2256 -55794
rect 2320 -55950 2354 -55794
rect 2418 -55902 2452 -55794
rect 2516 -55950 2550 -55794
rect 2729 -55908 2790 -55759
rect 2929 -55908 2963 -55564
rect 3125 -55908 3159 -55564
rect 2729 -55938 3159 -55908
rect 3349 -55915 3385 -55165
rect 2740 -55946 3159 -55938
rect 3207 -55923 3385 -55915
rect 1071 -56004 2027 -55970
rect 1071 -56011 1206 -56004
rect 2075 -56036 2690 -55950
rect 3207 -55959 3394 -55923
rect 3207 -55963 3372 -55959
rect 3207 -55969 3342 -55963
rect 2803 -56019 2877 -55993
rect 3430 -56017 3470 -55081
rect 3729 -55737 3763 -55565
rect 3925 -55673 3959 -55565
rect 4121 -55673 4155 -55565
rect 3288 -56019 3470 -56017
rect 804 -56094 1037 -56060
rect 1210 -56094 1653 -56060
rect 489 -56654 523 -56258
rect 804 -56466 838 -56094
rect 902 -56564 936 -56158
rect 1000 -56466 1034 -56094
rect 1210 -56095 1457 -56094
rect 1210 -56158 1245 -56095
rect 1113 -56455 1147 -56158
rect 1112 -56561 1147 -56455
rect 1211 -56466 1245 -56158
rect 1309 -56457 1343 -56158
rect 1308 -56561 1343 -56457
rect 1423 -56465 1457 -56095
rect 1112 -56564 1343 -56561
rect 902 -56598 1343 -56564
rect 1521 -56654 1555 -56157
rect 1619 -56465 1653 -56094
rect 2385 -56443 2446 -56036
rect 2803 -56057 3470 -56019
rect 3565 -55807 3763 -55737
rect 4200 -55720 4273 -55707
rect 4200 -55748 4373 -55720
rect 4200 -55761 4395 -55748
rect 4200 -55767 4273 -55761
rect 2803 -56058 3289 -56057
rect 2803 -56064 2877 -56058
rect 3218 -56059 3289 -56058
rect 2831 -56409 2865 -56101
rect 2929 -56409 2963 -56101
rect 3027 -56409 3061 -56101
rect 3125 -56409 3159 -56101
rect 3223 -56409 3257 -56101
rect 2385 -56461 2835 -56443
rect 3125 -56461 3160 -56409
rect 2385 -56504 3277 -56461
rect 379 -56719 1653 -56654
rect 392 -56984 522 -56719
rect 698 -56984 828 -56719
rect 1015 -56984 1145 -56719
rect 1461 -56984 1591 -56719
rect 2385 -56984 2536 -56504
rect 2762 -56522 3277 -56504
rect 2762 -56984 2886 -56522
rect 3092 -56984 3216 -56522
rect 3565 -56542 3635 -55807
rect 3827 -55904 3861 -55796
rect 3925 -55952 3959 -55796
rect 4023 -55904 4057 -55796
rect 4121 -55952 4155 -55796
rect 4334 -55910 4395 -55761
rect 4534 -55910 4568 -55566
rect 4730 -55910 4764 -55566
rect 4334 -55940 4764 -55910
rect 4345 -55948 4764 -55940
rect 4812 -55923 4947 -55917
rect 4983 -55923 5019 -54596
rect 3680 -56038 4295 -55952
rect 4812 -55961 5019 -55923
rect 4812 -55963 4999 -55961
rect 4812 -55971 4947 -55963
rect 4408 -56021 4482 -55995
rect 5058 -56019 5098 -54526
rect 4893 -56021 5098 -56019
rect 3499 -56588 3635 -56542
rect 3990 -56445 4051 -56038
rect 4408 -56059 5098 -56021
rect 4408 -56060 4894 -56059
rect 4408 -56066 4482 -56060
rect 4823 -56061 4894 -56060
rect 4436 -56411 4470 -56103
rect 4534 -56411 4568 -56103
rect 4632 -56411 4666 -56103
rect 4730 -56411 4764 -56103
rect 4828 -56411 4862 -56103
rect 5353 -56141 5387 -55541
rect 6091 -55785 6125 -55541
rect 6287 -55785 6321 -55541
rect 6483 -55785 6517 -55541
rect 5962 -55822 6517 -55785
rect 6557 -55796 6692 -55788
rect 5422 -55960 5557 -55950
rect 5962 -55960 5999 -55822
rect 6556 -55833 6711 -55796
rect 6556 -55842 6692 -55833
rect 6221 -55879 6356 -55870
rect 6748 -55879 6782 -54510
rect 6221 -55917 6782 -55879
rect 6221 -55924 6356 -55917
rect 5422 -55997 5999 -55960
rect 5422 -56004 5557 -55997
rect 5962 -56051 5999 -55997
rect 6033 -55961 6168 -55948
rect 6818 -55961 6852 -54418
rect 6966 -55448 7694 -55414
rect 6966 -55760 7000 -55448
rect 7064 -55796 7098 -55552
rect 7162 -55760 7196 -55448
rect 7282 -55517 7624 -55483
rect 7282 -55760 7316 -55517
rect 7380 -55796 7414 -55552
rect 7478 -55760 7512 -55517
rect 6915 -55830 7529 -55796
rect 6033 -55995 6852 -55961
rect 6965 -55964 7104 -55910
rect 7495 -55945 7529 -55830
rect 7590 -55869 7624 -55517
rect 7660 -55795 7694 -55448
rect 7840 -55795 7874 -55552
rect 7660 -55829 7874 -55795
rect 8036 -55869 8070 -55552
rect 8346 -55745 8380 -55552
rect 7590 -55903 8070 -55869
rect 8123 -55920 8262 -55866
rect 7495 -55979 7641 -55945
rect 6033 -56002 6168 -55995
rect 5137 -56199 5387 -56141
rect 3990 -56463 4440 -56445
rect 4730 -56463 4765 -56411
rect 3990 -56506 4882 -56463
rect 3990 -56984 4141 -56506
rect 4432 -56524 4882 -56506
rect 4432 -56984 4583 -56524
rect 4725 -56984 4876 -56524
rect 5137 -56654 5202 -56199
rect 5353 -56457 5387 -56199
rect 5766 -56085 5999 -56051
rect 6172 -56085 6615 -56051
rect 5451 -56645 5485 -56249
rect 5766 -56457 5800 -56085
rect 5864 -56555 5898 -56149
rect 5962 -56457 5996 -56085
rect 6172 -56086 6419 -56085
rect 6172 -56149 6207 -56086
rect 6075 -56446 6109 -56149
rect 6074 -56552 6109 -56446
rect 6173 -56457 6207 -56149
rect 6271 -56448 6305 -56149
rect 6270 -56552 6305 -56448
rect 6385 -56456 6419 -56086
rect 6074 -56555 6305 -56552
rect 5864 -56589 6305 -56555
rect 6483 -56645 6517 -56148
rect 6581 -56456 6615 -56085
rect 6964 -56082 7295 -56045
rect 7607 -56041 7641 -55979
rect 7714 -55994 7853 -55940
rect 7607 -56075 8168 -56041
rect 6964 -56165 7001 -56082
rect 7258 -56106 7295 -56082
rect 7258 -56143 7414 -56106
rect 6966 -56354 7000 -56165
rect 6962 -56477 7001 -56354
rect 7064 -56403 7098 -56158
rect 7377 -56164 7414 -56143
rect 7380 -56366 7414 -56164
rect 7476 -56167 7776 -56128
rect 7478 -56366 7512 -56167
rect 7742 -56366 7776 -56167
rect 7840 -56366 7874 -56075
rect 8036 -56349 8070 -56158
rect 8036 -56403 8072 -56349
rect 8134 -56366 8168 -56075
rect 8341 -56084 8384 -55745
rect 8655 -55743 8689 -55552
rect 8651 -55940 8694 -55743
rect 8738 -55926 8877 -55872
rect 8551 -55986 8694 -55940
rect 8245 -56130 8384 -56084
rect 8341 -56175 8384 -56130
rect 8346 -56366 8380 -56175
rect 8444 -56359 8478 -56158
rect 8651 -56177 8694 -55986
rect 7064 -56439 8072 -56403
rect 8439 -56443 8482 -56359
rect 8655 -56366 8689 -56177
rect 8753 -56357 8787 -56158
rect 8748 -56443 8791 -56357
rect 8163 -56477 8795 -56443
rect 6962 -56530 8795 -56477
rect 5067 -56700 5203 -56654
rect 5341 -56710 6615 -56645
rect 5365 -56984 5511 -56710
rect 5810 -56984 5956 -56710
rect 6076 -56984 6222 -56710
rect 6436 -56984 6582 -56710
rect 7000 -56984 7197 -56530
rect 7533 -56984 7730 -56530
rect 8046 -56539 8795 -56530
rect 8046 -56984 8243 -56539
rect 8549 -56984 8746 -56539
rect 8944 -56984 9205 -54301
rect 9641 -54352 16907 -54213
rect 16582 -55232 16849 -55196
rect 11237 -55467 16849 -55232
rect 16582 -55494 16849 -55467
rect 9669 -55826 9887 -55818
rect 16845 -55826 16998 -55787
rect 9669 -55901 16998 -55826
rect 9669 -55907 9887 -55901
rect 16845 -55938 16998 -55901
rect 10651 -56047 10701 -56041
rect 16163 -56047 16261 -56033
rect 10642 -56170 16261 -56047
rect 10651 -56174 10701 -56170
rect 16163 -56197 16261 -56170
rect 17080 -56452 17208 -53540
rect 17333 -56363 17465 -53112
rect 17575 -55787 17664 -52637
rect 19667 -53851 20212 -52313
rect 19084 -54357 85057 -53851
rect 17575 -55938 17672 -55787
rect 19667 -55821 20212 -54357
rect 29413 -54818 29696 -54357
rect 29169 -54846 29834 -54818
rect 34781 -54833 35138 -54766
rect 35959 -54833 36316 -54800
rect 37812 -54829 38095 -54357
rect 29169 -54904 30204 -54846
rect 29169 -54985 29255 -54904
rect 29429 -54941 29464 -54904
rect 29754 -54907 30204 -54904
rect 28317 -55071 29255 -54985
rect 28165 -55361 28295 -55269
rect 28457 -55327 28491 -55071
rect 28555 -55327 28589 -55119
rect 28653 -55327 28687 -55071
rect 28751 -55293 28785 -55119
rect 29332 -55249 29366 -54941
rect 29430 -55249 29464 -54941
rect 29528 -55249 29562 -54941
rect 29626 -55249 29660 -54941
rect 29724 -55249 29758 -54941
rect 29300 -55292 29371 -55291
rect 29712 -55292 29786 -55286
rect 29300 -55293 29786 -55292
rect 28751 -55327 29786 -55293
rect 30143 -55314 30204 -54907
rect 34781 -55022 36316 -54833
rect 37609 -54857 38274 -54829
rect 37609 -54915 38644 -54857
rect 46724 -54868 47007 -54357
rect 55943 -54834 56226 -54357
rect 61292 -54802 61668 -54707
rect 64738 -54768 65045 -54357
rect 62893 -54802 63143 -54775
rect 37609 -54996 37695 -54915
rect 37869 -54952 37904 -54915
rect 38194 -54918 38644 -54915
rect 34781 -55033 35138 -55022
rect 35959 -55067 36316 -55022
rect 36757 -55082 37695 -54996
rect 28752 -55331 29786 -55327
rect 28752 -55333 29301 -55331
rect 28339 -55361 28412 -55355
rect 29712 -55357 29786 -55331
rect 28165 -55402 28412 -55361
rect 28165 -55419 28295 -55402
rect 28339 -55415 28412 -55402
rect 29899 -55400 30684 -55314
rect 36605 -55372 36735 -55280
rect 36897 -55338 36931 -55082
rect 36995 -55338 37029 -55130
rect 37093 -55338 37127 -55082
rect 37191 -55304 37225 -55130
rect 37772 -55260 37806 -54952
rect 37870 -55260 37904 -54952
rect 37968 -55260 38002 -54952
rect 38066 -55260 38100 -54952
rect 38164 -55260 38198 -54952
rect 37740 -55303 37811 -55302
rect 38152 -55303 38226 -55297
rect 37740 -55304 38226 -55303
rect 37191 -55338 38226 -55304
rect 38583 -55325 38644 -54918
rect 43337 -54922 43602 -54891
rect 44863 -54922 45160 -54889
rect 43337 -55089 45160 -54922
rect 46472 -54896 47137 -54868
rect 46472 -54954 47507 -54896
rect 46472 -55035 46558 -54954
rect 46732 -54991 46767 -54954
rect 47057 -54957 47507 -54954
rect 43337 -55156 43602 -55089
rect 44863 -55111 45160 -55089
rect 45620 -55121 46558 -55035
rect 37192 -55342 38226 -55338
rect 37192 -55344 37741 -55342
rect 36779 -55372 36852 -55366
rect 38152 -55368 38226 -55342
rect 29430 -55412 29849 -55404
rect 29430 -55442 29860 -55412
rect 28457 -55657 28491 -55449
rect 28653 -55657 28687 -55449
rect 28849 -55657 28883 -55449
rect 21077 -55783 21705 -55749
rect 17575 -56271 17664 -55938
rect 18769 -55927 20539 -55821
rect 20984 -55917 21018 -55817
rect 21077 -55834 21119 -55783
rect 18873 -56073 18921 -55927
rect 18878 -56244 18912 -56073
rect 18976 -56227 19010 -56036
rect 19067 -56076 19115 -55927
rect 18692 -56271 18837 -56264
rect 17575 -56312 18837 -56271
rect 18692 -56320 18837 -56312
rect 18972 -56278 19014 -56227
rect 19074 -56244 19108 -56076
rect 19172 -56227 19206 -56036
rect 19168 -56278 19210 -56227
rect 18972 -56320 19758 -56278
rect 19619 -56338 19758 -56320
rect 19021 -56363 19166 -56359
rect 17333 -56404 19166 -56363
rect 19021 -56415 19166 -56404
rect 19341 -56447 19486 -56391
rect 19341 -56452 19401 -56447
rect 17080 -56493 19401 -56452
rect 19619 -56520 19661 -56338
rect 18874 -56566 19323 -56529
rect -1619 -57112 -991 -57078
rect -11819 -57239 -11664 -57237
rect -11799 -57247 -11664 -57239
rect -12294 -57297 -11745 -57295
rect -11334 -57297 -11260 -57271
rect -12294 -57301 -11260 -57297
rect -12589 -57557 -12555 -57301
rect -12491 -57509 -12457 -57301
rect -12393 -57557 -12359 -57301
rect -12295 -57335 -11260 -57301
rect -11147 -57314 -10362 -57228
rect -12295 -57509 -12261 -57335
rect -11746 -57336 -11260 -57335
rect -11746 -57337 -11675 -57336
rect -11334 -57342 -11260 -57336
rect -12729 -57643 -11791 -57557
rect -11877 -57724 -11791 -57643
rect -11714 -57687 -11680 -57379
rect -11616 -57687 -11582 -57379
rect -11518 -57687 -11484 -57379
rect -11420 -57687 -11386 -57379
rect -11322 -57687 -11288 -57379
rect -11617 -57724 -11582 -57687
rect -10903 -57721 -10842 -57314
rect -11292 -57724 -10842 -57721
rect -11877 -57782 -10842 -57724
rect -11877 -57810 -11212 -57782
rect -27236 -60993 -26896 -60851
rect -23096 -62272 -22910 -57887
rect -15693 -57919 -15425 -57887
rect -13640 -58026 -13606 -58022
rect -13646 -58279 -13600 -58026
rect -13444 -58214 -13410 -58022
rect -13450 -58279 -13404 -58214
rect -13248 -58214 -13214 -58022
rect -13024 -58108 -12967 -58044
rect -13167 -58157 -12967 -58108
rect -13254 -58279 -13208 -58214
rect -13646 -58287 -13208 -58279
rect -13167 -58287 -13121 -58157
rect -13024 -58208 -12967 -58157
rect -12803 -58026 -12769 -58022
rect -13850 -58324 -13682 -58294
rect -13857 -58368 -13682 -58324
rect -13646 -58325 -13121 -58287
rect -12809 -58279 -12763 -58026
rect -12607 -58214 -12573 -58022
rect -12613 -58279 -12567 -58214
rect -12193 -58003 -11565 -57969
rect -12411 -58214 -12377 -58022
rect -12193 -58048 -12157 -58003
rect -12417 -58279 -12371 -58214
rect -12809 -58287 -12371 -58279
rect -12316 -58263 -12242 -58095
rect -12192 -58122 -12158 -58048
rect -12316 -58287 -12243 -58263
rect -13013 -58305 -12845 -58294
rect -13048 -58306 -12845 -58305
rect -21117 -59698 -21083 -59107
rect -20817 -59071 -20354 -59037
rect -21121 -59749 -21080 -59698
rect -20905 -59705 -20871 -59107
rect -20817 -59113 -20764 -59071
rect -20910 -59749 -20868 -59705
rect -20807 -59715 -20773 -59113
rect -20709 -59704 -20675 -59107
rect -20608 -59113 -20552 -59071
rect -20714 -59749 -20672 -59704
rect -20596 -59715 -20562 -59113
rect -20498 -59697 -20464 -59107
rect -20410 -59113 -20354 -59071
rect -21121 -59786 -20672 -59749
rect -20502 -59753 -20460 -59697
rect -20400 -59715 -20366 -59113
rect -19911 -59439 -19877 -59036
rect -19707 -59000 -19463 -58962
rect -19912 -59478 -19876 -59439
rect -19707 -59064 -19661 -59000
rect -19700 -59444 -19666 -59064
rect -19602 -59434 -19568 -59036
rect -19509 -59064 -19463 -59000
rect -19504 -59398 -19470 -59064
rect -19609 -59478 -19564 -59434
rect -19912 -59514 -19564 -59478
rect -19507 -59630 -19457 -59398
rect -19006 -59440 -18972 -59037
rect -18802 -59001 -18558 -58963
rect -19273 -59561 -19215 -59466
rect -19007 -59479 -18971 -59440
rect -18802 -59065 -18756 -59001
rect -18795 -59445 -18761 -59065
rect -18697 -59435 -18663 -59037
rect -18604 -59065 -18558 -59001
rect -16891 -59039 -15414 -58926
rect -18599 -59399 -18565 -59065
rect -17722 -59334 -17273 -59316
rect -16891 -59334 -16830 -59039
rect -16164 -59157 -16117 -59039
rect -18234 -59395 -16830 -59334
rect -18704 -59479 -18659 -59435
rect -19007 -59515 -18659 -59479
rect -18877 -59561 -18734 -59554
rect -19273 -59597 -18734 -59561
rect -19273 -59603 -19215 -59597
rect -18877 -59614 -18734 -59597
rect -20114 -59649 -20056 -59636
rect -20005 -59649 -19859 -59633
rect -19507 -59643 -19361 -59630
rect -18602 -59631 -18552 -59399
rect -20114 -59685 -19859 -59649
rect -19563 -59652 -19361 -59643
rect -20502 -59795 -20334 -59753
rect -20114 -59773 -20056 -59685
rect -20005 -59693 -19859 -59685
rect -19818 -59688 -19361 -59652
rect -19196 -59650 -19138 -59638
rect -19100 -59650 -18954 -59634
rect -18602 -59644 -18430 -59631
rect -19196 -59686 -18954 -59650
rect -18658 -59653 -18430 -59644
rect -20376 -59979 -20334 -59795
rect -19911 -59887 -19877 -59728
rect -19818 -59737 -19773 -59688
rect -20385 -59995 -20248 -59979
rect -21023 -60037 -20248 -59995
rect -21117 -60242 -21083 -60071
rect -21023 -60088 -20981 -60037
rect -21122 -60371 -21074 -60242
rect -21019 -60279 -20985 -60088
rect -20921 -60239 -20887 -60071
rect -20827 -60088 -20785 -60037
rect -19915 -60039 -19871 -59887
rect -19813 -59936 -19779 -59737
rect -19715 -59888 -19681 -59728
rect -19196 -59775 -19138 -59686
rect -19100 -59694 -18954 -59686
rect -18913 -59689 -18430 -59653
rect -19006 -59888 -18972 -59729
rect -18913 -59738 -18868 -59689
rect -19721 -60039 -19677 -59888
rect -20044 -60074 -19447 -60039
rect -19010 -60040 -18966 -59888
rect -18908 -59937 -18874 -59738
rect -18810 -59889 -18776 -59729
rect -18234 -59753 -18173 -59395
rect -17605 -59429 -17570 -59395
rect -17702 -59737 -17668 -59429
rect -17604 -59737 -17570 -59429
rect -17506 -59737 -17472 -59429
rect -17408 -59737 -17374 -59429
rect -17310 -59737 -17276 -59429
rect -18621 -59814 -18173 -59753
rect -17734 -59780 -17663 -59779
rect -17322 -59780 -17248 -59774
rect -17734 -59781 -17248 -59780
rect -18816 -60040 -18772 -59889
rect -18621 -60040 -18560 -59814
rect -17960 -59819 -17248 -59781
rect -16891 -59802 -16830 -59395
rect -16157 -59451 -16123 -59157
rect -16059 -59435 -16025 -59143
rect -15968 -59158 -15921 -59039
rect -16266 -59497 -16111 -59485
rect -16303 -59531 -16111 -59497
rect -16266 -59540 -16111 -59531
rect -16065 -59505 -16020 -59435
rect -15961 -59451 -15927 -59158
rect -15726 -59168 -15679 -59039
rect -15719 -59451 -15685 -59168
rect -15621 -59442 -15587 -59143
rect -15625 -59482 -15581 -59442
rect -14733 -59482 -14596 -59412
rect -15625 -59485 -14596 -59482
rect -16065 -59545 -15711 -59505
rect -15673 -59525 -14596 -59485
rect -16401 -59602 -16331 -59600
rect -15996 -59602 -15841 -59593
rect -16401 -59638 -15841 -59602
rect -17960 -59821 -17733 -59819
rect -17322 -59845 -17248 -59819
rect -18306 -59879 -18189 -59864
rect -17787 -59877 -17652 -59869
rect -17807 -59879 -17652 -59877
rect -18306 -59915 -17652 -59879
rect -17135 -59888 -16520 -59802
rect -18306 -59987 -18189 -59915
rect -17807 -59917 -17652 -59915
rect -17787 -59923 -17652 -59917
rect -17604 -59900 -17185 -59892
rect -17604 -59930 -17174 -59900
rect -19139 -60074 -18542 -60040
rect -20928 -60371 -20880 -60239
rect -20823 -60279 -20789 -60088
rect -20599 -60129 -18542 -60074
rect -20599 -60190 -18758 -60129
rect -20599 -60371 -20483 -60190
rect -21257 -60388 -20453 -60371
rect -17604 -60274 -17570 -59930
rect -17408 -60274 -17374 -59930
rect -17235 -60079 -17174 -59930
rect -16995 -60044 -16961 -59888
rect -16897 -60044 -16863 -59936
rect -16799 -60044 -16765 -59888
rect -16701 -60044 -16667 -59936
rect -16401 -60033 -16331 -59638
rect -15996 -59648 -15841 -59638
rect -15754 -59615 -15711 -59545
rect -15754 -59670 -15573 -59615
rect -15754 -59682 -15711 -59670
rect -16161 -59720 -15907 -59684
rect -17113 -60079 -17040 -60073
rect -17235 -60092 -17040 -60079
rect -17213 -60120 -17040 -60092
rect -17113 -60133 -17040 -60120
rect -16603 -60103 -16325 -60033
rect -16995 -60275 -16961 -60167
rect -16799 -60275 -16765 -60167
rect -16603 -60275 -16569 -60103
rect -16161 -59779 -16119 -59720
rect -21257 -60494 -20369 -60388
rect -16157 -60363 -16123 -59779
rect -15949 -59773 -15907 -59720
rect -15852 -59721 -15711 -59682
rect -15946 -60355 -15912 -59773
rect -15852 -59775 -15810 -59721
rect -15950 -60397 -15908 -60355
rect -15848 -60363 -15814 -59775
rect -15750 -60353 -15716 -59755
rect -15539 -59769 -15496 -59525
rect -14733 -59578 -14596 -59525
rect -15313 -59700 -15208 -59628
rect -13857 -58740 -13809 -58368
rect -13738 -58561 -13704 -58402
rect -13646 -58418 -13600 -58325
rect -13640 -58510 -13606 -58418
rect -13542 -58561 -13508 -58402
rect -13450 -58418 -13404 -58325
rect -13254 -58357 -13121 -58325
rect -13444 -58510 -13410 -58418
rect -13346 -58561 -13312 -58402
rect -13254 -58418 -13208 -58357
rect -13085 -58368 -12845 -58306
rect -12809 -58325 -12243 -58287
rect -13248 -58510 -13214 -58418
rect -13085 -58512 -13025 -58368
rect -12901 -58561 -12867 -58402
rect -12809 -58418 -12763 -58325
rect -12803 -58510 -12769 -58418
rect -12705 -58561 -12671 -58402
rect -12613 -58418 -12567 -58325
rect -12417 -58357 -12243 -58325
rect -12198 -58269 -12151 -58122
rect -12094 -58129 -12060 -58037
rect -11997 -58058 -11955 -58003
rect -12095 -58181 -12059 -58129
rect -11996 -58145 -11962 -58058
rect -11898 -58127 -11864 -58037
rect -11803 -58059 -11761 -58003
rect -11898 -58145 -11861 -58127
rect -11800 -58145 -11766 -58059
rect -11702 -58127 -11668 -58037
rect -11607 -58054 -11565 -58003
rect -11897 -58181 -11861 -58145
rect -11703 -58181 -11667 -58127
rect -11604 -58145 -11570 -58054
rect -11506 -58137 -11472 -58037
rect -11509 -58181 -11467 -58137
rect -12095 -58215 -11467 -58181
rect -12198 -58343 -12026 -58269
rect -11642 -58322 -11467 -58215
rect -10940 -58026 -10906 -58022
rect -10946 -58279 -10900 -58026
rect -10744 -58214 -10710 -58022
rect -10750 -58279 -10704 -58214
rect -10548 -58214 -10514 -58022
rect -10324 -58096 -10267 -58044
rect -10472 -58158 -10267 -58096
rect -10554 -58279 -10508 -58214
rect -10946 -58287 -10508 -58279
rect -10472 -58287 -10410 -58158
rect -10324 -58208 -10267 -58158
rect -10103 -58026 -10069 -58022
rect -11150 -58301 -10982 -58294
rect -12607 -58510 -12573 -58418
rect -12509 -58561 -12475 -58402
rect -12417 -58418 -12371 -58357
rect -12411 -58510 -12377 -58418
rect -12198 -58478 -12151 -58343
rect -11642 -58382 -11376 -58322
rect -11172 -58361 -10982 -58301
rect -11150 -58368 -10982 -58361
rect -10946 -58325 -10410 -58287
rect -10109 -58279 -10063 -58026
rect -9907 -58214 -9873 -58022
rect -9913 -58279 -9867 -58214
rect -9493 -58003 -8865 -57969
rect -9711 -58214 -9677 -58022
rect -9493 -58048 -9457 -58003
rect -9717 -58279 -9671 -58214
rect -10109 -58287 -9671 -58279
rect -9616 -58263 -9542 -58095
rect -9492 -58122 -9458 -58048
rect -9616 -58287 -9543 -58263
rect -10313 -58305 -10145 -58294
rect -12098 -58416 -11467 -58382
rect -12098 -58457 -12057 -58416
rect -12192 -58548 -12158 -58478
rect -13747 -58629 -12376 -58561
rect -12197 -58606 -12153 -58548
rect -12094 -58560 -12060 -58457
rect -11996 -58537 -11962 -58452
rect -11900 -58465 -11859 -58416
rect -12001 -58606 -11957 -58537
rect -11898 -58560 -11864 -58465
rect -11800 -58537 -11766 -58452
rect -11706 -58465 -11665 -58416
rect -11509 -58423 -11467 -58416
rect -11805 -58606 -11761 -58537
rect -11702 -58560 -11668 -58465
rect -11604 -58548 -11570 -58452
rect -11509 -58466 -11468 -58423
rect -11608 -58606 -11564 -58548
rect -11506 -58560 -11472 -58466
rect -11038 -58561 -11004 -58402
rect -10946 -58418 -10900 -58325
rect -10940 -58510 -10906 -58418
rect -10842 -58561 -10808 -58402
rect -10750 -58418 -10704 -58325
rect -10554 -58357 -10410 -58325
rect -10744 -58510 -10710 -58418
rect -10646 -58561 -10612 -58402
rect -10554 -58418 -10508 -58357
rect -10373 -58368 -10145 -58305
rect -10109 -58325 -9543 -58287
rect -10548 -58510 -10514 -58418
rect -10373 -58527 -10313 -58368
rect -10201 -58561 -10167 -58402
rect -10109 -58418 -10063 -58325
rect -10103 -58510 -10069 -58418
rect -10005 -58561 -9971 -58402
rect -9913 -58418 -9867 -58325
rect -9717 -58357 -9543 -58325
rect -9498 -58269 -9451 -58122
rect -9394 -58129 -9360 -58037
rect -9297 -58058 -9255 -58003
rect -9395 -58181 -9359 -58129
rect -9296 -58145 -9262 -58058
rect -9198 -58127 -9164 -58037
rect -9103 -58059 -9061 -58003
rect -9198 -58145 -9161 -58127
rect -9100 -58145 -9066 -58059
rect -9002 -58127 -8968 -58037
rect -8907 -58054 -8865 -58003
rect -9197 -58181 -9161 -58145
rect -9003 -58181 -8967 -58127
rect -8904 -58145 -8870 -58054
rect -8806 -58137 -8772 -58037
rect -8809 -58181 -8767 -58137
rect -9395 -58215 -8767 -58181
rect -9498 -58343 -9326 -58269
rect -8942 -58324 -8767 -58215
rect -9907 -58510 -9873 -58418
rect -9809 -58561 -9775 -58402
rect -9717 -58418 -9671 -58357
rect -9711 -58510 -9677 -58418
rect -9498 -58478 -9451 -58343
rect -8942 -58382 -8692 -58324
rect -9398 -58384 -8692 -58382
rect -9398 -58416 -8767 -58384
rect -9398 -58457 -9357 -58416
rect -9492 -58548 -9458 -58478
rect -13499 -58669 -13388 -58629
rect -13510 -58677 -13373 -58669
rect -12688 -58677 -12577 -58629
rect -12197 -58640 -11564 -58606
rect -11047 -58563 -10513 -58561
rect -10210 -58563 -9676 -58561
rect -11047 -58629 -9676 -58563
rect -9497 -58606 -9453 -58548
rect -9394 -58560 -9360 -58457
rect -9296 -58537 -9262 -58452
rect -9200 -58465 -9159 -58416
rect -9301 -58606 -9257 -58537
rect -9198 -58560 -9164 -58465
rect -9100 -58537 -9066 -58452
rect -9006 -58465 -8965 -58416
rect -8809 -58423 -8767 -58416
rect -9105 -58606 -9061 -58537
rect -9002 -58560 -8968 -58465
rect -8904 -58548 -8870 -58452
rect -8809 -58466 -8768 -58423
rect -8908 -58606 -8864 -58548
rect -8806 -58560 -8772 -58466
rect -10890 -58675 -10779 -58629
rect -10707 -58631 -10187 -58629
rect -10913 -58677 -10776 -58675
rect -10012 -58677 -9901 -58629
rect -9497 -58640 -8864 -58606
rect -7447 -58633 -7413 -58039
rect -7241 -58005 -7001 -57971
rect -7241 -58049 -7199 -58005
rect -8275 -58677 -8143 -58675
rect -13527 -58716 -8142 -58677
rect -13510 -58729 -13373 -58716
rect -10913 -58735 -10776 -58716
rect -8275 -58735 -8143 -58716
rect -13858 -58877 -13798 -58740
rect -11348 -58769 -11211 -58758
rect -10402 -58769 -10270 -58759
rect -13527 -58808 -7797 -58769
rect -11348 -58818 -11211 -58808
rect -10402 -58819 -10270 -58808
rect -13121 -58855 -12989 -58847
rect -8598 -58855 -8466 -58845
rect -13857 -59235 -13809 -58877
rect -13527 -58894 -8466 -58855
rect -13121 -58907 -12989 -58894
rect -8598 -58905 -8466 -58894
rect -7836 -58877 -7797 -58808
rect -7455 -58877 -7412 -58633
rect -7235 -58647 -7201 -58049
rect -7137 -58627 -7103 -58039
rect -7043 -58047 -7001 -58005
rect -7141 -58681 -7099 -58627
rect -7039 -58629 -7005 -58047
rect -7240 -58720 -7099 -58681
rect -7044 -58682 -7002 -58629
rect -6828 -58623 -6794 -58039
rect -6832 -58682 -6790 -58623
rect -654 -57245 9205 -56984
rect 18874 -56617 18915 -56566
rect -654 -58103 -356 -57245
rect 955 -58103 1216 -57245
rect 1792 -58103 2053 -57245
rect 2832 -58103 3093 -57245
rect 4290 -58103 4551 -57245
rect 5504 -58103 5765 -57245
rect 7450 -58103 7711 -57245
rect 8944 -58103 9205 -57245
rect 18878 -57208 18912 -56617
rect 19085 -56610 19127 -56566
rect 19090 -57208 19124 -56610
rect 19188 -57202 19222 -56600
rect 19281 -56611 19323 -56566
rect 19493 -56562 19661 -56520
rect 19178 -57244 19231 -57202
rect 19286 -57208 19320 -56611
rect 19399 -57202 19433 -56600
rect 19493 -56618 19535 -56562
rect 19387 -57244 19443 -57202
rect 19497 -57208 19531 -56618
rect 19595 -57202 19629 -56600
rect 19585 -57244 19641 -57202
rect 19178 -57278 19641 -57244
rect -7044 -58718 -6790 -58682
rect -7240 -58732 -7197 -58720
rect -7378 -58787 -7197 -58732
rect -7240 -58857 -7197 -58787
rect -7110 -58764 -6955 -58754
rect -6597 -58764 -6465 -58712
rect -7110 -58800 -6465 -58764
rect -7110 -58809 -6955 -58800
rect -7836 -58917 -7278 -58877
rect -7240 -58897 -6886 -58857
rect -7836 -58920 -7326 -58917
rect -13739 -59009 -13205 -58941
rect -12808 -58964 -12175 -58930
rect -13738 -59152 -13704 -59060
rect -13744 -59213 -13698 -59152
rect -13640 -59168 -13606 -59009
rect -13542 -59152 -13508 -59060
rect -13774 -59235 -13698 -59213
rect -13857 -59245 -13698 -59235
rect -13548 -59245 -13502 -59152
rect -13444 -59168 -13410 -59009
rect -13346 -59152 -13312 -59060
rect -13352 -59245 -13306 -59152
rect -13248 -59168 -13214 -59009
rect -12900 -59104 -12866 -59010
rect -12808 -59022 -12764 -58964
rect -12904 -59147 -12863 -59104
rect -12802 -59118 -12768 -59022
rect -12704 -59105 -12670 -59010
rect -12611 -59033 -12567 -58964
rect -12905 -59154 -12863 -59147
rect -12707 -59154 -12666 -59105
rect -12606 -59118 -12572 -59033
rect -12508 -59105 -12474 -59010
rect -12415 -59033 -12371 -58964
rect -12513 -59154 -12472 -59105
rect -12410 -59118 -12376 -59033
rect -12312 -59113 -12278 -59010
rect -12219 -59022 -12175 -58964
rect -11996 -59009 -10505 -58941
rect -10108 -58964 -9475 -58930
rect -12214 -59092 -12180 -59022
rect -12315 -59154 -12274 -59113
rect -12905 -59188 -12274 -59154
rect -13857 -59272 -13306 -59245
rect -13856 -59274 -13306 -59272
rect -13774 -59283 -13306 -59274
rect -13270 -59217 -13102 -59202
rect -12905 -59217 -12730 -59188
rect -13270 -59270 -12730 -59217
rect -12221 -59227 -12174 -59092
rect -11995 -59152 -11961 -59060
rect -12001 -59213 -11955 -59152
rect -11897 -59168 -11863 -59009
rect -11799 -59152 -11765 -59060
rect -13270 -59276 -13102 -59270
rect -13744 -59291 -13306 -59283
rect -13744 -59356 -13698 -59291
rect -13738 -59548 -13704 -59356
rect -13548 -59356 -13502 -59291
rect -13542 -59548 -13508 -59356
rect -13352 -59544 -13306 -59291
rect -13346 -59548 -13312 -59544
rect -12905 -59355 -12730 -59270
rect -12346 -59301 -12174 -59227
rect -12905 -59389 -12277 -59355
rect -12905 -59433 -12863 -59389
rect -12900 -59533 -12866 -59433
rect -12802 -59516 -12768 -59425
rect -12705 -59443 -12669 -59389
rect -12511 -59425 -12475 -59389
rect -12807 -59567 -12765 -59516
rect -12704 -59533 -12670 -59443
rect -12606 -59511 -12572 -59425
rect -12511 -59443 -12474 -59425
rect -12611 -59567 -12569 -59511
rect -12508 -59533 -12474 -59443
rect -12410 -59512 -12376 -59425
rect -12313 -59441 -12277 -59389
rect -12417 -59567 -12375 -59512
rect -12312 -59533 -12278 -59441
rect -12221 -59448 -12174 -59301
rect -12129 -59245 -11955 -59213
rect -11805 -59245 -11759 -59152
rect -11701 -59168 -11667 -59009
rect -11603 -59152 -11569 -59060
rect -11609 -59245 -11563 -59152
rect -11505 -59168 -11471 -59009
rect -12129 -59283 -11563 -59245
rect -11527 -59207 -11359 -59202
rect -11299 -59207 -11239 -59134
rect -11527 -59265 -11239 -59207
rect -11184 -59224 -11124 -59109
rect -11038 -59152 -11004 -59060
rect -11044 -59213 -10998 -59152
rect -10940 -59168 -10906 -59009
rect -10842 -59152 -10808 -59060
rect -11074 -59224 -10998 -59213
rect -11527 -59276 -11359 -59265
rect -11299 -59266 -11239 -59265
rect -11189 -59245 -10998 -59224
rect -10848 -59245 -10802 -59152
rect -10744 -59168 -10710 -59009
rect -10646 -59152 -10612 -59060
rect -10652 -59245 -10606 -59152
rect -10548 -59168 -10514 -59009
rect -10203 -59104 -10157 -58982
rect -10108 -59022 -10064 -58964
rect -10204 -59114 -10157 -59104
rect -10204 -59147 -10163 -59114
rect -10102 -59118 -10068 -59022
rect -10004 -59105 -9970 -59010
rect -9911 -59033 -9867 -58964
rect -10205 -59154 -10163 -59147
rect -10007 -59154 -9966 -59105
rect -9906 -59118 -9872 -59033
rect -9808 -59105 -9774 -59010
rect -9715 -59033 -9671 -58964
rect -9813 -59154 -9772 -59105
rect -9710 -59118 -9676 -59033
rect -9612 -59113 -9578 -59010
rect -9519 -59022 -9475 -58964
rect -9296 -59009 -7880 -58941
rect -9514 -59092 -9480 -59022
rect -9615 -59154 -9574 -59113
rect -10205 -59188 -9574 -59154
rect -11189 -59269 -10606 -59245
rect -12129 -59307 -12056 -59283
rect -12214 -59522 -12180 -59448
rect -12130 -59475 -12056 -59307
rect -12001 -59291 -11563 -59283
rect -12001 -59356 -11955 -59291
rect -12215 -59567 -12179 -59522
rect -11995 -59548 -11961 -59356
rect -12807 -59601 -12179 -59567
rect -11805 -59356 -11759 -59291
rect -11799 -59548 -11765 -59356
rect -11609 -59544 -11563 -59291
rect -11603 -59548 -11569 -59544
rect -11405 -59403 -11348 -59362
rect -11189 -59403 -11144 -59269
rect -11074 -59283 -10606 -59269
rect -10570 -59210 -10402 -59202
rect -10205 -59210 -10030 -59188
rect -10570 -59267 -10030 -59210
rect -9521 -59227 -9474 -59092
rect -9295 -59152 -9261 -59060
rect -9301 -59213 -9255 -59152
rect -9197 -59168 -9163 -59009
rect -9099 -59152 -9065 -59060
rect -10570 -59276 -10402 -59267
rect -11044 -59291 -10606 -59283
rect -11044 -59356 -10998 -59291
rect -11405 -59448 -11144 -59403
rect -11405 -59526 -11348 -59448
rect -11038 -59548 -11004 -59356
rect -10848 -59356 -10802 -59291
rect -10842 -59548 -10808 -59356
rect -10652 -59544 -10606 -59291
rect -10646 -59548 -10612 -59544
rect -10205 -59355 -10030 -59267
rect -9646 -59301 -9474 -59227
rect -10205 -59389 -9577 -59355
rect -10205 -59433 -10163 -59389
rect -10200 -59533 -10166 -59433
rect -10102 -59516 -10068 -59425
rect -10005 -59443 -9969 -59389
rect -9811 -59425 -9775 -59389
rect -10107 -59567 -10065 -59516
rect -10004 -59533 -9970 -59443
rect -9906 -59511 -9872 -59425
rect -9811 -59443 -9774 -59425
rect -9911 -59567 -9869 -59511
rect -9808 -59533 -9774 -59443
rect -9710 -59512 -9676 -59425
rect -9613 -59441 -9577 -59389
rect -9717 -59567 -9675 -59512
rect -9612 -59533 -9578 -59441
rect -9521 -59448 -9474 -59301
rect -9429 -59245 -9255 -59213
rect -9105 -59245 -9059 -59152
rect -9001 -59168 -8967 -59009
rect -8903 -59152 -8869 -59060
rect -8909 -59245 -8863 -59152
rect -8805 -59168 -8771 -59009
rect -9429 -59283 -8863 -59245
rect -8827 -59207 -8659 -59202
rect -8827 -59219 -8624 -59207
rect -8567 -59219 -8507 -59133
rect -8413 -59152 -8379 -59060
rect -8419 -59213 -8373 -59152
rect -8315 -59168 -8281 -59009
rect -8217 -59152 -8183 -59060
rect -8449 -59219 -8373 -59213
rect -8827 -59245 -8373 -59219
rect -8223 -59245 -8177 -59152
rect -8119 -59168 -8085 -59009
rect -8021 -59152 -7987 -59060
rect -8027 -59245 -7981 -59152
rect -7923 -59168 -7889 -59009
rect -7836 -59202 -7797 -58920
rect -7370 -58960 -7326 -58920
rect -8827 -59261 -7981 -59245
rect -8827 -59265 -8624 -59261
rect -8567 -59265 -8507 -59261
rect -8827 -59276 -8659 -59265
rect -8449 -59283 -7981 -59261
rect -7945 -59276 -7777 -59202
rect -7364 -59259 -7330 -58960
rect -7266 -59234 -7232 -58951
rect -9429 -59307 -9356 -59283
rect -9514 -59522 -9480 -59448
rect -9430 -59475 -9356 -59307
rect -9301 -59291 -8863 -59283
rect -9301 -59356 -9255 -59291
rect -9515 -59567 -9479 -59522
rect -9295 -59548 -9261 -59356
rect -10107 -59601 -9479 -59567
rect -9105 -59356 -9059 -59291
rect -9099 -59548 -9065 -59356
rect -8909 -59544 -8863 -59291
rect -8419 -59291 -7981 -59283
rect -8903 -59548 -8869 -59544
rect -8419 -59356 -8373 -59291
rect -8705 -59526 -8648 -59362
rect -8413 -59548 -8379 -59356
rect -8223 -59356 -8177 -59291
rect -8217 -59548 -8183 -59356
rect -8027 -59544 -7981 -59291
rect -8021 -59548 -7987 -59544
rect -7272 -59364 -7225 -59234
rect -7024 -59244 -6990 -58951
rect -6931 -58967 -6886 -58897
rect -6840 -58871 -6685 -58862
rect -6322 -58871 -6180 -58854
rect -6840 -58905 -6180 -58871
rect -6840 -58917 -6685 -58905
rect -6322 -58918 -6180 -58905
rect -7030 -59364 -6983 -59244
rect -6926 -59259 -6892 -58967
rect -6828 -59245 -6794 -58951
rect -6834 -59364 -6787 -59245
rect -6323 -59364 -6218 -59358
rect -7452 -59446 -6218 -59364
rect -6323 -59453 -6218 -59446
rect -15752 -60397 -15710 -60353
rect -15950 -60431 -15710 -60397
rect -15538 -60363 -15504 -59769
rect -21257 -60521 -20453 -60494
rect -21971 -60686 -21913 -60683
rect -20116 -60686 -20058 -60590
rect -21971 -60727 -20058 -60686
rect -21971 -60820 -21913 -60727
rect -21857 -60765 -21799 -60764
rect -19295 -60765 -19237 -60669
rect -21857 -60806 -19237 -60765
rect -21857 -60901 -21799 -60806
rect -19202 -60842 -19144 -60746
rect -21712 -60883 -19144 -60842
rect -21712 -60979 -21654 -60883
rect -21470 -60964 -20487 -60933
rect -21470 -61029 -20192 -60964
rect -21470 -61048 -20487 -61029
rect -21454 -62133 -21420 -61217
rect -21356 -61425 -21322 -61048
rect -20943 -61119 -20502 -61085
rect -21041 -61589 -21007 -61217
rect -20943 -61525 -20909 -61119
rect -20733 -61122 -20502 -61119
rect -20845 -61589 -20811 -61217
rect -20733 -61228 -20698 -61122
rect -20732 -61525 -20698 -61228
rect -20634 -61525 -20600 -61217
rect -20537 -61226 -20502 -61122
rect -20536 -61525 -20502 -61226
rect -20635 -61588 -20600 -61525
rect -20422 -61588 -20388 -61218
rect -20324 -61526 -20290 -61029
rect -20635 -61589 -20388 -61588
rect -20226 -61589 -20192 -61218
rect -21041 -61623 -20808 -61589
rect -20635 -61623 -20192 -61589
rect -21385 -61677 -21250 -61670
rect -20845 -61677 -20808 -61623
rect -21385 -61714 -20808 -61677
rect -21385 -61724 -21250 -61714
rect -20845 -61852 -20808 -61714
rect -20774 -61679 -20639 -61672
rect -20145 -61679 -20087 -61576
rect -20774 -61713 -20087 -61679
rect -20774 -61726 -20639 -61713
rect -20586 -61757 -20451 -61750
rect -19415 -61757 -19357 -61658
rect -17578 -61203 -17544 -60995
rect -17382 -61203 -17348 -60995
rect -17186 -61203 -17152 -60995
rect -16605 -61210 -16571 -60866
rect -16409 -61210 -16375 -60866
rect -15996 -60973 -15962 -60865
rect -15800 -60973 -15766 -60865
rect -16114 -61020 -16041 -61007
rect -16214 -61048 -16041 -61020
rect -16236 -61061 -16041 -61048
rect -16236 -61210 -16175 -61061
rect -16114 -61067 -16041 -61061
rect -15604 -61037 -15570 -60865
rect -15302 -61037 -15232 -59700
rect -5766 -58293 -5732 -58289
rect -5772 -58546 -5726 -58293
rect -5570 -58481 -5536 -58289
rect -5576 -58546 -5530 -58481
rect -5374 -58481 -5340 -58289
rect -5150 -58375 -5093 -58311
rect -5293 -58424 -5093 -58375
rect -5380 -58546 -5334 -58481
rect -5772 -58554 -5334 -58546
rect -5293 -58554 -5247 -58424
rect -5150 -58475 -5093 -58424
rect -4929 -58293 -4895 -58289
rect -5976 -58591 -5808 -58561
rect -5983 -58635 -5808 -58591
rect -5772 -58592 -5247 -58554
rect -4935 -58546 -4889 -58293
rect -4733 -58481 -4699 -58289
rect -4739 -58546 -4693 -58481
rect -4319 -58270 -3691 -58236
rect -4537 -58481 -4503 -58289
rect -4319 -58315 -4283 -58270
rect -4543 -58546 -4497 -58481
rect -4935 -58554 -4497 -58546
rect -4442 -58530 -4368 -58362
rect -4318 -58389 -4284 -58315
rect -4442 -58554 -4369 -58530
rect -5139 -58572 -4971 -58561
rect -5174 -58573 -4971 -58572
rect -5983 -59007 -5935 -58635
rect -5864 -58828 -5830 -58669
rect -5772 -58685 -5726 -58592
rect -5766 -58777 -5732 -58685
rect -5668 -58828 -5634 -58669
rect -5576 -58685 -5530 -58592
rect -5380 -58624 -5247 -58592
rect -5570 -58777 -5536 -58685
rect -5472 -58828 -5438 -58669
rect -5380 -58685 -5334 -58624
rect -5211 -58635 -4971 -58573
rect -4935 -58592 -4369 -58554
rect -5374 -58777 -5340 -58685
rect -5211 -58779 -5151 -58635
rect -5027 -58828 -4993 -58669
rect -4935 -58685 -4889 -58592
rect -4929 -58777 -4895 -58685
rect -4831 -58828 -4797 -58669
rect -4739 -58685 -4693 -58592
rect -4543 -58624 -4369 -58592
rect -4324 -58536 -4277 -58389
rect -4220 -58396 -4186 -58304
rect -4123 -58325 -4081 -58270
rect -4221 -58448 -4185 -58396
rect -4122 -58412 -4088 -58325
rect -4024 -58394 -3990 -58304
rect -3929 -58326 -3887 -58270
rect -4024 -58412 -3987 -58394
rect -3926 -58412 -3892 -58326
rect -3828 -58394 -3794 -58304
rect -3733 -58321 -3691 -58270
rect -4023 -58448 -3987 -58412
rect -3829 -58448 -3793 -58394
rect -3730 -58412 -3696 -58321
rect -3632 -58404 -3598 -58304
rect -3635 -58448 -3593 -58404
rect -4221 -58482 -3593 -58448
rect -4324 -58610 -4152 -58536
rect -3768 -58589 -3593 -58482
rect -3066 -58293 -3032 -58289
rect -3072 -58546 -3026 -58293
rect -2870 -58481 -2836 -58289
rect -2876 -58546 -2830 -58481
rect -2674 -58481 -2640 -58289
rect -2450 -58363 -2393 -58311
rect -2598 -58425 -2393 -58363
rect -2680 -58546 -2634 -58481
rect -3072 -58554 -2634 -58546
rect -2598 -58554 -2536 -58425
rect -2450 -58475 -2393 -58425
rect -2229 -58293 -2195 -58289
rect -3276 -58568 -3108 -58561
rect -4733 -58777 -4699 -58685
rect -4635 -58828 -4601 -58669
rect -4543 -58685 -4497 -58624
rect -4537 -58777 -4503 -58685
rect -4324 -58745 -4277 -58610
rect -3768 -58649 -3502 -58589
rect -3298 -58628 -3108 -58568
rect -3276 -58635 -3108 -58628
rect -3072 -58592 -2536 -58554
rect -2235 -58546 -2189 -58293
rect -2033 -58481 -1999 -58289
rect -2039 -58546 -1993 -58481
rect -1619 -58270 -991 -58236
rect -1837 -58481 -1803 -58289
rect -1619 -58315 -1583 -58270
rect -1843 -58546 -1797 -58481
rect -2235 -58554 -1797 -58546
rect -1742 -58530 -1668 -58362
rect -1618 -58389 -1584 -58315
rect -1742 -58554 -1669 -58530
rect -4224 -58683 -3593 -58649
rect -4224 -58724 -4183 -58683
rect -4318 -58815 -4284 -58745
rect -5873 -58896 -4502 -58828
rect -4323 -58873 -4279 -58815
rect -4220 -58827 -4186 -58724
rect -4122 -58804 -4088 -58719
rect -4026 -58732 -3985 -58683
rect -4127 -58873 -4083 -58804
rect -4024 -58827 -3990 -58732
rect -3926 -58804 -3892 -58719
rect -3832 -58732 -3791 -58683
rect -3635 -58690 -3593 -58683
rect -3931 -58873 -3887 -58804
rect -3828 -58827 -3794 -58732
rect -3730 -58815 -3696 -58719
rect -3635 -58733 -3594 -58690
rect -3734 -58873 -3690 -58815
rect -3632 -58827 -3598 -58733
rect -3164 -58828 -3130 -58669
rect -3072 -58685 -3026 -58592
rect -3066 -58777 -3032 -58685
rect -2968 -58828 -2934 -58669
rect -2876 -58685 -2830 -58592
rect -2680 -58624 -2536 -58592
rect -2870 -58777 -2836 -58685
rect -2772 -58828 -2738 -58669
rect -2680 -58685 -2634 -58624
rect -2235 -58592 -1669 -58554
rect -2674 -58777 -2640 -58685
rect -2327 -58828 -2293 -58669
rect -2235 -58685 -2189 -58592
rect -2229 -58777 -2195 -58685
rect -2131 -58828 -2097 -58669
rect -2039 -58685 -1993 -58592
rect -1843 -58624 -1669 -58592
rect -1624 -58536 -1577 -58389
rect -1520 -58396 -1486 -58304
rect -1423 -58325 -1381 -58270
rect -1521 -58448 -1485 -58396
rect -1422 -58412 -1388 -58325
rect -1324 -58394 -1290 -58304
rect -1229 -58326 -1187 -58270
rect -1324 -58412 -1287 -58394
rect -1226 -58412 -1192 -58326
rect -1128 -58394 -1094 -58304
rect -1033 -58321 -991 -58270
rect -1323 -58448 -1287 -58412
rect -1129 -58448 -1093 -58394
rect -1030 -58412 -996 -58321
rect -932 -58404 -898 -58304
rect -654 -58364 9205 -58103
rect 14951 -57976 15465 -57813
rect 16711 -57976 16932 -57948
rect 14951 -58106 16932 -57976
rect 14951 -58238 15465 -58106
rect -935 -58448 -893 -58404
rect -1521 -58482 -893 -58448
rect -1624 -58610 -1452 -58536
rect -1068 -58591 -893 -58482
rect -2033 -58777 -1999 -58685
rect -1935 -58828 -1901 -58669
rect -1843 -58685 -1797 -58624
rect -1837 -58777 -1803 -58685
rect -1624 -58745 -1577 -58610
rect -1068 -58649 -818 -58591
rect -1524 -58651 -818 -58649
rect -1524 -58683 -893 -58651
rect -1524 -58724 -1483 -58683
rect -1618 -58815 -1584 -58745
rect -5625 -58936 -5514 -58896
rect -5636 -58944 -5499 -58936
rect -4814 -58944 -4703 -58896
rect -4323 -58907 -3690 -58873
rect -3173 -58830 -2639 -58828
rect -2336 -58830 -1802 -58828
rect -3173 -58896 -1802 -58830
rect -1623 -58873 -1579 -58815
rect -1520 -58827 -1486 -58724
rect -1422 -58804 -1388 -58719
rect -1326 -58732 -1285 -58683
rect -1427 -58873 -1383 -58804
rect -1324 -58827 -1290 -58732
rect -1226 -58804 -1192 -58719
rect -1132 -58732 -1091 -58683
rect -935 -58690 -893 -58683
rect -1231 -58873 -1187 -58804
rect -1128 -58827 -1094 -58732
rect -1030 -58815 -996 -58719
rect -935 -58733 -894 -58690
rect -1034 -58873 -990 -58815
rect -932 -58827 -898 -58733
rect -3016 -58942 -2905 -58896
rect -2833 -58898 -2313 -58896
rect -3039 -58944 -2902 -58942
rect -2138 -58944 -2027 -58896
rect -1623 -58907 -990 -58873
rect -654 -58942 -356 -58364
rect 392 -58629 522 -58364
rect 698 -58629 828 -58364
rect 1015 -58629 1145 -58364
rect 1461 -58629 1591 -58364
rect 379 -58694 1653 -58629
rect -654 -58944 -269 -58942
rect -5653 -58983 -268 -58944
rect -5636 -58996 -5499 -58983
rect -3039 -59002 -2902 -58983
rect -401 -59002 -269 -58983
rect -5984 -59144 -5924 -59007
rect -5247 -59122 -5115 -59114
rect -724 -59122 -592 -59112
rect -5983 -59502 -5935 -59144
rect -5653 -59161 -592 -59122
rect -5247 -59174 -5115 -59161
rect -724 -59172 -592 -59161
rect -5865 -59276 -5331 -59208
rect -4934 -59231 -4301 -59197
rect -5864 -59419 -5830 -59327
rect -5870 -59480 -5824 -59419
rect -5766 -59435 -5732 -59276
rect -5668 -59419 -5634 -59327
rect -5900 -59502 -5824 -59480
rect -5983 -59512 -5824 -59502
rect -5674 -59512 -5628 -59419
rect -5570 -59435 -5536 -59276
rect -5472 -59419 -5438 -59327
rect -5478 -59512 -5432 -59419
rect -5374 -59435 -5340 -59276
rect -5026 -59371 -4992 -59277
rect -4934 -59289 -4890 -59231
rect -5030 -59414 -4989 -59371
rect -4928 -59385 -4894 -59289
rect -4830 -59372 -4796 -59277
rect -4737 -59300 -4693 -59231
rect -5031 -59421 -4989 -59414
rect -4833 -59421 -4792 -59372
rect -4732 -59385 -4698 -59300
rect -4634 -59372 -4600 -59277
rect -4541 -59300 -4497 -59231
rect -4639 -59421 -4598 -59372
rect -4536 -59385 -4502 -59300
rect -4438 -59380 -4404 -59277
rect -4345 -59289 -4301 -59231
rect -4122 -59276 -2631 -59208
rect -2234 -59231 -1601 -59197
rect -4340 -59359 -4306 -59289
rect -4441 -59421 -4400 -59380
rect -5031 -59455 -4400 -59421
rect -5983 -59539 -5432 -59512
rect -5982 -59541 -5432 -59539
rect -5900 -59550 -5432 -59541
rect -5396 -59484 -5228 -59469
rect -5031 -59484 -4856 -59455
rect -5396 -59537 -4856 -59484
rect -4347 -59494 -4300 -59359
rect -4121 -59419 -4087 -59327
rect -4127 -59480 -4081 -59419
rect -4023 -59435 -3989 -59276
rect -3925 -59419 -3891 -59327
rect -5396 -59543 -5228 -59537
rect -5870 -59558 -5432 -59550
rect -5870 -59623 -5824 -59558
rect -5864 -59815 -5830 -59623
rect -5674 -59623 -5628 -59558
rect -5668 -59815 -5634 -59623
rect -5478 -59811 -5432 -59558
rect -5472 -59815 -5438 -59811
rect -5031 -59622 -4856 -59537
rect -4472 -59568 -4300 -59494
rect -5031 -59656 -4403 -59622
rect -5031 -59700 -4989 -59656
rect -5026 -59800 -4992 -59700
rect -4928 -59783 -4894 -59692
rect -4831 -59710 -4795 -59656
rect -4637 -59692 -4601 -59656
rect -4933 -59834 -4891 -59783
rect -4830 -59800 -4796 -59710
rect -4732 -59778 -4698 -59692
rect -4637 -59710 -4600 -59692
rect -4737 -59834 -4695 -59778
rect -4634 -59800 -4600 -59710
rect -4536 -59779 -4502 -59692
rect -4439 -59708 -4403 -59656
rect -4543 -59834 -4501 -59779
rect -4438 -59800 -4404 -59708
rect -4347 -59715 -4300 -59568
rect -4255 -59512 -4081 -59480
rect -3931 -59512 -3885 -59419
rect -3827 -59435 -3793 -59276
rect -3729 -59419 -3695 -59327
rect -3735 -59512 -3689 -59419
rect -3631 -59435 -3597 -59276
rect -4255 -59550 -3689 -59512
rect -3310 -59491 -3250 -59376
rect -3164 -59419 -3130 -59327
rect -3170 -59480 -3124 -59419
rect -3066 -59435 -3032 -59276
rect -2968 -59419 -2934 -59327
rect -3200 -59491 -3124 -59480
rect -3315 -59512 -3124 -59491
rect -2974 -59512 -2928 -59419
rect -2870 -59435 -2836 -59276
rect -2772 -59419 -2738 -59327
rect -2778 -59512 -2732 -59419
rect -2674 -59435 -2640 -59276
rect -2329 -59371 -2283 -59249
rect -2234 -59289 -2190 -59231
rect -2330 -59381 -2283 -59371
rect -2330 -59414 -2289 -59381
rect -2228 -59385 -2194 -59289
rect -2130 -59372 -2096 -59277
rect -2037 -59300 -1993 -59231
rect -2331 -59421 -2289 -59414
rect -2133 -59421 -2092 -59372
rect -2032 -59385 -1998 -59300
rect -1934 -59372 -1900 -59277
rect -1841 -59300 -1797 -59231
rect -1939 -59421 -1898 -59372
rect -1836 -59385 -1802 -59300
rect -1738 -59380 -1704 -59277
rect -1645 -59289 -1601 -59231
rect -1422 -59276 -6 -59208
rect -1640 -59359 -1606 -59289
rect -1741 -59421 -1700 -59380
rect -2331 -59455 -1700 -59421
rect -3315 -59536 -2732 -59512
rect -4255 -59574 -4182 -59550
rect -4340 -59789 -4306 -59715
rect -4256 -59742 -4182 -59574
rect -4127 -59558 -3689 -59550
rect -4127 -59623 -4081 -59558
rect -4341 -59834 -4305 -59789
rect -4121 -59815 -4087 -59623
rect -4933 -59868 -4305 -59834
rect -3931 -59623 -3885 -59558
rect -3925 -59815 -3891 -59623
rect -3735 -59811 -3689 -59558
rect -3729 -59815 -3695 -59811
rect -3531 -59670 -3474 -59629
rect -3315 -59670 -3270 -59536
rect -3200 -59550 -2732 -59536
rect -2696 -59477 -2528 -59469
rect -2331 -59477 -2156 -59455
rect -2696 -59534 -2156 -59477
rect -1647 -59494 -1600 -59359
rect -1421 -59419 -1387 -59327
rect -1427 -59480 -1381 -59419
rect -1323 -59435 -1289 -59276
rect -1225 -59419 -1191 -59327
rect -2696 -59543 -2528 -59534
rect -3170 -59558 -2732 -59550
rect -3170 -59623 -3124 -59558
rect -3531 -59715 -3270 -59670
rect -3531 -59793 -3474 -59715
rect -3164 -59815 -3130 -59623
rect -2974 -59623 -2928 -59558
rect -2968 -59815 -2934 -59623
rect -2778 -59811 -2732 -59558
rect -2772 -59815 -2738 -59811
rect -2331 -59622 -2156 -59534
rect -1772 -59568 -1600 -59494
rect -2331 -59656 -1703 -59622
rect -2331 -59700 -2289 -59656
rect -2326 -59800 -2292 -59700
rect -2228 -59783 -2194 -59692
rect -2131 -59710 -2095 -59656
rect -1937 -59692 -1901 -59656
rect -2233 -59834 -2191 -59783
rect -2130 -59800 -2096 -59710
rect -2032 -59778 -1998 -59692
rect -1937 -59710 -1900 -59692
rect -2037 -59834 -1995 -59778
rect -1934 -59800 -1900 -59710
rect -1836 -59779 -1802 -59692
rect -1739 -59708 -1703 -59656
rect -1843 -59834 -1801 -59779
rect -1738 -59800 -1704 -59708
rect -1647 -59715 -1600 -59568
rect -1555 -59512 -1381 -59480
rect -1231 -59512 -1185 -59419
rect -1127 -59435 -1093 -59276
rect -1029 -59419 -995 -59327
rect -1035 -59512 -989 -59419
rect -931 -59435 -897 -59276
rect -1555 -59550 -989 -59512
rect -953 -59474 -785 -59469
rect -953 -59486 -750 -59474
rect -693 -59486 -633 -59400
rect -539 -59419 -505 -59327
rect -545 -59480 -499 -59419
rect -441 -59435 -407 -59276
rect -343 -59419 -309 -59327
rect -575 -59486 -499 -59480
rect -953 -59512 -499 -59486
rect -349 -59512 -303 -59419
rect -245 -59435 -211 -59276
rect -147 -59419 -113 -59327
rect -153 -59512 -107 -59419
rect -49 -59435 -15 -59276
rect 391 -59335 425 -58882
rect 489 -59090 523 -58694
rect 902 -58784 1343 -58750
rect 804 -59254 838 -58882
rect 902 -59190 936 -58784
rect 1112 -58787 1343 -58784
rect 1000 -59254 1034 -58882
rect 1112 -58893 1147 -58787
rect 1113 -59190 1147 -58893
rect 1211 -59190 1245 -58882
rect 1308 -58891 1343 -58787
rect 1309 -59190 1343 -58891
rect 1210 -59253 1245 -59190
rect 1423 -59253 1457 -58883
rect 1521 -59191 1555 -58694
rect 2385 -58844 2536 -58364
rect 2762 -58826 2886 -58364
rect 3092 -58826 3216 -58364
rect 3499 -58806 3635 -58760
rect 2762 -58844 3277 -58826
rect 1210 -59254 1457 -59253
rect 1619 -59254 1653 -58883
rect 804 -59288 1037 -59254
rect 1210 -59288 1653 -59254
rect 2385 -58887 3277 -58844
rect 2385 -58905 2835 -58887
rect 240 -59388 425 -59335
rect -953 -59528 -107 -59512
rect -953 -59532 -750 -59528
rect -693 -59532 -633 -59528
rect -953 -59543 -785 -59532
rect -575 -59550 -107 -59528
rect -1555 -59574 -1482 -59550
rect -1640 -59789 -1606 -59715
rect -1556 -59742 -1482 -59574
rect -1427 -59558 -989 -59550
rect -1427 -59623 -1381 -59558
rect -1641 -59834 -1605 -59789
rect -1421 -59815 -1387 -59623
rect -2233 -59868 -1605 -59834
rect -1231 -59623 -1185 -59558
rect -1225 -59815 -1191 -59623
rect -1035 -59811 -989 -59558
rect -545 -59558 -107 -59550
rect -1029 -59815 -995 -59811
rect -545 -59623 -499 -59558
rect -831 -59793 -774 -59629
rect -539 -59815 -505 -59623
rect -349 -59623 -303 -59558
rect -343 -59815 -309 -59623
rect -153 -59811 -107 -59558
rect -147 -59815 -113 -59811
rect -6195 -60238 -6059 -60192
rect -16788 -61223 -16653 -61217
rect -16808 -61225 -16653 -61223
rect -17870 -61250 -17740 -61233
rect -17696 -61250 -17623 -61237
rect -18405 -61256 -18347 -61255
rect -17870 -61256 -17623 -61250
rect -18405 -61291 -17623 -61256
rect -17015 -61261 -16653 -61225
rect -16605 -61240 -16175 -61210
rect -16605 -61248 -16186 -61240
rect -15996 -61252 -15962 -61096
rect -15898 -61204 -15864 -61096
rect -15800 -61252 -15766 -61096
rect -15702 -61204 -15668 -61096
rect -15604 -61107 -15232 -61037
rect -16808 -61263 -16653 -61261
rect -16788 -61271 -16653 -61263
rect -18405 -61324 -17740 -61291
rect -17696 -61297 -17623 -61291
rect -18405 -61392 -18347 -61324
rect -17870 -61383 -17740 -61324
rect -17283 -61321 -16734 -61319
rect -16323 -61321 -16249 -61295
rect -17283 -61325 -16249 -61321
rect -17578 -61581 -17544 -61325
rect -17480 -61533 -17446 -61325
rect -17382 -61581 -17348 -61325
rect -17284 -61359 -16249 -61325
rect -16136 -61338 -15351 -61252
rect -17284 -61533 -17250 -61359
rect -16735 -61360 -16249 -61359
rect -16735 -61361 -16664 -61360
rect -16323 -61366 -16249 -61360
rect -17718 -61667 -16780 -61581
rect -20586 -61795 -19357 -61757
rect -20586 -61804 -20451 -61795
rect -20250 -61841 -20115 -61832
rect -18490 -61841 -18432 -61744
rect -16866 -61748 -16780 -61667
rect -16703 -61711 -16669 -61403
rect -16605 -61711 -16571 -61403
rect -16507 -61711 -16473 -61403
rect -16409 -61711 -16375 -61403
rect -16311 -61711 -16277 -61403
rect -16606 -61748 -16571 -61711
rect -15892 -61745 -15831 -61338
rect -16281 -61748 -15831 -61745
rect -16866 -61806 -15831 -61748
rect -6155 -61769 -6121 -60238
rect -3715 -60311 -3579 -60265
rect -3715 -60564 -3675 -60311
rect -3718 -60700 -3672 -60564
rect 391 -59798 425 -59388
rect 460 -59342 595 -59335
rect 1000 -59342 1037 -59288
rect 2385 -59312 2446 -58905
rect 3125 -58939 3160 -58887
rect 2831 -59247 2865 -58939
rect 2929 -59247 2963 -58939
rect 3027 -59247 3061 -58939
rect 3125 -59247 3159 -58939
rect 3223 -59247 3257 -58939
rect 2803 -59290 2877 -59284
rect 3218 -59290 3289 -59289
rect 2803 -59291 3289 -59290
rect 460 -59379 1037 -59342
rect 460 -59389 595 -59379
rect 1000 -59517 1037 -59379
rect 1071 -59344 1206 -59337
rect 1071 -59378 2027 -59344
rect 1071 -59391 1206 -59378
rect 1259 -59422 1394 -59415
rect 1822 -59422 1958 -59415
rect 1259 -59460 1958 -59422
rect 1259 -59469 1394 -59460
rect 1822 -59461 1958 -59460
rect 1000 -59554 1555 -59517
rect 1595 -59551 1787 -59497
rect 1993 -59543 2027 -59378
rect 2075 -59398 2690 -59312
rect 2803 -59329 3470 -59291
rect 2803 -59355 2877 -59329
rect 3288 -59331 3470 -59329
rect 3207 -59385 3342 -59379
rect 3207 -59389 3372 -59385
rect 1129 -59798 1163 -59554
rect 1325 -59798 1359 -59554
rect 1521 -59798 1555 -59554
rect 1741 -59635 1787 -59551
rect 1987 -59613 2158 -59543
rect 2222 -59554 2256 -59446
rect 2320 -59554 2354 -59398
rect 2418 -59554 2452 -59446
rect 2516 -59554 2550 -59398
rect 2740 -59410 3159 -59402
rect 2729 -59440 3159 -59410
rect 3207 -59425 3394 -59389
rect 3207 -59433 3385 -59425
rect 2124 -59785 2158 -59613
rect 2595 -59589 2668 -59583
rect 2729 -59589 2790 -59440
rect 2595 -59602 2790 -59589
rect 2595 -59630 2768 -59602
rect 2595 -59643 2668 -59630
rect 2320 -59785 2354 -59677
rect 2516 -59785 2550 -59677
rect 2929 -59784 2963 -59440
rect 3125 -59784 3159 -59440
rect 3349 -60183 3385 -59433
rect 3230 -60229 3385 -60183
rect 3430 -60267 3470 -59331
rect 3565 -59541 3635 -58806
rect 3990 -58842 4141 -58364
rect 4432 -58824 4583 -58364
rect 4725 -58824 4876 -58364
rect 5365 -58638 5511 -58364
rect 5810 -58638 5956 -58364
rect 6076 -58638 6222 -58364
rect 6436 -58638 6582 -58364
rect 5067 -58694 5203 -58648
rect 4432 -58842 4882 -58824
rect 3990 -58885 4882 -58842
rect 3990 -58903 4440 -58885
rect 3990 -59310 4051 -58903
rect 4730 -58937 4765 -58885
rect 4436 -59245 4470 -58937
rect 4534 -59245 4568 -58937
rect 4632 -59245 4666 -58937
rect 4730 -59245 4764 -58937
rect 4828 -59245 4862 -58937
rect 5137 -59149 5202 -58694
rect 5341 -58703 6615 -58638
rect 5353 -59149 5387 -58891
rect 5451 -59099 5485 -58703
rect 5864 -58793 6305 -58759
rect 5137 -59207 5387 -59149
rect 4408 -59288 4482 -59282
rect 4823 -59288 4894 -59287
rect 4408 -59289 4894 -59288
rect 3680 -59396 4295 -59310
rect 4408 -59327 5098 -59289
rect 4408 -59353 4482 -59327
rect 4893 -59329 5098 -59327
rect 4812 -59385 4947 -59377
rect 4812 -59387 4999 -59385
rect 3565 -59611 3763 -59541
rect 3827 -59552 3861 -59444
rect 3925 -59552 3959 -59396
rect 4023 -59552 4057 -59444
rect 4121 -59552 4155 -59396
rect 4345 -59408 4764 -59400
rect 4334 -59438 4764 -59408
rect 4812 -59425 5019 -59387
rect 4812 -59431 4947 -59425
rect 3729 -59783 3763 -59611
rect 4200 -59587 4273 -59581
rect 4334 -59587 4395 -59438
rect 4200 -59600 4395 -59587
rect 4200 -59628 4373 -59600
rect 4200 -59641 4273 -59628
rect 3925 -59783 3959 -59675
rect 4121 -59783 4155 -59675
rect 4534 -59782 4568 -59438
rect 4730 -59782 4764 -59438
rect 3334 -60313 3470 -60267
rect 4983 -60752 5019 -59425
rect 3498 -60788 5019 -60752
rect 3498 -60900 3534 -60788
rect 5058 -60822 5098 -59329
rect 5353 -59807 5387 -59207
rect 5766 -59263 5800 -58891
rect 5864 -59199 5898 -58793
rect 6074 -58796 6305 -58793
rect 5962 -59263 5996 -58891
rect 6074 -58902 6109 -58796
rect 6075 -59199 6109 -58902
rect 6173 -59199 6207 -58891
rect 6270 -58900 6305 -58796
rect 6271 -59199 6305 -58900
rect 6172 -59262 6207 -59199
rect 6385 -59262 6419 -58892
rect 6483 -59200 6517 -58703
rect 7000 -58818 7197 -58364
rect 7533 -58818 7730 -58364
rect 8046 -58809 8243 -58364
rect 8549 -58809 8746 -58364
rect 8944 -58791 9205 -58364
rect 10489 -58301 10553 -58278
rect 15854 -58301 15937 -58106
rect 16711 -58128 16932 -58106
rect 10489 -58384 15937 -58301
rect 10489 -58396 10553 -58384
rect 19794 -58462 19943 -55927
rect 20355 -56457 20539 -55927
rect 20979 -55961 21021 -55917
rect 21082 -55925 21116 -55834
rect 21180 -55907 21214 -55817
rect 21273 -55839 21315 -55783
rect 21179 -55961 21215 -55907
rect 21278 -55925 21312 -55839
rect 21376 -55907 21410 -55817
rect 21467 -55838 21509 -55783
rect 21373 -55925 21410 -55907
rect 21474 -55925 21508 -55838
rect 21572 -55909 21606 -55817
rect 21669 -55828 21705 -55783
rect 21670 -55902 21704 -55828
rect 21373 -55961 21409 -55925
rect 21571 -55961 21607 -55909
rect 20979 -55995 21607 -55961
rect 20979 -56104 21154 -55995
rect 21663 -56049 21710 -55902
rect 21754 -56043 21828 -55875
rect 21889 -55994 21923 -55802
rect 20904 -56162 21154 -56104
rect 21538 -56123 21710 -56049
rect 20904 -56164 21610 -56162
rect 20979 -56196 21610 -56164
rect 20979 -56203 21021 -56196
rect 20980 -56246 21021 -56203
rect 20984 -56340 21018 -56246
rect 21082 -56328 21116 -56232
rect 21177 -56245 21218 -56196
rect 21076 -56386 21120 -56328
rect 21180 -56340 21214 -56245
rect 21278 -56317 21312 -56232
rect 21371 -56245 21412 -56196
rect 21273 -56386 21317 -56317
rect 21376 -56340 21410 -56245
rect 21474 -56317 21508 -56232
rect 21569 -56237 21610 -56196
rect 21469 -56386 21513 -56317
rect 21572 -56340 21606 -56237
rect 21663 -56258 21710 -56123
rect 21755 -56067 21828 -56043
rect 21883 -56059 21929 -55994
rect 22085 -55994 22119 -55802
rect 22079 -56059 22125 -55994
rect 22281 -55806 22315 -55802
rect 22275 -56059 22321 -55806
rect 22479 -55876 22536 -55824
rect 22479 -55938 22684 -55876
rect 22479 -55988 22536 -55938
rect 21883 -56067 22321 -56059
rect 21755 -56105 22321 -56067
rect 22622 -56067 22684 -55938
rect 22726 -55994 22760 -55802
rect 22720 -56059 22766 -55994
rect 22922 -55994 22956 -55802
rect 22916 -56059 22962 -55994
rect 23118 -55806 23152 -55802
rect 23112 -56059 23158 -55806
rect 23777 -55783 24405 -55749
rect 23684 -55917 23718 -55817
rect 23777 -55834 23819 -55783
rect 23679 -55961 23721 -55917
rect 23782 -55925 23816 -55834
rect 23880 -55907 23914 -55817
rect 23973 -55839 24015 -55783
rect 23879 -55961 23915 -55907
rect 23978 -55925 24012 -55839
rect 24076 -55907 24110 -55817
rect 24167 -55838 24209 -55783
rect 24073 -55925 24110 -55907
rect 24174 -55925 24208 -55838
rect 24272 -55909 24306 -55817
rect 24369 -55828 24405 -55783
rect 24370 -55902 24404 -55828
rect 24073 -55961 24109 -55925
rect 24271 -55961 24307 -55909
rect 23679 -55995 24307 -55961
rect 22720 -56067 23158 -56059
rect 21755 -56137 21929 -56105
rect 21883 -56198 21929 -56137
rect 21670 -56328 21704 -56258
rect 21889 -56290 21923 -56198
rect 21665 -56386 21709 -56328
rect 21987 -56341 22021 -56182
rect 22079 -56198 22125 -56105
rect 22085 -56290 22119 -56198
rect 22183 -56341 22217 -56182
rect 22275 -56198 22321 -56105
rect 22622 -56105 23158 -56067
rect 22622 -56137 22766 -56105
rect 22281 -56290 22315 -56198
rect 22379 -56341 22413 -56182
rect 22720 -56198 22766 -56137
rect 22726 -56290 22760 -56198
rect 22824 -56341 22858 -56182
rect 22916 -56198 22962 -56105
rect 22922 -56290 22956 -56198
rect 23020 -56341 23054 -56182
rect 23112 -56198 23158 -56105
rect 23194 -56081 23362 -56074
rect 23194 -56141 23384 -56081
rect 23679 -56102 23854 -55995
rect 24363 -56049 24410 -55902
rect 24454 -56043 24528 -55875
rect 24589 -55994 24623 -55802
rect 23194 -56148 23362 -56141
rect 23588 -56162 23854 -56102
rect 24238 -56123 24410 -56049
rect 23118 -56290 23152 -56198
rect 23216 -56341 23250 -56182
rect 23679 -56196 24310 -56162
rect 23679 -56203 23721 -56196
rect 23680 -56246 23721 -56203
rect 23684 -56340 23718 -56246
rect 23782 -56328 23816 -56232
rect 23877 -56245 23918 -56196
rect 21076 -56420 21709 -56386
rect 21888 -56343 22422 -56341
rect 22725 -56343 23259 -56341
rect 21888 -56409 23259 -56343
rect 23776 -56386 23820 -56328
rect 23880 -56340 23914 -56245
rect 23978 -56317 24012 -56232
rect 24071 -56245 24112 -56196
rect 23973 -56386 24017 -56317
rect 24076 -56340 24110 -56245
rect 24174 -56317 24208 -56232
rect 24269 -56237 24310 -56196
rect 24169 -56386 24213 -56317
rect 24272 -56340 24306 -56237
rect 24363 -56258 24410 -56123
rect 24455 -56067 24528 -56043
rect 24583 -56059 24629 -55994
rect 24785 -55994 24819 -55802
rect 24779 -56059 24825 -55994
rect 24981 -55806 25015 -55802
rect 24975 -56059 25021 -55806
rect 25179 -55888 25236 -55824
rect 25179 -55937 25379 -55888
rect 25179 -55988 25236 -55937
rect 24583 -56067 25021 -56059
rect 24455 -56105 25021 -56067
rect 25333 -56067 25379 -55937
rect 25426 -55994 25460 -55802
rect 25420 -56059 25466 -55994
rect 25622 -55994 25656 -55802
rect 25616 -56059 25662 -55994
rect 25818 -55806 25852 -55802
rect 25812 -56059 25858 -55806
rect 29430 -55786 29464 -55442
rect 29626 -55786 29660 -55442
rect 29799 -55591 29860 -55442
rect 30039 -55556 30073 -55400
rect 30137 -55556 30171 -55448
rect 30235 -55556 30269 -55400
rect 36605 -55413 36852 -55372
rect 37687 -55400 37822 -55392
rect 37667 -55402 37822 -55400
rect 36605 -55430 36735 -55413
rect 36779 -55426 36852 -55413
rect 37460 -55438 37822 -55402
rect 38339 -55411 39124 -55325
rect 45468 -55411 45598 -55319
rect 45760 -55377 45794 -55121
rect 45858 -55377 45892 -55169
rect 45956 -55377 45990 -55121
rect 46054 -55343 46088 -55169
rect 46635 -55299 46669 -54991
rect 46733 -55299 46767 -54991
rect 46831 -55299 46865 -54991
rect 46929 -55299 46963 -54991
rect 47027 -55299 47061 -54991
rect 46603 -55342 46674 -55341
rect 47015 -55342 47089 -55336
rect 46603 -55343 47089 -55342
rect 46054 -55377 47089 -55343
rect 47446 -55364 47507 -54957
rect 52201 -54925 52427 -54916
rect 53854 -54925 54100 -54845
rect 52201 -55058 54100 -54925
rect 55670 -54862 56335 -54834
rect 55670 -54920 56705 -54862
rect 55670 -55001 55756 -54920
rect 55930 -54957 55965 -54920
rect 56255 -54923 56705 -54920
rect 52201 -55150 52427 -55058
rect 53854 -55065 54100 -55058
rect 54818 -55087 55756 -55001
rect 46055 -55381 47089 -55377
rect 46055 -55383 46604 -55381
rect 45642 -55411 45715 -55405
rect 47015 -55407 47089 -55381
rect 37667 -55440 37822 -55438
rect 37687 -55446 37822 -55440
rect 37870 -55423 38289 -55415
rect 30333 -55556 30367 -55448
rect 37870 -55453 38300 -55423
rect 29921 -55591 29994 -55585
rect 29799 -55604 29994 -55591
rect 29821 -55632 29994 -55604
rect 29921 -55645 29994 -55632
rect 30431 -55615 30803 -55545
rect 30039 -55787 30073 -55679
rect 30235 -55787 30269 -55679
rect 30431 -55787 30465 -55615
rect 25420 -56067 25858 -56059
rect 24455 -56137 24629 -56105
rect 24583 -56198 24629 -56137
rect 24370 -56328 24404 -56258
rect 24589 -56290 24623 -56198
rect 24365 -56386 24409 -56328
rect 24687 -56341 24721 -56182
rect 24779 -56198 24825 -56105
rect 24785 -56290 24819 -56198
rect 24883 -56341 24917 -56182
rect 24975 -56198 25021 -56105
rect 25057 -56085 25225 -56074
rect 25057 -56086 25260 -56085
rect 25057 -56148 25297 -56086
rect 25333 -56105 25858 -56067
rect 25333 -56137 25466 -56105
rect 24981 -56290 25015 -56198
rect 25079 -56341 25113 -56182
rect 25237 -56292 25297 -56148
rect 25420 -56198 25466 -56137
rect 25426 -56290 25460 -56198
rect 25524 -56341 25558 -56182
rect 25616 -56198 25662 -56105
rect 25622 -56290 25656 -56198
rect 25720 -56341 25754 -56182
rect 25812 -56198 25858 -56105
rect 25894 -56104 26062 -56074
rect 25894 -56148 26069 -56104
rect 25818 -56290 25852 -56198
rect 25916 -56341 25950 -56182
rect 22113 -56457 22224 -56409
rect 22399 -56411 22919 -56409
rect 22991 -56455 23102 -56409
rect 23776 -56420 24409 -56386
rect 24588 -56409 25959 -56341
rect 22988 -56457 23125 -56455
rect 24789 -56457 24900 -56409
rect 25600 -56449 25711 -56409
rect 25585 -56457 25722 -56449
rect 20354 -56496 25739 -56457
rect 20355 -56515 20487 -56496
rect 22988 -56515 23125 -56496
rect 25585 -56509 25722 -56496
rect 26021 -56520 26069 -56148
rect 20678 -56635 20810 -56625
rect 25201 -56635 25333 -56627
rect 20678 -56674 25739 -56635
rect 26010 -56657 26070 -56520
rect 20678 -56685 20810 -56674
rect 25201 -56687 25333 -56674
rect 20092 -56789 21508 -56721
rect 21687 -56744 22320 -56710
rect 20101 -56948 20135 -56789
rect 20199 -56932 20233 -56840
rect 20193 -57025 20239 -56932
rect 20297 -56948 20331 -56789
rect 20395 -56932 20429 -56840
rect 20389 -57025 20435 -56932
rect 20493 -56948 20527 -56789
rect 20591 -56932 20625 -56840
rect 20585 -56993 20631 -56932
rect 20585 -56999 20661 -56993
rect 20719 -56999 20779 -56913
rect 20983 -56948 21017 -56789
rect 21081 -56932 21115 -56840
rect 20871 -56987 21039 -56982
rect 20836 -56999 21039 -56987
rect 20585 -57025 21039 -56999
rect 20193 -57041 21039 -57025
rect 20193 -57063 20661 -57041
rect 20719 -57045 20779 -57041
rect 20836 -57045 21039 -57041
rect 20871 -57056 21039 -57045
rect 21075 -57025 21121 -56932
rect 21179 -56948 21213 -56789
rect 21277 -56932 21311 -56840
rect 21271 -57025 21317 -56932
rect 21375 -56948 21409 -56789
rect 21687 -56802 21731 -56744
rect 21473 -56932 21507 -56840
rect 21692 -56872 21726 -56802
rect 21467 -56993 21513 -56932
rect 21467 -57025 21641 -56993
rect 21075 -57063 21641 -57025
rect 20193 -57071 20631 -57063
rect 20193 -57324 20239 -57071
rect 20199 -57328 20233 -57324
rect 20389 -57136 20435 -57071
rect 20395 -57328 20429 -57136
rect 20585 -57136 20631 -57071
rect 21075 -57071 21513 -57063
rect 20591 -57328 20625 -57136
rect 20860 -57306 20917 -57142
rect 21075 -57324 21121 -57071
rect 21081 -57328 21115 -57324
rect 21271 -57136 21317 -57071
rect 21277 -57328 21311 -57136
rect 21467 -57136 21513 -57071
rect 21568 -57087 21641 -57063
rect 21686 -57007 21733 -56872
rect 21790 -56893 21824 -56790
rect 21883 -56813 21927 -56744
rect 21786 -56934 21827 -56893
rect 21888 -56898 21922 -56813
rect 21986 -56885 22020 -56790
rect 22079 -56813 22123 -56744
rect 21984 -56934 22025 -56885
rect 22084 -56898 22118 -56813
rect 22182 -56885 22216 -56790
rect 22276 -56802 22320 -56744
rect 22178 -56934 22219 -56885
rect 22280 -56898 22314 -56802
rect 22369 -56884 22415 -56762
rect 22717 -56789 24208 -56721
rect 24387 -56744 25020 -56710
rect 22369 -56894 22416 -56884
rect 22375 -56927 22416 -56894
rect 22375 -56934 22417 -56927
rect 21786 -56968 22417 -56934
rect 22726 -56948 22760 -56789
rect 22824 -56932 22858 -56840
rect 22242 -56990 22417 -56968
rect 22614 -56990 22782 -56982
rect 21686 -57081 21858 -57007
rect 22242 -57047 22782 -56990
rect 21473 -57328 21507 -57136
rect 21568 -57255 21642 -57087
rect 21686 -57228 21733 -57081
rect 22242 -57135 22417 -57047
rect 22614 -57056 22782 -57047
rect 22818 -57025 22864 -56932
rect 22922 -56948 22956 -56789
rect 23020 -56932 23054 -56840
rect 23014 -57025 23060 -56932
rect 23118 -56948 23152 -56789
rect 23216 -56932 23250 -56840
rect 23210 -56993 23256 -56932
rect 23210 -57004 23286 -56993
rect 23336 -57004 23396 -56889
rect 23683 -56948 23717 -56789
rect 23781 -56932 23815 -56840
rect 23210 -57025 23401 -57004
rect 22818 -57049 23401 -57025
rect 22818 -57063 23286 -57049
rect 22818 -57071 23256 -57063
rect 21789 -57169 22417 -57135
rect 21789 -57221 21825 -57169
rect 21987 -57205 22023 -57169
rect 21692 -57302 21726 -57228
rect 21691 -57347 21727 -57302
rect 21790 -57313 21824 -57221
rect 21888 -57292 21922 -57205
rect 21986 -57223 22023 -57205
rect 21887 -57347 21929 -57292
rect 21986 -57313 22020 -57223
rect 22084 -57291 22118 -57205
rect 22181 -57223 22217 -57169
rect 22081 -57347 22123 -57291
rect 22182 -57313 22216 -57223
rect 22280 -57296 22314 -57205
rect 22375 -57213 22417 -57169
rect 22277 -57347 22319 -57296
rect 22378 -57313 22412 -57213
rect 21691 -57381 22319 -57347
rect 22818 -57324 22864 -57071
rect 22824 -57328 22858 -57324
rect 23014 -57136 23060 -57071
rect 23020 -57328 23054 -57136
rect 23210 -57136 23256 -57071
rect 23216 -57328 23250 -57136
rect 23356 -57183 23401 -57049
rect 23775 -57025 23821 -56932
rect 23879 -56948 23913 -56789
rect 23977 -56932 24011 -56840
rect 23971 -57025 24017 -56932
rect 24075 -56948 24109 -56789
rect 24387 -56802 24431 -56744
rect 24173 -56932 24207 -56840
rect 24392 -56872 24426 -56802
rect 24167 -56993 24213 -56932
rect 24167 -57025 24341 -56993
rect 23775 -57063 24341 -57025
rect 23775 -57071 24213 -57063
rect 23560 -57183 23617 -57142
rect 23356 -57228 23617 -57183
rect 23560 -57306 23617 -57228
rect 23775 -57324 23821 -57071
rect 23781 -57328 23815 -57324
rect 23971 -57136 24017 -57071
rect 23977 -57328 24011 -57136
rect 24167 -57136 24213 -57071
rect 24268 -57087 24341 -57063
rect 24386 -57007 24433 -56872
rect 24490 -56893 24524 -56790
rect 24583 -56813 24627 -56744
rect 24486 -56934 24527 -56893
rect 24588 -56898 24622 -56813
rect 24686 -56885 24720 -56790
rect 24779 -56813 24823 -56744
rect 24684 -56934 24725 -56885
rect 24784 -56898 24818 -56813
rect 24882 -56885 24916 -56790
rect 24976 -56802 25020 -56744
rect 25417 -56789 25951 -56721
rect 24878 -56934 24919 -56885
rect 24980 -56898 25014 -56802
rect 25078 -56884 25112 -56790
rect 25075 -56927 25116 -56884
rect 25075 -56934 25117 -56927
rect 24486 -56968 25117 -56934
rect 25426 -56948 25460 -56789
rect 25524 -56932 25558 -56840
rect 24942 -56997 25117 -56968
rect 25314 -56997 25482 -56982
rect 24386 -57081 24558 -57007
rect 24942 -57050 25482 -56997
rect 24173 -57328 24207 -57136
rect 24268 -57255 24342 -57087
rect 24386 -57228 24433 -57081
rect 24942 -57135 25117 -57050
rect 25314 -57056 25482 -57050
rect 25518 -57025 25564 -56932
rect 25622 -56948 25656 -56789
rect 25720 -56932 25754 -56840
rect 25714 -57025 25760 -56932
rect 25818 -56948 25852 -56789
rect 25916 -56932 25950 -56840
rect 25910 -56993 25956 -56932
rect 25910 -57015 25986 -56993
rect 26021 -57015 26069 -56657
rect 25910 -57025 26069 -57015
rect 25518 -57052 26069 -57025
rect 25518 -57054 26068 -57052
rect 25518 -57063 25986 -57054
rect 25518 -57071 25956 -57063
rect 24489 -57169 25117 -57135
rect 24489 -57221 24525 -57169
rect 24687 -57205 24723 -57169
rect 24392 -57302 24426 -57228
rect 24391 -57347 24427 -57302
rect 24490 -57313 24524 -57221
rect 24588 -57292 24622 -57205
rect 24686 -57223 24723 -57205
rect 24587 -57347 24629 -57292
rect 24686 -57313 24720 -57223
rect 24784 -57291 24818 -57205
rect 24881 -57223 24917 -57169
rect 24781 -57347 24823 -57291
rect 24882 -57313 24916 -57223
rect 24980 -57296 25014 -57205
rect 25075 -57213 25117 -57169
rect 24977 -57347 25019 -57296
rect 25078 -57313 25112 -57213
rect 24391 -57381 25019 -57347
rect 25518 -57324 25564 -57071
rect 25524 -57328 25558 -57324
rect 25714 -57136 25760 -57071
rect 25720 -57328 25754 -57136
rect 25910 -57136 25956 -57071
rect 25916 -57328 25950 -57136
rect 28431 -56722 28465 -56378
rect 28627 -56722 28661 -56378
rect 29040 -56485 29074 -56377
rect 29236 -56485 29270 -56377
rect 28922 -56532 28995 -56519
rect 28822 -56560 28995 -56532
rect 28800 -56573 28995 -56560
rect 28800 -56722 28861 -56573
rect 28922 -56579 28995 -56573
rect 29432 -56549 29466 -56377
rect 28431 -56752 28861 -56722
rect 28431 -56760 28850 -56752
rect 29040 -56764 29074 -56608
rect 29138 -56716 29172 -56608
rect 29236 -56764 29270 -56608
rect 29334 -56716 29368 -56608
rect 29432 -56619 29710 -56549
rect 28075 -56833 28302 -56831
rect 28713 -56833 28787 -56807
rect 28075 -56871 28787 -56833
rect 28900 -56850 29515 -56764
rect 22124 -57682 22284 -57550
rect 22131 -57865 22266 -57682
rect 22121 -57997 22281 -57865
rect 22644 -58316 22678 -57872
rect 22840 -58316 22874 -57872
rect 23082 -57804 26006 -57707
rect 22644 -58317 22874 -58316
rect 22018 -58330 22150 -58320
rect 22461 -58329 22596 -58323
rect 22441 -58330 22596 -58329
rect 22018 -58366 22596 -58330
rect 22644 -58354 22888 -58317
rect 22018 -58380 22150 -58366
rect 22441 -58369 22596 -58366
rect 22461 -58377 22596 -58369
rect 22854 -58389 22888 -58354
rect 22984 -58389 23044 -58329
rect 20589 -58462 22185 -58419
rect 18740 -58484 22185 -58462
rect 22371 -58422 22530 -58421
rect 22371 -58427 22531 -58422
rect 22679 -58427 22814 -58421
rect 22371 -58466 22814 -58427
rect 22371 -58467 22585 -58466
rect 22371 -58480 22531 -58467
rect 22679 -58475 22814 -58466
rect 22854 -58450 23044 -58389
rect 22371 -58481 22530 -58480
rect 18740 -58551 20769 -58484
rect 10168 -58605 10227 -58598
rect 10168 -58688 14144 -58605
rect 10168 -58693 10227 -58688
rect 8046 -58818 8795 -58809
rect 6962 -58871 8795 -58818
rect 6172 -59263 6419 -59262
rect 6581 -59263 6615 -58892
rect 6962 -58994 7001 -58871
rect 8163 -58905 8795 -58871
rect 7064 -58945 8072 -58909
rect 6966 -59183 7000 -58994
rect 5766 -59297 5999 -59263
rect 6172 -59297 6615 -59263
rect 6964 -59266 7001 -59183
rect 7064 -59190 7098 -58945
rect 7380 -59184 7414 -58982
rect 7478 -59181 7512 -58982
rect 7742 -59181 7776 -58982
rect 7377 -59205 7414 -59184
rect 7258 -59242 7414 -59205
rect 7476 -59220 7776 -59181
rect 7258 -59266 7295 -59242
rect 5422 -59351 5557 -59344
rect 5962 -59351 5999 -59297
rect 6964 -59303 7295 -59266
rect 7840 -59273 7874 -58982
rect 8036 -58999 8072 -58945
rect 8036 -59190 8070 -58999
rect 8134 -59273 8168 -58982
rect 8346 -59173 8380 -58982
rect 8439 -58989 8482 -58905
rect 8341 -59218 8384 -59173
rect 8444 -59190 8478 -58989
rect 8655 -59171 8689 -58982
rect 8748 -58991 8791 -58905
rect 8245 -59264 8384 -59218
rect 7607 -59307 8168 -59273
rect 5422 -59388 5999 -59351
rect 5422 -59398 5557 -59388
rect 5962 -59526 5999 -59388
rect 6033 -59353 6168 -59346
rect 6033 -59387 6852 -59353
rect 7607 -59369 7641 -59307
rect 6033 -59400 6168 -59387
rect 6221 -59431 6356 -59424
rect 6221 -59469 6782 -59431
rect 6221 -59478 6356 -59469
rect 6556 -59515 6692 -59506
rect 5962 -59563 6517 -59526
rect 6556 -59552 6711 -59515
rect 6557 -59560 6692 -59552
rect 6091 -59807 6125 -59563
rect 6287 -59807 6321 -59563
rect 6483 -59807 6517 -59563
rect -918 -60936 3534 -60900
rect 3596 -60856 5098 -60822
rect 6748 -60838 6782 -59469
rect -918 -60984 -869 -60936
rect 1492 -60980 1628 -60971
rect 3596 -60980 3630 -60856
rect 6442 -60872 6782 -60838
rect 3675 -60911 3811 -60908
rect 6442 -60911 6476 -60872
rect 3675 -60945 6476 -60911
rect 6580 -60930 6716 -60924
rect 6818 -60930 6852 -59387
rect 6965 -59438 7104 -59384
rect 7495 -59403 7641 -59369
rect 7495 -59518 7529 -59403
rect 7714 -59408 7853 -59354
rect 6915 -59552 7529 -59518
rect 7590 -59479 8070 -59445
rect 6966 -59900 7000 -59588
rect 7064 -59796 7098 -59552
rect 7162 -59900 7196 -59588
rect 7282 -59831 7316 -59588
rect 7380 -59796 7414 -59552
rect 7478 -59831 7512 -59588
rect 7590 -59831 7624 -59479
rect 7282 -59865 7624 -59831
rect 7660 -59553 7874 -59519
rect 7660 -59900 7694 -59553
rect 7840 -59796 7874 -59553
rect 6966 -59934 7694 -59900
rect 8036 -59796 8070 -59479
rect 8123 -59482 8262 -59428
rect 8341 -59603 8384 -59264
rect 8651 -59362 8694 -59171
rect 8753 -59190 8787 -58991
rect 8944 -59052 10099 -58791
rect 13481 -58877 13766 -58819
rect 14061 -58877 14144 -58688
rect 18869 -58703 18913 -58551
rect 18873 -58862 18907 -58703
rect 18971 -58853 19005 -58654
rect 19063 -58702 19107 -58551
rect 13481 -58905 18441 -58877
rect 18779 -58905 18925 -58897
rect 13481 -58941 18925 -58905
rect 18966 -58902 19011 -58853
rect 19069 -58862 19103 -58702
rect 19815 -58703 19859 -58551
rect 19819 -58862 19853 -58703
rect 19917 -58853 19951 -58654
rect 20009 -58702 20053 -58551
rect 18966 -58903 19360 -58902
rect 18966 -58938 19409 -58903
rect 19725 -58905 19871 -58897
rect 13481 -58971 18441 -58941
rect 18779 -58957 18925 -58941
rect 19221 -58947 19409 -58938
rect 19666 -58941 19871 -58905
rect 19912 -58902 19957 -58853
rect 20015 -58862 20049 -58702
rect 19912 -58938 20582 -58902
rect 19277 -58963 19409 -58947
rect 19725 -58957 19871 -58941
rect 20167 -58947 20582 -58938
rect 13481 -59038 13766 -58971
rect 19002 -58994 19145 -58977
rect 18544 -59030 19145 -58994
rect 8551 -59408 8694 -59362
rect 8346 -59796 8380 -59603
rect 8651 -59605 8694 -59408
rect 8738 -59476 8877 -59422
rect 8655 -59796 8689 -59605
rect 3675 -60954 3811 -60945
rect 6580 -60964 6852 -60930
rect 6580 -60970 6716 -60964
rect -1005 -61030 -869 -60984
rect 1459 -61014 3630 -60980
rect 1492 -61017 1628 -61014
rect 8944 -61047 9205 -59052
rect -4847 -61069 -4215 -61060
rect -2347 -61069 -1715 -61060
rect 153 -61069 785 -61060
rect 2653 -61069 3285 -61060
rect 5153 -61069 5785 -61060
rect 8137 -61069 9205 -61047
rect -6048 -61070 -4215 -61069
rect -3548 -61070 9205 -61069
rect -6048 -61122 9205 -61070
rect -6048 -61245 -6009 -61122
rect -4847 -61156 -3509 -61122
rect -2347 -61156 -1715 -61122
rect -5946 -61196 -4938 -61160
rect -6044 -61434 -6010 -61245
rect -6046 -61517 -6009 -61434
rect -5946 -61441 -5912 -61196
rect -5630 -61435 -5596 -61233
rect -5532 -61432 -5498 -61233
rect -5268 -61432 -5234 -61233
rect -5633 -61456 -5596 -61435
rect -5752 -61493 -5596 -61456
rect -5534 -61471 -5234 -61432
rect -5752 -61517 -5715 -61493
rect -6046 -61554 -5715 -61517
rect -5170 -61524 -5136 -61233
rect -4974 -61250 -4938 -61196
rect -4974 -61441 -4940 -61250
rect -4876 -61524 -4842 -61233
rect -4664 -61424 -4630 -61233
rect -4571 -61240 -4528 -61156
rect -4336 -61157 -3509 -61156
rect -4669 -61469 -4626 -61424
rect -4566 -61441 -4532 -61240
rect -4355 -61422 -4321 -61233
rect -4262 -61242 -4219 -61157
rect -4765 -61515 -4626 -61469
rect -5403 -61558 -4842 -61524
rect -5403 -61620 -5369 -61558
rect -6045 -61689 -5906 -61635
rect -5515 -61654 -5369 -61620
rect -5515 -61769 -5481 -61654
rect -5296 -61659 -5157 -61605
rect -6155 -61803 -5481 -61769
rect -5420 -61730 -4940 -61696
rect -16866 -61834 -16201 -61806
rect -20845 -61889 -20290 -61852
rect -20250 -61876 -18432 -61841
rect -20250 -61878 -20096 -61876
rect -20250 -61886 -20115 -61878
rect -18490 -61881 -18432 -61876
rect -20716 -62133 -20682 -61889
rect -20520 -62133 -20486 -61889
rect -20324 -62133 -20290 -61889
rect -7745 -61997 -7545 -61973
rect -18126 -62133 -7545 -61997
rect -7745 -62144 -7545 -62133
rect -6044 -62151 -6010 -61839
rect -5946 -62047 -5912 -61803
rect -5848 -62151 -5814 -61839
rect -5728 -62082 -5694 -61839
rect -5630 -62047 -5596 -61803
rect -5532 -62082 -5498 -61839
rect -5420 -62082 -5386 -61730
rect -5728 -62116 -5386 -62082
rect -5350 -61804 -5136 -61770
rect -5350 -62151 -5316 -61804
rect -6044 -62185 -5316 -62151
rect -5170 -62047 -5136 -61804
rect -4974 -62047 -4940 -61730
rect -4887 -61733 -4748 -61679
rect -4669 -61854 -4626 -61515
rect -4359 -61613 -4316 -61422
rect -4257 -61441 -4223 -61242
rect -3548 -61245 -3509 -61157
rect -3446 -61196 -2438 -61160
rect -3718 -61406 -3672 -61270
rect -4459 -61659 -4316 -61613
rect -4664 -62047 -4630 -61854
rect -4359 -61856 -4316 -61659
rect -4272 -61727 -4133 -61673
rect -4355 -62047 -4321 -61856
rect -23449 -62311 -22910 -62272
rect -6608 -62251 -6445 -62231
rect -28147 -62448 -22910 -62311
rect -18303 -62387 -6445 -62251
rect -3712 -61769 -3678 -61406
rect -3544 -61434 -3510 -61245
rect -3546 -61517 -3509 -61434
rect -3446 -61441 -3412 -61196
rect -3130 -61435 -3096 -61233
rect -3032 -61432 -2998 -61233
rect -2768 -61432 -2734 -61233
rect -3133 -61456 -3096 -61435
rect -3252 -61493 -3096 -61456
rect -3034 -61471 -2734 -61432
rect -3252 -61517 -3215 -61493
rect -3546 -61554 -3215 -61517
rect -2670 -61524 -2636 -61233
rect -2474 -61250 -2438 -61196
rect -2474 -61441 -2440 -61250
rect -2376 -61524 -2342 -61233
rect -2164 -61424 -2130 -61233
rect -2071 -61240 -2028 -61156
rect -2169 -61469 -2126 -61424
rect -2066 -61441 -2032 -61240
rect -1855 -61422 -1821 -61233
rect -1762 -61242 -1719 -61156
rect -2265 -61515 -2126 -61469
rect -3163 -61585 -3024 -61531
rect -2903 -61558 -2342 -61524
rect -2903 -61620 -2869 -61558
rect -3545 -61689 -3406 -61635
rect -3015 -61654 -2869 -61620
rect -3015 -61769 -2981 -61654
rect -2796 -61659 -2657 -61605
rect -3712 -61803 -2981 -61769
rect -2920 -61730 -2440 -61696
rect -3544 -62151 -3510 -61839
rect -3446 -62047 -3412 -61803
rect -3348 -62151 -3314 -61839
rect -3228 -62082 -3194 -61839
rect -3130 -62047 -3096 -61803
rect -3032 -62082 -2998 -61839
rect -2920 -62082 -2886 -61730
rect -3228 -62116 -2886 -62082
rect -2850 -61804 -2636 -61770
rect -2850 -62151 -2816 -61804
rect -3544 -62185 -2816 -62151
rect -2670 -62047 -2636 -61804
rect -2474 -62047 -2440 -61730
rect -2387 -61733 -2248 -61679
rect -2169 -61854 -2126 -61515
rect -2085 -61579 -1946 -61525
rect -1859 -61613 -1816 -61422
rect -1757 -61441 -1723 -61242
rect -1048 -61245 -1009 -61122
rect 153 -61156 785 -61122
rect -946 -61196 62 -61160
rect -1959 -61659 -1816 -61613
rect -2164 -62047 -2130 -61854
rect -1859 -61856 -1816 -61659
rect -1772 -61727 -1633 -61673
rect -1855 -62047 -1821 -61856
rect -1170 -61402 -1124 -61266
rect -1164 -61769 -1130 -61402
rect -1044 -61434 -1010 -61245
rect -1046 -61517 -1009 -61434
rect -946 -61441 -912 -61196
rect -630 -61435 -596 -61233
rect -532 -61432 -498 -61233
rect -268 -61432 -234 -61233
rect -633 -61456 -596 -61435
rect -752 -61493 -596 -61456
rect -534 -61471 -234 -61432
rect -752 -61517 -715 -61493
rect -1046 -61554 -715 -61517
rect -170 -61524 -136 -61233
rect 26 -61250 62 -61196
rect 26 -61441 60 -61250
rect 124 -61524 158 -61233
rect 336 -61424 370 -61233
rect 429 -61240 472 -61156
rect 331 -61469 374 -61424
rect 434 -61441 468 -61240
rect 645 -61422 679 -61233
rect 738 -61242 781 -61156
rect 235 -61515 374 -61469
rect -663 -61585 -524 -61531
rect -403 -61558 158 -61524
rect -403 -61620 -369 -61558
rect -1045 -61689 -906 -61635
rect -515 -61654 -369 -61620
rect -515 -61769 -481 -61654
rect -296 -61659 -157 -61605
rect -1164 -61803 -481 -61769
rect -420 -61730 60 -61696
rect -1044 -62151 -1010 -61839
rect -946 -62047 -912 -61803
rect -848 -62151 -814 -61839
rect -728 -62082 -694 -61839
rect -630 -62047 -596 -61803
rect -532 -62082 -498 -61839
rect -420 -62082 -386 -61730
rect -728 -62116 -386 -62082
rect -350 -61804 -136 -61770
rect -350 -62151 -316 -61804
rect -1044 -62185 -316 -62151
rect -170 -62047 -136 -61804
rect 26 -62047 60 -61730
rect 113 -61733 252 -61679
rect 331 -61854 374 -61515
rect 415 -61579 554 -61525
rect 641 -61613 684 -61422
rect 743 -61441 777 -61242
rect 1452 -61245 1491 -61122
rect 2653 -61156 3285 -61122
rect 1554 -61196 2562 -61160
rect 541 -61659 684 -61613
rect 336 -62047 370 -61854
rect 641 -61856 684 -61659
rect 728 -61727 867 -61673
rect 645 -62047 679 -61856
rect 1310 -61402 1356 -61266
rect 1316 -61769 1350 -61402
rect 1456 -61434 1490 -61245
rect 1454 -61517 1491 -61434
rect 1554 -61441 1588 -61196
rect 1870 -61435 1904 -61233
rect 1968 -61432 2002 -61233
rect 2232 -61432 2266 -61233
rect 1867 -61456 1904 -61435
rect 1748 -61493 1904 -61456
rect 1966 -61471 2266 -61432
rect 1748 -61517 1785 -61493
rect 1454 -61554 1785 -61517
rect 2330 -61524 2364 -61233
rect 2526 -61250 2562 -61196
rect 2526 -61441 2560 -61250
rect 2624 -61524 2658 -61233
rect 2836 -61424 2870 -61233
rect 2929 -61240 2972 -61156
rect 2831 -61469 2874 -61424
rect 2934 -61441 2968 -61240
rect 3145 -61422 3179 -61233
rect 3238 -61242 3281 -61156
rect 2735 -61515 2874 -61469
rect 1837 -61585 1976 -61531
rect 2097 -61558 2658 -61524
rect 2097 -61620 2131 -61558
rect 1455 -61689 1594 -61635
rect 1985 -61654 2131 -61620
rect 1985 -61769 2019 -61654
rect 2204 -61659 2343 -61605
rect 1316 -61803 2019 -61769
rect 2080 -61730 2560 -61696
rect 1316 -61804 1350 -61803
rect 1456 -62151 1490 -61839
rect 1554 -62047 1588 -61803
rect 1652 -62151 1686 -61839
rect 1772 -62082 1806 -61839
rect 1870 -62047 1904 -61803
rect 1968 -62082 2002 -61839
rect 2080 -62082 2114 -61730
rect 1772 -62116 2114 -62082
rect 2150 -61804 2364 -61770
rect 2150 -62151 2184 -61804
rect 1456 -62185 2184 -62151
rect 2330 -62047 2364 -61804
rect 2526 -62047 2560 -61730
rect 2613 -61733 2752 -61679
rect 2831 -61854 2874 -61515
rect 2915 -61579 3054 -61525
rect 3141 -61613 3184 -61422
rect 3243 -61441 3277 -61242
rect 3952 -61245 3991 -61122
rect 5153 -61156 5785 -61122
rect 4054 -61196 5062 -61160
rect 3727 -61402 3773 -61266
rect 3732 -61403 3767 -61402
rect 3041 -61659 3184 -61613
rect 2836 -62047 2870 -61854
rect 3141 -61856 3184 -61659
rect 3228 -61727 3367 -61673
rect 3732 -61769 3766 -61403
rect 3956 -61434 3990 -61245
rect 3954 -61517 3991 -61434
rect 4054 -61441 4088 -61196
rect 4370 -61435 4404 -61233
rect 4468 -61432 4502 -61233
rect 4732 -61432 4766 -61233
rect 4367 -61456 4404 -61435
rect 4248 -61493 4404 -61456
rect 4466 -61471 4766 -61432
rect 4248 -61517 4285 -61493
rect 3954 -61554 4285 -61517
rect 4830 -61524 4864 -61233
rect 5026 -61250 5062 -61196
rect 5026 -61441 5060 -61250
rect 5124 -61524 5158 -61233
rect 5336 -61424 5370 -61233
rect 5429 -61240 5472 -61156
rect 5331 -61469 5374 -61424
rect 5434 -61441 5468 -61240
rect 5645 -61422 5679 -61233
rect 5738 -61242 5781 -61156
rect 5235 -61515 5374 -61469
rect 4597 -61558 5158 -61524
rect 4597 -61620 4631 -61558
rect 3955 -61689 4094 -61635
rect 4485 -61654 4631 -61620
rect 4485 -61769 4519 -61654
rect 4704 -61659 4843 -61605
rect 3732 -61803 4519 -61769
rect 4580 -61730 5060 -61696
rect 3145 -62047 3179 -61856
rect 3956 -62151 3990 -61839
rect 4054 -62047 4088 -61803
rect 4152 -62151 4186 -61839
rect 4272 -62082 4306 -61839
rect 4370 -62047 4404 -61803
rect 4468 -62082 4502 -61839
rect 4580 -62082 4614 -61730
rect 4272 -62116 4614 -62082
rect 4650 -61804 4864 -61770
rect 4650 -62151 4684 -61804
rect 3956 -62185 4684 -62151
rect 4830 -62047 4864 -61804
rect 5026 -62047 5060 -61730
rect 5113 -61733 5252 -61679
rect 5331 -61854 5374 -61515
rect 5641 -61613 5684 -61422
rect 5743 -61441 5777 -61242
rect 6952 -61245 6991 -61122
rect 7054 -61196 8062 -61160
rect 8137 -61174 9205 -61122
rect 6632 -61402 6678 -61266
rect 5541 -61659 5684 -61613
rect 5336 -62047 5370 -61854
rect 5641 -61856 5684 -61659
rect 5728 -61727 5867 -61673
rect 6638 -61769 6672 -61402
rect 6956 -61434 6990 -61245
rect 6954 -61517 6991 -61434
rect 7054 -61441 7088 -61196
rect 7370 -61435 7404 -61233
rect 7468 -61432 7502 -61233
rect 7732 -61432 7766 -61233
rect 7367 -61456 7404 -61435
rect 7248 -61493 7404 -61456
rect 7466 -61471 7766 -61432
rect 7248 -61517 7285 -61493
rect 6954 -61554 7285 -61517
rect 7830 -61524 7864 -61233
rect 8026 -61250 8062 -61196
rect 8026 -61441 8060 -61250
rect 8124 -61524 8158 -61233
rect 8336 -61424 8370 -61233
rect 8429 -61240 8472 -61174
rect 8331 -61469 8374 -61424
rect 8434 -61441 8468 -61240
rect 8645 -61422 8679 -61233
rect 8738 -61242 8781 -61174
rect 8235 -61515 8374 -61469
rect 7597 -61558 8158 -61524
rect 7597 -61620 7631 -61558
rect 6955 -61689 7094 -61635
rect 7485 -61654 7631 -61620
rect 7485 -61769 7519 -61654
rect 7704 -61659 7843 -61605
rect 6638 -61803 7519 -61769
rect 7580 -61730 8060 -61696
rect 5645 -62047 5679 -61856
rect 6956 -62151 6990 -61839
rect 7054 -62047 7088 -61803
rect 7152 -62151 7186 -61839
rect 7272 -62082 7306 -61839
rect 7370 -62047 7404 -61803
rect 7468 -62082 7502 -61839
rect 7580 -62082 7614 -61730
rect 7272 -62116 7614 -62082
rect 7650 -61804 7864 -61770
rect 7650 -62151 7684 -61804
rect 6956 -62185 7684 -62151
rect 7830 -62047 7864 -61804
rect 8026 -62047 8060 -61730
rect 8113 -61733 8252 -61679
rect 8331 -61854 8374 -61515
rect 8641 -61613 8684 -61422
rect 8743 -61441 8777 -61242
rect 8541 -61659 8684 -61613
rect 8336 -62047 8370 -61854
rect 8641 -61856 8684 -61659
rect 8728 -61727 8867 -61673
rect 8645 -62047 8679 -61856
rect -18303 -62388 -18165 -62387
rect -23449 -62458 -22910 -62448
rect -21509 -62433 -21351 -62400
rect -6608 -62406 -6445 -62387
rect -18441 -62433 -18304 -62428
rect -21509 -62485 -18304 -62433
rect -21509 -62516 -21351 -62485
rect -18441 -62486 -18304 -62485
rect 9838 -59846 10099 -59052
rect 18544 -59083 18580 -59030
rect 19002 -59037 19145 -59030
rect 14463 -59245 18580 -59083
rect 18872 -59112 19220 -59076
rect 10321 -59408 10390 -59390
rect 15534 -59408 15645 -59245
rect 10321 -59519 15645 -59408
rect 10321 -59529 10390 -59519
rect 18872 -59151 18908 -59112
rect 18873 -59554 18907 -59151
rect 19084 -59526 19118 -59146
rect 19175 -59156 19220 -59112
rect 19077 -59590 19123 -59526
rect 19182 -59554 19216 -59156
rect 19277 -59192 19327 -58963
rect 19948 -58994 20091 -58977
rect 19665 -59030 20091 -58994
rect 19948 -59037 20091 -59030
rect 19818 -59112 20166 -59076
rect 19280 -59526 19314 -59192
rect 19275 -59590 19321 -59526
rect 19818 -59151 19854 -59112
rect 19077 -59628 19321 -59590
rect 19819 -59554 19853 -59151
rect 20030 -59526 20064 -59146
rect 20121 -59156 20166 -59112
rect 20023 -59590 20069 -59526
rect 20128 -59554 20162 -59156
rect 20223 -59192 20273 -58947
rect 20226 -59526 20260 -59192
rect 20313 -59212 20373 -59046
rect 20548 -59134 20582 -58947
rect 20637 -59044 20671 -58673
rect 20735 -58981 20769 -58551
rect 20947 -58574 21388 -58540
rect 20947 -58577 21178 -58574
rect 20833 -59043 20867 -58673
rect 20947 -58681 20982 -58577
rect 20947 -58980 20981 -58681
rect 21045 -58980 21079 -58672
rect 21143 -58683 21178 -58577
rect 21143 -58980 21177 -58683
rect 21045 -59043 21080 -58980
rect 20833 -59044 21080 -59043
rect 21256 -59044 21290 -58672
rect 21354 -58980 21388 -58574
rect 21452 -59044 21486 -58672
rect 21767 -58880 21801 -58484
rect 21869 -58500 22185 -58484
rect 21869 -58535 22184 -58500
rect 20637 -59078 21080 -59044
rect 21253 -59078 21486 -59044
rect 21865 -59065 21899 -58672
rect 22103 -58841 22184 -58535
rect 22546 -58838 22580 -58526
rect 22644 -58754 22678 -58526
rect 22756 -58754 22790 -58526
rect 22854 -58734 22888 -58450
rect 22984 -58463 23044 -58450
rect 22644 -58789 22790 -58754
rect 22513 -58841 22992 -58838
rect 23082 -58841 23152 -57804
rect 22103 -58999 23152 -58841
rect 22487 -59042 23152 -58999
rect 23209 -58683 23279 -57949
rect 23376 -58625 23410 -57804
rect 23474 -58681 23508 -57917
rect 23776 -58625 23810 -57804
rect 23706 -58681 23840 -58668
rect 23209 -58737 23438 -58683
rect 23474 -58715 23840 -58681
rect 21084 -59134 21219 -59127
rect 20543 -59168 21219 -59134
rect 21084 -59181 21219 -59168
rect 21253 -59132 21290 -59078
rect 21865 -59101 22142 -59065
rect 21695 -59132 21830 -59125
rect 21253 -59169 21830 -59132
rect 20896 -59212 21031 -59205
rect 20313 -59250 21031 -59212
rect 20896 -59259 21031 -59250
rect 20560 -59296 20695 -59287
rect 20428 -59331 20695 -59296
rect 21253 -59307 21290 -59169
rect 21695 -59179 21830 -59169
rect 20428 -59428 20488 -59331
rect 20541 -59333 20695 -59331
rect 20560 -59341 20695 -59333
rect 20735 -59344 21290 -59307
rect 20221 -59590 20267 -59526
rect 20023 -59628 20267 -59590
rect 20735 -59588 20769 -59344
rect 20931 -59588 20965 -59344
rect 21127 -59588 21161 -59344
rect 21865 -59588 21899 -59101
rect 22011 -59125 22142 -59101
rect 22496 -59201 22530 -59042
rect 22594 -59185 22628 -59093
rect 22384 -59309 22552 -59235
rect 22588 -59278 22634 -59185
rect 22692 -59201 22726 -59042
rect 22790 -59185 22824 -59093
rect 22784 -59278 22830 -59185
rect 22888 -59201 22922 -59042
rect 22986 -59185 23020 -59093
rect 22980 -59246 23026 -59185
rect 23209 -59246 23279 -58737
rect 22980 -59278 23279 -59246
rect 22588 -59316 23279 -59278
rect 22588 -59324 23026 -59316
rect 22588 -59577 22634 -59324
rect 22594 -59581 22628 -59577
rect 22784 -59389 22830 -59324
rect 22790 -59581 22824 -59389
rect 22980 -59389 23026 -59324
rect 22986 -59581 23020 -59389
rect 23474 -59510 23508 -58715
rect 23706 -58722 23840 -58715
rect 23874 -58671 23908 -57917
rect 23982 -58671 24100 -58659
rect 23874 -58705 24100 -58671
rect 23874 -59510 23908 -58705
rect 23982 -58717 24100 -58705
rect 24253 -58681 24323 -58500
rect 24376 -58625 24410 -57804
rect 24253 -58735 24427 -58681
rect 24474 -58691 24508 -57917
rect 24776 -58625 24810 -57804
rect 24706 -58691 24840 -58683
rect 24474 -58730 24840 -58691
rect 24474 -59510 24508 -58730
rect 24706 -58737 24840 -58730
rect 24874 -58698 24908 -57917
rect 25059 -58698 25177 -58686
rect 24874 -58732 25177 -58698
rect 24874 -59510 24908 -58732
rect 25059 -58744 25177 -58732
rect 25244 -58688 25314 -58501
rect 25376 -58625 25410 -57804
rect 25244 -58742 25427 -58688
rect 25474 -58692 25508 -57917
rect 25776 -58625 25810 -57804
rect 25874 -58682 25908 -57917
rect 25955 -58682 26073 -58674
rect 25699 -58692 25833 -58685
rect 25474 -58731 25833 -58692
rect 25474 -59510 25508 -58731
rect 25699 -58739 25833 -58731
rect 25874 -58716 26076 -58682
rect 25874 -59510 25908 -58716
rect 25955 -58732 26073 -58716
rect 28086 -57943 28162 -56871
rect 28301 -56872 28787 -56871
rect 28301 -56873 28372 -56872
rect 28713 -56878 28787 -56872
rect 28333 -57223 28367 -56915
rect 28431 -57223 28465 -56915
rect 28529 -57223 28563 -56915
rect 28627 -57223 28661 -56915
rect 28725 -57223 28759 -56915
rect 28430 -57275 28465 -57223
rect 29144 -57257 29205 -56850
rect 29634 -57014 29704 -56619
rect 29878 -56873 29912 -56289
rect 30085 -56255 30325 -56221
rect 30085 -56297 30127 -56255
rect 29874 -56932 29916 -56873
rect 30089 -56879 30123 -56297
rect 30187 -56877 30221 -56289
rect 30283 -56299 30325 -56255
rect 30086 -56932 30128 -56879
rect 29874 -56968 30128 -56932
rect 30183 -56931 30225 -56877
rect 30285 -56897 30319 -56299
rect 30497 -56883 30531 -56289
rect 30183 -56970 30324 -56931
rect 30281 -56982 30324 -56970
rect 30039 -57014 30194 -57004
rect 29634 -57050 30194 -57014
rect 29634 -57052 29704 -57050
rect 30039 -57059 30194 -57050
rect 30281 -57037 30462 -56982
rect 30281 -57107 30324 -57037
rect 29769 -57121 29924 -57112
rect 29732 -57155 29924 -57121
rect 29769 -57167 29924 -57155
rect 29970 -57147 30324 -57107
rect 30496 -57127 30539 -56883
rect 30733 -56952 30803 -55615
rect 36897 -55668 36931 -55460
rect 37093 -55668 37127 -55460
rect 37289 -55668 37323 -55460
rect 31870 -56647 31904 -56147
rect 32049 -56111 32370 -56077
rect 31869 -56693 31904 -56647
rect 32049 -56693 32089 -56111
rect 32138 -56151 32173 -56111
rect 32139 -56655 32173 -56151
rect 32237 -56648 32271 -56147
rect 32335 -56150 32370 -56111
rect 31869 -56733 32089 -56693
rect 32234 -56768 32272 -56648
rect 32335 -56655 32369 -56150
rect 32465 -56731 32499 -56147
rect 32791 -56661 32825 -56147
rect 33019 -56437 33053 -56147
rect 37870 -55797 37904 -55453
rect 38066 -55797 38100 -55453
rect 38239 -55602 38300 -55453
rect 38479 -55567 38513 -55411
rect 38577 -55567 38611 -55459
rect 38675 -55567 38709 -55411
rect 45468 -55452 45715 -55411
rect 46550 -55439 46685 -55431
rect 46530 -55441 46685 -55439
rect 38773 -55567 38807 -55459
rect 45468 -55469 45598 -55452
rect 45642 -55465 45715 -55452
rect 46323 -55477 46685 -55441
rect 47202 -55450 47987 -55364
rect 54666 -55377 54796 -55285
rect 54958 -55343 54992 -55087
rect 55056 -55343 55090 -55135
rect 55154 -55343 55188 -55087
rect 55252 -55309 55286 -55135
rect 55833 -55265 55867 -54957
rect 55931 -55265 55965 -54957
rect 56029 -55265 56063 -54957
rect 56127 -55265 56161 -54957
rect 56225 -55265 56259 -54957
rect 55801 -55308 55872 -55307
rect 56213 -55308 56287 -55302
rect 55801 -55309 56287 -55308
rect 55252 -55343 56287 -55309
rect 56644 -55330 56705 -54923
rect 61292 -54953 63143 -54802
rect 64424 -54796 65089 -54768
rect 64424 -54854 65459 -54796
rect 64424 -54935 64510 -54854
rect 64684 -54891 64719 -54854
rect 65009 -54857 65459 -54854
rect 61292 -55021 61668 -54953
rect 62893 -55004 63143 -54953
rect 63572 -55021 64510 -54935
rect 63420 -55311 63550 -55219
rect 63712 -55277 63746 -55021
rect 63810 -55277 63844 -55069
rect 63908 -55277 63942 -55021
rect 64006 -55243 64040 -55069
rect 64587 -55199 64621 -54891
rect 64685 -55199 64719 -54891
rect 64783 -55199 64817 -54891
rect 64881 -55199 64915 -54891
rect 64979 -55199 65013 -54891
rect 64555 -55242 64626 -55241
rect 64967 -55242 65041 -55236
rect 64555 -55243 65041 -55242
rect 64006 -55277 65041 -55243
rect 65398 -55264 65459 -54857
rect 70068 -54808 70406 -54712
rect 73844 -54751 74184 -54357
rect 79298 -54747 79568 -54626
rect 81311 -54747 81606 -54705
rect 83180 -54713 83391 -54357
rect 72056 -54808 72324 -54767
rect 70068 -54939 72324 -54808
rect 73577 -54779 74242 -54751
rect 73577 -54837 74612 -54779
rect 73577 -54918 73663 -54837
rect 73837 -54874 73872 -54837
rect 74162 -54840 74612 -54837
rect 70068 -55003 70406 -54939
rect 72056 -55007 72324 -54939
rect 72725 -55004 73663 -54918
rect 64007 -55281 65041 -55277
rect 64007 -55283 64556 -55281
rect 63594 -55311 63667 -55305
rect 64967 -55307 65041 -55281
rect 55253 -55347 56287 -55343
rect 55253 -55349 55802 -55347
rect 54840 -55377 54913 -55371
rect 56213 -55373 56287 -55347
rect 54666 -55418 54913 -55377
rect 55748 -55405 55883 -55397
rect 55728 -55407 55883 -55405
rect 54666 -55435 54796 -55418
rect 54840 -55431 54913 -55418
rect 55521 -55443 55883 -55407
rect 56400 -55416 57185 -55330
rect 63420 -55352 63667 -55311
rect 64502 -55339 64637 -55331
rect 64482 -55341 64637 -55339
rect 63420 -55369 63550 -55352
rect 63594 -55365 63667 -55352
rect 64275 -55377 64637 -55341
rect 65154 -55350 65939 -55264
rect 72573 -55294 72703 -55202
rect 72865 -55260 72899 -55004
rect 72963 -55260 72997 -55052
rect 73061 -55260 73095 -55004
rect 73159 -55226 73193 -55052
rect 73740 -55182 73774 -54874
rect 73838 -55182 73872 -54874
rect 73936 -55182 73970 -54874
rect 74034 -55182 74068 -54874
rect 74132 -55182 74166 -54874
rect 73708 -55225 73779 -55224
rect 74120 -55225 74194 -55219
rect 73708 -55226 74194 -55225
rect 73159 -55260 74194 -55226
rect 74551 -55247 74612 -54840
rect 79298 -54886 81606 -54747
rect 82941 -54741 83606 -54713
rect 82941 -54799 83976 -54741
rect 82941 -54880 83027 -54799
rect 83201 -54836 83236 -54799
rect 83526 -54802 83976 -54799
rect 79298 -54911 79568 -54886
rect 81311 -54978 81606 -54886
rect 82089 -54966 83027 -54880
rect 73160 -55264 74194 -55260
rect 73160 -55266 73709 -55264
rect 72747 -55294 72820 -55288
rect 74120 -55290 74194 -55264
rect 72573 -55335 72820 -55294
rect 73655 -55322 73790 -55314
rect 73635 -55324 73790 -55322
rect 64482 -55379 64637 -55377
rect 64502 -55385 64637 -55379
rect 64685 -55362 65104 -55354
rect 64685 -55392 65115 -55362
rect 55728 -55445 55883 -55443
rect 46530 -55479 46685 -55477
rect 46550 -55485 46685 -55479
rect 46733 -55462 47152 -55454
rect 46733 -55492 47163 -55462
rect 38361 -55602 38434 -55596
rect 38239 -55615 38434 -55602
rect 38261 -55643 38434 -55615
rect 38361 -55656 38434 -55643
rect 38871 -55626 39243 -55556
rect 38479 -55798 38513 -55690
rect 38675 -55798 38709 -55690
rect 38871 -55798 38905 -55626
rect 33018 -56530 33055 -56437
rect 33018 -56567 33155 -56530
rect 32791 -56695 32950 -56661
rect 32614 -56731 32752 -56720
rect 31870 -56806 32272 -56768
rect 32339 -56765 32752 -56731
rect 31633 -56817 31771 -56807
rect 31243 -56851 31771 -56817
rect 30722 -57024 30827 -56952
rect 31243 -57127 31286 -56851
rect 31633 -56861 31771 -56851
rect 31689 -56952 31827 -56943
rect 31479 -56986 31827 -56952
rect 31479 -57113 31551 -56986
rect 31689 -56997 31827 -56986
rect 31479 -57122 31563 -57113
rect 28755 -57275 29205 -57257
rect 28313 -57318 29205 -57275
rect 28313 -57336 28762 -57318
rect 29144 -57613 29205 -57318
rect 29878 -57495 29912 -57201
rect 29970 -57217 30015 -57147
rect 30362 -57167 31286 -57127
rect 30410 -57170 31286 -57167
rect 29871 -57613 29918 -57495
rect 29976 -57509 30010 -57217
rect 30074 -57494 30108 -57201
rect 30316 -57484 30350 -57201
rect 30410 -57210 30454 -57170
rect 31484 -57192 31563 -57122
rect 30067 -57613 30114 -57494
rect 30309 -57613 30356 -57484
rect 30414 -57509 30448 -57210
rect 31772 -57434 31806 -57143
rect 31770 -57545 31807 -57434
rect 31870 -57451 31904 -56806
rect 32099 -56876 32137 -56806
rect 32339 -56844 32373 -56765
rect 32614 -56774 32752 -56765
rect 32089 -57014 32143 -56876
rect 32242 -56878 32373 -56844
rect 32439 -56861 32577 -56807
rect 32824 -56876 32878 -56738
rect 32916 -56739 32950 -56695
rect 32916 -56793 33082 -56739
rect 32242 -57451 32276 -56878
rect 32916 -56908 32950 -56793
rect 33002 -56908 33056 -56891
rect 32340 -56947 32499 -56912
rect 32916 -56913 33056 -56908
rect 32888 -56942 33056 -56913
rect 32340 -57451 32374 -56947
rect 32465 -57451 32499 -56947
rect 32563 -57434 32597 -56943
rect 32693 -57433 32727 -56943
rect 31233 -57549 31844 -57545
rect 32562 -57549 32599 -57434
rect 32690 -57549 32727 -57433
rect 32791 -57451 32825 -56943
rect 32888 -56947 32950 -56942
rect 32889 -57451 32923 -56947
rect 33002 -56950 33056 -56942
rect 33117 -57060 33155 -56567
rect 33117 -57098 33409 -57060
rect 33019 -57432 33053 -57143
rect 33117 -57148 33155 -57098
rect 33017 -57549 33054 -57432
rect 33117 -57451 33151 -57148
rect 31233 -57613 33167 -57549
rect 29144 -57658 33167 -57613
rect 29144 -57726 31346 -57658
rect 31694 -57710 33167 -57658
rect 9838 -60107 10808 -59846
rect 9986 -60550 10134 -60502
rect 9830 -60685 9953 -60641
rect 9671 -60812 9828 -60772
rect 9671 -62343 9725 -60812
rect 9885 -61116 9939 -60685
rect 9786 -61170 9939 -61116
rect 9786 -62343 9840 -61170
rect 9930 -62248 9984 -62218
rect 10028 -62248 10082 -60550
rect 10547 -61887 10808 -60107
rect 27290 -57999 28162 -57943
rect 33371 -57993 33409 -57098
rect 27290 -58075 31396 -57999
rect 27290 -58089 28162 -58075
rect 12071 -60362 12105 -60358
rect 12065 -60615 12111 -60362
rect 12267 -60550 12301 -60358
rect 12261 -60615 12307 -60550
rect 12463 -60550 12497 -60358
rect 12732 -60544 12789 -60380
rect 12457 -60615 12503 -60550
rect 12953 -60362 12987 -60358
rect 12065 -60623 12503 -60615
rect 12947 -60615 12993 -60362
rect 13149 -60550 13183 -60358
rect 13143 -60615 13189 -60550
rect 13563 -60339 14191 -60305
rect 13345 -60550 13379 -60358
rect 13563 -60384 13599 -60339
rect 13339 -60615 13385 -60550
rect 12947 -60623 13385 -60615
rect 13440 -60599 13514 -60431
rect 13564 -60458 13598 -60384
rect 13440 -60623 13513 -60599
rect 12065 -60645 12533 -60623
rect 12743 -60641 12911 -60630
rect 12591 -60645 12651 -60641
rect 12708 -60645 12911 -60641
rect 12065 -60661 12911 -60645
rect 11973 -60897 12007 -60738
rect 12065 -60754 12111 -60661
rect 12071 -60846 12105 -60754
rect 12169 -60897 12203 -60738
rect 12261 -60754 12307 -60661
rect 12457 -60687 12911 -60661
rect 12457 -60693 12533 -60687
rect 12267 -60846 12301 -60754
rect 12365 -60897 12399 -60738
rect 12457 -60754 12503 -60693
rect 12463 -60846 12497 -60754
rect 12591 -60773 12651 -60687
rect 12708 -60699 12911 -60687
rect 12743 -60704 12911 -60699
rect 12947 -60661 13513 -60623
rect 12855 -60897 12889 -60738
rect 12947 -60754 12993 -60661
rect 12953 -60846 12987 -60754
rect 13051 -60897 13085 -60738
rect 13143 -60754 13189 -60661
rect 13339 -60693 13513 -60661
rect 13558 -60605 13605 -60458
rect 13662 -60465 13696 -60373
rect 13759 -60394 13801 -60339
rect 13661 -60517 13697 -60465
rect 13760 -60481 13794 -60394
rect 13858 -60463 13892 -60373
rect 13953 -60395 13995 -60339
rect 13858 -60481 13895 -60463
rect 13956 -60481 13990 -60395
rect 14054 -60463 14088 -60373
rect 14149 -60390 14191 -60339
rect 13859 -60517 13895 -60481
rect 14053 -60517 14089 -60463
rect 14152 -60481 14186 -60390
rect 14250 -60473 14284 -60373
rect 14247 -60517 14289 -60473
rect 13661 -60551 14289 -60517
rect 13558 -60679 13730 -60605
rect 14114 -60639 14289 -60551
rect 14696 -60362 14730 -60358
rect 14690 -60615 14736 -60362
rect 14892 -60550 14926 -60358
rect 14886 -60615 14932 -60550
rect 15088 -60550 15122 -60358
rect 15432 -60458 15489 -60380
rect 15228 -60503 15489 -60458
rect 15082 -60615 15128 -60550
rect 14690 -60623 15128 -60615
rect 14486 -60639 14654 -60630
rect 13149 -60846 13183 -60754
rect 13247 -60897 13281 -60738
rect 13339 -60754 13385 -60693
rect 13345 -60846 13379 -60754
rect 13558 -60814 13605 -60679
rect 14114 -60696 14654 -60639
rect 14114 -60718 14289 -60696
rect 14486 -60704 14654 -60696
rect 14690 -60637 15158 -60623
rect 15228 -60637 15273 -60503
rect 15432 -60544 15489 -60503
rect 15653 -60362 15687 -60358
rect 15647 -60615 15693 -60362
rect 15849 -60550 15883 -60358
rect 15843 -60615 15889 -60550
rect 16263 -60339 16891 -60305
rect 16045 -60550 16079 -60358
rect 16263 -60384 16299 -60339
rect 16039 -60615 16085 -60550
rect 15647 -60623 16085 -60615
rect 16140 -60599 16214 -60431
rect 16264 -60458 16298 -60384
rect 16140 -60623 16213 -60599
rect 14690 -60661 15273 -60637
rect 13658 -60752 14289 -60718
rect 13658 -60793 13699 -60752
rect 13564 -60884 13598 -60814
rect 11964 -60965 13380 -60897
rect 13559 -60942 13603 -60884
rect 13662 -60896 13696 -60793
rect 13760 -60873 13794 -60788
rect 13856 -60801 13897 -60752
rect 13755 -60942 13799 -60873
rect 13858 -60896 13892 -60801
rect 13956 -60873 13990 -60788
rect 14050 -60801 14091 -60752
rect 14247 -60759 14289 -60752
rect 13951 -60942 13995 -60873
rect 14054 -60896 14088 -60801
rect 14152 -60884 14186 -60788
rect 14247 -60792 14288 -60759
rect 14241 -60802 14288 -60792
rect 14148 -60942 14192 -60884
rect 14241 -60924 14287 -60802
rect 14598 -60897 14632 -60738
rect 14690 -60754 14736 -60661
rect 14696 -60846 14730 -60754
rect 14794 -60897 14828 -60738
rect 14886 -60754 14932 -60661
rect 15082 -60682 15273 -60661
rect 15082 -60693 15158 -60682
rect 14892 -60846 14926 -60754
rect 14990 -60897 15024 -60738
rect 15082 -60754 15128 -60693
rect 15088 -60846 15122 -60754
rect 15208 -60797 15268 -60682
rect 15647 -60661 16213 -60623
rect 15555 -60897 15589 -60738
rect 15647 -60754 15693 -60661
rect 15653 -60846 15687 -60754
rect 15751 -60897 15785 -60738
rect 15843 -60754 15889 -60661
rect 16039 -60693 16213 -60661
rect 16258 -60605 16305 -60458
rect 16362 -60465 16396 -60373
rect 16459 -60394 16501 -60339
rect 16361 -60517 16397 -60465
rect 16460 -60481 16494 -60394
rect 16558 -60463 16592 -60373
rect 16653 -60395 16695 -60339
rect 16558 -60481 16595 -60463
rect 16656 -60481 16690 -60395
rect 16754 -60463 16788 -60373
rect 16849 -60390 16891 -60339
rect 16559 -60517 16595 -60481
rect 16753 -60517 16789 -60463
rect 16852 -60481 16886 -60390
rect 16950 -60473 16984 -60373
rect 16947 -60517 16989 -60473
rect 16361 -60551 16989 -60517
rect 16258 -60679 16430 -60605
rect 16814 -60636 16989 -60551
rect 17396 -60362 17430 -60358
rect 17390 -60615 17436 -60362
rect 17592 -60550 17626 -60358
rect 17586 -60615 17632 -60550
rect 17788 -60550 17822 -60358
rect 17782 -60615 17828 -60550
rect 17390 -60623 17828 -60615
rect 17186 -60636 17354 -60630
rect 15849 -60846 15883 -60754
rect 15947 -60897 15981 -60738
rect 16039 -60754 16085 -60693
rect 16045 -60846 16079 -60754
rect 16258 -60814 16305 -60679
rect 16814 -60689 17354 -60636
rect 16814 -60718 16989 -60689
rect 17186 -60704 17354 -60689
rect 17390 -60632 17858 -60623
rect 17390 -60634 17940 -60632
rect 17390 -60661 17941 -60634
rect 16358 -60752 16989 -60718
rect 16358 -60793 16399 -60752
rect 16264 -60884 16298 -60814
rect 13559 -60976 14192 -60942
rect 14589 -60965 16080 -60897
rect 16259 -60942 16303 -60884
rect 16362 -60896 16396 -60793
rect 16460 -60873 16494 -60788
rect 16556 -60801 16597 -60752
rect 16455 -60942 16499 -60873
rect 16558 -60896 16592 -60801
rect 16656 -60873 16690 -60788
rect 16750 -60801 16791 -60752
rect 16947 -60759 16989 -60752
rect 16651 -60942 16695 -60873
rect 16754 -60896 16788 -60801
rect 16852 -60884 16886 -60788
rect 16947 -60802 16988 -60759
rect 16848 -60942 16892 -60884
rect 16950 -60896 16984 -60802
rect 17298 -60897 17332 -60738
rect 17390 -60754 17436 -60661
rect 17396 -60846 17430 -60754
rect 17494 -60897 17528 -60738
rect 17586 -60754 17632 -60661
rect 17782 -60671 17941 -60661
rect 17782 -60693 17858 -60671
rect 17592 -60846 17626 -60754
rect 17690 -60897 17724 -60738
rect 17782 -60754 17828 -60693
rect 17788 -60846 17822 -60754
rect 16259 -60976 16892 -60942
rect 17289 -60965 17823 -60897
rect 12550 -61012 12682 -61001
rect 17073 -61012 17205 -60999
rect 12550 -61051 17611 -61012
rect 17893 -61029 17941 -60671
rect 12550 -61061 12682 -61051
rect 17073 -61059 17205 -61051
rect 17882 -61166 17942 -61029
rect 12227 -61190 12359 -61171
rect 14860 -61190 14997 -61171
rect 17457 -61190 17594 -61177
rect 12226 -61229 17611 -61190
rect 12227 -61231 12592 -61229
rect 12331 -61887 12592 -61231
rect 12948 -61300 13581 -61266
rect 13985 -61277 14096 -61229
rect 14860 -61231 14997 -61229
rect 14271 -61277 14791 -61275
rect 14863 -61277 14974 -61231
rect 12856 -61440 12890 -61346
rect 12948 -61358 12992 -61300
rect 12852 -61483 12893 -61440
rect 12954 -61454 12988 -61358
rect 13052 -61441 13086 -61346
rect 13145 -61369 13189 -61300
rect 12851 -61490 12893 -61483
rect 13049 -61490 13090 -61441
rect 13150 -61454 13184 -61369
rect 13248 -61441 13282 -61346
rect 13341 -61369 13385 -61300
rect 13243 -61490 13284 -61441
rect 13346 -61454 13380 -61369
rect 13444 -61449 13478 -61346
rect 13537 -61358 13581 -61300
rect 13760 -61343 15131 -61277
rect 13760 -61345 14294 -61343
rect 14597 -61345 15131 -61343
rect 15648 -61300 16281 -61266
rect 16661 -61277 16772 -61229
rect 17457 -61237 17594 -61229
rect 17472 -61277 17583 -61237
rect 13542 -61428 13576 -61358
rect 13441 -61490 13482 -61449
rect 12851 -61522 13482 -61490
rect 12776 -61524 13482 -61522
rect 12776 -61582 13026 -61524
rect 13535 -61563 13582 -61428
rect 13761 -61488 13795 -61396
rect 13755 -61549 13801 -61488
rect 13859 -61504 13893 -61345
rect 13957 -61488 13991 -61396
rect 12851 -61691 13026 -61582
rect 13410 -61637 13582 -61563
rect 12851 -61725 13479 -61691
rect 12851 -61769 12893 -61725
rect 12856 -61869 12890 -61769
rect 12954 -61852 12988 -61761
rect 13051 -61779 13087 -61725
rect 13245 -61761 13281 -61725
rect 10547 -62148 12592 -61887
rect 12949 -61903 12991 -61852
rect 13052 -61869 13086 -61779
rect 13150 -61847 13184 -61761
rect 13245 -61779 13282 -61761
rect 13145 -61903 13187 -61847
rect 13248 -61869 13282 -61779
rect 13346 -61848 13380 -61761
rect 13443 -61777 13479 -61725
rect 13339 -61903 13381 -61848
rect 13444 -61869 13478 -61777
rect 13535 -61784 13582 -61637
rect 13627 -61581 13801 -61549
rect 13951 -61581 13997 -61488
rect 14055 -61504 14089 -61345
rect 14153 -61488 14187 -61396
rect 14147 -61581 14193 -61488
rect 14251 -61504 14285 -61345
rect 14598 -61488 14632 -61396
rect 13627 -61619 14193 -61581
rect 14592 -61549 14638 -61488
rect 14696 -61504 14730 -61345
rect 14794 -61488 14828 -61396
rect 14494 -61581 14638 -61549
rect 14788 -61581 14834 -61488
rect 14892 -61504 14926 -61345
rect 14990 -61488 15024 -61396
rect 14984 -61581 15030 -61488
rect 15088 -61504 15122 -61345
rect 15556 -61440 15590 -61346
rect 15648 -61358 15692 -61300
rect 15552 -61483 15593 -61440
rect 15654 -61454 15688 -61358
rect 15752 -61441 15786 -61346
rect 15845 -61369 15889 -61300
rect 15551 -61490 15593 -61483
rect 15749 -61490 15790 -61441
rect 15850 -61454 15884 -61369
rect 15948 -61441 15982 -61346
rect 16041 -61369 16085 -61300
rect 15943 -61490 15984 -61441
rect 16046 -61454 16080 -61369
rect 16144 -61449 16178 -61346
rect 16237 -61358 16281 -61300
rect 16460 -61345 17831 -61277
rect 16242 -61428 16276 -61358
rect 16141 -61490 16182 -61449
rect 15551 -61524 16182 -61490
rect 13627 -61643 13700 -61619
rect 13542 -61858 13576 -61784
rect 13626 -61811 13700 -61643
rect 13755 -61627 14193 -61619
rect 13755 -61692 13801 -61627
rect 13541 -61903 13577 -61858
rect 13761 -61884 13795 -61692
rect 12949 -61937 13577 -61903
rect 13951 -61692 13997 -61627
rect 13957 -61884 13991 -61692
rect 14147 -61880 14193 -61627
rect 14494 -61619 15030 -61581
rect 15066 -61545 15234 -61538
rect 15066 -61605 15256 -61545
rect 15460 -61584 15726 -61524
rect 16235 -61563 16282 -61428
rect 16461 -61488 16495 -61396
rect 16455 -61549 16501 -61488
rect 16559 -61504 16593 -61345
rect 16657 -61488 16691 -61396
rect 15066 -61612 15234 -61605
rect 14153 -61884 14187 -61880
rect 14351 -61748 14408 -61698
rect 14494 -61748 14556 -61619
rect 14592 -61627 15030 -61619
rect 14592 -61692 14638 -61627
rect 14351 -61810 14556 -61748
rect 14351 -61862 14408 -61810
rect 14598 -61884 14632 -61692
rect 14788 -61692 14834 -61627
rect 14794 -61884 14828 -61692
rect 14984 -61880 15030 -61627
rect 14990 -61884 15024 -61880
rect 15551 -61691 15726 -61584
rect 16110 -61637 16282 -61563
rect 15551 -61725 16179 -61691
rect 15551 -61769 15593 -61725
rect 15556 -61869 15590 -61769
rect 15654 -61852 15688 -61761
rect 15751 -61779 15787 -61725
rect 15945 -61761 15981 -61725
rect 15649 -61903 15691 -61852
rect 15752 -61869 15786 -61779
rect 15850 -61847 15884 -61761
rect 15945 -61779 15982 -61761
rect 15845 -61903 15887 -61847
rect 15948 -61869 15982 -61779
rect 16046 -61848 16080 -61761
rect 16143 -61777 16179 -61725
rect 16039 -61903 16081 -61848
rect 16144 -61869 16178 -61777
rect 16235 -61784 16282 -61637
rect 16327 -61581 16501 -61549
rect 16651 -61581 16697 -61488
rect 16755 -61504 16789 -61345
rect 16853 -61488 16887 -61396
rect 16847 -61581 16893 -61488
rect 16951 -61504 16985 -61345
rect 17109 -61538 17169 -61394
rect 17298 -61488 17332 -61396
rect 16327 -61619 16893 -61581
rect 16929 -61600 17169 -61538
rect 17292 -61549 17338 -61488
rect 17396 -61504 17430 -61345
rect 17494 -61488 17528 -61396
rect 17205 -61581 17338 -61549
rect 17488 -61581 17534 -61488
rect 17592 -61504 17626 -61345
rect 17690 -61488 17724 -61396
rect 17684 -61581 17730 -61488
rect 17788 -61504 17822 -61345
rect 17893 -61538 17941 -61166
rect 16929 -61601 17132 -61600
rect 16929 -61612 17097 -61601
rect 16327 -61643 16400 -61619
rect 16242 -61858 16276 -61784
rect 16326 -61811 16400 -61643
rect 16455 -61627 16893 -61619
rect 16455 -61692 16501 -61627
rect 16241 -61903 16277 -61858
rect 16461 -61884 16495 -61692
rect 15649 -61937 16277 -61903
rect 16651 -61692 16697 -61627
rect 16657 -61884 16691 -61692
rect 16847 -61880 16893 -61627
rect 17205 -61619 17730 -61581
rect 17766 -61582 17941 -61538
rect 17766 -61612 17934 -61582
rect 16853 -61884 16887 -61880
rect 17051 -61749 17108 -61698
rect 17205 -61749 17251 -61619
rect 17292 -61627 17730 -61619
rect 17292 -61692 17338 -61627
rect 17051 -61798 17251 -61749
rect 17051 -61862 17108 -61798
rect 17298 -61884 17332 -61692
rect 17488 -61692 17534 -61627
rect 17494 -61884 17528 -61692
rect 17684 -61880 17730 -61627
rect 17690 -61884 17724 -61880
rect 27290 -61839 27436 -58089
rect 28086 -58257 28162 -58089
rect 28086 -58333 28228 -58257
rect 28152 -58722 28228 -58333
rect 29161 -58299 29826 -58271
rect 29161 -58357 30196 -58299
rect 29161 -58438 29247 -58357
rect 29421 -58394 29456 -58357
rect 29746 -58360 30196 -58357
rect 28309 -58524 29247 -58438
rect 28152 -58814 28287 -58722
rect 28449 -58780 28483 -58524
rect 28547 -58780 28581 -58572
rect 28645 -58780 28679 -58524
rect 28743 -58746 28777 -58572
rect 29324 -58702 29358 -58394
rect 29422 -58702 29456 -58394
rect 29520 -58702 29554 -58394
rect 29618 -58702 29652 -58394
rect 29716 -58702 29750 -58394
rect 29292 -58745 29363 -58744
rect 29704 -58745 29778 -58739
rect 29292 -58746 29778 -58745
rect 28743 -58780 29778 -58746
rect 30135 -58767 30196 -58360
rect 28744 -58784 29778 -58780
rect 28744 -58786 29293 -58784
rect 28331 -58814 28404 -58808
rect 29704 -58810 29778 -58784
rect 28152 -58831 28404 -58814
rect 28157 -58855 28404 -58831
rect 29239 -58842 29374 -58834
rect 29219 -58844 29374 -58842
rect 28157 -58872 28287 -58855
rect 28331 -58868 28404 -58855
rect 29012 -58880 29374 -58844
rect 29891 -58853 30676 -58767
rect 29219 -58882 29374 -58880
rect 29239 -58888 29374 -58882
rect 29422 -58865 29841 -58857
rect 29422 -58895 29852 -58865
rect 28449 -59110 28483 -58902
rect 28645 -59110 28679 -58902
rect 28841 -59110 28875 -58902
rect 29422 -59239 29456 -58895
rect 29618 -59239 29652 -58895
rect 29791 -59044 29852 -58895
rect 30031 -59009 30065 -58853
rect 30129 -59009 30163 -58901
rect 30227 -59009 30261 -58853
rect 30325 -59009 30359 -58901
rect 29913 -59044 29986 -59038
rect 29791 -59057 29986 -59044
rect 29813 -59085 29986 -59057
rect 29913 -59098 29986 -59085
rect 30423 -59068 30795 -58998
rect 30031 -59240 30065 -59132
rect 30227 -59240 30261 -59132
rect 30423 -59240 30457 -59068
rect 28423 -60175 28457 -59831
rect 28619 -60175 28653 -59831
rect 29032 -59938 29066 -59830
rect 29228 -59938 29262 -59830
rect 28914 -59985 28987 -59972
rect 28814 -60013 28987 -59985
rect 28792 -60026 28987 -60013
rect 28792 -60175 28853 -60026
rect 28914 -60032 28987 -60026
rect 29424 -60002 29458 -59830
rect 28423 -60205 28853 -60175
rect 28423 -60213 28842 -60205
rect 29032 -60217 29066 -60061
rect 29130 -60169 29164 -60061
rect 29228 -60217 29262 -60061
rect 29326 -60169 29360 -60061
rect 29424 -60072 29702 -60002
rect 25424 -61841 27436 -61839
rect 28067 -60286 28294 -60284
rect 28705 -60286 28779 -60260
rect 28067 -60324 28779 -60286
rect 28892 -60303 29507 -60217
rect 28293 -60325 28779 -60324
rect 28293 -60326 28364 -60325
rect 28705 -60331 28779 -60325
rect 28325 -60676 28359 -60368
rect 28423 -60676 28457 -60368
rect 28521 -60676 28555 -60368
rect 28619 -60676 28653 -60368
rect 28717 -60676 28751 -60368
rect 28422 -60728 28457 -60676
rect 29136 -60710 29197 -60303
rect 29626 -60467 29696 -60072
rect 29870 -60326 29904 -59742
rect 30077 -59708 30317 -59674
rect 30077 -59750 30119 -59708
rect 29866 -60385 29908 -60326
rect 30081 -60332 30115 -59750
rect 30179 -60330 30213 -59742
rect 30275 -59752 30317 -59708
rect 30078 -60385 30120 -60332
rect 29866 -60421 30120 -60385
rect 30175 -60384 30217 -60330
rect 30277 -60350 30311 -59752
rect 30489 -60336 30523 -59742
rect 30175 -60423 30316 -60384
rect 30273 -60435 30316 -60423
rect 30031 -60467 30186 -60457
rect 29626 -60503 30186 -60467
rect 29626 -60505 29696 -60503
rect 30031 -60512 30186 -60503
rect 30273 -60490 30454 -60435
rect 30273 -60560 30316 -60490
rect 29761 -60574 29916 -60565
rect 29724 -60608 29916 -60574
rect 29761 -60620 29916 -60608
rect 29962 -60600 30316 -60560
rect 30488 -60580 30531 -60336
rect 30725 -60405 30795 -59068
rect 30970 -58356 31062 -58271
rect 30993 -60331 31036 -58356
rect 31320 -58779 31396 -58075
rect 31622 -58031 33409 -57993
rect 31622 -58409 31660 -58031
rect 32829 -58330 33494 -58302
rect 32829 -58388 33864 -58330
rect 31599 -58463 31672 -58409
rect 32829 -58469 32915 -58388
rect 33089 -58425 33124 -58388
rect 33414 -58391 33864 -58388
rect 31977 -58555 32915 -58469
rect 31825 -58779 31955 -58753
rect 31320 -58845 31955 -58779
rect 32117 -58811 32151 -58555
rect 32215 -58811 32249 -58603
rect 32313 -58811 32347 -58555
rect 32411 -58777 32445 -58603
rect 32992 -58733 33026 -58425
rect 33090 -58733 33124 -58425
rect 33188 -58733 33222 -58425
rect 33286 -58733 33320 -58425
rect 33384 -58733 33418 -58425
rect 32960 -58776 33031 -58775
rect 33372 -58776 33446 -58770
rect 32960 -58777 33446 -58776
rect 32411 -58811 33446 -58777
rect 33803 -58798 33864 -58391
rect 36871 -56733 36905 -56389
rect 37067 -56733 37101 -56389
rect 37480 -56496 37514 -56388
rect 37676 -56496 37710 -56388
rect 37362 -56543 37435 -56530
rect 37262 -56571 37435 -56543
rect 37240 -56584 37435 -56571
rect 37240 -56733 37301 -56584
rect 37362 -56590 37435 -56584
rect 37872 -56560 37906 -56388
rect 36871 -56763 37301 -56733
rect 36871 -56771 37290 -56763
rect 37480 -56775 37514 -56619
rect 37578 -56727 37612 -56619
rect 37676 -56775 37710 -56619
rect 37774 -56727 37808 -56619
rect 37872 -56630 38150 -56560
rect 32412 -58815 33446 -58811
rect 32412 -58817 32961 -58815
rect 31999 -58845 32072 -58839
rect 33372 -58841 33446 -58815
rect 31320 -58855 32072 -58845
rect 31825 -58886 32072 -58855
rect 32907 -58873 33042 -58865
rect 32887 -58875 33042 -58873
rect 31825 -58903 31955 -58886
rect 31999 -58899 32072 -58886
rect 31852 -58953 31928 -58903
rect 32680 -58911 33042 -58875
rect 33559 -58884 34344 -58798
rect 32887 -58913 33042 -58911
rect 32907 -58919 33042 -58913
rect 33090 -58896 33509 -58888
rect 33090 -58926 33520 -58896
rect 32117 -59141 32151 -58933
rect 32313 -59141 32347 -58933
rect 32509 -59141 32543 -58933
rect 33090 -59270 33124 -58926
rect 33286 -59270 33320 -58926
rect 33459 -59075 33520 -58926
rect 33699 -59040 33733 -58884
rect 33797 -59040 33831 -58932
rect 33895 -59040 33929 -58884
rect 33993 -59040 34027 -58932
rect 33581 -59075 33654 -59069
rect 33459 -59088 33654 -59075
rect 33481 -59116 33654 -59088
rect 33581 -59129 33654 -59116
rect 34091 -59099 34463 -59029
rect 33699 -59271 33733 -59163
rect 33895 -59271 33929 -59163
rect 34091 -59271 34125 -59099
rect 32091 -60206 32125 -59862
rect 32287 -60206 32321 -59862
rect 32700 -59969 32734 -59861
rect 32896 -59969 32930 -59861
rect 32582 -60016 32655 -60003
rect 32482 -60044 32655 -60016
rect 32460 -60057 32655 -60044
rect 32460 -60206 32521 -60057
rect 32582 -60063 32655 -60057
rect 33092 -60033 33126 -59861
rect 32091 -60236 32521 -60206
rect 32091 -60244 32510 -60236
rect 32700 -60248 32734 -60092
rect 32798 -60200 32832 -60092
rect 32896 -60248 32930 -60092
rect 32994 -60200 33028 -60092
rect 33092 -60103 33370 -60033
rect 30993 -60374 31278 -60331
rect 30714 -60477 30819 -60405
rect 31235 -60580 31278 -60374
rect 28747 -60728 29197 -60710
rect 28305 -60771 29197 -60728
rect 28305 -60789 28754 -60771
rect 29136 -61066 29197 -60771
rect 29870 -60948 29904 -60654
rect 29962 -60670 30007 -60600
rect 30354 -60620 31278 -60580
rect 30402 -60623 31278 -60620
rect 29863 -61066 29910 -60948
rect 29968 -60962 30002 -60670
rect 30066 -60947 30100 -60654
rect 30308 -60937 30342 -60654
rect 30402 -60663 30446 -60623
rect 30059 -61066 30106 -60947
rect 30301 -61066 30348 -60937
rect 30406 -60962 30440 -60663
rect 29136 -61179 30613 -61066
rect 31735 -60317 31962 -60315
rect 32373 -60317 32447 -60291
rect 31735 -60355 32447 -60317
rect 32560 -60334 33175 -60248
rect 31961 -60356 32447 -60355
rect 31961 -60357 32032 -60356
rect 32373 -60362 32447 -60356
rect 31993 -60707 32027 -60399
rect 32091 -60707 32125 -60399
rect 32189 -60707 32223 -60399
rect 32287 -60707 32321 -60399
rect 32385 -60707 32419 -60399
rect 32090 -60759 32125 -60707
rect 32804 -60741 32865 -60334
rect 33294 -60498 33364 -60103
rect 33538 -60357 33572 -59773
rect 33745 -59739 33985 -59705
rect 33745 -59781 33787 -59739
rect 33534 -60416 33576 -60357
rect 33749 -60363 33783 -59781
rect 33847 -60361 33881 -59773
rect 33943 -59783 33985 -59739
rect 33746 -60416 33788 -60363
rect 33534 -60452 33788 -60416
rect 33843 -60415 33885 -60361
rect 33945 -60381 33979 -59783
rect 34157 -60367 34191 -59773
rect 33843 -60454 33984 -60415
rect 33941 -60466 33984 -60454
rect 33699 -60498 33854 -60488
rect 33294 -60534 33854 -60498
rect 33294 -60536 33364 -60534
rect 33699 -60543 33854 -60534
rect 33941 -60521 34122 -60466
rect 33941 -60591 33984 -60521
rect 33429 -60605 33584 -60596
rect 33392 -60639 33584 -60605
rect 33429 -60651 33584 -60639
rect 33630 -60631 33984 -60591
rect 34156 -60611 34199 -60367
rect 34393 -60436 34463 -59099
rect 34382 -60508 34487 -60436
rect 34888 -60611 35111 -60521
rect 32415 -60759 32865 -60741
rect 31973 -60802 32865 -60759
rect 31973 -60820 32422 -60802
rect 32804 -61097 32865 -60802
rect 33538 -60979 33572 -60685
rect 33630 -60701 33675 -60631
rect 34022 -60651 35224 -60611
rect 34070 -60654 35224 -60651
rect 33531 -61097 33578 -60979
rect 33636 -60993 33670 -60701
rect 33734 -60978 33768 -60685
rect 33976 -60968 34010 -60685
rect 34070 -60694 34114 -60654
rect 34888 -60691 35111 -60654
rect 33727 -61097 33774 -60978
rect 33969 -61097 34016 -60968
rect 34074 -60993 34108 -60694
rect 32804 -61210 34281 -61097
rect 25424 -62009 27455 -61841
rect 25424 -62010 27379 -62009
rect 9930 -62302 10082 -62248
rect 9930 -62343 9984 -62302
rect 36515 -56844 36742 -56842
rect 37153 -56844 37227 -56818
rect 36515 -56882 37227 -56844
rect 37340 -56861 37955 -56775
rect 36526 -57732 36602 -56882
rect 36741 -56883 37227 -56882
rect 36741 -56884 36812 -56883
rect 37153 -56889 37227 -56883
rect 36773 -57234 36807 -56926
rect 36871 -57234 36905 -56926
rect 36969 -57234 37003 -56926
rect 37067 -57234 37101 -56926
rect 37165 -57234 37199 -56926
rect 36870 -57286 36905 -57234
rect 37584 -57268 37645 -56861
rect 38074 -57025 38144 -56630
rect 38318 -56884 38352 -56300
rect 38525 -56266 38765 -56232
rect 38525 -56308 38567 -56266
rect 38314 -56943 38356 -56884
rect 38529 -56890 38563 -56308
rect 38627 -56888 38661 -56300
rect 38723 -56310 38765 -56266
rect 38526 -56943 38568 -56890
rect 38314 -56979 38568 -56943
rect 38623 -56942 38665 -56888
rect 38725 -56908 38759 -56310
rect 38937 -56894 38971 -56300
rect 38623 -56981 38764 -56942
rect 38721 -56993 38764 -56981
rect 38479 -57025 38634 -57015
rect 38074 -57061 38634 -57025
rect 38074 -57063 38144 -57061
rect 38479 -57070 38634 -57061
rect 38721 -57048 38902 -56993
rect 38721 -57118 38764 -57048
rect 38209 -57132 38364 -57123
rect 38172 -57166 38364 -57132
rect 38209 -57178 38364 -57166
rect 38410 -57158 38764 -57118
rect 38936 -57138 38979 -56894
rect 39173 -56963 39243 -55626
rect 45760 -55707 45794 -55499
rect 45956 -55707 45990 -55499
rect 46152 -55707 46186 -55499
rect 46733 -55836 46767 -55492
rect 46929 -55836 46963 -55492
rect 47102 -55641 47163 -55492
rect 47342 -55606 47376 -55450
rect 47440 -55606 47474 -55498
rect 47538 -55606 47572 -55450
rect 55748 -55451 55883 -55445
rect 55931 -55428 56350 -55420
rect 55931 -55458 56361 -55428
rect 47636 -55606 47670 -55498
rect 47224 -55641 47297 -55635
rect 47102 -55654 47297 -55641
rect 47124 -55682 47297 -55654
rect 47224 -55695 47297 -55682
rect 47734 -55665 48106 -55595
rect 47342 -55837 47376 -55729
rect 47538 -55837 47572 -55729
rect 47734 -55837 47768 -55665
rect 40310 -56658 40344 -56158
rect 40489 -56122 40810 -56088
rect 40309 -56704 40344 -56658
rect 40489 -56704 40529 -56122
rect 40578 -56162 40613 -56122
rect 40579 -56666 40613 -56162
rect 40677 -56659 40711 -56158
rect 40775 -56161 40810 -56122
rect 40309 -56744 40529 -56704
rect 40674 -56779 40712 -56659
rect 40775 -56666 40809 -56161
rect 40905 -56742 40939 -56158
rect 41231 -56672 41265 -56158
rect 41459 -56448 41493 -56158
rect 41458 -56541 41495 -56448
rect 41458 -56578 41595 -56541
rect 41231 -56706 41390 -56672
rect 41054 -56742 41192 -56731
rect 40310 -56817 40712 -56779
rect 40779 -56776 41192 -56742
rect 40073 -56828 40211 -56818
rect 39683 -56862 40211 -56828
rect 39162 -57035 39267 -56963
rect 39683 -57138 39726 -56862
rect 40073 -56872 40211 -56862
rect 40129 -56963 40267 -56954
rect 39919 -56997 40267 -56963
rect 39919 -57124 39991 -56997
rect 40129 -57008 40267 -56997
rect 39919 -57133 40003 -57124
rect 37195 -57286 37645 -57268
rect 36753 -57329 37645 -57286
rect 36753 -57347 37202 -57329
rect 35870 -57878 36602 -57732
rect 37584 -57624 37645 -57329
rect 38318 -57506 38352 -57212
rect 38410 -57228 38455 -57158
rect 38802 -57178 39726 -57138
rect 38850 -57181 39726 -57178
rect 38311 -57624 38358 -57506
rect 38416 -57520 38450 -57228
rect 38514 -57505 38548 -57212
rect 38756 -57495 38790 -57212
rect 38850 -57221 38894 -57181
rect 39924 -57203 40003 -57133
rect 38507 -57624 38554 -57505
rect 38749 -57624 38796 -57495
rect 38854 -57520 38888 -57221
rect 40212 -57445 40246 -57154
rect 40210 -57556 40247 -57445
rect 40310 -57462 40344 -56817
rect 40539 -56887 40577 -56817
rect 40779 -56855 40813 -56776
rect 41054 -56785 41192 -56776
rect 40529 -57025 40583 -56887
rect 40682 -56889 40813 -56855
rect 40879 -56872 41017 -56818
rect 41264 -56887 41318 -56749
rect 41356 -56750 41390 -56706
rect 41356 -56804 41522 -56750
rect 40682 -57462 40716 -56889
rect 41356 -56919 41390 -56804
rect 41442 -56919 41496 -56902
rect 40780 -56958 40939 -56923
rect 41356 -56924 41496 -56919
rect 41328 -56953 41496 -56924
rect 40780 -57462 40814 -56958
rect 40905 -57462 40939 -56958
rect 41003 -57445 41037 -56954
rect 41133 -57444 41167 -56954
rect 39673 -57560 40284 -57556
rect 41002 -57560 41039 -57445
rect 41130 -57560 41167 -57444
rect 41231 -57462 41265 -56954
rect 41328 -56958 41390 -56953
rect 41329 -57462 41363 -56958
rect 41442 -56961 41496 -56953
rect 41557 -57071 41595 -56578
rect 41557 -57109 41849 -57071
rect 41459 -57443 41493 -57154
rect 41557 -57159 41595 -57109
rect 41457 -57560 41494 -57443
rect 41557 -57462 41591 -57159
rect 39673 -57624 41607 -57560
rect 37584 -57669 41607 -57624
rect 37584 -57737 39786 -57669
rect 40134 -57721 41607 -57669
rect 35870 -61861 36016 -57878
rect 36526 -58010 36602 -57878
rect 41811 -58004 41849 -57109
rect 36526 -58086 39836 -58010
rect 36526 -58268 36602 -58086
rect 36526 -58344 36668 -58268
rect 36592 -58733 36668 -58344
rect 37601 -58310 38266 -58282
rect 37601 -58368 38636 -58310
rect 37601 -58449 37687 -58368
rect 37861 -58405 37896 -58368
rect 38186 -58371 38636 -58368
rect 36749 -58535 37687 -58449
rect 36592 -58825 36727 -58733
rect 36889 -58791 36923 -58535
rect 36987 -58791 37021 -58583
rect 37085 -58791 37119 -58535
rect 37183 -58757 37217 -58583
rect 37764 -58713 37798 -58405
rect 37862 -58713 37896 -58405
rect 37960 -58713 37994 -58405
rect 38058 -58713 38092 -58405
rect 38156 -58713 38190 -58405
rect 37732 -58756 37803 -58755
rect 38144 -58756 38218 -58750
rect 37732 -58757 38218 -58756
rect 37183 -58791 38218 -58757
rect 38575 -58778 38636 -58371
rect 37184 -58795 38218 -58791
rect 37184 -58797 37733 -58795
rect 36771 -58825 36844 -58819
rect 38144 -58821 38218 -58795
rect 36592 -58842 36844 -58825
rect 36597 -58866 36844 -58842
rect 37679 -58853 37814 -58845
rect 37659 -58855 37814 -58853
rect 36597 -58883 36727 -58866
rect 36771 -58879 36844 -58866
rect 37452 -58891 37814 -58855
rect 38331 -58864 39116 -58778
rect 37659 -58893 37814 -58891
rect 37679 -58899 37814 -58893
rect 37862 -58876 38281 -58868
rect 37862 -58906 38292 -58876
rect 36889 -59121 36923 -58913
rect 37085 -59121 37119 -58913
rect 37281 -59121 37315 -58913
rect 37862 -59250 37896 -58906
rect 38058 -59250 38092 -58906
rect 38231 -59055 38292 -58906
rect 38471 -59020 38505 -58864
rect 38569 -59020 38603 -58912
rect 38667 -59020 38701 -58864
rect 38765 -59020 38799 -58912
rect 38353 -59055 38426 -59049
rect 38231 -59068 38426 -59055
rect 38253 -59096 38426 -59068
rect 38353 -59109 38426 -59096
rect 38863 -59079 39235 -59009
rect 38471 -59251 38505 -59143
rect 38667 -59251 38701 -59143
rect 38863 -59251 38897 -59079
rect 36863 -60186 36897 -59842
rect 37059 -60186 37093 -59842
rect 37472 -59949 37506 -59841
rect 37668 -59949 37702 -59841
rect 37354 -59996 37427 -59983
rect 37254 -60024 37427 -59996
rect 37232 -60037 37427 -60024
rect 37232 -60186 37293 -60037
rect 37354 -60043 37427 -60037
rect 37864 -60013 37898 -59841
rect 36863 -60216 37293 -60186
rect 36863 -60224 37282 -60216
rect 37472 -60228 37506 -60072
rect 37570 -60180 37604 -60072
rect 37668 -60228 37702 -60072
rect 37766 -60180 37800 -60072
rect 37864 -60083 38142 -60013
rect 36507 -60297 36734 -60295
rect 37145 -60297 37219 -60271
rect 36507 -60335 37219 -60297
rect 37332 -60314 37947 -60228
rect 36733 -60336 37219 -60335
rect 36733 -60337 36804 -60336
rect 37145 -60342 37219 -60336
rect 36765 -60687 36799 -60379
rect 36863 -60687 36897 -60379
rect 36961 -60687 36995 -60379
rect 37059 -60687 37093 -60379
rect 37157 -60687 37191 -60379
rect 36862 -60739 36897 -60687
rect 37576 -60721 37637 -60314
rect 38066 -60478 38136 -60083
rect 38310 -60337 38344 -59753
rect 38517 -59719 38757 -59685
rect 38517 -59761 38559 -59719
rect 38306 -60396 38348 -60337
rect 38521 -60343 38555 -59761
rect 38619 -60341 38653 -59753
rect 38715 -59763 38757 -59719
rect 38518 -60396 38560 -60343
rect 38306 -60432 38560 -60396
rect 38615 -60395 38657 -60341
rect 38717 -60361 38751 -59763
rect 38929 -60347 38963 -59753
rect 38615 -60434 38756 -60395
rect 38713 -60446 38756 -60434
rect 38471 -60478 38626 -60468
rect 38066 -60514 38626 -60478
rect 38066 -60516 38136 -60514
rect 38471 -60523 38626 -60514
rect 38713 -60501 38894 -60446
rect 38713 -60571 38756 -60501
rect 38201 -60585 38356 -60576
rect 38164 -60619 38356 -60585
rect 38201 -60631 38356 -60619
rect 38402 -60611 38756 -60571
rect 38928 -60591 38971 -60347
rect 39165 -60416 39235 -59079
rect 39410 -58367 39502 -58282
rect 39433 -60342 39476 -58367
rect 39760 -58790 39836 -58086
rect 40062 -58042 41849 -58004
rect 40062 -58420 40100 -58042
rect 41269 -58341 41934 -58313
rect 41269 -58399 42304 -58341
rect 40039 -58474 40112 -58420
rect 41269 -58480 41355 -58399
rect 41529 -58436 41564 -58399
rect 41854 -58402 42304 -58399
rect 40417 -58566 41355 -58480
rect 40265 -58790 40395 -58764
rect 39760 -58856 40395 -58790
rect 40557 -58822 40591 -58566
rect 40655 -58822 40689 -58614
rect 40753 -58822 40787 -58566
rect 40851 -58788 40885 -58614
rect 41432 -58744 41466 -58436
rect 41530 -58744 41564 -58436
rect 41628 -58744 41662 -58436
rect 41726 -58744 41760 -58436
rect 41824 -58744 41858 -58436
rect 41400 -58787 41471 -58786
rect 41812 -58787 41886 -58781
rect 41400 -58788 41886 -58787
rect 40851 -58822 41886 -58788
rect 42243 -58809 42304 -58402
rect 45734 -56772 45768 -56428
rect 45930 -56772 45964 -56428
rect 46343 -56535 46377 -56427
rect 46539 -56535 46573 -56427
rect 46225 -56582 46298 -56569
rect 46125 -56610 46298 -56582
rect 46103 -56623 46298 -56610
rect 46103 -56772 46164 -56623
rect 46225 -56629 46298 -56623
rect 46735 -56599 46769 -56427
rect 45734 -56802 46164 -56772
rect 45734 -56810 46153 -56802
rect 46343 -56814 46377 -56658
rect 46441 -56766 46475 -56658
rect 46539 -56814 46573 -56658
rect 46637 -56766 46671 -56658
rect 46735 -56669 47013 -56599
rect 45378 -56883 45605 -56881
rect 46016 -56883 46090 -56857
rect 45378 -56921 46090 -56883
rect 46203 -56900 46818 -56814
rect 40852 -58826 41886 -58822
rect 40852 -58828 41401 -58826
rect 40439 -58856 40512 -58850
rect 41812 -58852 41886 -58826
rect 39760 -58866 40512 -58856
rect 40265 -58897 40512 -58866
rect 41347 -58884 41482 -58876
rect 41327 -58886 41482 -58884
rect 40265 -58914 40395 -58897
rect 40439 -58910 40512 -58897
rect 40292 -58964 40368 -58914
rect 41120 -58922 41482 -58886
rect 41999 -58895 42784 -58809
rect 41327 -58924 41482 -58922
rect 41347 -58930 41482 -58924
rect 41530 -58907 41949 -58899
rect 41530 -58937 41960 -58907
rect 40557 -59152 40591 -58944
rect 40753 -59152 40787 -58944
rect 40949 -59152 40983 -58944
rect 41530 -59281 41564 -58937
rect 41726 -59281 41760 -58937
rect 41899 -59086 41960 -58937
rect 42139 -59051 42173 -58895
rect 42237 -59051 42271 -58943
rect 42335 -59051 42369 -58895
rect 42433 -59051 42467 -58943
rect 42021 -59086 42094 -59080
rect 41899 -59099 42094 -59086
rect 41921 -59127 42094 -59099
rect 42021 -59140 42094 -59127
rect 42531 -59110 42903 -59040
rect 42139 -59282 42173 -59174
rect 42335 -59282 42369 -59174
rect 42531 -59282 42565 -59110
rect 40531 -60217 40565 -59873
rect 40727 -60217 40761 -59873
rect 41140 -59980 41174 -59872
rect 41336 -59980 41370 -59872
rect 41022 -60027 41095 -60014
rect 40922 -60055 41095 -60027
rect 40900 -60068 41095 -60055
rect 40900 -60217 40961 -60068
rect 41022 -60074 41095 -60068
rect 41532 -60044 41566 -59872
rect 40531 -60247 40961 -60217
rect 40531 -60255 40950 -60247
rect 41140 -60259 41174 -60103
rect 41238 -60211 41272 -60103
rect 41336 -60259 41370 -60103
rect 41434 -60211 41468 -60103
rect 41532 -60114 41810 -60044
rect 39433 -60385 39718 -60342
rect 39154 -60488 39259 -60416
rect 39675 -60591 39718 -60385
rect 37187 -60739 37637 -60721
rect 36745 -60782 37637 -60739
rect 36745 -60800 37194 -60782
rect 37576 -61077 37637 -60782
rect 38310 -60959 38344 -60665
rect 38402 -60681 38447 -60611
rect 38794 -60631 39718 -60591
rect 38842 -60634 39718 -60631
rect 38303 -61077 38350 -60959
rect 38408 -60973 38442 -60681
rect 38506 -60958 38540 -60665
rect 38748 -60948 38782 -60665
rect 38842 -60674 38886 -60634
rect 38499 -61077 38546 -60958
rect 38741 -61077 38788 -60948
rect 38846 -60973 38880 -60674
rect 37576 -61190 39053 -61077
rect 40175 -60328 40402 -60326
rect 40813 -60328 40887 -60302
rect 40175 -60366 40887 -60328
rect 41000 -60345 41615 -60259
rect 40401 -60367 40887 -60366
rect 40401 -60368 40472 -60367
rect 40813 -60373 40887 -60367
rect 40433 -60718 40467 -60410
rect 40531 -60718 40565 -60410
rect 40629 -60718 40663 -60410
rect 40727 -60718 40761 -60410
rect 40825 -60718 40859 -60410
rect 40530 -60770 40565 -60718
rect 41244 -60752 41305 -60345
rect 41734 -60509 41804 -60114
rect 41978 -60368 42012 -59784
rect 42185 -59750 42425 -59716
rect 42185 -59792 42227 -59750
rect 41974 -60427 42016 -60368
rect 42189 -60374 42223 -59792
rect 42287 -60372 42321 -59784
rect 42383 -59794 42425 -59750
rect 42186 -60427 42228 -60374
rect 41974 -60463 42228 -60427
rect 42283 -60426 42325 -60372
rect 42385 -60392 42419 -59794
rect 42597 -60378 42631 -59784
rect 42283 -60465 42424 -60426
rect 42381 -60477 42424 -60465
rect 42139 -60509 42294 -60499
rect 41734 -60545 42294 -60509
rect 41734 -60547 41804 -60545
rect 42139 -60554 42294 -60545
rect 42381 -60532 42562 -60477
rect 42381 -60602 42424 -60532
rect 41869 -60616 42024 -60607
rect 41832 -60650 42024 -60616
rect 41869 -60662 42024 -60650
rect 42070 -60642 42424 -60602
rect 42596 -60622 42639 -60378
rect 42833 -60447 42903 -59110
rect 42822 -60519 42927 -60447
rect 43337 -60622 43674 -60459
rect 40855 -60770 41305 -60752
rect 40413 -60813 41305 -60770
rect 40413 -60831 40862 -60813
rect 41244 -61108 41305 -60813
rect 41978 -60990 42012 -60696
rect 42070 -60712 42115 -60642
rect 42462 -60662 43674 -60622
rect 42510 -60665 43674 -60662
rect 41971 -61108 42018 -60990
rect 42076 -61004 42110 -60712
rect 42174 -60989 42208 -60696
rect 42416 -60979 42450 -60696
rect 42510 -60705 42554 -60665
rect 42167 -61108 42214 -60989
rect 42409 -61108 42456 -60979
rect 42514 -61004 42548 -60705
rect 43337 -60790 43674 -60665
rect 41244 -61221 42721 -61108
rect 35847 -62008 36050 -61861
rect 42978 -62042 43295 -61751
rect 42995 -62822 43261 -62042
rect 45389 -57859 45465 -56921
rect 45604 -56922 46090 -56921
rect 45604 -56923 45675 -56922
rect 46016 -56928 46090 -56922
rect 45636 -57273 45670 -56965
rect 45734 -57273 45768 -56965
rect 45832 -57273 45866 -56965
rect 45930 -57273 45964 -56965
rect 46028 -57273 46062 -56965
rect 45733 -57325 45768 -57273
rect 46447 -57307 46508 -56900
rect 46937 -57064 47007 -56669
rect 47181 -56923 47215 -56339
rect 47388 -56305 47628 -56271
rect 47388 -56347 47430 -56305
rect 47177 -56982 47219 -56923
rect 47392 -56929 47426 -56347
rect 47490 -56927 47524 -56339
rect 47586 -56349 47628 -56305
rect 47389 -56982 47431 -56929
rect 47177 -57018 47431 -56982
rect 47486 -56981 47528 -56927
rect 47588 -56947 47622 -56349
rect 47800 -56933 47834 -56339
rect 47486 -57020 47627 -56981
rect 47584 -57032 47627 -57020
rect 47342 -57064 47497 -57054
rect 46937 -57100 47497 -57064
rect 46937 -57102 47007 -57100
rect 47342 -57109 47497 -57100
rect 47584 -57087 47765 -57032
rect 47584 -57157 47627 -57087
rect 47072 -57171 47227 -57162
rect 47035 -57205 47227 -57171
rect 47072 -57217 47227 -57205
rect 47273 -57197 47627 -57157
rect 47799 -57177 47842 -56933
rect 48036 -57002 48106 -55665
rect 54958 -55673 54992 -55465
rect 55154 -55673 55188 -55465
rect 55350 -55673 55384 -55465
rect 55931 -55802 55965 -55458
rect 56127 -55802 56161 -55458
rect 56300 -55607 56361 -55458
rect 56540 -55572 56574 -55416
rect 56638 -55572 56672 -55464
rect 56736 -55572 56770 -55416
rect 56834 -55572 56868 -55464
rect 56422 -55607 56495 -55601
rect 56300 -55620 56495 -55607
rect 56322 -55648 56495 -55620
rect 56422 -55661 56495 -55648
rect 56932 -55631 57304 -55561
rect 56540 -55803 56574 -55695
rect 56736 -55803 56770 -55695
rect 56932 -55803 56966 -55631
rect 49173 -56697 49207 -56197
rect 49352 -56161 49673 -56127
rect 49172 -56743 49207 -56697
rect 49352 -56743 49392 -56161
rect 49441 -56201 49476 -56161
rect 49442 -56705 49476 -56201
rect 49540 -56698 49574 -56197
rect 49638 -56200 49673 -56161
rect 49172 -56783 49392 -56743
rect 49537 -56818 49575 -56698
rect 49638 -56705 49672 -56200
rect 49768 -56781 49802 -56197
rect 50094 -56711 50128 -56197
rect 50322 -56487 50356 -56197
rect 50321 -56580 50358 -56487
rect 50321 -56617 50458 -56580
rect 50094 -56745 50253 -56711
rect 49917 -56781 50055 -56770
rect 49173 -56856 49575 -56818
rect 49642 -56815 50055 -56781
rect 48936 -56867 49074 -56857
rect 48546 -56901 49074 -56867
rect 48025 -57074 48130 -57002
rect 48546 -57177 48589 -56901
rect 48936 -56911 49074 -56901
rect 48992 -57002 49130 -56993
rect 48782 -57036 49130 -57002
rect 48782 -57163 48854 -57036
rect 48992 -57047 49130 -57036
rect 48782 -57172 48866 -57163
rect 46058 -57325 46508 -57307
rect 45616 -57368 46508 -57325
rect 45616 -57386 46065 -57368
rect 46447 -57663 46508 -57368
rect 47181 -57545 47215 -57251
rect 47273 -57267 47318 -57197
rect 47665 -57217 48589 -57177
rect 47713 -57220 48589 -57217
rect 47174 -57663 47221 -57545
rect 47279 -57559 47313 -57267
rect 47377 -57544 47411 -57251
rect 47619 -57534 47653 -57251
rect 47713 -57260 47757 -57220
rect 48787 -57242 48866 -57172
rect 47370 -57663 47417 -57544
rect 47612 -57663 47659 -57534
rect 47717 -57559 47751 -57260
rect 49075 -57484 49109 -57193
rect 49073 -57595 49110 -57484
rect 49173 -57501 49207 -56856
rect 49402 -56926 49440 -56856
rect 49642 -56894 49676 -56815
rect 49917 -56824 50055 -56815
rect 49392 -57064 49446 -56926
rect 49545 -56928 49676 -56894
rect 49742 -56911 49880 -56857
rect 50127 -56926 50181 -56788
rect 50219 -56789 50253 -56745
rect 50219 -56843 50385 -56789
rect 49545 -57501 49579 -56928
rect 50219 -56958 50253 -56843
rect 50305 -56958 50359 -56941
rect 49643 -56997 49802 -56962
rect 50219 -56963 50359 -56958
rect 50191 -56992 50359 -56963
rect 49643 -57501 49677 -56997
rect 49768 -57501 49802 -56997
rect 49866 -57484 49900 -56993
rect 49996 -57483 50030 -56993
rect 48536 -57599 49147 -57595
rect 49865 -57599 49902 -57484
rect 49993 -57599 50030 -57483
rect 50094 -57501 50128 -56993
rect 50191 -56997 50253 -56992
rect 50192 -57501 50226 -56997
rect 50305 -57000 50359 -56992
rect 50420 -57110 50458 -56617
rect 50420 -57148 50712 -57110
rect 50322 -57482 50356 -57193
rect 50420 -57198 50458 -57148
rect 50320 -57599 50357 -57482
rect 50420 -57501 50454 -57198
rect 48536 -57663 50470 -57599
rect 46447 -57708 50470 -57663
rect 46447 -57776 48649 -57708
rect 48997 -57760 50470 -57708
rect 44739 -58005 45465 -57859
rect 44739 -62006 44885 -58005
rect 45389 -58049 45465 -58005
rect 50674 -58043 50712 -57148
rect 45389 -58125 48699 -58049
rect 45389 -58307 45465 -58125
rect 45389 -58383 45531 -58307
rect 45455 -58772 45531 -58383
rect 46464 -58349 47129 -58321
rect 46464 -58407 47499 -58349
rect 46464 -58488 46550 -58407
rect 46724 -58444 46759 -58407
rect 47049 -58410 47499 -58407
rect 45612 -58574 46550 -58488
rect 45455 -58864 45590 -58772
rect 45752 -58830 45786 -58574
rect 45850 -58830 45884 -58622
rect 45948 -58830 45982 -58574
rect 46046 -58796 46080 -58622
rect 46627 -58752 46661 -58444
rect 46725 -58752 46759 -58444
rect 46823 -58752 46857 -58444
rect 46921 -58752 46955 -58444
rect 47019 -58752 47053 -58444
rect 46595 -58795 46666 -58794
rect 47007 -58795 47081 -58789
rect 46595 -58796 47081 -58795
rect 46046 -58830 47081 -58796
rect 47438 -58817 47499 -58410
rect 46047 -58834 47081 -58830
rect 46047 -58836 46596 -58834
rect 45634 -58864 45707 -58858
rect 47007 -58860 47081 -58834
rect 45455 -58881 45707 -58864
rect 45460 -58905 45707 -58881
rect 46542 -58892 46677 -58884
rect 46522 -58894 46677 -58892
rect 45460 -58922 45590 -58905
rect 45634 -58918 45707 -58905
rect 46315 -58930 46677 -58894
rect 47194 -58903 47979 -58817
rect 46522 -58932 46677 -58930
rect 46542 -58938 46677 -58932
rect 46725 -58915 47144 -58907
rect 46725 -58945 47155 -58915
rect 45752 -59160 45786 -58952
rect 45948 -59160 45982 -58952
rect 46144 -59160 46178 -58952
rect 46725 -59289 46759 -58945
rect 46921 -59289 46955 -58945
rect 47094 -59094 47155 -58945
rect 47334 -59059 47368 -58903
rect 47432 -59059 47466 -58951
rect 47530 -59059 47564 -58903
rect 47628 -59059 47662 -58951
rect 47216 -59094 47289 -59088
rect 47094 -59107 47289 -59094
rect 47116 -59135 47289 -59107
rect 47216 -59148 47289 -59135
rect 47726 -59118 48098 -59048
rect 47334 -59290 47368 -59182
rect 47530 -59290 47564 -59182
rect 47726 -59290 47760 -59118
rect 45726 -60225 45760 -59881
rect 45922 -60225 45956 -59881
rect 46335 -59988 46369 -59880
rect 46531 -59988 46565 -59880
rect 46217 -60035 46290 -60022
rect 46117 -60063 46290 -60035
rect 46095 -60076 46290 -60063
rect 46095 -60225 46156 -60076
rect 46217 -60082 46290 -60076
rect 46727 -60052 46761 -59880
rect 45726 -60255 46156 -60225
rect 45726 -60263 46145 -60255
rect 46335 -60267 46369 -60111
rect 46433 -60219 46467 -60111
rect 46531 -60267 46565 -60111
rect 46629 -60219 46663 -60111
rect 46727 -60122 47005 -60052
rect 45370 -60336 45597 -60334
rect 46008 -60336 46082 -60310
rect 45370 -60374 46082 -60336
rect 46195 -60353 46810 -60267
rect 45596 -60375 46082 -60374
rect 45596 -60376 45667 -60375
rect 46008 -60381 46082 -60375
rect 45628 -60726 45662 -60418
rect 45726 -60726 45760 -60418
rect 45824 -60726 45858 -60418
rect 45922 -60726 45956 -60418
rect 46020 -60726 46054 -60418
rect 45725 -60778 45760 -60726
rect 46439 -60760 46500 -60353
rect 46929 -60517 46999 -60122
rect 47173 -60376 47207 -59792
rect 47380 -59758 47620 -59724
rect 47380 -59800 47422 -59758
rect 47169 -60435 47211 -60376
rect 47384 -60382 47418 -59800
rect 47482 -60380 47516 -59792
rect 47578 -59802 47620 -59758
rect 47381 -60435 47423 -60382
rect 47169 -60471 47423 -60435
rect 47478 -60434 47520 -60380
rect 47580 -60400 47614 -59802
rect 47792 -60386 47826 -59792
rect 47478 -60473 47619 -60434
rect 47576 -60485 47619 -60473
rect 47334 -60517 47489 -60507
rect 46929 -60553 47489 -60517
rect 46929 -60555 46999 -60553
rect 47334 -60562 47489 -60553
rect 47576 -60540 47757 -60485
rect 47576 -60610 47619 -60540
rect 47064 -60624 47219 -60615
rect 47027 -60658 47219 -60624
rect 47064 -60670 47219 -60658
rect 47265 -60650 47619 -60610
rect 47791 -60630 47834 -60386
rect 48028 -60455 48098 -59118
rect 48273 -58406 48365 -58321
rect 48296 -60381 48339 -58406
rect 48623 -58829 48699 -58125
rect 48925 -58081 50712 -58043
rect 48925 -58459 48963 -58081
rect 50132 -58380 50797 -58352
rect 50132 -58438 51167 -58380
rect 48902 -58513 48975 -58459
rect 50132 -58519 50218 -58438
rect 50392 -58475 50427 -58438
rect 50717 -58441 51167 -58438
rect 49280 -58605 50218 -58519
rect 49128 -58829 49258 -58803
rect 48623 -58895 49258 -58829
rect 49420 -58861 49454 -58605
rect 49518 -58861 49552 -58653
rect 49616 -58861 49650 -58605
rect 49714 -58827 49748 -58653
rect 50295 -58783 50329 -58475
rect 50393 -58783 50427 -58475
rect 50491 -58783 50525 -58475
rect 50589 -58783 50623 -58475
rect 50687 -58783 50721 -58475
rect 50263 -58826 50334 -58825
rect 50675 -58826 50749 -58820
rect 50263 -58827 50749 -58826
rect 49714 -58861 50749 -58827
rect 51106 -58848 51167 -58441
rect 54932 -56738 54966 -56394
rect 55128 -56738 55162 -56394
rect 55541 -56501 55575 -56393
rect 55737 -56501 55771 -56393
rect 55423 -56548 55496 -56535
rect 55323 -56576 55496 -56548
rect 55301 -56589 55496 -56576
rect 55301 -56738 55362 -56589
rect 55423 -56595 55496 -56589
rect 55933 -56565 55967 -56393
rect 54932 -56768 55362 -56738
rect 54932 -56776 55351 -56768
rect 55541 -56780 55575 -56624
rect 55639 -56732 55673 -56624
rect 55737 -56780 55771 -56624
rect 55835 -56732 55869 -56624
rect 55933 -56635 56211 -56565
rect 49715 -58865 50749 -58861
rect 49715 -58867 50264 -58865
rect 49302 -58895 49375 -58889
rect 50675 -58891 50749 -58865
rect 48623 -58905 49375 -58895
rect 49128 -58936 49375 -58905
rect 50210 -58923 50345 -58915
rect 50190 -58925 50345 -58923
rect 49128 -58953 49258 -58936
rect 49302 -58949 49375 -58936
rect 49155 -59003 49231 -58953
rect 49983 -58961 50345 -58925
rect 50862 -58934 51647 -58848
rect 50190 -58963 50345 -58961
rect 50210 -58969 50345 -58963
rect 50393 -58946 50812 -58938
rect 50393 -58976 50823 -58946
rect 49420 -59191 49454 -58983
rect 49616 -59191 49650 -58983
rect 49812 -59191 49846 -58983
rect 50393 -59320 50427 -58976
rect 50589 -59320 50623 -58976
rect 50762 -59125 50823 -58976
rect 51002 -59090 51036 -58934
rect 51100 -59090 51134 -58982
rect 51198 -59090 51232 -58934
rect 51296 -59090 51330 -58982
rect 50884 -59125 50957 -59119
rect 50762 -59138 50957 -59125
rect 50784 -59166 50957 -59138
rect 50884 -59179 50957 -59166
rect 51394 -59149 51766 -59079
rect 51002 -59321 51036 -59213
rect 51198 -59321 51232 -59213
rect 51394 -59321 51428 -59149
rect 49394 -60256 49428 -59912
rect 49590 -60256 49624 -59912
rect 50003 -60019 50037 -59911
rect 50199 -60019 50233 -59911
rect 49885 -60066 49958 -60053
rect 49785 -60094 49958 -60066
rect 49763 -60107 49958 -60094
rect 49763 -60256 49824 -60107
rect 49885 -60113 49958 -60107
rect 50395 -60083 50429 -59911
rect 49394 -60286 49824 -60256
rect 49394 -60294 49813 -60286
rect 50003 -60298 50037 -60142
rect 50101 -60250 50135 -60142
rect 50199 -60298 50233 -60142
rect 50297 -60250 50331 -60142
rect 50395 -60153 50673 -60083
rect 48296 -60424 48581 -60381
rect 48017 -60527 48122 -60455
rect 48538 -60630 48581 -60424
rect 46050 -60778 46500 -60760
rect 45608 -60821 46500 -60778
rect 45608 -60839 46057 -60821
rect 46439 -61116 46500 -60821
rect 47173 -60998 47207 -60704
rect 47265 -60720 47310 -60650
rect 47657 -60670 48581 -60630
rect 47705 -60673 48581 -60670
rect 47166 -61116 47213 -60998
rect 47271 -61012 47305 -60720
rect 47369 -60997 47403 -60704
rect 47611 -60987 47645 -60704
rect 47705 -60713 47749 -60673
rect 47362 -61116 47409 -60997
rect 47604 -61116 47651 -60987
rect 47709 -61012 47743 -60713
rect 46439 -61229 47916 -61116
rect 49038 -60367 49265 -60365
rect 49676 -60367 49750 -60341
rect 49038 -60405 49750 -60367
rect 49863 -60384 50478 -60298
rect 49264 -60406 49750 -60405
rect 49264 -60407 49335 -60406
rect 49676 -60412 49750 -60406
rect 49296 -60757 49330 -60449
rect 49394 -60757 49428 -60449
rect 49492 -60757 49526 -60449
rect 49590 -60757 49624 -60449
rect 49688 -60757 49722 -60449
rect 49393 -60809 49428 -60757
rect 50107 -60791 50168 -60384
rect 50597 -60548 50667 -60153
rect 50841 -60407 50875 -59823
rect 51048 -59789 51288 -59755
rect 51048 -59831 51090 -59789
rect 50837 -60466 50879 -60407
rect 51052 -60413 51086 -59831
rect 51150 -60411 51184 -59823
rect 51246 -59833 51288 -59789
rect 51049 -60466 51091 -60413
rect 50837 -60502 51091 -60466
rect 51146 -60465 51188 -60411
rect 51248 -60431 51282 -59833
rect 51460 -60417 51494 -59823
rect 51146 -60504 51287 -60465
rect 51244 -60516 51287 -60504
rect 51002 -60548 51157 -60538
rect 50597 -60584 51157 -60548
rect 50597 -60586 50667 -60584
rect 51002 -60593 51157 -60584
rect 51244 -60571 51425 -60516
rect 51244 -60641 51287 -60571
rect 50732 -60655 50887 -60646
rect 50695 -60689 50887 -60655
rect 50732 -60701 50887 -60689
rect 50933 -60681 51287 -60641
rect 51459 -60661 51502 -60417
rect 51696 -60486 51766 -59149
rect 51685 -60558 51790 -60486
rect 52215 -60661 52429 -60546
rect 49718 -60809 50168 -60791
rect 49276 -60852 50168 -60809
rect 49276 -60870 49725 -60852
rect 50107 -61147 50168 -60852
rect 50841 -61029 50875 -60735
rect 50933 -60751 50978 -60681
rect 51325 -60701 52527 -60661
rect 51373 -60704 52527 -60701
rect 50834 -61147 50881 -61029
rect 50939 -61043 50973 -60751
rect 51037 -61028 51071 -60735
rect 51279 -61018 51313 -60735
rect 51373 -60744 51417 -60704
rect 51030 -61147 51077 -61028
rect 51272 -61147 51319 -61018
rect 51377 -61043 51411 -60744
rect 52215 -60766 52429 -60704
rect 50107 -61260 51584 -61147
rect 43012 -62831 43252 -62822
rect 54576 -56849 54803 -56847
rect 55214 -56849 55288 -56823
rect 54576 -56887 55288 -56849
rect 55401 -56866 56016 -56780
rect 54587 -57758 54663 -56887
rect 54802 -56888 55288 -56887
rect 54802 -56889 54873 -56888
rect 55214 -56894 55288 -56888
rect 54834 -57239 54868 -56931
rect 54932 -57239 54966 -56931
rect 55030 -57239 55064 -56931
rect 55128 -57239 55162 -56931
rect 55226 -57239 55260 -56931
rect 54931 -57291 54966 -57239
rect 55645 -57273 55706 -56866
rect 56135 -57030 56205 -56635
rect 56379 -56889 56413 -56305
rect 56586 -56271 56826 -56237
rect 56586 -56313 56628 -56271
rect 56375 -56948 56417 -56889
rect 56590 -56895 56624 -56313
rect 56688 -56893 56722 -56305
rect 56784 -56315 56826 -56271
rect 56587 -56948 56629 -56895
rect 56375 -56984 56629 -56948
rect 56684 -56947 56726 -56893
rect 56786 -56913 56820 -56315
rect 56998 -56899 57032 -56305
rect 56684 -56986 56825 -56947
rect 56782 -56998 56825 -56986
rect 56540 -57030 56695 -57020
rect 56135 -57066 56695 -57030
rect 56135 -57068 56205 -57066
rect 56540 -57075 56695 -57066
rect 56782 -57053 56963 -56998
rect 56782 -57123 56825 -57053
rect 56270 -57137 56425 -57128
rect 56233 -57171 56425 -57137
rect 56270 -57183 56425 -57171
rect 56471 -57163 56825 -57123
rect 56997 -57143 57040 -56899
rect 57234 -56968 57304 -55631
rect 63712 -55607 63746 -55399
rect 63908 -55607 63942 -55399
rect 64104 -55607 64138 -55399
rect 64685 -55736 64719 -55392
rect 64881 -55736 64915 -55392
rect 65054 -55541 65115 -55392
rect 65294 -55506 65328 -55350
rect 65392 -55506 65426 -55398
rect 65490 -55506 65524 -55350
rect 72573 -55352 72703 -55335
rect 72747 -55348 72820 -55335
rect 73428 -55360 73790 -55324
rect 74307 -55333 75092 -55247
rect 81937 -55256 82067 -55164
rect 82229 -55222 82263 -54966
rect 82327 -55222 82361 -55014
rect 82425 -55222 82459 -54966
rect 82523 -55188 82557 -55014
rect 83104 -55144 83138 -54836
rect 83202 -55144 83236 -54836
rect 83300 -55144 83334 -54836
rect 83398 -55144 83432 -54836
rect 83496 -55144 83530 -54836
rect 83072 -55187 83143 -55186
rect 83484 -55187 83558 -55181
rect 83072 -55188 83558 -55187
rect 82523 -55222 83558 -55188
rect 83915 -55209 83976 -54802
rect 82524 -55226 83558 -55222
rect 82524 -55228 83073 -55226
rect 82111 -55256 82184 -55250
rect 83484 -55252 83558 -55226
rect 81937 -55297 82184 -55256
rect 83019 -55284 83154 -55276
rect 82999 -55286 83154 -55284
rect 81937 -55314 82067 -55297
rect 82111 -55310 82184 -55297
rect 82792 -55322 83154 -55286
rect 83671 -55295 84456 -55209
rect 82999 -55324 83154 -55322
rect 83019 -55330 83154 -55324
rect 83202 -55307 83621 -55299
rect 73635 -55362 73790 -55360
rect 73655 -55368 73790 -55362
rect 73838 -55345 74257 -55337
rect 73838 -55375 74268 -55345
rect 65588 -55506 65622 -55398
rect 65176 -55541 65249 -55535
rect 65054 -55554 65249 -55541
rect 65076 -55582 65249 -55554
rect 65176 -55595 65249 -55582
rect 65686 -55565 66058 -55495
rect 65294 -55737 65328 -55629
rect 65490 -55737 65524 -55629
rect 65686 -55737 65720 -55565
rect 58371 -56663 58405 -56163
rect 58550 -56127 58871 -56093
rect 58370 -56709 58405 -56663
rect 58550 -56709 58590 -56127
rect 58639 -56167 58674 -56127
rect 58640 -56671 58674 -56167
rect 58738 -56664 58772 -56163
rect 58836 -56166 58871 -56127
rect 58370 -56749 58590 -56709
rect 58735 -56784 58773 -56664
rect 58836 -56671 58870 -56166
rect 58966 -56747 59000 -56163
rect 59292 -56677 59326 -56163
rect 59520 -56453 59554 -56163
rect 59519 -56546 59556 -56453
rect 59519 -56583 59656 -56546
rect 59292 -56711 59451 -56677
rect 59115 -56747 59253 -56736
rect 58371 -56822 58773 -56784
rect 58840 -56781 59253 -56747
rect 58134 -56833 58272 -56823
rect 57744 -56867 58272 -56833
rect 57223 -57040 57328 -56968
rect 57744 -57143 57787 -56867
rect 58134 -56877 58272 -56867
rect 58190 -56968 58328 -56959
rect 57980 -57002 58328 -56968
rect 57980 -57129 58052 -57002
rect 58190 -57013 58328 -57002
rect 57980 -57138 58064 -57129
rect 55256 -57291 55706 -57273
rect 54814 -57334 55706 -57291
rect 54814 -57352 55263 -57334
rect 55645 -57629 55706 -57334
rect 56379 -57511 56413 -57217
rect 56471 -57233 56516 -57163
rect 56863 -57183 57787 -57143
rect 56911 -57186 57787 -57183
rect 56372 -57629 56419 -57511
rect 56477 -57525 56511 -57233
rect 56575 -57510 56609 -57217
rect 56817 -57500 56851 -57217
rect 56911 -57226 56955 -57186
rect 57985 -57208 58064 -57138
rect 56568 -57629 56615 -57510
rect 56810 -57629 56857 -57500
rect 56915 -57525 56949 -57226
rect 58273 -57450 58307 -57159
rect 58271 -57561 58308 -57450
rect 58371 -57467 58405 -56822
rect 58600 -56892 58638 -56822
rect 58840 -56860 58874 -56781
rect 59115 -56790 59253 -56781
rect 58590 -57030 58644 -56892
rect 58743 -56894 58874 -56860
rect 58940 -56877 59078 -56823
rect 59325 -56892 59379 -56754
rect 59417 -56755 59451 -56711
rect 59417 -56809 59583 -56755
rect 58743 -57467 58777 -56894
rect 59417 -56924 59451 -56809
rect 59503 -56924 59557 -56907
rect 58841 -56963 59000 -56928
rect 59417 -56929 59557 -56924
rect 59389 -56958 59557 -56929
rect 58841 -57467 58875 -56963
rect 58966 -57467 59000 -56963
rect 59064 -57450 59098 -56959
rect 59194 -57449 59228 -56959
rect 57734 -57565 58345 -57561
rect 59063 -57565 59100 -57450
rect 59191 -57565 59228 -57449
rect 59292 -57467 59326 -56959
rect 59389 -56963 59451 -56958
rect 59390 -57467 59424 -56963
rect 59503 -56966 59557 -56958
rect 59618 -57076 59656 -56583
rect 59618 -57114 59910 -57076
rect 59520 -57448 59554 -57159
rect 59618 -57164 59656 -57114
rect 59518 -57565 59555 -57448
rect 59618 -57467 59652 -57164
rect 57734 -57629 59668 -57565
rect 55645 -57674 59668 -57629
rect 55645 -57742 57847 -57674
rect 58195 -57726 59668 -57674
rect 53876 -57919 54663 -57758
rect 53876 -61840 54037 -57919
rect 54587 -58015 54663 -57919
rect 59872 -58009 59910 -57114
rect 54587 -58091 57897 -58015
rect 54587 -58273 54663 -58091
rect 54587 -58349 54729 -58273
rect 54653 -58738 54729 -58349
rect 55662 -58315 56327 -58287
rect 55662 -58373 56697 -58315
rect 55662 -58454 55748 -58373
rect 55922 -58410 55957 -58373
rect 56247 -58376 56697 -58373
rect 54810 -58540 55748 -58454
rect 54653 -58830 54788 -58738
rect 54950 -58796 54984 -58540
rect 55048 -58796 55082 -58588
rect 55146 -58796 55180 -58540
rect 55244 -58762 55278 -58588
rect 55825 -58718 55859 -58410
rect 55923 -58718 55957 -58410
rect 56021 -58718 56055 -58410
rect 56119 -58718 56153 -58410
rect 56217 -58718 56251 -58410
rect 55793 -58761 55864 -58760
rect 56205 -58761 56279 -58755
rect 55793 -58762 56279 -58761
rect 55244 -58796 56279 -58762
rect 56636 -58783 56697 -58376
rect 55245 -58800 56279 -58796
rect 55245 -58802 55794 -58800
rect 54832 -58830 54905 -58824
rect 56205 -58826 56279 -58800
rect 54653 -58847 54905 -58830
rect 54658 -58871 54905 -58847
rect 55740 -58858 55875 -58850
rect 55720 -58860 55875 -58858
rect 54658 -58888 54788 -58871
rect 54832 -58884 54905 -58871
rect 55513 -58896 55875 -58860
rect 56392 -58869 57177 -58783
rect 55720 -58898 55875 -58896
rect 55740 -58904 55875 -58898
rect 55923 -58881 56342 -58873
rect 55923 -58911 56353 -58881
rect 54950 -59126 54984 -58918
rect 55146 -59126 55180 -58918
rect 55342 -59126 55376 -58918
rect 55923 -59255 55957 -58911
rect 56119 -59255 56153 -58911
rect 56292 -59060 56353 -58911
rect 56532 -59025 56566 -58869
rect 56630 -59025 56664 -58917
rect 56728 -59025 56762 -58869
rect 56826 -59025 56860 -58917
rect 56414 -59060 56487 -59054
rect 56292 -59073 56487 -59060
rect 56314 -59101 56487 -59073
rect 56414 -59114 56487 -59101
rect 56924 -59084 57296 -59014
rect 56532 -59256 56566 -59148
rect 56728 -59256 56762 -59148
rect 56924 -59256 56958 -59084
rect 54924 -60191 54958 -59847
rect 55120 -60191 55154 -59847
rect 55533 -59954 55567 -59846
rect 55729 -59954 55763 -59846
rect 55415 -60001 55488 -59988
rect 55315 -60029 55488 -60001
rect 55293 -60042 55488 -60029
rect 55293 -60191 55354 -60042
rect 55415 -60048 55488 -60042
rect 55925 -60018 55959 -59846
rect 54924 -60221 55354 -60191
rect 54924 -60229 55343 -60221
rect 55533 -60233 55567 -60077
rect 55631 -60185 55665 -60077
rect 55729 -60233 55763 -60077
rect 55827 -60185 55861 -60077
rect 55925 -60088 56203 -60018
rect 54568 -60302 54795 -60300
rect 55206 -60302 55280 -60276
rect 54568 -60340 55280 -60302
rect 55393 -60319 56008 -60233
rect 54794 -60341 55280 -60340
rect 54794 -60342 54865 -60341
rect 55206 -60347 55280 -60341
rect 54826 -60692 54860 -60384
rect 54924 -60692 54958 -60384
rect 55022 -60692 55056 -60384
rect 55120 -60692 55154 -60384
rect 55218 -60692 55252 -60384
rect 54923 -60744 54958 -60692
rect 55637 -60726 55698 -60319
rect 56127 -60483 56197 -60088
rect 56371 -60342 56405 -59758
rect 56578 -59724 56818 -59690
rect 56578 -59766 56620 -59724
rect 56367 -60401 56409 -60342
rect 56582 -60348 56616 -59766
rect 56680 -60346 56714 -59758
rect 56776 -59768 56818 -59724
rect 56579 -60401 56621 -60348
rect 56367 -60437 56621 -60401
rect 56676 -60400 56718 -60346
rect 56778 -60366 56812 -59768
rect 56990 -60352 57024 -59758
rect 56676 -60439 56817 -60400
rect 56774 -60451 56817 -60439
rect 56532 -60483 56687 -60473
rect 56127 -60519 56687 -60483
rect 56127 -60521 56197 -60519
rect 56532 -60528 56687 -60519
rect 56774 -60506 56955 -60451
rect 56774 -60576 56817 -60506
rect 56262 -60590 56417 -60581
rect 56225 -60624 56417 -60590
rect 56262 -60636 56417 -60624
rect 56463 -60616 56817 -60576
rect 56989 -60596 57032 -60352
rect 57226 -60421 57296 -59084
rect 57471 -58372 57563 -58287
rect 57494 -60347 57537 -58372
rect 57821 -58795 57897 -58091
rect 58123 -58047 59910 -58009
rect 58123 -58425 58161 -58047
rect 59330 -58346 59995 -58318
rect 59330 -58404 60365 -58346
rect 58100 -58479 58173 -58425
rect 59330 -58485 59416 -58404
rect 59590 -58441 59625 -58404
rect 59915 -58407 60365 -58404
rect 58478 -58571 59416 -58485
rect 58326 -58795 58456 -58769
rect 57821 -58861 58456 -58795
rect 58618 -58827 58652 -58571
rect 58716 -58827 58750 -58619
rect 58814 -58827 58848 -58571
rect 58912 -58793 58946 -58619
rect 59493 -58749 59527 -58441
rect 59591 -58749 59625 -58441
rect 59689 -58749 59723 -58441
rect 59787 -58749 59821 -58441
rect 59885 -58749 59919 -58441
rect 59461 -58792 59532 -58791
rect 59873 -58792 59947 -58786
rect 59461 -58793 59947 -58792
rect 58912 -58827 59947 -58793
rect 60304 -58814 60365 -58407
rect 63686 -56672 63720 -56328
rect 63882 -56672 63916 -56328
rect 64295 -56435 64329 -56327
rect 64491 -56435 64525 -56327
rect 64177 -56482 64250 -56469
rect 64077 -56510 64250 -56482
rect 64055 -56523 64250 -56510
rect 64055 -56672 64116 -56523
rect 64177 -56529 64250 -56523
rect 64687 -56499 64721 -56327
rect 63686 -56702 64116 -56672
rect 63686 -56710 64105 -56702
rect 64295 -56714 64329 -56558
rect 64393 -56666 64427 -56558
rect 64491 -56714 64525 -56558
rect 64589 -56666 64623 -56558
rect 64687 -56569 64965 -56499
rect 63330 -56783 63557 -56781
rect 63968 -56783 64042 -56757
rect 58913 -58831 59947 -58827
rect 58913 -58833 59462 -58831
rect 58500 -58861 58573 -58855
rect 59873 -58857 59947 -58831
rect 57821 -58871 58573 -58861
rect 58326 -58902 58573 -58871
rect 59408 -58889 59543 -58881
rect 59388 -58891 59543 -58889
rect 58326 -58919 58456 -58902
rect 58500 -58915 58573 -58902
rect 58353 -58969 58429 -58919
rect 59181 -58927 59543 -58891
rect 60060 -58900 60845 -58814
rect 59388 -58929 59543 -58927
rect 59408 -58935 59543 -58929
rect 59591 -58912 60010 -58904
rect 59591 -58942 60021 -58912
rect 58618 -59157 58652 -58949
rect 58814 -59157 58848 -58949
rect 59010 -59157 59044 -58949
rect 59591 -59286 59625 -58942
rect 59787 -59286 59821 -58942
rect 59960 -59091 60021 -58942
rect 60200 -59056 60234 -58900
rect 60298 -59056 60332 -58948
rect 60396 -59056 60430 -58900
rect 60494 -59056 60528 -58948
rect 60082 -59091 60155 -59085
rect 59960 -59104 60155 -59091
rect 59982 -59132 60155 -59104
rect 60082 -59145 60155 -59132
rect 60592 -59115 60964 -59045
rect 60200 -59287 60234 -59179
rect 60396 -59287 60430 -59179
rect 60592 -59287 60626 -59115
rect 58592 -60222 58626 -59878
rect 58788 -60222 58822 -59878
rect 59201 -59985 59235 -59877
rect 59397 -59985 59431 -59877
rect 59083 -60032 59156 -60019
rect 58983 -60060 59156 -60032
rect 58961 -60073 59156 -60060
rect 58961 -60222 59022 -60073
rect 59083 -60079 59156 -60073
rect 59593 -60049 59627 -59877
rect 58592 -60252 59022 -60222
rect 58592 -60260 59011 -60252
rect 59201 -60264 59235 -60108
rect 59299 -60216 59333 -60108
rect 59397 -60264 59431 -60108
rect 59495 -60216 59529 -60108
rect 59593 -60119 59871 -60049
rect 57494 -60390 57779 -60347
rect 57215 -60493 57320 -60421
rect 57736 -60596 57779 -60390
rect 55248 -60744 55698 -60726
rect 54806 -60787 55698 -60744
rect 54806 -60805 55255 -60787
rect 55637 -61082 55698 -60787
rect 56371 -60964 56405 -60670
rect 56463 -60686 56508 -60616
rect 56855 -60636 57779 -60596
rect 56903 -60639 57779 -60636
rect 56364 -61082 56411 -60964
rect 56469 -60978 56503 -60686
rect 56567 -60963 56601 -60670
rect 56809 -60953 56843 -60670
rect 56903 -60679 56947 -60639
rect 56560 -61082 56607 -60963
rect 56802 -61082 56849 -60953
rect 56907 -60978 56941 -60679
rect 55637 -61195 57114 -61082
rect 58236 -60333 58463 -60331
rect 58874 -60333 58948 -60307
rect 58236 -60371 58948 -60333
rect 59061 -60350 59676 -60264
rect 58462 -60372 58948 -60371
rect 58462 -60373 58533 -60372
rect 58874 -60378 58948 -60372
rect 58494 -60723 58528 -60415
rect 58592 -60723 58626 -60415
rect 58690 -60723 58724 -60415
rect 58788 -60723 58822 -60415
rect 58886 -60723 58920 -60415
rect 58591 -60775 58626 -60723
rect 59305 -60757 59366 -60350
rect 59795 -60514 59865 -60119
rect 60039 -60373 60073 -59789
rect 60246 -59755 60486 -59721
rect 60246 -59797 60288 -59755
rect 60035 -60432 60077 -60373
rect 60250 -60379 60284 -59797
rect 60348 -60377 60382 -59789
rect 60444 -59799 60486 -59755
rect 60247 -60432 60289 -60379
rect 60035 -60468 60289 -60432
rect 60344 -60431 60386 -60377
rect 60446 -60397 60480 -59799
rect 60658 -60383 60692 -59789
rect 60344 -60470 60485 -60431
rect 60442 -60482 60485 -60470
rect 60200 -60514 60355 -60504
rect 59795 -60550 60355 -60514
rect 59795 -60552 59865 -60550
rect 60200 -60559 60355 -60550
rect 60442 -60537 60623 -60482
rect 60442 -60607 60485 -60537
rect 59930 -60621 60085 -60612
rect 59893 -60655 60085 -60621
rect 59930 -60667 60085 -60655
rect 60131 -60647 60485 -60607
rect 60657 -60627 60700 -60383
rect 60894 -60452 60964 -59115
rect 60883 -60524 60988 -60452
rect 61341 -60627 61633 -60458
rect 58916 -60775 59366 -60757
rect 58474 -60818 59366 -60775
rect 58474 -60836 58923 -60818
rect 59305 -61113 59366 -60818
rect 60039 -60995 60073 -60701
rect 60131 -60717 60176 -60647
rect 60523 -60667 61725 -60627
rect 60571 -60670 61725 -60667
rect 60032 -61113 60079 -60995
rect 60137 -61009 60171 -60717
rect 60235 -60994 60269 -60701
rect 60477 -60984 60511 -60701
rect 60571 -60710 60615 -60670
rect 60228 -61113 60275 -60994
rect 60470 -61113 60517 -60984
rect 60575 -61009 60609 -60710
rect 61341 -60757 61633 -60670
rect 59305 -61226 60782 -61113
rect 53858 -62007 54052 -61840
rect 63330 -56821 64042 -56783
rect 64155 -56800 64770 -56714
rect 63341 -57785 63417 -56821
rect 63556 -56822 64042 -56821
rect 63556 -56823 63627 -56822
rect 63968 -56828 64042 -56822
rect 63588 -57173 63622 -56865
rect 63686 -57173 63720 -56865
rect 63784 -57173 63818 -56865
rect 63882 -57173 63916 -56865
rect 63980 -57173 64014 -56865
rect 63685 -57225 63720 -57173
rect 64399 -57207 64460 -56800
rect 64889 -56964 64959 -56569
rect 65133 -56823 65167 -56239
rect 65340 -56205 65580 -56171
rect 65340 -56247 65382 -56205
rect 65129 -56882 65171 -56823
rect 65344 -56829 65378 -56247
rect 65442 -56827 65476 -56239
rect 65538 -56249 65580 -56205
rect 65341 -56882 65383 -56829
rect 65129 -56918 65383 -56882
rect 65438 -56881 65480 -56827
rect 65540 -56847 65574 -56249
rect 65752 -56833 65786 -56239
rect 65438 -56920 65579 -56881
rect 65536 -56932 65579 -56920
rect 65294 -56964 65449 -56954
rect 64889 -57000 65449 -56964
rect 64889 -57002 64959 -57000
rect 65294 -57009 65449 -57000
rect 65536 -56987 65717 -56932
rect 65536 -57057 65579 -56987
rect 65024 -57071 65179 -57062
rect 64987 -57105 65179 -57071
rect 65024 -57117 65179 -57105
rect 65225 -57097 65579 -57057
rect 65751 -57077 65794 -56833
rect 65988 -56902 66058 -55565
rect 72865 -55590 72899 -55382
rect 73061 -55590 73095 -55382
rect 73257 -55590 73291 -55382
rect 73838 -55719 73872 -55375
rect 74034 -55719 74068 -55375
rect 74207 -55524 74268 -55375
rect 74447 -55489 74481 -55333
rect 74545 -55489 74579 -55381
rect 74643 -55489 74677 -55333
rect 83202 -55337 83632 -55307
rect 74741 -55489 74775 -55381
rect 74329 -55524 74402 -55518
rect 74207 -55537 74402 -55524
rect 74229 -55565 74402 -55537
rect 74329 -55578 74402 -55565
rect 74839 -55548 75211 -55478
rect 74447 -55720 74481 -55612
rect 74643 -55720 74677 -55612
rect 74839 -55720 74873 -55548
rect 67125 -56597 67159 -56097
rect 67304 -56061 67625 -56027
rect 67124 -56643 67159 -56597
rect 67304 -56643 67344 -56061
rect 67393 -56101 67428 -56061
rect 67394 -56605 67428 -56101
rect 67492 -56598 67526 -56097
rect 67590 -56100 67625 -56061
rect 67124 -56683 67344 -56643
rect 67489 -56718 67527 -56598
rect 67590 -56605 67624 -56100
rect 67720 -56681 67754 -56097
rect 68046 -56611 68080 -56097
rect 68274 -56387 68308 -56097
rect 68273 -56480 68310 -56387
rect 68273 -56517 68410 -56480
rect 68046 -56645 68205 -56611
rect 67869 -56681 68007 -56670
rect 67125 -56756 67527 -56718
rect 67594 -56715 68007 -56681
rect 66888 -56767 67026 -56757
rect 66498 -56801 67026 -56767
rect 65977 -56974 66082 -56902
rect 66498 -57077 66541 -56801
rect 66888 -56811 67026 -56801
rect 66944 -56902 67082 -56893
rect 66734 -56936 67082 -56902
rect 66734 -57063 66806 -56936
rect 66944 -56947 67082 -56936
rect 66734 -57072 66818 -57063
rect 64010 -57225 64460 -57207
rect 63568 -57268 64460 -57225
rect 63568 -57286 64017 -57268
rect 64399 -57563 64460 -57268
rect 65133 -57445 65167 -57151
rect 65225 -57167 65270 -57097
rect 65617 -57117 66541 -57077
rect 65665 -57120 66541 -57117
rect 65126 -57563 65173 -57445
rect 65231 -57459 65265 -57167
rect 65329 -57444 65363 -57151
rect 65571 -57434 65605 -57151
rect 65665 -57160 65709 -57120
rect 66739 -57142 66818 -57072
rect 65322 -57563 65369 -57444
rect 65564 -57563 65611 -57434
rect 65669 -57459 65703 -57160
rect 67027 -57384 67061 -57093
rect 67025 -57495 67062 -57384
rect 67125 -57401 67159 -56756
rect 67354 -56826 67392 -56756
rect 67594 -56794 67628 -56715
rect 67869 -56724 68007 -56715
rect 67344 -56964 67398 -56826
rect 67497 -56828 67628 -56794
rect 67694 -56811 67832 -56757
rect 68079 -56826 68133 -56688
rect 68171 -56689 68205 -56645
rect 68171 -56743 68337 -56689
rect 67497 -57401 67531 -56828
rect 68171 -56858 68205 -56743
rect 68257 -56858 68311 -56841
rect 67595 -56897 67754 -56862
rect 68171 -56863 68311 -56858
rect 68143 -56892 68311 -56863
rect 67595 -57401 67629 -56897
rect 67720 -57401 67754 -56897
rect 67818 -57384 67852 -56893
rect 67948 -57383 67982 -56893
rect 66488 -57499 67099 -57495
rect 67817 -57499 67854 -57384
rect 67945 -57499 67982 -57383
rect 68046 -57401 68080 -56893
rect 68143 -56897 68205 -56892
rect 68144 -57401 68178 -56897
rect 68257 -56900 68311 -56892
rect 68372 -57010 68410 -56517
rect 68372 -57048 68664 -57010
rect 68274 -57382 68308 -57093
rect 68372 -57098 68410 -57048
rect 68272 -57499 68309 -57382
rect 68372 -57401 68406 -57098
rect 66488 -57563 68422 -57499
rect 64399 -57608 68422 -57563
rect 64399 -57676 66601 -57608
rect 66949 -57660 68422 -57608
rect 62628 -57949 63417 -57785
rect 68626 -57943 68664 -57048
rect 62628 -58002 66651 -57949
rect 62628 -62572 62845 -58002
rect 63341 -58025 66651 -58002
rect 63341 -58207 63417 -58025
rect 63341 -58283 63483 -58207
rect 63407 -58672 63483 -58283
rect 64416 -58249 65081 -58221
rect 64416 -58307 65451 -58249
rect 64416 -58388 64502 -58307
rect 64676 -58344 64711 -58307
rect 65001 -58310 65451 -58307
rect 63564 -58474 64502 -58388
rect 63407 -58764 63542 -58672
rect 63704 -58730 63738 -58474
rect 63802 -58730 63836 -58522
rect 63900 -58730 63934 -58474
rect 63998 -58696 64032 -58522
rect 64579 -58652 64613 -58344
rect 64677 -58652 64711 -58344
rect 64775 -58652 64809 -58344
rect 64873 -58652 64907 -58344
rect 64971 -58652 65005 -58344
rect 64547 -58695 64618 -58694
rect 64959 -58695 65033 -58689
rect 64547 -58696 65033 -58695
rect 63998 -58730 65033 -58696
rect 65390 -58717 65451 -58310
rect 63999 -58734 65033 -58730
rect 63999 -58736 64548 -58734
rect 63586 -58764 63659 -58758
rect 64959 -58760 65033 -58734
rect 63407 -58781 63659 -58764
rect 63412 -58805 63659 -58781
rect 64494 -58792 64629 -58784
rect 64474 -58794 64629 -58792
rect 63412 -58822 63542 -58805
rect 63586 -58818 63659 -58805
rect 64267 -58830 64629 -58794
rect 65146 -58803 65931 -58717
rect 64474 -58832 64629 -58830
rect 64494 -58838 64629 -58832
rect 64677 -58815 65096 -58807
rect 64677 -58845 65107 -58815
rect 63704 -59060 63738 -58852
rect 63900 -59060 63934 -58852
rect 64096 -59060 64130 -58852
rect 64677 -59189 64711 -58845
rect 64873 -59189 64907 -58845
rect 65046 -58994 65107 -58845
rect 65286 -58959 65320 -58803
rect 65384 -58959 65418 -58851
rect 65482 -58959 65516 -58803
rect 65580 -58959 65614 -58851
rect 65168 -58994 65241 -58988
rect 65046 -59007 65241 -58994
rect 65068 -59035 65241 -59007
rect 65168 -59048 65241 -59035
rect 65678 -59018 66050 -58948
rect 65286 -59190 65320 -59082
rect 65482 -59190 65516 -59082
rect 65678 -59190 65712 -59018
rect 63678 -60125 63712 -59781
rect 63874 -60125 63908 -59781
rect 64287 -59888 64321 -59780
rect 64483 -59888 64517 -59780
rect 64169 -59935 64242 -59922
rect 64069 -59963 64242 -59935
rect 64047 -59976 64242 -59963
rect 64047 -60125 64108 -59976
rect 64169 -59982 64242 -59976
rect 64679 -59952 64713 -59780
rect 63495 -60138 63630 -60132
rect 63475 -60140 63630 -60138
rect 62947 -60176 63630 -60140
rect 63678 -60155 64108 -60125
rect 63678 -60163 64097 -60155
rect 64287 -60167 64321 -60011
rect 64385 -60119 64419 -60011
rect 64483 -60167 64517 -60011
rect 64581 -60119 64615 -60011
rect 64679 -60022 64957 -59952
rect 63130 -61203 63266 -60176
rect 63475 -60178 63630 -60176
rect 63495 -60186 63630 -60178
rect 63322 -60236 63549 -60234
rect 63960 -60236 64034 -60210
rect 63322 -60274 64034 -60236
rect 64147 -60253 64762 -60167
rect 63548 -60275 64034 -60274
rect 63548 -60276 63619 -60275
rect 63960 -60281 64034 -60275
rect 63580 -60626 63614 -60318
rect 63678 -60626 63712 -60318
rect 63776 -60626 63810 -60318
rect 63874 -60626 63908 -60318
rect 63972 -60626 64006 -60318
rect 63677 -60678 63712 -60626
rect 64391 -60660 64452 -60253
rect 64881 -60417 64951 -60022
rect 65125 -60276 65159 -59692
rect 65332 -59658 65572 -59624
rect 65332 -59700 65374 -59658
rect 65121 -60335 65163 -60276
rect 65336 -60282 65370 -59700
rect 65434 -60280 65468 -59692
rect 65530 -59702 65572 -59658
rect 65333 -60335 65375 -60282
rect 65121 -60371 65375 -60335
rect 65430 -60334 65472 -60280
rect 65532 -60300 65566 -59702
rect 65744 -60286 65778 -59692
rect 65430 -60373 65571 -60334
rect 65528 -60385 65571 -60373
rect 65286 -60417 65441 -60407
rect 64881 -60453 65441 -60417
rect 64881 -60455 64951 -60453
rect 65286 -60462 65441 -60453
rect 65528 -60440 65709 -60385
rect 65528 -60510 65571 -60440
rect 65016 -60524 65171 -60515
rect 64979 -60558 65171 -60524
rect 65016 -60570 65171 -60558
rect 65217 -60550 65571 -60510
rect 65743 -60530 65786 -60286
rect 65980 -60355 66050 -59018
rect 66225 -58306 66317 -58221
rect 66248 -60281 66291 -58306
rect 66575 -58729 66651 -58025
rect 66877 -57981 68664 -57943
rect 66877 -58359 66915 -57981
rect 68084 -58280 68749 -58252
rect 68084 -58338 69119 -58280
rect 66854 -58413 66927 -58359
rect 68084 -58419 68170 -58338
rect 68344 -58375 68379 -58338
rect 68669 -58341 69119 -58338
rect 67232 -58505 68170 -58419
rect 67080 -58729 67210 -58703
rect 66575 -58795 67210 -58729
rect 67372 -58761 67406 -58505
rect 67470 -58761 67504 -58553
rect 67568 -58761 67602 -58505
rect 67666 -58727 67700 -58553
rect 68247 -58683 68281 -58375
rect 68345 -58683 68379 -58375
rect 68443 -58683 68477 -58375
rect 68541 -58683 68575 -58375
rect 68639 -58683 68673 -58375
rect 68215 -58726 68286 -58725
rect 68627 -58726 68701 -58720
rect 68215 -58727 68701 -58726
rect 67666 -58761 68701 -58727
rect 69058 -58748 69119 -58341
rect 72839 -56655 72873 -56311
rect 73035 -56655 73069 -56311
rect 73448 -56418 73482 -56310
rect 73644 -56418 73678 -56310
rect 73330 -56465 73403 -56452
rect 73230 -56493 73403 -56465
rect 73208 -56506 73403 -56493
rect 73208 -56655 73269 -56506
rect 73330 -56512 73403 -56506
rect 73840 -56482 73874 -56310
rect 72839 -56685 73269 -56655
rect 72839 -56693 73258 -56685
rect 73448 -56697 73482 -56541
rect 73546 -56649 73580 -56541
rect 73644 -56697 73678 -56541
rect 73742 -56649 73776 -56541
rect 73840 -56552 74118 -56482
rect 72483 -56766 72710 -56764
rect 73121 -56766 73195 -56740
rect 67667 -58765 68701 -58761
rect 67667 -58767 68216 -58765
rect 67254 -58795 67327 -58789
rect 68627 -58791 68701 -58765
rect 66575 -58805 67327 -58795
rect 67080 -58836 67327 -58805
rect 68162 -58823 68297 -58815
rect 68142 -58825 68297 -58823
rect 67080 -58853 67210 -58836
rect 67254 -58849 67327 -58836
rect 67107 -58903 67183 -58853
rect 67935 -58861 68297 -58825
rect 68814 -58834 69599 -58748
rect 68142 -58863 68297 -58861
rect 68162 -58869 68297 -58863
rect 68345 -58846 68764 -58838
rect 68345 -58876 68775 -58846
rect 67372 -59091 67406 -58883
rect 67568 -59091 67602 -58883
rect 67764 -59091 67798 -58883
rect 68345 -59220 68379 -58876
rect 68541 -59220 68575 -58876
rect 68714 -59025 68775 -58876
rect 68954 -58990 68988 -58834
rect 69052 -58990 69086 -58882
rect 69150 -58990 69184 -58834
rect 69248 -58990 69282 -58882
rect 68836 -59025 68909 -59019
rect 68714 -59038 68909 -59025
rect 68736 -59066 68909 -59038
rect 68836 -59079 68909 -59066
rect 69346 -59049 69718 -58979
rect 68954 -59221 68988 -59113
rect 69150 -59221 69184 -59113
rect 69346 -59221 69380 -59049
rect 67346 -60156 67380 -59812
rect 67542 -60156 67576 -59812
rect 67955 -59919 67989 -59811
rect 68151 -59919 68185 -59811
rect 67837 -59966 67910 -59953
rect 67737 -59994 67910 -59966
rect 67715 -60007 67910 -59994
rect 67715 -60156 67776 -60007
rect 67837 -60013 67910 -60007
rect 68347 -59983 68381 -59811
rect 67163 -60169 67298 -60163
rect 67143 -60171 67298 -60169
rect 66729 -60207 67298 -60171
rect 67346 -60186 67776 -60156
rect 67346 -60194 67765 -60186
rect 67955 -60198 67989 -60042
rect 68053 -60150 68087 -60042
rect 68151 -60198 68185 -60042
rect 68249 -60150 68283 -60042
rect 68347 -60053 68625 -59983
rect 66248 -60324 66533 -60281
rect 65969 -60427 66074 -60355
rect 66490 -60530 66533 -60324
rect 64002 -60678 64452 -60660
rect 63560 -60721 64452 -60678
rect 63560 -60739 64009 -60721
rect 64391 -61016 64452 -60721
rect 65125 -60898 65159 -60604
rect 65217 -60620 65262 -60550
rect 65609 -60570 66533 -60530
rect 65657 -60573 66533 -60570
rect 65118 -61016 65165 -60898
rect 65223 -60912 65257 -60620
rect 65321 -60897 65355 -60604
rect 65563 -60887 65597 -60604
rect 65657 -60613 65701 -60573
rect 65314 -61016 65361 -60897
rect 65556 -61016 65603 -60887
rect 65661 -60912 65695 -60613
rect 64391 -61129 65868 -61016
rect 66729 -61203 66865 -60207
rect 67143 -60209 67298 -60207
rect 67163 -60217 67298 -60209
rect 66990 -60267 67217 -60265
rect 67628 -60267 67702 -60241
rect 66990 -60305 67702 -60267
rect 67815 -60284 68430 -60198
rect 67216 -60306 67702 -60305
rect 67216 -60307 67287 -60306
rect 67628 -60312 67702 -60306
rect 67248 -60657 67282 -60349
rect 67346 -60657 67380 -60349
rect 67444 -60657 67478 -60349
rect 67542 -60657 67576 -60349
rect 67640 -60657 67674 -60349
rect 67345 -60709 67380 -60657
rect 68059 -60691 68120 -60284
rect 68549 -60448 68619 -60053
rect 68793 -60307 68827 -59723
rect 69000 -59689 69240 -59655
rect 69000 -59731 69042 -59689
rect 68789 -60366 68831 -60307
rect 69004 -60313 69038 -59731
rect 69102 -60311 69136 -59723
rect 69198 -59733 69240 -59689
rect 69001 -60366 69043 -60313
rect 68789 -60402 69043 -60366
rect 69098 -60365 69140 -60311
rect 69200 -60331 69234 -59733
rect 69412 -60317 69446 -59723
rect 69098 -60404 69239 -60365
rect 69196 -60416 69239 -60404
rect 68954 -60448 69109 -60438
rect 68549 -60484 69109 -60448
rect 68549 -60486 68619 -60484
rect 68954 -60493 69109 -60484
rect 69196 -60471 69377 -60416
rect 69196 -60541 69239 -60471
rect 68684 -60555 68839 -60546
rect 68647 -60589 68839 -60555
rect 68684 -60601 68839 -60589
rect 68885 -60581 69239 -60541
rect 69411 -60561 69454 -60317
rect 69648 -60386 69718 -59049
rect 69637 -60458 69742 -60386
rect 70106 -60561 70367 -60400
rect 67670 -60709 68120 -60691
rect 67228 -60752 68120 -60709
rect 67228 -60770 67677 -60752
rect 68059 -61047 68120 -60752
rect 68793 -60929 68827 -60635
rect 68885 -60651 68930 -60581
rect 69277 -60601 70479 -60561
rect 69325 -60604 70479 -60601
rect 68786 -61047 68833 -60929
rect 68891 -60943 68925 -60651
rect 68989 -60928 69023 -60635
rect 69231 -60918 69265 -60635
rect 69325 -60644 69369 -60604
rect 68982 -61047 69029 -60928
rect 69224 -61047 69271 -60918
rect 69329 -60943 69363 -60644
rect 70106 -60704 70367 -60604
rect 68059 -61160 69536 -61047
rect 63130 -61339 66865 -61203
rect 62571 -62855 62915 -62572
rect 9690 -63588 9826 -63586
rect 63130 -63588 63266 -61339
rect 72483 -56804 73195 -56766
rect 73308 -56783 73923 -56697
rect 72494 -57826 72570 -56804
rect 72709 -56805 73195 -56804
rect 72709 -56806 72780 -56805
rect 73121 -56811 73195 -56805
rect 72741 -57156 72775 -56848
rect 72839 -57156 72873 -56848
rect 72937 -57156 72971 -56848
rect 73035 -57156 73069 -56848
rect 73133 -57156 73167 -56848
rect 72838 -57208 72873 -57156
rect 73552 -57190 73613 -56783
rect 74042 -56947 74112 -56552
rect 74286 -56806 74320 -56222
rect 74493 -56188 74733 -56154
rect 74493 -56230 74535 -56188
rect 74282 -56865 74324 -56806
rect 74497 -56812 74531 -56230
rect 74595 -56810 74629 -56222
rect 74691 -56232 74733 -56188
rect 74494 -56865 74536 -56812
rect 74282 -56901 74536 -56865
rect 74591 -56864 74633 -56810
rect 74693 -56830 74727 -56232
rect 74905 -56816 74939 -56222
rect 74591 -56903 74732 -56864
rect 74689 -56915 74732 -56903
rect 74447 -56947 74602 -56937
rect 74042 -56983 74602 -56947
rect 74042 -56985 74112 -56983
rect 74447 -56992 74602 -56983
rect 74689 -56970 74870 -56915
rect 74689 -57040 74732 -56970
rect 74177 -57054 74332 -57045
rect 74140 -57088 74332 -57054
rect 74177 -57100 74332 -57088
rect 74378 -57080 74732 -57040
rect 74904 -57060 74947 -56816
rect 75141 -56885 75211 -55548
rect 82229 -55552 82263 -55344
rect 82425 -55552 82459 -55344
rect 82621 -55552 82655 -55344
rect 83202 -55681 83236 -55337
rect 83398 -55681 83432 -55337
rect 83571 -55486 83632 -55337
rect 83811 -55451 83845 -55295
rect 83909 -55451 83943 -55343
rect 84007 -55451 84041 -55295
rect 84105 -55451 84139 -55343
rect 83693 -55486 83766 -55480
rect 83571 -55499 83766 -55486
rect 83593 -55527 83766 -55499
rect 83693 -55540 83766 -55527
rect 84203 -55510 84575 -55440
rect 83811 -55682 83845 -55574
rect 84007 -55682 84041 -55574
rect 84203 -55682 84237 -55510
rect 76278 -56580 76312 -56080
rect 76457 -56044 76778 -56010
rect 76277 -56626 76312 -56580
rect 76457 -56626 76497 -56044
rect 76546 -56084 76581 -56044
rect 76547 -56588 76581 -56084
rect 76645 -56581 76679 -56080
rect 76743 -56083 76778 -56044
rect 76277 -56666 76497 -56626
rect 76642 -56701 76680 -56581
rect 76743 -56588 76777 -56083
rect 76873 -56664 76907 -56080
rect 77199 -56594 77233 -56080
rect 77427 -56370 77461 -56080
rect 77426 -56463 77463 -56370
rect 77426 -56500 77563 -56463
rect 77199 -56628 77358 -56594
rect 77022 -56664 77160 -56653
rect 76278 -56739 76680 -56701
rect 76747 -56698 77160 -56664
rect 76041 -56750 76179 -56740
rect 75651 -56784 76179 -56750
rect 75130 -56957 75235 -56885
rect 75651 -57060 75694 -56784
rect 76041 -56794 76179 -56784
rect 76097 -56885 76235 -56876
rect 75887 -56919 76235 -56885
rect 75887 -57046 75959 -56919
rect 76097 -56930 76235 -56919
rect 75887 -57055 75971 -57046
rect 73163 -57208 73613 -57190
rect 72721 -57251 73613 -57208
rect 72721 -57269 73170 -57251
rect 73552 -57546 73613 -57251
rect 74286 -57428 74320 -57134
rect 74378 -57150 74423 -57080
rect 74770 -57100 75694 -57060
rect 74818 -57103 75694 -57100
rect 74279 -57546 74326 -57428
rect 74384 -57442 74418 -57150
rect 74482 -57427 74516 -57134
rect 74724 -57417 74758 -57134
rect 74818 -57143 74862 -57103
rect 75892 -57125 75971 -57055
rect 74475 -57546 74522 -57427
rect 74717 -57546 74764 -57417
rect 74822 -57442 74856 -57143
rect 76180 -57367 76214 -57076
rect 76178 -57478 76215 -57367
rect 76278 -57384 76312 -56739
rect 76507 -56809 76545 -56739
rect 76747 -56777 76781 -56698
rect 77022 -56707 77160 -56698
rect 76497 -56947 76551 -56809
rect 76650 -56811 76781 -56777
rect 76847 -56794 76985 -56740
rect 77232 -56809 77286 -56671
rect 77324 -56672 77358 -56628
rect 77324 -56726 77490 -56672
rect 76650 -57384 76684 -56811
rect 77324 -56841 77358 -56726
rect 77410 -56841 77464 -56824
rect 76748 -56880 76907 -56845
rect 77324 -56846 77464 -56841
rect 77296 -56875 77464 -56846
rect 76748 -57384 76782 -56880
rect 76873 -57384 76907 -56880
rect 76971 -57367 77005 -56876
rect 77101 -57366 77135 -56876
rect 75641 -57482 76252 -57478
rect 76970 -57482 77007 -57367
rect 77098 -57482 77135 -57366
rect 77199 -57384 77233 -56876
rect 77296 -56880 77358 -56875
rect 77297 -57384 77331 -56880
rect 77410 -56883 77464 -56875
rect 77525 -56993 77563 -56500
rect 77525 -57031 77817 -56993
rect 77427 -57365 77461 -57076
rect 77525 -57081 77563 -57031
rect 77425 -57482 77462 -57365
rect 77525 -57384 77559 -57081
rect 75641 -57546 77575 -57482
rect 73552 -57591 77575 -57546
rect 73552 -57659 75754 -57591
rect 76102 -57643 77575 -57591
rect 71819 -57932 72570 -57826
rect 77779 -57926 77817 -57031
rect 71819 -57996 75804 -57932
rect 71819 -61832 71989 -57996
rect 72494 -58008 75804 -57996
rect 72494 -58190 72570 -58008
rect 72494 -58266 72636 -58190
rect 72560 -58655 72636 -58266
rect 73569 -58232 74234 -58204
rect 73569 -58290 74604 -58232
rect 73569 -58371 73655 -58290
rect 73829 -58327 73864 -58290
rect 74154 -58293 74604 -58290
rect 72717 -58457 73655 -58371
rect 72560 -58747 72695 -58655
rect 72857 -58713 72891 -58457
rect 72955 -58713 72989 -58505
rect 73053 -58713 73087 -58457
rect 73151 -58679 73185 -58505
rect 73732 -58635 73766 -58327
rect 73830 -58635 73864 -58327
rect 73928 -58635 73962 -58327
rect 74026 -58635 74060 -58327
rect 74124 -58635 74158 -58327
rect 73700 -58678 73771 -58677
rect 74112 -58678 74186 -58672
rect 73700 -58679 74186 -58678
rect 73151 -58713 74186 -58679
rect 74543 -58700 74604 -58293
rect 73152 -58717 74186 -58713
rect 73152 -58719 73701 -58717
rect 72739 -58747 72812 -58741
rect 74112 -58743 74186 -58717
rect 72560 -58764 72812 -58747
rect 72565 -58788 72812 -58764
rect 73647 -58775 73782 -58767
rect 73627 -58777 73782 -58775
rect 72565 -58805 72695 -58788
rect 72739 -58801 72812 -58788
rect 73420 -58813 73782 -58777
rect 74299 -58786 75084 -58700
rect 73627 -58815 73782 -58813
rect 73647 -58821 73782 -58815
rect 73830 -58798 74249 -58790
rect 73830 -58828 74260 -58798
rect 72857 -59043 72891 -58835
rect 73053 -59043 73087 -58835
rect 73249 -59043 73283 -58835
rect 73830 -59172 73864 -58828
rect 74026 -59172 74060 -58828
rect 74199 -58977 74260 -58828
rect 74439 -58942 74473 -58786
rect 74537 -58942 74571 -58834
rect 74635 -58942 74669 -58786
rect 74733 -58942 74767 -58834
rect 74321 -58977 74394 -58971
rect 74199 -58990 74394 -58977
rect 74221 -59018 74394 -58990
rect 74321 -59031 74394 -59018
rect 74831 -59001 75203 -58931
rect 74439 -59173 74473 -59065
rect 74635 -59173 74669 -59065
rect 74831 -59173 74865 -59001
rect 72831 -60108 72865 -59764
rect 73027 -60108 73061 -59764
rect 73440 -59871 73474 -59763
rect 73636 -59871 73670 -59763
rect 73322 -59918 73395 -59905
rect 73222 -59946 73395 -59918
rect 73200 -59959 73395 -59946
rect 73200 -60108 73261 -59959
rect 73322 -59965 73395 -59959
rect 73832 -59935 73866 -59763
rect 72648 -60121 72783 -60115
rect 72628 -60123 72783 -60121
rect 72100 -60159 72783 -60123
rect 72831 -60138 73261 -60108
rect 72831 -60146 73250 -60138
rect 73440 -60150 73474 -59994
rect 73538 -60102 73572 -59994
rect 73636 -60150 73670 -59994
rect 73734 -60102 73768 -59994
rect 73832 -60005 74110 -59935
rect 72283 -61186 72419 -60159
rect 72628 -60161 72783 -60159
rect 72648 -60169 72783 -60161
rect 72475 -60219 72702 -60217
rect 73113 -60219 73187 -60193
rect 72475 -60257 73187 -60219
rect 73300 -60236 73915 -60150
rect 72701 -60258 73187 -60257
rect 72701 -60259 72772 -60258
rect 73113 -60264 73187 -60258
rect 72733 -60609 72767 -60301
rect 72831 -60609 72865 -60301
rect 72929 -60609 72963 -60301
rect 73027 -60609 73061 -60301
rect 73125 -60609 73159 -60301
rect 72830 -60661 72865 -60609
rect 73544 -60643 73605 -60236
rect 74034 -60400 74104 -60005
rect 74278 -60259 74312 -59675
rect 74485 -59641 74725 -59607
rect 74485 -59683 74527 -59641
rect 74274 -60318 74316 -60259
rect 74489 -60265 74523 -59683
rect 74587 -60263 74621 -59675
rect 74683 -59685 74725 -59641
rect 74486 -60318 74528 -60265
rect 74274 -60354 74528 -60318
rect 74583 -60317 74625 -60263
rect 74685 -60283 74719 -59685
rect 74897 -60269 74931 -59675
rect 74583 -60356 74724 -60317
rect 74681 -60368 74724 -60356
rect 74439 -60400 74594 -60390
rect 74034 -60436 74594 -60400
rect 74034 -60438 74104 -60436
rect 74439 -60445 74594 -60436
rect 74681 -60423 74862 -60368
rect 74681 -60493 74724 -60423
rect 74169 -60507 74324 -60498
rect 74132 -60541 74324 -60507
rect 74169 -60553 74324 -60541
rect 74370 -60533 74724 -60493
rect 74896 -60513 74939 -60269
rect 75133 -60338 75203 -59001
rect 75378 -58289 75470 -58204
rect 75401 -60264 75444 -58289
rect 75728 -58712 75804 -58008
rect 76030 -57964 77817 -57926
rect 76030 -58342 76068 -57964
rect 77237 -58263 77902 -58235
rect 77237 -58321 78272 -58263
rect 76007 -58396 76080 -58342
rect 77237 -58402 77323 -58321
rect 77497 -58358 77532 -58321
rect 77822 -58324 78272 -58321
rect 76385 -58488 77323 -58402
rect 76233 -58712 76363 -58686
rect 75728 -58778 76363 -58712
rect 76525 -58744 76559 -58488
rect 76623 -58744 76657 -58536
rect 76721 -58744 76755 -58488
rect 76819 -58710 76853 -58536
rect 77400 -58666 77434 -58358
rect 77498 -58666 77532 -58358
rect 77596 -58666 77630 -58358
rect 77694 -58666 77728 -58358
rect 77792 -58666 77826 -58358
rect 77368 -58709 77439 -58708
rect 77780 -58709 77854 -58703
rect 77368 -58710 77854 -58709
rect 76819 -58744 77854 -58710
rect 78211 -58731 78272 -58324
rect 82203 -56617 82237 -56273
rect 82399 -56617 82433 -56273
rect 82812 -56380 82846 -56272
rect 83008 -56380 83042 -56272
rect 82694 -56427 82767 -56414
rect 82594 -56455 82767 -56427
rect 82572 -56468 82767 -56455
rect 82572 -56617 82633 -56468
rect 82694 -56474 82767 -56468
rect 83204 -56444 83238 -56272
rect 82203 -56647 82633 -56617
rect 82203 -56655 82622 -56647
rect 82812 -56659 82846 -56503
rect 82910 -56611 82944 -56503
rect 83008 -56659 83042 -56503
rect 83106 -56611 83140 -56503
rect 83204 -56514 83482 -56444
rect 81847 -56728 82074 -56726
rect 82485 -56728 82559 -56702
rect 76820 -58748 77854 -58744
rect 76820 -58750 77369 -58748
rect 76407 -58778 76480 -58772
rect 77780 -58774 77854 -58748
rect 75728 -58788 76480 -58778
rect 76233 -58819 76480 -58788
rect 77315 -58806 77450 -58798
rect 77295 -58808 77450 -58806
rect 76233 -58836 76363 -58819
rect 76407 -58832 76480 -58819
rect 76260 -58886 76336 -58836
rect 77088 -58844 77450 -58808
rect 77967 -58817 78752 -58731
rect 77295 -58846 77450 -58844
rect 77315 -58852 77450 -58846
rect 77498 -58829 77917 -58821
rect 77498 -58859 77928 -58829
rect 76525 -59074 76559 -58866
rect 76721 -59074 76755 -58866
rect 76917 -59074 76951 -58866
rect 77498 -59203 77532 -58859
rect 77694 -59203 77728 -58859
rect 77867 -59008 77928 -58859
rect 78107 -58973 78141 -58817
rect 78205 -58973 78239 -58865
rect 78303 -58973 78337 -58817
rect 78401 -58973 78435 -58865
rect 77989 -59008 78062 -59002
rect 77867 -59021 78062 -59008
rect 77889 -59049 78062 -59021
rect 77989 -59062 78062 -59049
rect 78499 -59032 78871 -58962
rect 78107 -59204 78141 -59096
rect 78303 -59204 78337 -59096
rect 78499 -59204 78533 -59032
rect 76499 -60139 76533 -59795
rect 76695 -60139 76729 -59795
rect 77108 -59902 77142 -59794
rect 77304 -59902 77338 -59794
rect 76990 -59949 77063 -59936
rect 76890 -59977 77063 -59949
rect 76868 -59990 77063 -59977
rect 76868 -60139 76929 -59990
rect 76990 -59996 77063 -59990
rect 77500 -59966 77534 -59794
rect 76316 -60152 76451 -60146
rect 76296 -60154 76451 -60152
rect 75882 -60190 76451 -60154
rect 76499 -60169 76929 -60139
rect 76499 -60177 76918 -60169
rect 77108 -60181 77142 -60025
rect 77206 -60133 77240 -60025
rect 77304 -60181 77338 -60025
rect 77402 -60133 77436 -60025
rect 77500 -60036 77778 -59966
rect 75401 -60307 75686 -60264
rect 75122 -60410 75227 -60338
rect 75643 -60513 75686 -60307
rect 73155 -60661 73605 -60643
rect 72713 -60704 73605 -60661
rect 72713 -60722 73162 -60704
rect 73544 -60999 73605 -60704
rect 74278 -60881 74312 -60587
rect 74370 -60603 74415 -60533
rect 74762 -60553 75686 -60513
rect 74810 -60556 75686 -60553
rect 74271 -60999 74318 -60881
rect 74376 -60895 74410 -60603
rect 74474 -60880 74508 -60587
rect 74716 -60870 74750 -60587
rect 74810 -60596 74854 -60556
rect 74467 -60999 74514 -60880
rect 74709 -60999 74756 -60870
rect 74814 -60895 74848 -60596
rect 73544 -61112 75021 -60999
rect 75882 -61186 76018 -60190
rect 76296 -60192 76451 -60190
rect 76316 -60200 76451 -60192
rect 76143 -60250 76370 -60248
rect 76781 -60250 76855 -60224
rect 76143 -60288 76855 -60250
rect 76968 -60267 77583 -60181
rect 76369 -60289 76855 -60288
rect 76369 -60290 76440 -60289
rect 76781 -60295 76855 -60289
rect 76401 -60640 76435 -60332
rect 76499 -60640 76533 -60332
rect 76597 -60640 76631 -60332
rect 76695 -60640 76729 -60332
rect 76793 -60640 76827 -60332
rect 76498 -60692 76533 -60640
rect 77212 -60674 77273 -60267
rect 77702 -60431 77772 -60036
rect 77946 -60290 77980 -59706
rect 78153 -59672 78393 -59638
rect 78153 -59714 78195 -59672
rect 77942 -60349 77984 -60290
rect 78157 -60296 78191 -59714
rect 78255 -60294 78289 -59706
rect 78351 -59716 78393 -59672
rect 78154 -60349 78196 -60296
rect 77942 -60385 78196 -60349
rect 78251 -60348 78293 -60294
rect 78353 -60314 78387 -59716
rect 78565 -60300 78599 -59706
rect 78251 -60387 78392 -60348
rect 78349 -60399 78392 -60387
rect 78107 -60431 78262 -60421
rect 77702 -60467 78262 -60431
rect 77702 -60469 77772 -60467
rect 78107 -60476 78262 -60467
rect 78349 -60454 78530 -60399
rect 78349 -60524 78392 -60454
rect 77837 -60538 77992 -60529
rect 77800 -60572 77992 -60538
rect 77837 -60584 77992 -60572
rect 78038 -60564 78392 -60524
rect 78564 -60544 78607 -60300
rect 78801 -60369 78871 -59032
rect 78790 -60441 78895 -60369
rect 79392 -60544 79494 -60506
rect 76823 -60692 77273 -60674
rect 76381 -60735 77273 -60692
rect 76381 -60753 76830 -60735
rect 77212 -61030 77273 -60735
rect 77946 -60912 77980 -60618
rect 78038 -60634 78083 -60564
rect 78430 -60584 79632 -60544
rect 78478 -60587 79632 -60584
rect 77939 -61030 77986 -60912
rect 78044 -60926 78078 -60634
rect 78142 -60911 78176 -60618
rect 78384 -60901 78418 -60618
rect 78478 -60627 78522 -60587
rect 79392 -60617 79494 -60587
rect 78135 -61030 78182 -60911
rect 78377 -61030 78424 -60901
rect 78482 -60926 78516 -60627
rect 77212 -61143 78689 -61030
rect 72283 -61322 76018 -61186
rect 71780 -62012 72026 -61832
rect -23846 -63724 63266 -63588
rect -23846 -63729 -21540 -63724
rect -23846 -63887 -23710 -63729
rect 72283 -63887 72419 -61322
rect 81847 -56766 82559 -56728
rect 82672 -56745 83287 -56659
rect 81858 -57747 81934 -56766
rect 82073 -56767 82559 -56766
rect 82073 -56768 82144 -56767
rect 82485 -56773 82559 -56767
rect 82105 -57118 82139 -56810
rect 82203 -57118 82237 -56810
rect 82301 -57118 82335 -56810
rect 82399 -57118 82433 -56810
rect 82497 -57118 82531 -56810
rect 82202 -57170 82237 -57118
rect 82916 -57152 82977 -56745
rect 83406 -56909 83476 -56514
rect 83650 -56768 83684 -56184
rect 83857 -56150 84097 -56116
rect 83857 -56192 83899 -56150
rect 83646 -56827 83688 -56768
rect 83861 -56774 83895 -56192
rect 83959 -56772 83993 -56184
rect 84055 -56194 84097 -56150
rect 83858 -56827 83900 -56774
rect 83646 -56863 83900 -56827
rect 83955 -56826 83997 -56772
rect 84057 -56792 84091 -56194
rect 84269 -56778 84303 -56184
rect 83955 -56865 84096 -56826
rect 84053 -56877 84096 -56865
rect 83811 -56909 83966 -56899
rect 83406 -56945 83966 -56909
rect 83406 -56947 83476 -56945
rect 83811 -56954 83966 -56945
rect 84053 -56932 84234 -56877
rect 84053 -57002 84096 -56932
rect 83541 -57016 83696 -57007
rect 83504 -57050 83696 -57016
rect 83541 -57062 83696 -57050
rect 83742 -57042 84096 -57002
rect 84268 -57022 84311 -56778
rect 84505 -56847 84575 -55510
rect 85642 -56542 85676 -56042
rect 85821 -56006 86142 -55972
rect 85641 -56588 85676 -56542
rect 85821 -56588 85861 -56006
rect 85910 -56046 85945 -56006
rect 85911 -56550 85945 -56046
rect 86009 -56543 86043 -56042
rect 86107 -56045 86142 -56006
rect 85641 -56628 85861 -56588
rect 86006 -56663 86044 -56543
rect 86107 -56550 86141 -56045
rect 86237 -56626 86271 -56042
rect 86563 -56556 86597 -56042
rect 86791 -56332 86825 -56042
rect 86790 -56425 86827 -56332
rect 86790 -56462 86927 -56425
rect 86563 -56590 86722 -56556
rect 86386 -56626 86524 -56615
rect 85642 -56701 86044 -56663
rect 86111 -56660 86524 -56626
rect 85405 -56712 85543 -56702
rect 85015 -56746 85543 -56712
rect 84494 -56919 84599 -56847
rect 85015 -57022 85058 -56746
rect 85405 -56756 85543 -56746
rect 85461 -56847 85599 -56838
rect 85251 -56881 85599 -56847
rect 85251 -57008 85323 -56881
rect 85461 -56892 85599 -56881
rect 85251 -57017 85335 -57008
rect 82527 -57170 82977 -57152
rect 82085 -57213 82977 -57170
rect 82085 -57231 82534 -57213
rect 82916 -57508 82977 -57213
rect 83650 -57390 83684 -57096
rect 83742 -57112 83787 -57042
rect 84134 -57062 85058 -57022
rect 84182 -57065 85058 -57062
rect 83643 -57508 83690 -57390
rect 83748 -57404 83782 -57112
rect 83846 -57389 83880 -57096
rect 84088 -57379 84122 -57096
rect 84182 -57105 84226 -57065
rect 85256 -57087 85335 -57017
rect 83839 -57508 83886 -57389
rect 84081 -57508 84128 -57379
rect 84186 -57404 84220 -57105
rect 85544 -57329 85578 -57038
rect 85542 -57440 85579 -57329
rect 85642 -57346 85676 -56701
rect 85871 -56771 85909 -56701
rect 86111 -56739 86145 -56660
rect 86386 -56669 86524 -56660
rect 85861 -56909 85915 -56771
rect 86014 -56773 86145 -56739
rect 86211 -56756 86349 -56702
rect 86596 -56771 86650 -56633
rect 86688 -56634 86722 -56590
rect 86688 -56688 86854 -56634
rect 86014 -57346 86048 -56773
rect 86688 -56803 86722 -56688
rect 86774 -56803 86828 -56786
rect 86112 -56842 86271 -56807
rect 86688 -56808 86828 -56803
rect 86660 -56837 86828 -56808
rect 86112 -57346 86146 -56842
rect 86237 -57346 86271 -56842
rect 86335 -57329 86369 -56838
rect 86465 -57328 86499 -56838
rect 85005 -57444 85616 -57440
rect 86334 -57444 86371 -57329
rect 86462 -57444 86499 -57328
rect 86563 -57346 86597 -56838
rect 86660 -56842 86722 -56837
rect 86661 -57346 86695 -56842
rect 86774 -56845 86828 -56837
rect 86889 -56955 86927 -56462
rect 86889 -56993 87181 -56955
rect 86791 -57327 86825 -57038
rect 86889 -57043 86927 -56993
rect 86789 -57444 86826 -57327
rect 86889 -57346 86923 -57043
rect 85005 -57508 86939 -57444
rect 82916 -57553 86939 -57508
rect 82916 -57621 85118 -57553
rect 85466 -57605 86939 -57553
rect 81095 -57894 81976 -57747
rect 87143 -57888 87181 -56993
rect 81095 -57970 85168 -57894
rect 81095 -57973 81976 -57970
rect 81095 -62575 81321 -57973
rect 81858 -58152 81934 -57973
rect 81858 -58228 82000 -58152
rect 81924 -58617 82000 -58228
rect 82933 -58194 83598 -58166
rect 82933 -58252 83968 -58194
rect 82933 -58333 83019 -58252
rect 83193 -58289 83228 -58252
rect 83518 -58255 83968 -58252
rect 82081 -58419 83019 -58333
rect 81924 -58709 82059 -58617
rect 82221 -58675 82255 -58419
rect 82319 -58675 82353 -58467
rect 82417 -58675 82451 -58419
rect 82515 -58641 82549 -58467
rect 83096 -58597 83130 -58289
rect 83194 -58597 83228 -58289
rect 83292 -58597 83326 -58289
rect 83390 -58597 83424 -58289
rect 83488 -58597 83522 -58289
rect 83064 -58640 83135 -58639
rect 83476 -58640 83550 -58634
rect 83064 -58641 83550 -58640
rect 82515 -58675 83550 -58641
rect 83907 -58662 83968 -58255
rect 82516 -58679 83550 -58675
rect 82516 -58681 83065 -58679
rect 82103 -58709 82176 -58703
rect 83476 -58705 83550 -58679
rect 81924 -58726 82176 -58709
rect 81929 -58750 82176 -58726
rect 83011 -58737 83146 -58729
rect 82991 -58739 83146 -58737
rect 81929 -58767 82059 -58750
rect 82103 -58763 82176 -58750
rect 82784 -58775 83146 -58739
rect 83663 -58748 84448 -58662
rect 82991 -58777 83146 -58775
rect 83011 -58783 83146 -58777
rect 83194 -58760 83613 -58752
rect 83194 -58790 83624 -58760
rect 82221 -59005 82255 -58797
rect 82417 -59005 82451 -58797
rect 82613 -59005 82647 -58797
rect 83194 -59134 83228 -58790
rect 83390 -59134 83424 -58790
rect 83563 -58939 83624 -58790
rect 83803 -58904 83837 -58748
rect 83901 -58904 83935 -58796
rect 83999 -58904 84033 -58748
rect 84097 -58904 84131 -58796
rect 83685 -58939 83758 -58933
rect 83563 -58952 83758 -58939
rect 83585 -58980 83758 -58952
rect 83685 -58993 83758 -58980
rect 84195 -58963 84567 -58893
rect 83803 -59135 83837 -59027
rect 83999 -59135 84033 -59027
rect 84195 -59135 84229 -58963
rect 82195 -60070 82229 -59726
rect 82391 -60070 82425 -59726
rect 82804 -59833 82838 -59725
rect 83000 -59833 83034 -59725
rect 82686 -59880 82759 -59867
rect 82586 -59908 82759 -59880
rect 82564 -59921 82759 -59908
rect 82564 -60070 82625 -59921
rect 82686 -59927 82759 -59921
rect 83196 -59897 83230 -59725
rect 82012 -60083 82147 -60077
rect 81992 -60085 82147 -60083
rect 81464 -60121 82147 -60085
rect 82195 -60100 82625 -60070
rect 82195 -60108 82614 -60100
rect 82804 -60112 82838 -59956
rect 82902 -60064 82936 -59956
rect 83000 -60112 83034 -59956
rect 83098 -60064 83132 -59956
rect 83196 -59967 83474 -59897
rect 81647 -61148 81783 -60121
rect 81992 -60123 82147 -60121
rect 82012 -60131 82147 -60123
rect 81839 -60181 82066 -60179
rect 82477 -60181 82551 -60155
rect 81839 -60219 82551 -60181
rect 82664 -60198 83279 -60112
rect 82065 -60220 82551 -60219
rect 82065 -60221 82136 -60220
rect 82477 -60226 82551 -60220
rect 82097 -60571 82131 -60263
rect 82195 -60571 82229 -60263
rect 82293 -60571 82327 -60263
rect 82391 -60571 82425 -60263
rect 82489 -60571 82523 -60263
rect 82194 -60623 82229 -60571
rect 82908 -60605 82969 -60198
rect 83398 -60362 83468 -59967
rect 83642 -60221 83676 -59637
rect 83849 -59603 84089 -59569
rect 83849 -59645 83891 -59603
rect 83638 -60280 83680 -60221
rect 83853 -60227 83887 -59645
rect 83951 -60225 83985 -59637
rect 84047 -59647 84089 -59603
rect 83850 -60280 83892 -60227
rect 83638 -60316 83892 -60280
rect 83947 -60279 83989 -60225
rect 84049 -60245 84083 -59647
rect 84261 -60231 84295 -59637
rect 83947 -60318 84088 -60279
rect 84045 -60330 84088 -60318
rect 83803 -60362 83958 -60352
rect 83398 -60398 83958 -60362
rect 83398 -60400 83468 -60398
rect 83803 -60407 83958 -60398
rect 84045 -60385 84226 -60330
rect 84045 -60455 84088 -60385
rect 83533 -60469 83688 -60460
rect 83496 -60503 83688 -60469
rect 83533 -60515 83688 -60503
rect 83734 -60495 84088 -60455
rect 84260 -60475 84303 -60231
rect 84497 -60300 84567 -58963
rect 84742 -58251 84834 -58166
rect 84765 -60226 84808 -58251
rect 85092 -58674 85168 -57970
rect 85394 -57926 87181 -57888
rect 85394 -58304 85432 -57926
rect 86601 -58225 87266 -58197
rect 86601 -58283 87636 -58225
rect 85371 -58358 85444 -58304
rect 86601 -58364 86687 -58283
rect 86861 -58320 86896 -58283
rect 87186 -58286 87636 -58283
rect 85749 -58450 86687 -58364
rect 85597 -58674 85727 -58648
rect 85092 -58740 85727 -58674
rect 85889 -58706 85923 -58450
rect 85987 -58706 86021 -58498
rect 86085 -58706 86119 -58450
rect 86183 -58672 86217 -58498
rect 86764 -58628 86798 -58320
rect 86862 -58628 86896 -58320
rect 86960 -58628 86994 -58320
rect 87058 -58628 87092 -58320
rect 87156 -58628 87190 -58320
rect 86732 -58671 86803 -58670
rect 87144 -58671 87218 -58665
rect 86732 -58672 87218 -58671
rect 86183 -58706 87218 -58672
rect 87575 -58693 87636 -58286
rect 86184 -58710 87218 -58706
rect 86184 -58712 86733 -58710
rect 85771 -58740 85844 -58734
rect 87144 -58736 87218 -58710
rect 85092 -58750 85844 -58740
rect 85597 -58781 85844 -58750
rect 86679 -58768 86814 -58760
rect 86659 -58770 86814 -58768
rect 85597 -58798 85727 -58781
rect 85771 -58794 85844 -58781
rect 85624 -58848 85700 -58798
rect 86452 -58806 86814 -58770
rect 87331 -58779 88116 -58693
rect 86659 -58808 86814 -58806
rect 86679 -58814 86814 -58808
rect 86862 -58791 87281 -58783
rect 86862 -58821 87292 -58791
rect 85889 -59036 85923 -58828
rect 86085 -59036 86119 -58828
rect 86281 -59036 86315 -58828
rect 86862 -59165 86896 -58821
rect 87058 -59165 87092 -58821
rect 87231 -58970 87292 -58821
rect 87471 -58935 87505 -58779
rect 87569 -58935 87603 -58827
rect 87667 -58935 87701 -58779
rect 87765 -58935 87799 -58827
rect 87353 -58970 87426 -58964
rect 87231 -58983 87426 -58970
rect 87253 -59011 87426 -58983
rect 87353 -59024 87426 -59011
rect 87863 -58994 88235 -58924
rect 87471 -59166 87505 -59058
rect 87667 -59166 87701 -59058
rect 87863 -59166 87897 -58994
rect 85863 -60101 85897 -59757
rect 86059 -60101 86093 -59757
rect 86472 -59864 86506 -59756
rect 86668 -59864 86702 -59756
rect 86354 -59911 86427 -59898
rect 86254 -59939 86427 -59911
rect 86232 -59952 86427 -59939
rect 86232 -60101 86293 -59952
rect 86354 -59958 86427 -59952
rect 86864 -59928 86898 -59756
rect 85680 -60114 85815 -60108
rect 85660 -60116 85815 -60114
rect 85246 -60152 85815 -60116
rect 85863 -60131 86293 -60101
rect 85863 -60139 86282 -60131
rect 86472 -60143 86506 -59987
rect 86570 -60095 86604 -59987
rect 86668 -60143 86702 -59987
rect 86766 -60095 86800 -59987
rect 86864 -59998 87142 -59928
rect 84765 -60269 85050 -60226
rect 84486 -60372 84591 -60300
rect 85007 -60475 85050 -60269
rect 82519 -60623 82969 -60605
rect 82077 -60666 82969 -60623
rect 82077 -60684 82526 -60666
rect 82908 -60961 82969 -60666
rect 83642 -60843 83676 -60549
rect 83734 -60565 83779 -60495
rect 84126 -60515 85050 -60475
rect 84174 -60518 85050 -60515
rect 83635 -60961 83682 -60843
rect 83740 -60857 83774 -60565
rect 83838 -60842 83872 -60549
rect 84080 -60832 84114 -60549
rect 84174 -60558 84218 -60518
rect 83831 -60961 83878 -60842
rect 84073 -60961 84120 -60832
rect 84178 -60857 84212 -60558
rect 82908 -61074 84385 -60961
rect 85246 -61148 85382 -60152
rect 85660 -60154 85815 -60152
rect 85680 -60162 85815 -60154
rect 85507 -60212 85734 -60210
rect 86145 -60212 86219 -60186
rect 85507 -60250 86219 -60212
rect 86332 -60229 86947 -60143
rect 85733 -60251 86219 -60250
rect 85733 -60252 85804 -60251
rect 86145 -60257 86219 -60251
rect 85765 -60602 85799 -60294
rect 85863 -60602 85897 -60294
rect 85961 -60602 85995 -60294
rect 86059 -60602 86093 -60294
rect 86157 -60602 86191 -60294
rect 85862 -60654 85897 -60602
rect 86576 -60636 86637 -60229
rect 87066 -60393 87136 -59998
rect 87310 -60252 87344 -59668
rect 87517 -59634 87757 -59600
rect 87517 -59676 87559 -59634
rect 87306 -60311 87348 -60252
rect 87521 -60258 87555 -59676
rect 87619 -60256 87653 -59668
rect 87715 -59678 87757 -59634
rect 87518 -60311 87560 -60258
rect 87306 -60347 87560 -60311
rect 87615 -60310 87657 -60256
rect 87717 -60276 87751 -59678
rect 87929 -60262 87963 -59668
rect 87615 -60349 87756 -60310
rect 87713 -60361 87756 -60349
rect 87471 -60393 87626 -60383
rect 87066 -60429 87626 -60393
rect 87066 -60431 87136 -60429
rect 87471 -60438 87626 -60429
rect 87713 -60416 87894 -60361
rect 87713 -60486 87756 -60416
rect 87201 -60500 87356 -60491
rect 87164 -60534 87356 -60500
rect 87201 -60546 87356 -60534
rect 87402 -60526 87756 -60486
rect 87928 -60506 87971 -60262
rect 88165 -60331 88235 -58994
rect 88154 -60403 88259 -60331
rect 88783 -60506 89142 -60356
rect 86187 -60654 86637 -60636
rect 85745 -60697 86637 -60654
rect 85745 -60715 86194 -60697
rect 86576 -60992 86637 -60697
rect 87310 -60874 87344 -60580
rect 87402 -60596 87447 -60526
rect 87794 -60546 89142 -60506
rect 87842 -60549 89142 -60546
rect 87303 -60992 87350 -60874
rect 87408 -60888 87442 -60596
rect 87506 -60873 87540 -60580
rect 87748 -60863 87782 -60580
rect 87842 -60589 87886 -60549
rect 87499 -60992 87546 -60873
rect 87741 -60992 87788 -60863
rect 87846 -60888 87880 -60589
rect 88783 -60699 89142 -60549
rect 86576 -61105 88053 -60992
rect 81647 -61284 85382 -61148
rect 81006 -62851 81393 -62575
rect -23846 -64023 72419 -63887
rect -23846 -64257 -23710 -64023
rect 81671 -64257 81807 -61284
rect -23846 -64393 81807 -64257
rect -6606 -64897 18338 -64761
rect -23356 -65134 11812 -64999
<< metal1 >>
rect -12872 120359 -10450 120472
rect -12872 116804 -12759 120359
rect -11358 120177 -11167 120328
rect -12651 119654 -12351 119700
rect -12651 119412 -12351 119458
rect -12651 119216 -12351 119262
rect -11333 120018 -11194 120177
rect -11345 119927 -11182 120018
rect -10929 119867 -10829 119913
rect -12039 119737 -11439 119783
rect -10563 119764 -10450 120359
rect -10929 119671 -10829 119717
rect -10698 119573 -10598 119619
rect -10929 119475 -10829 119521
rect -10698 119377 -10598 119423
rect -12039 119314 -11439 119360
rect -10929 119279 -10829 119325
rect -12039 119118 -11439 119164
rect -10928 119062 -10628 119108
rect -11627 118868 -11527 118914
rect -10928 118866 -10628 118912
rect -10391 118768 -10091 118814
rect -11627 118672 -11527 118718
rect -10928 118670 -10628 118716
rect -8113 118795 -7813 118841
rect -9109 118697 -8809 118743
rect -11858 118574 -11758 118620
rect -11627 118476 -11527 118522
rect -11858 118378 -11758 118424
rect -11627 118280 -11527 118326
rect -10799 118285 -10599 118331
rect -8113 118599 -7813 118645
rect -9109 118371 -8609 118417
rect -11828 118063 -11528 118109
rect -10799 118089 -10599 118135
rect -10469 117991 -10269 118037
rect -11828 117867 -11528 117913
rect -10799 117893 -10599 117939
rect -12365 117769 -12065 117815
rect -10469 117795 -10269 117841
rect -11828 117671 -11528 117717
rect -10799 117697 -10599 117743
rect -9109 118241 -8609 118287
rect -8313 118371 -7813 118417
rect -8313 118241 -7813 118287
rect -9109 117450 -8809 117496
rect -8313 117646 -7813 117692
rect -8313 117450 -7813 117496
rect -12872 116691 -10419 116804
rect -12872 116131 -12728 116691
rect -11280 116507 -11143 116603
rect -12841 116127 -12728 116131
rect -12620 115986 -12320 116032
rect -12620 115744 -12320 115790
rect -12620 115548 -12320 115594
rect -12008 116069 -11408 116115
rect -12008 115646 -11408 115692
rect -12008 115450 -11408 115496
rect -11254 115387 -11172 116507
rect -10532 116438 -10419 116691
rect -9388 116699 -6966 116812
rect -9388 116438 -9275 116699
rect -7874 116517 -7724 116627
rect -10898 116199 -10798 116245
rect -10532 116325 -9274 116438
rect -10532 116096 -10419 116325
rect -9388 116135 -9275 116325
rect -10898 116003 -10798 116049
rect -9167 115994 -8867 116040
rect -10667 115905 -10567 115951
rect -10898 115807 -10798 115853
rect -10667 115709 -10567 115755
rect -9167 115752 -8867 115798
rect -10898 115611 -10798 115657
rect -9167 115556 -8867 115602
rect -7856 116363 -7760 116517
rect -7862 116289 -7744 116363
rect -7445 116207 -7345 116253
rect -8555 116077 -7955 116123
rect -7079 116104 -6966 116699
rect -7445 116011 -7345 116057
rect -7214 115913 -7114 115959
rect -7445 115815 -7345 115861
rect -7214 115717 -7114 115763
rect -8555 115654 -7955 115700
rect -7445 115619 -7345 115665
rect -8555 115458 -7955 115504
rect -10897 115394 -10597 115440
rect -7444 115402 -7144 115448
rect -11596 115200 -11496 115246
rect -11261 115204 -11131 115387
rect -10897 115198 -10597 115244
rect -10360 115100 -10060 115146
rect -11596 115004 -11496 115050
rect -10897 115002 -10597 115048
rect -8143 115208 -8043 115254
rect -7444 115206 -7144 115252
rect -6907 115108 -6607 115154
rect -8143 115012 -8043 115058
rect -11827 114906 -11727 114952
rect -7444 115010 -7144 115056
rect -11596 114808 -11496 114854
rect -11827 114710 -11727 114756
rect -14196 58887 -13951 114640
rect -11596 114612 -11496 114658
rect -10768 114617 -10568 114663
rect -8374 114914 -8274 114960
rect -8143 114816 -8043 114862
rect -8374 114718 -8274 114764
rect -11797 114395 -11497 114441
rect -10768 114421 -10568 114467
rect -10438 114323 -10238 114369
rect -11797 114199 -11497 114245
rect -10768 114225 -10568 114271
rect -12334 114101 -12034 114147
rect -10438 114127 -10238 114173
rect -11797 114003 -11497 114049
rect -10768 114029 -10568 114075
rect -8143 114620 -8043 114666
rect -7315 114625 -7115 114671
rect -8344 114403 -8044 114449
rect -7315 114429 -7115 114475
rect -6985 114331 -6785 114377
rect -8344 114207 -8044 114253
rect -7315 114233 -7115 114279
rect -8881 114109 -8581 114155
rect -6985 114135 -6785 114181
rect -8344 114011 -8044 114057
rect -7315 114037 -7115 114083
rect -12910 110995 -10488 111108
rect -12910 107440 -12797 110995
rect -11396 110813 -11205 110964
rect -12689 110290 -12389 110336
rect -12689 110048 -12389 110094
rect -12689 109852 -12389 109898
rect -11371 110654 -11232 110813
rect -11383 110563 -11220 110654
rect -10967 110503 -10867 110549
rect -12077 110373 -11477 110419
rect -10601 110400 -10488 110995
rect -10967 110307 -10867 110353
rect -10736 110209 -10636 110255
rect -10967 110111 -10867 110157
rect -10736 110013 -10636 110059
rect -12077 109950 -11477 109996
rect -10967 109915 -10867 109961
rect -12077 109754 -11477 109800
rect -10966 109698 -10666 109744
rect -11665 109504 -11565 109550
rect -10966 109502 -10666 109548
rect -10429 109404 -10129 109450
rect -11665 109308 -11565 109354
rect -10966 109306 -10666 109352
rect -8151 109431 -7851 109477
rect -9147 109333 -8847 109379
rect -11896 109210 -11796 109256
rect -11665 109112 -11565 109158
rect -11896 109014 -11796 109060
rect -11665 108916 -11565 108962
rect -10837 108921 -10637 108967
rect -8151 109235 -7851 109281
rect -9147 109007 -8647 109053
rect -11866 108699 -11566 108745
rect -10837 108725 -10637 108771
rect -10507 108627 -10307 108673
rect -11866 108503 -11566 108549
rect -10837 108529 -10637 108575
rect -12403 108405 -12103 108451
rect -10507 108431 -10307 108477
rect -11866 108307 -11566 108353
rect -10837 108333 -10637 108379
rect -9147 108877 -8647 108923
rect -8351 109007 -7851 109053
rect -8351 108877 -7851 108923
rect -9147 108086 -8847 108132
rect -8351 108282 -7851 108328
rect -8351 108086 -7851 108132
rect -12910 107327 -10457 107440
rect -12910 106767 -12766 107327
rect -11318 107143 -11181 107239
rect -12879 106763 -12766 106767
rect -12658 106622 -12358 106668
rect -12658 106380 -12358 106426
rect -12658 106184 -12358 106230
rect -12046 106705 -11446 106751
rect -12046 106282 -11446 106328
rect -12046 106086 -11446 106132
rect -11292 106023 -11210 107143
rect -10570 107074 -10457 107327
rect -9426 107335 -7004 107448
rect -9426 107074 -9313 107335
rect -7912 107153 -7762 107263
rect -10936 106835 -10836 106881
rect -10570 106961 -9312 107074
rect -10570 106732 -10457 106961
rect -9426 106771 -9313 106961
rect -10936 106639 -10836 106685
rect -9205 106630 -8905 106676
rect -10705 106541 -10605 106587
rect -10936 106443 -10836 106489
rect -10705 106345 -10605 106391
rect -9205 106388 -8905 106434
rect -10936 106247 -10836 106293
rect -9205 106192 -8905 106238
rect -7894 106999 -7798 107153
rect -7900 106925 -7782 106999
rect -7483 106843 -7383 106889
rect -8593 106713 -7993 106759
rect -7117 106740 -7004 107335
rect -7483 106647 -7383 106693
rect -7252 106549 -7152 106595
rect -7483 106451 -7383 106497
rect -7252 106353 -7152 106399
rect -8593 106290 -7993 106336
rect -7483 106255 -7383 106301
rect -8593 106094 -7993 106140
rect -10935 106030 -10635 106076
rect -7482 106038 -7182 106084
rect -11634 105836 -11534 105882
rect -11299 105840 -11169 106023
rect -10935 105834 -10635 105880
rect -10398 105736 -10098 105782
rect -11634 105640 -11534 105686
rect -10935 105638 -10635 105684
rect -8181 105844 -8081 105890
rect -7482 105842 -7182 105888
rect -6945 105744 -6645 105790
rect -8181 105648 -8081 105694
rect -11865 105542 -11765 105588
rect -7482 105646 -7182 105692
rect -11634 105444 -11534 105490
rect -11865 105346 -11765 105392
rect -11634 105248 -11534 105294
rect -10806 105253 -10606 105299
rect -8412 105550 -8312 105596
rect -8181 105452 -8081 105498
rect -8412 105354 -8312 105400
rect -11835 105031 -11535 105077
rect -10806 105057 -10606 105103
rect -10476 104959 -10276 105005
rect -11835 104835 -11535 104881
rect -10806 104861 -10606 104907
rect -12372 104737 -12072 104783
rect -10476 104763 -10276 104809
rect -11835 104639 -11535 104685
rect -10806 104665 -10606 104711
rect -8181 105256 -8081 105302
rect -7353 105261 -7153 105307
rect -8382 105039 -8082 105085
rect -7353 105065 -7153 105111
rect -7023 104967 -6823 105013
rect -8382 104843 -8082 104889
rect -7353 104869 -7153 104915
rect -8919 104745 -8619 104791
rect -7023 104771 -6823 104817
rect -8382 104647 -8082 104693
rect -7353 104673 -7153 104719
rect -12927 101842 -10505 101955
rect -12927 98287 -12814 101842
rect -11413 101660 -11222 101811
rect -12706 101137 -12406 101183
rect -12706 100895 -12406 100941
rect -12706 100699 -12406 100745
rect -11388 101501 -11249 101660
rect -11400 101410 -11237 101501
rect -10984 101350 -10884 101396
rect -12094 101220 -11494 101266
rect -10618 101247 -10505 101842
rect -10984 101154 -10884 101200
rect -10753 101056 -10653 101102
rect -10984 100958 -10884 101004
rect -10753 100860 -10653 100906
rect -12094 100797 -11494 100843
rect -10984 100762 -10884 100808
rect -12094 100601 -11494 100647
rect -10983 100545 -10683 100591
rect -11682 100351 -11582 100397
rect -10983 100349 -10683 100395
rect -10446 100251 -10146 100297
rect -11682 100155 -11582 100201
rect -10983 100153 -10683 100199
rect -8168 100278 -7868 100324
rect -9164 100180 -8864 100226
rect -11913 100057 -11813 100103
rect -11682 99959 -11582 100005
rect -11913 99861 -11813 99907
rect -11682 99763 -11582 99809
rect -10854 99768 -10654 99814
rect -8168 100082 -7868 100128
rect -9164 99854 -8664 99900
rect -11883 99546 -11583 99592
rect -10854 99572 -10654 99618
rect -10524 99474 -10324 99520
rect -11883 99350 -11583 99396
rect -10854 99376 -10654 99422
rect -12420 99252 -12120 99298
rect -10524 99278 -10324 99324
rect -11883 99154 -11583 99200
rect -10854 99180 -10654 99226
rect -9164 99724 -8664 99770
rect -8368 99854 -7868 99900
rect -8368 99724 -7868 99770
rect -9164 98933 -8864 98979
rect -8368 99129 -7868 99175
rect -8368 98933 -7868 98979
rect -12927 98174 -10474 98287
rect -12927 97614 -12783 98174
rect -11335 97990 -11198 98086
rect -12896 97610 -12783 97614
rect -12675 97469 -12375 97515
rect -12675 97227 -12375 97273
rect -12675 97031 -12375 97077
rect -12063 97552 -11463 97598
rect -12063 97129 -11463 97175
rect -12063 96933 -11463 96979
rect -11309 96870 -11227 97990
rect -10587 97921 -10474 98174
rect -9443 98182 -7021 98295
rect -9443 97921 -9330 98182
rect -7929 98000 -7779 98110
rect -10953 97682 -10853 97728
rect -10587 97808 -9329 97921
rect -10587 97579 -10474 97808
rect -9443 97618 -9330 97808
rect -10953 97486 -10853 97532
rect -9222 97477 -8922 97523
rect -10722 97388 -10622 97434
rect -10953 97290 -10853 97336
rect -10722 97192 -10622 97238
rect -9222 97235 -8922 97281
rect -10953 97094 -10853 97140
rect -9222 97039 -8922 97085
rect -7911 97846 -7815 98000
rect -7917 97772 -7799 97846
rect -7500 97690 -7400 97736
rect -8610 97560 -8010 97606
rect -7134 97587 -7021 98182
rect -7500 97494 -7400 97540
rect -7269 97396 -7169 97442
rect -7500 97298 -7400 97344
rect -7269 97200 -7169 97246
rect -8610 97137 -8010 97183
rect -7500 97102 -7400 97148
rect -8610 96941 -8010 96987
rect -10952 96877 -10652 96923
rect -7499 96885 -7199 96931
rect -11651 96683 -11551 96729
rect -11316 96687 -11186 96870
rect -10952 96681 -10652 96727
rect -10415 96583 -10115 96629
rect -11651 96487 -11551 96533
rect -10952 96485 -10652 96531
rect -8198 96691 -8098 96737
rect -7499 96689 -7199 96735
rect -6962 96591 -6662 96637
rect -8198 96495 -8098 96541
rect -11882 96389 -11782 96435
rect -7499 96493 -7199 96539
rect -11651 96291 -11551 96337
rect -11882 96193 -11782 96239
rect -11651 96095 -11551 96141
rect -10823 96100 -10623 96146
rect -8429 96397 -8329 96443
rect -8198 96299 -8098 96345
rect -8429 96201 -8329 96247
rect -11852 95878 -11552 95924
rect -10823 95904 -10623 95950
rect -10493 95806 -10293 95852
rect -11852 95682 -11552 95728
rect -10823 95708 -10623 95754
rect -12389 95584 -12089 95630
rect -10493 95610 -10293 95656
rect -11852 95486 -11552 95532
rect -10823 95512 -10623 95558
rect -8198 96103 -8098 96149
rect -7370 96108 -7170 96154
rect -8399 95886 -8099 95932
rect -7370 95912 -7170 95958
rect -7040 95814 -6840 95860
rect -8399 95690 -8099 95736
rect -7370 95716 -7170 95762
rect -8936 95592 -8636 95638
rect -7040 95618 -6840 95664
rect -8399 95494 -8099 95540
rect -7370 95520 -7170 95566
rect -12993 93088 -10571 93201
rect -12993 89533 -12880 93088
rect -11479 92906 -11288 93057
rect -12772 92383 -12472 92429
rect -12772 92141 -12472 92187
rect -12772 91945 -12472 91991
rect -11454 92747 -11315 92906
rect -11466 92656 -11303 92747
rect -11050 92596 -10950 92642
rect -12160 92466 -11560 92512
rect -10684 92493 -10571 93088
rect -11050 92400 -10950 92446
rect -10819 92302 -10719 92348
rect -11050 92204 -10950 92250
rect -10819 92106 -10719 92152
rect -12160 92043 -11560 92089
rect -11050 92008 -10950 92054
rect -12160 91847 -11560 91893
rect -11049 91791 -10749 91837
rect -11748 91597 -11648 91643
rect -11049 91595 -10749 91641
rect -10512 91497 -10212 91543
rect -11748 91401 -11648 91447
rect -11049 91399 -10749 91445
rect -8234 91524 -7934 91570
rect -9230 91426 -8930 91472
rect -11979 91303 -11879 91349
rect -11748 91205 -11648 91251
rect -11979 91107 -11879 91153
rect -11748 91009 -11648 91055
rect -10920 91014 -10720 91060
rect -8234 91328 -7934 91374
rect -9230 91100 -8730 91146
rect -11949 90792 -11649 90838
rect -10920 90818 -10720 90864
rect -10590 90720 -10390 90766
rect -11949 90596 -11649 90642
rect -10920 90622 -10720 90668
rect -12486 90498 -12186 90544
rect -10590 90524 -10390 90570
rect -11949 90400 -11649 90446
rect -10920 90426 -10720 90472
rect -9230 90970 -8730 91016
rect -8434 91100 -7934 91146
rect -8434 90970 -7934 91016
rect -9230 90179 -8930 90225
rect -8434 90375 -7934 90421
rect -8434 90179 -7934 90225
rect -12993 89420 -10540 89533
rect -12993 88860 -12849 89420
rect -11401 89236 -11264 89332
rect -12962 88856 -12849 88860
rect -12741 88715 -12441 88761
rect -12741 88473 -12441 88519
rect -12741 88277 -12441 88323
rect -12129 88798 -11529 88844
rect -12129 88375 -11529 88421
rect -12129 88179 -11529 88225
rect -11375 88116 -11293 89236
rect -10653 89167 -10540 89420
rect -9509 89428 -7087 89541
rect -9509 89167 -9396 89428
rect -7995 89246 -7845 89356
rect -11019 88928 -10919 88974
rect -10653 89054 -9395 89167
rect -10653 88825 -10540 89054
rect -9509 88864 -9396 89054
rect -11019 88732 -10919 88778
rect -9288 88723 -8988 88769
rect -10788 88634 -10688 88680
rect -11019 88536 -10919 88582
rect -10788 88438 -10688 88484
rect -9288 88481 -8988 88527
rect -11019 88340 -10919 88386
rect -9288 88285 -8988 88331
rect -7977 89092 -7881 89246
rect -7983 89018 -7865 89092
rect -7566 88936 -7466 88982
rect -8676 88806 -8076 88852
rect -7200 88833 -7087 89428
rect -7566 88740 -7466 88786
rect -7335 88642 -7235 88688
rect -7566 88544 -7466 88590
rect -7335 88446 -7235 88492
rect -8676 88383 -8076 88429
rect -7566 88348 -7466 88394
rect -8676 88187 -8076 88233
rect -11018 88123 -10718 88169
rect -7565 88131 -7265 88177
rect -11717 87929 -11617 87975
rect -11382 87933 -11252 88116
rect -11018 87927 -10718 87973
rect -10481 87829 -10181 87875
rect -11717 87733 -11617 87779
rect -11018 87731 -10718 87777
rect -8264 87937 -8164 87983
rect -7565 87935 -7265 87981
rect -7028 87837 -6728 87883
rect -8264 87741 -8164 87787
rect -11948 87635 -11848 87681
rect -7565 87739 -7265 87785
rect -11717 87537 -11617 87583
rect -11948 87439 -11848 87485
rect -11717 87341 -11617 87387
rect -10889 87346 -10689 87392
rect -8495 87643 -8395 87689
rect -8264 87545 -8164 87591
rect -8495 87447 -8395 87493
rect -11918 87124 -11618 87170
rect -10889 87150 -10689 87196
rect -10559 87052 -10359 87098
rect -11918 86928 -11618 86974
rect -10889 86954 -10689 87000
rect -12455 86830 -12155 86876
rect -10559 86856 -10359 86902
rect -11918 86732 -11618 86778
rect -10889 86758 -10689 86804
rect -8264 87349 -8164 87395
rect -7436 87354 -7236 87400
rect -8465 87132 -8165 87178
rect -7436 87158 -7236 87204
rect -7106 87060 -6906 87106
rect -8465 86936 -8165 86982
rect -7436 86962 -7236 87008
rect -9002 86838 -8702 86884
rect -7106 86864 -6906 86910
rect -8465 86740 -8165 86786
rect -7436 86766 -7236 86812
rect -13027 83890 -10605 84003
rect -13027 80335 -12914 83890
rect -11513 83708 -11322 83859
rect -12806 83185 -12506 83231
rect -12806 82943 -12506 82989
rect -12806 82747 -12506 82793
rect -11488 83549 -11349 83708
rect -11500 83458 -11337 83549
rect -11084 83398 -10984 83444
rect -12194 83268 -11594 83314
rect -10718 83295 -10605 83890
rect -11084 83202 -10984 83248
rect -10853 83104 -10753 83150
rect -11084 83006 -10984 83052
rect -10853 82908 -10753 82954
rect -12194 82845 -11594 82891
rect -11084 82810 -10984 82856
rect -12194 82649 -11594 82695
rect -11083 82593 -10783 82639
rect -11782 82399 -11682 82445
rect -11083 82397 -10783 82443
rect -10546 82299 -10246 82345
rect -11782 82203 -11682 82249
rect -11083 82201 -10783 82247
rect -8268 82326 -7968 82372
rect -9264 82228 -8964 82274
rect -12013 82105 -11913 82151
rect -11782 82007 -11682 82053
rect -12013 81909 -11913 81955
rect -11782 81811 -11682 81857
rect -10954 81816 -10754 81862
rect -8268 82130 -7968 82176
rect -9264 81902 -8764 81948
rect -11983 81594 -11683 81640
rect -10954 81620 -10754 81666
rect -10624 81522 -10424 81568
rect -11983 81398 -11683 81444
rect -10954 81424 -10754 81470
rect -12520 81300 -12220 81346
rect -10624 81326 -10424 81372
rect -11983 81202 -11683 81248
rect -10954 81228 -10754 81274
rect -9264 81772 -8764 81818
rect -8468 81902 -7968 81948
rect -8468 81772 -7968 81818
rect -9264 80981 -8964 81027
rect -8468 81177 -7968 81223
rect -8468 80981 -7968 81027
rect -13027 80222 -10574 80335
rect -13027 79662 -12883 80222
rect -11435 80038 -11298 80134
rect -12996 79658 -12883 79662
rect -12775 79517 -12475 79563
rect -12775 79275 -12475 79321
rect -12775 79079 -12475 79125
rect -12163 79600 -11563 79646
rect -12163 79177 -11563 79223
rect -12163 78981 -11563 79027
rect -11409 78918 -11327 80038
rect -10687 79969 -10574 80222
rect -9543 80230 -7121 80343
rect -9543 79969 -9430 80230
rect -8029 80048 -7879 80158
rect -11053 79730 -10953 79776
rect -10687 79856 -9429 79969
rect -10687 79627 -10574 79856
rect -9543 79666 -9430 79856
rect -11053 79534 -10953 79580
rect -9322 79525 -9022 79571
rect -10822 79436 -10722 79482
rect -11053 79338 -10953 79384
rect -10822 79240 -10722 79286
rect -9322 79283 -9022 79329
rect -11053 79142 -10953 79188
rect -9322 79087 -9022 79133
rect -8011 79894 -7915 80048
rect -8017 79820 -7899 79894
rect -7600 79738 -7500 79784
rect -8710 79608 -8110 79654
rect -7234 79635 -7121 80230
rect -7600 79542 -7500 79588
rect -7369 79444 -7269 79490
rect -7600 79346 -7500 79392
rect -7369 79248 -7269 79294
rect -8710 79185 -8110 79231
rect -7600 79150 -7500 79196
rect -8710 78989 -8110 79035
rect -11052 78925 -10752 78971
rect -7599 78933 -7299 78979
rect -11751 78731 -11651 78777
rect -11416 78735 -11286 78918
rect -11052 78729 -10752 78775
rect -10515 78631 -10215 78677
rect -11751 78535 -11651 78581
rect -11052 78533 -10752 78579
rect -8298 78739 -8198 78785
rect -7599 78737 -7299 78783
rect -7062 78639 -6762 78685
rect -8298 78543 -8198 78589
rect -11982 78437 -11882 78483
rect -7599 78541 -7299 78587
rect -11751 78339 -11651 78385
rect -11982 78241 -11882 78287
rect -11751 78143 -11651 78189
rect -10923 78148 -10723 78194
rect -8529 78445 -8429 78491
rect -8298 78347 -8198 78393
rect -8529 78249 -8429 78295
rect -11952 77926 -11652 77972
rect -10923 77952 -10723 77998
rect -10593 77854 -10393 77900
rect -11952 77730 -11652 77776
rect -10923 77756 -10723 77802
rect -12489 77632 -12189 77678
rect -10593 77658 -10393 77704
rect -11952 77534 -11652 77580
rect -10923 77560 -10723 77606
rect -8298 78151 -8198 78197
rect -7470 78156 -7270 78202
rect -8499 77934 -8199 77980
rect -7470 77960 -7270 78006
rect -7140 77862 -6940 77908
rect -8499 77738 -8199 77784
rect -7470 77764 -7270 77810
rect -9036 77640 -8736 77686
rect -7140 77666 -6940 77712
rect -8499 77542 -8199 77588
rect -7470 77568 -7270 77614
rect -12988 75027 -10566 75140
rect -12988 71472 -12875 75027
rect -11474 74845 -11283 74996
rect -12767 74322 -12467 74368
rect -12767 74080 -12467 74126
rect -12767 73884 -12467 73930
rect -11449 74686 -11310 74845
rect -11461 74595 -11298 74686
rect -11045 74535 -10945 74581
rect -12155 74405 -11555 74451
rect -10679 74432 -10566 75027
rect -11045 74339 -10945 74385
rect -10814 74241 -10714 74287
rect -11045 74143 -10945 74189
rect -10814 74045 -10714 74091
rect -12155 73982 -11555 74028
rect -11045 73947 -10945 73993
rect -12155 73786 -11555 73832
rect -11044 73730 -10744 73776
rect -11743 73536 -11643 73582
rect -11044 73534 -10744 73580
rect -10507 73436 -10207 73482
rect -11743 73340 -11643 73386
rect -11044 73338 -10744 73384
rect -8229 73463 -7929 73509
rect -9225 73365 -8925 73411
rect -11974 73242 -11874 73288
rect -11743 73144 -11643 73190
rect -11974 73046 -11874 73092
rect -11743 72948 -11643 72994
rect -10915 72953 -10715 72999
rect -8229 73267 -7929 73313
rect -9225 73039 -8725 73085
rect -11944 72731 -11644 72777
rect -10915 72757 -10715 72803
rect -10585 72659 -10385 72705
rect -11944 72535 -11644 72581
rect -10915 72561 -10715 72607
rect -12481 72437 -12181 72483
rect -10585 72463 -10385 72509
rect -11944 72339 -11644 72385
rect -10915 72365 -10715 72411
rect -9225 72909 -8725 72955
rect -8429 73039 -7929 73085
rect -8429 72909 -7929 72955
rect -9225 72118 -8925 72164
rect -8429 72314 -7929 72360
rect -8429 72118 -7929 72164
rect -12988 71359 -10535 71472
rect -12988 70799 -12844 71359
rect -11396 71175 -11259 71271
rect -12957 70795 -12844 70799
rect -12736 70654 -12436 70700
rect -12736 70412 -12436 70458
rect -12736 70216 -12436 70262
rect -12124 70737 -11524 70783
rect -12124 70314 -11524 70360
rect -12124 70118 -11524 70164
rect -11370 70055 -11288 71175
rect -10648 71106 -10535 71359
rect -9504 71367 -7082 71480
rect -9504 71106 -9391 71367
rect -7990 71185 -7840 71295
rect -11014 70867 -10914 70913
rect -10648 70993 -9390 71106
rect -10648 70764 -10535 70993
rect -9504 70803 -9391 70993
rect -11014 70671 -10914 70717
rect -9283 70662 -8983 70708
rect -10783 70573 -10683 70619
rect -11014 70475 -10914 70521
rect -10783 70377 -10683 70423
rect -9283 70420 -8983 70466
rect -11014 70279 -10914 70325
rect -9283 70224 -8983 70270
rect -7972 71031 -7876 71185
rect -7978 70957 -7860 71031
rect -7561 70875 -7461 70921
rect -8671 70745 -8071 70791
rect -7195 70772 -7082 71367
rect -7561 70679 -7461 70725
rect -7330 70581 -7230 70627
rect -7561 70483 -7461 70529
rect -7330 70385 -7230 70431
rect -8671 70322 -8071 70368
rect -7561 70287 -7461 70333
rect -8671 70126 -8071 70172
rect -11013 70062 -10713 70108
rect -7560 70070 -7260 70116
rect -11712 69868 -11612 69914
rect -11377 69872 -11247 70055
rect -11013 69866 -10713 69912
rect -10476 69768 -10176 69814
rect -11712 69672 -11612 69718
rect -11013 69670 -10713 69716
rect -8259 69876 -8159 69922
rect -7560 69874 -7260 69920
rect -7023 69776 -6723 69822
rect -8259 69680 -8159 69726
rect -11943 69574 -11843 69620
rect -7560 69678 -7260 69724
rect -11712 69476 -11612 69522
rect -11943 69378 -11843 69424
rect -11712 69280 -11612 69326
rect -10884 69285 -10684 69331
rect -8490 69582 -8390 69628
rect -8259 69484 -8159 69530
rect -8490 69386 -8390 69432
rect -11913 69063 -11613 69109
rect -10884 69089 -10684 69135
rect -10554 68991 -10354 69037
rect -11913 68867 -11613 68913
rect -10884 68893 -10684 68939
rect -12450 68769 -12150 68815
rect -10554 68795 -10354 68841
rect -11913 68671 -11613 68717
rect -10884 68697 -10684 68743
rect -8259 69288 -8159 69334
rect -7431 69293 -7231 69339
rect -8460 69071 -8160 69117
rect -7431 69097 -7231 69143
rect -7101 68999 -6901 69045
rect -8460 68875 -8160 68921
rect -7431 68901 -7231 68947
rect -8997 68777 -8697 68823
rect -7101 68803 -6901 68849
rect -8460 68679 -8160 68725
rect -7431 68705 -7231 68751
rect -12977 66587 -10555 66700
rect -12977 63032 -12864 66587
rect -11463 66405 -11272 66556
rect -12756 65882 -12456 65928
rect -12756 65640 -12456 65686
rect -12756 65444 -12456 65490
rect -11438 66246 -11299 66405
rect -11450 66155 -11287 66246
rect -11034 66095 -10934 66141
rect -12144 65965 -11544 66011
rect -10668 65992 -10555 66587
rect -11034 65899 -10934 65945
rect -10803 65801 -10703 65847
rect -11034 65703 -10934 65749
rect -10803 65605 -10703 65651
rect -12144 65542 -11544 65588
rect -11034 65507 -10934 65553
rect -12144 65346 -11544 65392
rect -11033 65290 -10733 65336
rect -11732 65096 -11632 65142
rect -11033 65094 -10733 65140
rect -10496 64996 -10196 65042
rect -11732 64900 -11632 64946
rect -11033 64898 -10733 64944
rect -8218 65023 -7918 65069
rect -9214 64925 -8914 64971
rect -11963 64802 -11863 64848
rect -11732 64704 -11632 64750
rect -11963 64606 -11863 64652
rect -11732 64508 -11632 64554
rect -10904 64513 -10704 64559
rect -8218 64827 -7918 64873
rect -9214 64599 -8714 64645
rect -11933 64291 -11633 64337
rect -10904 64317 -10704 64363
rect -10574 64219 -10374 64265
rect -11933 64095 -11633 64141
rect -10904 64121 -10704 64167
rect -12470 63997 -12170 64043
rect -10574 64023 -10374 64069
rect -11933 63899 -11633 63945
rect -10904 63925 -10704 63971
rect -9214 64469 -8714 64515
rect -8418 64599 -7918 64645
rect -8418 64469 -7918 64515
rect -9214 63678 -8914 63724
rect -8418 63874 -7918 63920
rect -8418 63678 -7918 63724
rect -12977 62919 -10524 63032
rect -12977 62359 -12833 62919
rect -11385 62735 -11248 62831
rect -12946 62355 -12833 62359
rect -12725 62214 -12425 62260
rect -12725 61972 -12425 62018
rect -12725 61776 -12425 61822
rect -12113 62297 -11513 62343
rect -12113 61874 -11513 61920
rect -12113 61678 -11513 61724
rect -11359 61615 -11277 62735
rect -10637 62666 -10524 62919
rect -9493 62927 -7071 63040
rect -9493 62666 -9380 62927
rect -7979 62745 -7829 62855
rect -11003 62427 -10903 62473
rect -10637 62553 -9379 62666
rect -10637 62324 -10524 62553
rect -9493 62363 -9380 62553
rect -11003 62231 -10903 62277
rect -9272 62222 -8972 62268
rect -10772 62133 -10672 62179
rect -11003 62035 -10903 62081
rect -10772 61937 -10672 61983
rect -9272 61980 -8972 62026
rect -11003 61839 -10903 61885
rect -9272 61784 -8972 61830
rect -7961 62591 -7865 62745
rect -7967 62517 -7849 62591
rect -7550 62435 -7450 62481
rect -8660 62305 -8060 62351
rect -7184 62332 -7071 62927
rect -7550 62239 -7450 62285
rect -7319 62141 -7219 62187
rect -7550 62043 -7450 62089
rect -7319 61945 -7219 61991
rect -8660 61882 -8060 61928
rect -7550 61847 -7450 61893
rect -8660 61686 -8060 61732
rect -11002 61622 -10702 61668
rect -7549 61630 -7249 61676
rect -11701 61428 -11601 61474
rect -11366 61432 -11236 61615
rect -11002 61426 -10702 61472
rect -10465 61328 -10165 61374
rect -11701 61232 -11601 61278
rect -11002 61230 -10702 61276
rect -8248 61436 -8148 61482
rect -7549 61434 -7249 61480
rect -7012 61336 -6712 61382
rect -8248 61240 -8148 61286
rect -11932 61134 -11832 61180
rect -7549 61238 -7249 61284
rect -7203 61222 -7145 61301
rect -11701 61036 -11601 61082
rect -11932 60938 -11832 60984
rect -11701 60840 -11601 60886
rect -10873 60845 -10673 60891
rect -8479 61142 -8379 61188
rect -7203 61168 -7036 61222
rect -7203 61142 -7145 61168
rect -8248 61044 -8148 61090
rect -8479 60946 -8379 60992
rect -11902 60623 -11602 60669
rect -10873 60649 -10673 60695
rect -10543 60551 -10343 60597
rect -11902 60427 -11602 60473
rect -10873 60453 -10673 60499
rect -12439 60329 -12139 60375
rect -10543 60355 -10343 60401
rect -11902 60231 -11602 60277
rect -10873 60257 -10673 60303
rect -8248 60848 -8148 60894
rect -7420 60853 -7220 60899
rect -7090 60948 -7036 61168
rect -7090 60894 -6692 60948
rect -8449 60631 -8149 60677
rect -7420 60657 -7220 60703
rect -7090 60559 -6890 60605
rect -8449 60435 -8149 60481
rect -7420 60461 -7220 60507
rect -8986 60337 -8686 60383
rect -7090 60363 -6890 60409
rect -8449 60239 -8149 60285
rect -7420 60265 -7220 60311
rect -8613 59511 -8350 59770
rect -6746 59723 -6692 60894
rect -6786 59510 -6653 59723
rect -6834 58887 -6540 58922
rect -14196 58742 -6540 58887
rect -14196 58642 -6500 58742
rect -11273 57878 -10573 57924
rect -11273 57682 -10573 57728
rect -10388 57682 -9688 57728
rect -11273 57478 -10573 57524
rect -11273 57282 -10573 57328
rect -10388 57282 -9688 57328
rect -11273 56878 -10573 56924
rect -11273 56682 -10573 56728
rect -10388 56682 -9688 56728
rect -11273 56478 -10573 56524
rect -11273 56282 -10573 56328
rect -10388 56282 -9688 56328
rect -11273 55878 -10573 55924
rect -11273 55682 -10573 55728
rect -10388 55682 -9688 55728
rect -11273 55478 -10573 55524
rect -11273 55282 -10573 55328
rect -10388 55282 -9688 55328
rect -10043 54844 -9643 54890
rect -11344 54794 -11144 54840
rect -10964 54794 -10864 54840
rect -10043 54648 -9643 54694
rect -11344 54598 -11144 54644
rect -10964 54598 -10864 54644
rect -10497 54452 -10297 54498
rect -10043 54452 -9643 54498
rect -11344 54402 -11144 54448
rect -10964 54402 -10864 54448
rect -11351 53869 -11151 53915
rect -11351 53673 -11151 53719
rect -10643 53673 -10443 53719
rect -11351 53131 -11151 53177
rect -11351 52935 -11151 52981
rect -11351 52739 -11151 52785
rect -10744 52641 -10444 52687
rect -11351 52543 -11151 52589
rect -11317 51823 -10917 51869
rect -11317 51627 -10917 51673
rect -10625 51921 -10425 51967
rect -10625 51725 -10425 51771
rect -8053 57822 -7953 57868
rect -7773 57822 -7573 57868
rect -9091 57724 -8891 57770
rect -8711 57724 -8611 57770
rect -8554 57619 -8494 57643
rect -8276 57619 -8216 57634
rect -8053 57626 -7953 57672
rect -7773 57626 -7573 57672
rect -9091 57528 -8891 57574
rect -8711 57528 -8611 57574
rect -8554 57524 -8216 57619
rect -8554 57511 -8494 57524
rect -8276 57497 -8216 57524
rect -8053 57430 -7953 57476
rect -7773 57430 -7573 57476
rect -9091 57332 -8891 57378
rect -8711 57332 -8611 57378
rect -8053 56985 -7953 57031
rect -8053 56789 -7953 56835
rect -8053 56593 -7953 56639
rect -9091 55981 -8891 56027
rect -9091 55785 -8891 55831
rect -9091 55589 -8891 55635
rect -8711 55981 -8611 56027
rect -8711 55785 -8611 55831
rect -8711 55589 -8611 55635
rect -7773 56985 -7573 57031
rect -7773 56789 -7573 56835
rect -7773 56593 -7573 56639
rect -8365 55423 -8305 55472
rect -8813 55363 -8305 55423
rect -8365 55335 -8305 55363
rect -8053 55122 -7953 55168
rect -7773 55122 -7573 55168
rect -9091 55024 -8891 55070
rect -8711 55024 -8611 55070
rect -8550 55026 -8490 55044
rect -8282 55026 -8222 55037
rect -8550 54931 -8222 55026
rect -8550 54907 -8490 54931
rect -8282 54900 -8222 54931
rect -8053 54926 -7953 54972
rect -7773 54926 -7573 54972
rect -9091 54828 -8891 54874
rect -8711 54828 -8611 54874
rect -8053 54730 -7953 54776
rect -7773 54730 -7573 54776
rect -9091 54632 -8891 54678
rect -8711 54632 -8611 54678
rect -8366 54497 -8306 54526
rect -8366 54437 -7942 54497
rect -8366 54394 -8306 54437
rect -8053 54285 -7953 54331
rect -8053 54089 -7953 54135
rect -8053 53893 -7953 53939
rect -9091 53281 -8891 53327
rect -9091 53085 -8891 53131
rect -9091 52889 -8891 52935
rect -7773 54285 -7573 54331
rect -7773 54089 -7573 54135
rect -7773 53893 -7573 53939
rect -8711 53281 -8611 53327
rect -8711 53085 -8611 53131
rect -8711 52889 -8611 52935
rect -9091 52399 -8891 52445
rect -8711 52399 -8611 52445
rect -8551 52382 -8491 52417
rect -8282 52382 -8222 52399
rect -8551 52287 -8222 52382
rect -8551 52280 -8491 52287
rect -8282 52267 -8222 52287
rect -9091 52203 -8891 52249
rect -8711 52203 -8611 52249
rect -9091 52007 -8891 52053
rect -8711 52007 -8611 52053
rect -7981 52023 -7846 52053
rect -7981 51948 -7696 52023
rect -7981 51921 -7846 51948
rect -10625 50975 -10425 51021
rect -11317 50877 -10917 50923
rect -10625 50779 -10425 50825
rect -11317 50681 -10917 50727
rect -8007 50980 -7807 51026
rect -8971 50882 -8371 50928
rect -8007 50784 -7807 50830
rect -8971 50686 -8371 50732
rect -13647 49694 -13447 49740
rect -13267 49694 -13167 49740
rect -12609 49596 -12509 49642
rect -12329 49596 -12129 49642
rect -13647 49498 -13447 49544
rect -13267 49498 -13167 49544
rect -13004 49491 -12944 49506
rect -12726 49491 -12666 49515
rect -13004 49396 -12666 49491
rect -12609 49400 -12509 49446
rect -12329 49400 -12129 49446
rect -13004 49369 -12944 49396
rect -12726 49383 -12666 49396
rect -13647 49302 -13447 49348
rect -13267 49302 -13167 49348
rect -12609 49204 -12509 49250
rect -12329 49204 -12129 49250
rect -13647 48857 -13447 48903
rect -13647 48661 -13447 48707
rect -13647 48465 -13447 48511
rect -13267 48857 -13167 48903
rect -13267 48661 -13167 48707
rect -13267 48465 -13167 48511
rect -12609 47853 -12509 47899
rect -12609 47657 -12509 47703
rect -12609 47461 -12509 47507
rect -7771 50532 -7696 51948
rect -7809 50353 -7620 50532
rect -6852 48509 -6500 58642
rect -12329 47853 -12129 47899
rect -12329 47657 -12129 47703
rect -12329 47461 -12129 47507
rect -12915 47295 -12855 47344
rect -12915 47235 -12407 47295
rect -12915 47207 -12855 47235
rect -13647 46994 -13447 47040
rect -13267 46994 -13167 47040
rect -12998 46898 -12938 46909
rect -12730 46898 -12670 46916
rect -13647 46798 -13447 46844
rect -13267 46798 -13167 46844
rect -12998 46803 -12670 46898
rect -12609 46896 -12509 46942
rect -12329 46896 -12129 46942
rect -12998 46772 -12938 46803
rect -12730 46779 -12670 46803
rect -12609 46700 -12509 46746
rect -12329 46700 -12129 46746
rect -13647 46602 -13447 46648
rect -13267 46602 -13167 46648
rect -12609 46504 -12509 46550
rect -12329 46504 -12129 46550
rect -12914 46369 -12854 46398
rect -13278 46309 -12854 46369
rect -12914 46266 -12854 46309
rect -13647 46157 -13447 46203
rect -13647 45961 -13447 46007
rect -13647 45765 -13447 45811
rect -13267 46157 -13167 46203
rect -13267 45961 -13167 46007
rect -13267 45765 -13167 45811
rect -12609 45153 -12509 45199
rect -12609 44957 -12509 45003
rect -12609 44761 -12509 44807
rect -12329 45153 -12129 45199
rect -12329 44957 -12129 45003
rect -12329 44761 -12129 44807
rect -12998 44254 -12938 44271
rect -12729 44254 -12669 44289
rect -12609 44271 -12509 44317
rect -12329 44271 -12129 44317
rect -12998 44159 -12669 44254
rect -12998 44139 -12938 44159
rect -12729 44152 -12669 44159
rect -12609 44075 -12509 44121
rect -12329 44075 -12129 44121
rect -4820 44054 -3786 44102
rect -1993 44054 -862 44070
rect -12609 43879 -12509 43925
rect -12329 43879 -12129 43925
rect -16404 43172 -6583 43467
rect -14142 42120 -13873 43172
rect -16152 41899 -16029 41945
rect -16152 41839 -13944 41899
rect -16152 41822 -16029 41839
rect -15785 41758 -15662 41794
rect -15785 41694 -13980 41758
rect -15785 41692 -15489 41694
rect -15785 41671 -15661 41692
rect -15480 41641 -15362 41642
rect -15480 41580 -13984 41641
rect -15480 41512 -15361 41580
rect -15395 41511 -15361 41512
rect -15200 41528 -15077 41529
rect -15200 41467 -14130 41528
rect -15200 41405 -15077 41467
rect -14943 41428 -14820 41435
rect -14943 41421 -13987 41428
rect -14943 41377 -13984 41421
rect -14943 41368 -13987 41377
rect -14943 41312 -14820 41368
rect -14710 41320 -14587 41329
rect -14710 41259 -13983 41320
rect -14710 41206 -14587 41259
rect -13345 42808 -5537 42836
rect -13345 41329 -13317 42808
rect -13350 41264 -13213 41329
rect -13810 40649 -13610 40695
rect -13810 40453 -13610 40499
rect -13810 40340 -13610 40386
rect -13810 40144 -13610 40190
rect -13345 40466 -13317 41264
rect -13204 40649 -13004 40695
rect -13810 40030 -13610 40076
rect -13810 39834 -13610 39880
rect -13346 40327 -13292 40466
rect -13204 40340 -13004 40386
rect -13345 40225 -13315 40327
rect -13810 39638 -13610 39684
rect -13343 39388 -13315 40225
rect -13352 39249 -13298 39388
rect -13204 39276 -13004 39322
rect -13204 38862 -13004 38908
rect -12719 42657 -6163 42685
rect -12719 41438 -12691 42657
rect -12572 42498 -6310 42526
rect -12723 41299 -12676 41438
rect -12719 38686 -12691 41299
rect -13345 38658 -12691 38686
rect -12572 41756 -12544 42498
rect -12584 41612 -12537 41756
rect -13810 37649 -13610 37695
rect -13810 37453 -13610 37499
rect -13810 37340 -13610 37386
rect -13810 37144 -13610 37190
rect -13345 37466 -13317 38658
rect -13204 37649 -13004 37695
rect -13810 37030 -13610 37076
rect -13810 36834 -13610 36880
rect -13346 37327 -13292 37466
rect -13204 37340 -13004 37386
rect -13810 36638 -13610 36684
rect -13343 36388 -13315 37327
rect -13352 36249 -13298 36388
rect -13204 36276 -13004 36322
rect -13204 35862 -13004 35908
rect -12572 35365 -12544 41612
rect -13345 35337 -12544 35365
rect -13810 35149 -13610 35195
rect -13810 34953 -13610 34999
rect -13810 34840 -13610 34886
rect -13810 34644 -13610 34690
rect -13345 34966 -13317 35337
rect -13204 35149 -13004 35195
rect -13810 34530 -13610 34576
rect -13810 34334 -13610 34380
rect -13346 34827 -13292 34966
rect -13204 34840 -13004 34886
rect -13810 34138 -13610 34184
rect -13343 33888 -13315 34827
rect -13352 33749 -13298 33888
rect -13204 33776 -13004 33822
rect -13204 33362 -13004 33408
rect -13153 33134 -13017 33139
rect -12599 33138 -12537 33321
rect -12600 33134 -12537 33138
rect -13153 33020 -12537 33134
rect -13153 33016 -13017 33020
rect -12600 33015 -12537 33020
rect -12452 42336 -6430 42364
rect -12452 41881 -12424 42336
rect -12313 42169 -6569 42205
rect -12313 42046 -12277 42169
rect -12453 41738 -12406 41881
rect -12452 32899 -12424 41738
rect -12317 41898 -12269 42046
rect -13345 32871 -12424 32899
rect -13810 32649 -13610 32695
rect -13810 32453 -13610 32499
rect -13810 32340 -13610 32386
rect -13810 32144 -13610 32190
rect -13345 32466 -13317 32871
rect -13204 32649 -13004 32695
rect -13810 32030 -13610 32076
rect -13810 31834 -13610 31880
rect -13346 32327 -13292 32466
rect -13204 32340 -13004 32386
rect -13810 31638 -13610 31684
rect -13343 31388 -13315 32327
rect -13352 31249 -13298 31388
rect -13204 31276 -13004 31322
rect -13204 30862 -13004 30908
rect -13153 30651 -13017 30656
rect -12565 30651 -12429 30655
rect -13153 30537 -12429 30651
rect -13153 30533 -13017 30537
rect -12565 30532 -12429 30537
rect -12313 30415 -12277 41898
rect -13345 30387 -12277 30415
rect -13810 30149 -13610 30195
rect -13810 29953 -13610 29999
rect -13810 29840 -13610 29886
rect -13810 29644 -13610 29690
rect -13345 29966 -13317 30387
rect -13204 30149 -13004 30195
rect -13810 29530 -13610 29576
rect -13810 29334 -13610 29380
rect -13346 29827 -13292 29966
rect -13204 29840 -13004 29886
rect -13810 29138 -13610 29184
rect -13343 28888 -13315 29827
rect -13352 28749 -13298 28888
rect -13204 28776 -13004 28822
rect -13204 28362 -13004 28408
rect -13188 28084 -13052 28089
rect -12421 28084 -12285 28088
rect -13188 27970 -12285 28084
rect -13188 27966 -13052 27970
rect -12421 27965 -12285 27970
rect -12167 41987 -6715 42038
rect -12167 27858 -12116 41987
rect -12088 41913 -11981 41933
rect -12088 41862 -6972 41913
rect -12088 41742 -11981 41862
rect -13345 27830 -12116 27858
rect -13810 27649 -13610 27695
rect -13810 27453 -13610 27499
rect -13810 27340 -13610 27386
rect -13810 27144 -13610 27190
rect -13345 27466 -13317 27830
rect -13204 27649 -13004 27695
rect -13810 27030 -13610 27076
rect -13810 26834 -13610 26880
rect -13346 27327 -13292 27466
rect -13204 27340 -13004 27386
rect -13810 26638 -13610 26684
rect -13343 26388 -13315 27327
rect -13352 26249 -13298 26388
rect -13204 26276 -13004 26322
rect -13204 25862 -13004 25908
rect -11910 31950 -11859 41862
rect -11094 41708 -11066 41710
rect -7831 41708 -7780 41718
rect -11094 41680 -7780 41708
rect -11094 41593 -11066 41680
rect -7831 41667 -7780 41680
rect -11106 41448 -10971 41593
rect -11559 40659 -11359 40705
rect -11559 40463 -11359 40509
rect -11559 40350 -11359 40396
rect -11559 40154 -11359 40200
rect -11094 40476 -11066 41448
rect -10953 40659 -10753 40705
rect -8129 40659 -7929 40705
rect -7816 40476 -7788 41667
rect -7523 40659 -7323 40705
rect -11559 40040 -11359 40086
rect -11559 39844 -11359 39890
rect -11763 39653 -11627 39776
rect -11095 40337 -11041 40476
rect -10953 40350 -10753 40396
rect -8129 40350 -7929 40396
rect -7841 40337 -7787 40476
rect -11751 38560 -11646 39653
rect -11559 39648 -11359 39694
rect -11092 39398 -11064 40337
rect -11101 39259 -11047 39398
rect -10953 39286 -10753 39332
rect -8129 39286 -7929 39332
rect -7818 39398 -7790 40337
rect -7523 40463 -7323 40509
rect -7523 40350 -7323 40396
rect -7523 40154 -7323 40200
rect -7523 40040 -7323 40086
rect -7523 39844 -7323 39890
rect -7523 39648 -7323 39694
rect -7255 39653 -7119 39776
rect -7835 39259 -7781 39398
rect -10953 38872 -10753 38918
rect -8129 38872 -7929 38918
rect -11764 38437 -11628 38560
rect -11570 38487 -11370 38533
rect -7236 38560 -7131 39653
rect -7512 38487 -7312 38533
rect -7254 38437 -7118 38560
rect -10963 38389 -10663 38435
rect -8219 38389 -7919 38435
rect -11570 38291 -11370 38337
rect -7512 38291 -7312 38337
rect -11570 38095 -11370 38141
rect -7512 38095 -7312 38141
rect -11570 37899 -11370 37945
rect -7512 37899 -7312 37945
rect -11570 37357 -11370 37403
rect -10862 37357 -10662 37403
rect -8220 37357 -8020 37403
rect -7512 37357 -7312 37403
rect -11769 37081 -11633 37204
rect -11570 37161 -11370 37207
rect -7512 37161 -7312 37207
rect -11758 36803 -11651 37081
rect -11767 36680 -11631 36803
rect -11545 36734 -11245 36780
rect -11008 36636 -10708 36682
rect -11545 36538 -11245 36584
rect -11545 36342 -11245 36388
rect -11546 36125 -11446 36171
rect -11315 36027 -11215 36073
rect -11546 35929 -11446 35975
rect -11315 35831 -11215 35877
rect -11546 35733 -11446 35779
rect -11744 35452 -11608 35575
rect -11546 35537 -11446 35583
rect -11728 35186 -11621 35452
rect -11743 35063 -11607 35186
rect -11547 35129 -11247 35175
rect -11010 35031 -10710 35077
rect -11547 34933 -11247 34979
rect -11547 34737 -11247 34783
rect -11548 34520 -11448 34566
rect -11317 34422 -11217 34468
rect -11548 34324 -11448 34370
rect -11317 34226 -11217 34272
rect -11548 34128 -11448 34174
rect -11548 33932 -11448 33978
rect -7249 37081 -7113 37204
rect -7231 36803 -7124 37081
rect -7637 36734 -7337 36780
rect -8174 36636 -7874 36682
rect -7251 36680 -7115 36803
rect -7637 36538 -7337 36584
rect -7637 36342 -7337 36388
rect -7436 36125 -7336 36171
rect -7667 36027 -7567 36073
rect -7436 35929 -7336 35975
rect -7667 35831 -7567 35877
rect -7436 35733 -7336 35779
rect -7436 35537 -7336 35583
rect -7274 35452 -7138 35575
rect -7261 35186 -7154 35452
rect -7635 35129 -7335 35175
rect -8172 35031 -7872 35077
rect -7275 35063 -7139 35186
rect -7635 34933 -7335 34979
rect -7635 34737 -7335 34783
rect -7434 34520 -7334 34566
rect -7665 34422 -7565 34468
rect -7434 34324 -7334 34370
rect -7665 34226 -7565 34272
rect -7434 34128 -7334 34174
rect -7434 33932 -7334 33978
rect -11561 33525 -11361 33571
rect -7521 33525 -7321 33571
rect -10954 33427 -10654 33473
rect -8228 33427 -7928 33473
rect -11561 33329 -11361 33375
rect -7521 33329 -7321 33375
rect -11561 33133 -11361 33179
rect -7521 33133 -7321 33179
rect -11561 32937 -11361 32983
rect -7521 32937 -7321 32983
rect -11561 32395 -11361 32441
rect -10853 32395 -10653 32441
rect -8229 32395 -8029 32441
rect -7521 32395 -7321 32441
rect -11756 32085 -11620 32208
rect -11561 32199 -11361 32245
rect -11743 31914 -11628 32085
rect -11755 31791 -11619 31914
rect -11578 31857 -11378 31903
rect -11198 31857 -11098 31903
rect -11578 31661 -11378 31707
rect -11198 31661 -11098 31707
rect -11038 31623 -10978 31630
rect -10769 31623 -10709 31643
rect -11038 31528 -10709 31623
rect -11578 31465 -11378 31511
rect -11198 31465 -11098 31511
rect -11038 31493 -10978 31528
rect -10769 31511 -10709 31528
rect -7521 32199 -7321 32245
rect -7262 32085 -7126 32208
rect -7254 31914 -7139 32085
rect -7023 31950 -6972 41862
rect -7784 31857 -7684 31903
rect -7504 31857 -7304 31903
rect -8173 31753 -8113 31773
rect -7904 31753 -7844 31760
rect -7263 31791 -7127 31914
rect -8173 31658 -7844 31753
rect -7784 31661 -7684 31707
rect -7504 31661 -7304 31707
rect -8173 31641 -8113 31658
rect -7904 31623 -7844 31658
rect -7784 31465 -7684 31511
rect -7504 31465 -7304 31511
rect -11578 30975 -11378 31021
rect -11578 30779 -11378 30825
rect -11578 30583 -11378 30629
rect -11198 30975 -11098 31021
rect -11198 30779 -11098 30825
rect -11198 30583 -11098 30629
rect -10540 29971 -10440 30017
rect -10540 29775 -10440 29821
rect -10540 29579 -10440 29625
rect -7784 30975 -7684 31021
rect -7784 30779 -7684 30825
rect -7784 30583 -7684 30629
rect -10260 29971 -10060 30017
rect -8822 29971 -8622 30017
rect -10260 29775 -10060 29821
rect -8822 29775 -8622 29821
rect -10260 29579 -10060 29625
rect -8822 29579 -8622 29625
rect -7504 30975 -7304 31021
rect -7504 30779 -7304 30825
rect -7504 30583 -7304 30629
rect -8442 29971 -8342 30017
rect -8442 29775 -8342 29821
rect -8442 29579 -8342 29625
rect -10853 29473 -10793 29516
rect -10853 29413 -10429 29473
rect -10853 29384 -10793 29413
rect -11578 29232 -11378 29278
rect -11198 29232 -11098 29278
rect -7784 29232 -7684 29278
rect -7504 29232 -7304 29278
rect -10540 29134 -10440 29180
rect -10260 29134 -10060 29180
rect -8822 29134 -8622 29180
rect -8442 29134 -8342 29180
rect -11578 29036 -11378 29082
rect -11198 29036 -11098 29082
rect -7784 29036 -7684 29082
rect -7504 29036 -7304 29082
rect -11037 28979 -10977 29003
rect -10769 28979 -10709 29010
rect -11578 28840 -11378 28886
rect -11198 28840 -11098 28886
rect -11037 28884 -10709 28979
rect -10540 28938 -10440 28984
rect -10260 28938 -10060 28984
rect -8822 28938 -8622 28984
rect -8442 28938 -8342 28984
rect -8173 28979 -8113 29010
rect -7905 28979 -7845 29003
rect -11037 28866 -10977 28884
rect -10769 28873 -10709 28884
rect -8173 28884 -7845 28979
rect -8173 28873 -8113 28884
rect -7905 28866 -7845 28884
rect -7784 28840 -7684 28886
rect -7504 28840 -7304 28886
rect -10540 28742 -10440 28788
rect -10260 28742 -10060 28788
rect -8822 28742 -8622 28788
rect -8442 28742 -8342 28788
rect -10852 28547 -10792 28575
rect -11300 28487 -10792 28547
rect -10852 28438 -10792 28487
rect -11578 28275 -11378 28321
rect -11578 28079 -11378 28125
rect -11578 27883 -11378 27929
rect -11198 28275 -11098 28321
rect -11198 28079 -11098 28125
rect -11198 27883 -11098 27929
rect -10540 27271 -10440 27317
rect -10540 27075 -10440 27121
rect -10540 26879 -10440 26925
rect -10260 27271 -10060 27317
rect -8822 27271 -8622 27317
rect -10260 27075 -10060 27121
rect -8822 27075 -8622 27121
rect -10260 26879 -10060 26925
rect -8822 26879 -8622 26925
rect -7784 28275 -7684 28321
rect -7784 28079 -7684 28125
rect -7784 27883 -7684 27929
rect -7504 28275 -7304 28321
rect -7504 28079 -7304 28125
rect -7504 27883 -7304 27929
rect -8442 27271 -8342 27317
rect -8442 27075 -8342 27121
rect -8442 26879 -8342 26925
rect -8001 26761 -7941 26797
rect -8468 26701 -7941 26761
rect -8001 26665 -7941 26701
rect -11578 26532 -11378 26578
rect -11198 26532 -11098 26578
rect -7784 26532 -7684 26578
rect -7504 26532 -7304 26578
rect -10540 26434 -10440 26480
rect -10260 26434 -10060 26480
rect -8822 26434 -8622 26480
rect -8442 26434 -8342 26480
rect -11041 26386 -10981 26399
rect -10763 26386 -10703 26413
rect -11578 26336 -11378 26382
rect -11198 26336 -11098 26382
rect -11046 26291 -10703 26386
rect -8179 26386 -8119 26413
rect -7901 26386 -7841 26399
rect -11578 26140 -11378 26186
rect -11198 26140 -11098 26186
rect -11046 25899 -10951 26291
rect -10763 26276 -10703 26291
rect -8179 26291 -7841 26386
rect -7784 26336 -7684 26382
rect -7504 26336 -7304 26382
rect -10540 26238 -10440 26284
rect -10260 26238 -10060 26284
rect -8822 26238 -8622 26284
rect -8442 26238 -8342 26284
rect -8179 26276 -8119 26291
rect -7901 26267 -7841 26291
rect -7784 26140 -7684 26186
rect -7504 26140 -7304 26186
rect -10540 26042 -10440 26088
rect -10260 26042 -10060 26088
rect -8822 26042 -8622 26088
rect -8442 26042 -8342 26088
rect -11220 25804 -10951 25899
rect -11220 25589 -11125 25804
rect -6766 26224 -6715 41987
rect -6605 30415 -6569 42169
rect -6458 32899 -6430 42336
rect -6338 35365 -6310 42498
rect -6191 38686 -6163 42657
rect -5878 40649 -5678 40695
rect -5565 40466 -5537 42808
rect -4820 42503 -797 44054
rect -4820 42470 -3786 42503
rect -1993 42470 -862 42503
rect -5272 40649 -5072 40695
rect -5878 40340 -5678 40386
rect -5590 40327 -5536 40466
rect -5567 40225 -5537 40327
rect -5878 39276 -5678 39322
rect -5567 39388 -5539 40225
rect -5272 40453 -5072 40499
rect -5272 40340 -5072 40386
rect -5272 40144 -5072 40190
rect -5272 40030 -5072 40076
rect -5272 39834 -5072 39880
rect -5272 39638 -5072 39684
rect -5584 39249 -5530 39388
rect -5878 38862 -5678 38908
rect -6191 38658 -5537 38686
rect -5878 37649 -5678 37695
rect -5565 37466 -5537 38658
rect -5272 37649 -5072 37695
rect -5878 37340 -5678 37386
rect -5590 37327 -5536 37466
rect -5878 36276 -5678 36322
rect -5567 36388 -5539 37327
rect -5272 37453 -5072 37499
rect -5272 37340 -5072 37386
rect -5272 37144 -5072 37190
rect -5272 37030 -5072 37076
rect -5272 36834 -5072 36880
rect -5272 36638 -5072 36684
rect -5584 36249 -5530 36388
rect -5878 35862 -5678 35908
rect -6338 35337 -5537 35365
rect -5878 35149 -5678 35195
rect -5565 34966 -5537 35337
rect -5272 35149 -5072 35195
rect -5878 34840 -5678 34886
rect -5590 34827 -5536 34966
rect -5878 33776 -5678 33822
rect -5567 33888 -5539 34827
rect -5272 34953 -5072 34999
rect -5272 34840 -5072 34886
rect -5272 34644 -5072 34690
rect -5272 34530 -5072 34576
rect -5272 34334 -5072 34380
rect -5272 34138 -5072 34184
rect -5584 33749 -5530 33888
rect -6345 33138 -6283 33321
rect -5878 33362 -5678 33408
rect -6345 33134 -6282 33138
rect -5865 33134 -5729 33139
rect -6345 33020 -5729 33134
rect -6345 33015 -6282 33020
rect -5865 33016 -5729 33020
rect -6458 32871 -5537 32899
rect -5878 32649 -5678 32695
rect -5565 32466 -5537 32871
rect -5272 32649 -5072 32695
rect -5878 32340 -5678 32386
rect -5590 32327 -5536 32466
rect -5878 31276 -5678 31322
rect -5567 31388 -5539 32327
rect -5272 32453 -5072 32499
rect -5272 32340 -5072 32386
rect -5272 32144 -5072 32190
rect -5272 32030 -5072 32076
rect -5272 31834 -5072 31880
rect -5272 31638 -5072 31684
rect -5584 31249 -5530 31388
rect -5878 30862 -5678 30908
rect -6453 30651 -6317 30655
rect -5865 30651 -5729 30656
rect -6453 30537 -5729 30651
rect -6453 30532 -6317 30537
rect -5865 30533 -5729 30537
rect -6605 30387 -5537 30415
rect -5878 30149 -5678 30195
rect -5565 29966 -5537 30387
rect -5272 30149 -5072 30195
rect -5878 29840 -5678 29886
rect -5590 29827 -5536 29966
rect -5878 28776 -5678 28822
rect -5567 28888 -5539 29827
rect -5272 29953 -5072 29999
rect -5272 29840 -5072 29886
rect -5272 29644 -5072 29690
rect -5272 29530 -5072 29576
rect -5272 29334 -5072 29380
rect -5272 29138 -5072 29184
rect -5584 28749 -5530 28888
rect -5878 28362 -5678 28408
rect -6597 28084 -6461 28088
rect -5830 28084 -5694 28089
rect -6597 27970 -5694 28084
rect -6597 27965 -6461 27970
rect -5830 27966 -5694 27970
rect -5878 27649 -5678 27695
rect -5272 27649 -5072 27695
rect -5878 27340 -5678 27386
rect -6601 26691 -6401 26737
rect -6221 26691 -6121 26737
rect -6601 26495 -6401 26541
rect -6221 26495 -6121 26541
rect -6601 26299 -6401 26345
rect -6333 26224 -6259 26309
rect -6221 26299 -6121 26345
rect -5878 26276 -5678 26322
rect -6766 26173 -6259 26224
rect -5272 27453 -5072 27499
rect -5272 27340 -5072 27386
rect -5272 27144 -5072 27190
rect -5272 27030 -5072 27076
rect -5272 26834 -5072 26880
rect -5272 26638 -5072 26684
rect -5878 25862 -5678 25908
rect -10410 25176 -9810 25222
rect -5476 25149 -4876 25195
rect -11022 25078 -10722 25124
rect -6088 25051 -5788 25097
rect -10410 24980 -9810 25026
rect -5476 24953 -4876 24999
rect -11022 24882 -10722 24928
rect -6088 24855 -5788 24901
rect -11022 24640 -10722 24686
rect -6088 24613 -5788 24659
rect -10410 24557 -9810 24603
rect -5476 24530 -4876 24576
rect -6782 24284 -6669 24285
rect -4604 24284 -4414 41117
rect -3742 40236 -2527 40571
rect -3742 39356 -2367 40236
rect -6782 24189 -4414 24284
rect -11311 23983 -11111 24029
rect -10931 23983 -10831 24029
rect -11311 23787 -11111 23833
rect -10931 23787 -10831 23833
rect -10771 23749 -10711 23756
rect -10502 23749 -10442 23769
rect -6782 23749 -6669 24189
rect -6384 23983 -6184 24029
rect -6004 23983 -5904 24029
rect -6384 23787 -6184 23833
rect -6004 23787 -5904 23833
rect -10771 23654 -6669 23749
rect -5844 23749 -5784 23756
rect -5735 23749 -5640 24189
rect -5575 23749 -5515 23769
rect -11311 23591 -11111 23637
rect -10931 23591 -10831 23637
rect -10771 23619 -10711 23654
rect -10502 23637 -10442 23654
rect -11311 23101 -11111 23147
rect -11311 22905 -11111 22951
rect -11311 22709 -11111 22755
rect -10931 23101 -10831 23147
rect -10931 22905 -10831 22951
rect -10931 22709 -10831 22755
rect -10273 22097 -10173 22143
rect -10273 21901 -10173 21947
rect -10273 21705 -10173 21751
rect -9993 22097 -9793 22143
rect -6782 21994 -6669 23654
rect -5844 23654 -5515 23749
rect -6384 23591 -6184 23637
rect -6004 23591 -5904 23637
rect -5844 23619 -5784 23654
rect -5575 23637 -5515 23654
rect -9993 21901 -9793 21947
rect -9091 21881 -6669 21994
rect -9993 21705 -9793 21751
rect -11311 21358 -11111 21404
rect -10931 21358 -10831 21404
rect -10273 21260 -10173 21306
rect -9993 21260 -9793 21306
rect -9091 21286 -8978 21881
rect -8712 21389 -8612 21435
rect -8102 21259 -7502 21305
rect -11311 21162 -11111 21208
rect -10931 21162 -10831 21208
rect -8712 21193 -8612 21239
rect -10770 21105 -10710 21129
rect -10502 21105 -10442 21136
rect -11311 20966 -11111 21012
rect -10931 20966 -10831 21012
rect -10770 21010 -10442 21105
rect -10273 21064 -10173 21110
rect -9993 21064 -9793 21110
rect -8943 21095 -8843 21141
rect -10770 20992 -10710 21010
rect -10502 20999 -10442 21010
rect -8712 20997 -8612 21043
rect -10273 20868 -10173 20914
rect -9993 20868 -9793 20914
rect -8943 20899 -8843 20945
rect -8712 20801 -8612 20847
rect -8102 20836 -7502 20882
rect -8102 20640 -7502 20686
rect -6782 21317 -6669 21881
rect -7190 21176 -6890 21222
rect -7190 20934 -6890 20980
rect -7190 20738 -6890 20784
rect -8913 20584 -8613 20630
rect -11311 20401 -11111 20447
rect -11311 20205 -11111 20251
rect -11311 20009 -11111 20055
rect -10931 20401 -10831 20447
rect -10931 20205 -10831 20251
rect -10931 20009 -10831 20055
rect -8913 20388 -8613 20434
rect -8014 20390 -7914 20436
rect -9450 20290 -9150 20336
rect -8913 20192 -8613 20238
rect -8014 20194 -7914 20240
rect -7783 20096 -7683 20142
rect -8014 19998 -7914 20044
rect -10273 19397 -10173 19443
rect -10273 19201 -10173 19247
rect -10273 19005 -10173 19051
rect -9993 19397 -9793 19443
rect -9993 19201 -9793 19247
rect -9993 19005 -9793 19051
rect -11311 18658 -11111 18704
rect -10931 18658 -10831 18704
rect -10273 18560 -10173 18606
rect -9993 18560 -9793 18606
rect -10774 18512 -10714 18525
rect -10496 18512 -10436 18539
rect -11311 18462 -11111 18508
rect -10931 18462 -10831 18508
rect -10774 18417 -10436 18512
rect -10774 18393 -10714 18417
rect -10496 18402 -10436 18417
rect -10273 18364 -10173 18410
rect -9993 18364 -9793 18410
rect -11311 18266 -11111 18312
rect -10931 18266 -10831 18312
rect -10273 18168 -10173 18214
rect -9993 18168 -9793 18214
rect -7783 19900 -7683 19946
rect -8942 19807 -8742 19853
rect -8014 19802 -7914 19848
rect -8942 19611 -8742 19657
rect -6384 23101 -6184 23147
rect -6384 22905 -6184 22951
rect -6384 22709 -6184 22755
rect -6004 23101 -5904 23147
rect -6004 22905 -5904 22951
rect -6004 22709 -5904 22755
rect -5346 22097 -5246 22143
rect -5346 21901 -5246 21947
rect -5346 21705 -5246 21751
rect -5066 22097 -4866 22143
rect -5066 21901 -4866 21947
rect -5066 21705 -4866 21751
rect -6384 21358 -6184 21404
rect -6004 21358 -5904 21404
rect -5346 21260 -5246 21306
rect -5066 21260 -4866 21306
rect -6384 21162 -6184 21208
rect -6004 21162 -5904 21208
rect -5843 21105 -5783 21129
rect -5575 21105 -5515 21136
rect -6384 20966 -6184 21012
rect -6004 20966 -5904 21012
rect -5843 21010 -5515 21105
rect -5346 21064 -5246 21110
rect -5066 21064 -4866 21110
rect -5843 20992 -5783 21010
rect -5575 20999 -5515 21010
rect -5346 20868 -5246 20914
rect -5066 20868 -4866 20914
rect -6384 20401 -6184 20447
rect -6384 20205 -6184 20251
rect -6384 20009 -6184 20055
rect -6004 20401 -5904 20447
rect -6004 20205 -5904 20251
rect -6004 20009 -5904 20055
rect -8013 19585 -7713 19631
rect -9272 19513 -9072 19559
rect -8942 19415 -8742 19461
rect -8013 19389 -7713 19435
rect -9272 19317 -9072 19363
rect -7476 19291 -7176 19337
rect -8942 19219 -8742 19265
rect -8013 19193 -7713 19239
rect -5346 19397 -5246 19443
rect -9126 19135 -8976 19161
rect -9126 19081 -7518 19135
rect -9126 19031 -8976 19081
rect -8779 17646 -8603 19081
rect -7572 18938 -7518 19081
rect -5346 19201 -5246 19247
rect -5346 19005 -5246 19051
rect -5066 19397 -4866 19443
rect -5066 19201 -4866 19247
rect -5066 19005 -4866 19051
rect -6384 18658 -6184 18704
rect -6004 18658 -5904 18704
rect -5346 18560 -5246 18606
rect -5066 18560 -4866 18606
rect -5847 18512 -5787 18525
rect -5569 18512 -5509 18539
rect -6384 18462 -6184 18508
rect -6004 18462 -5904 18508
rect -5847 18417 -5509 18512
rect -5847 18393 -5787 18417
rect -5569 18402 -5509 18417
rect -5346 18364 -5246 18410
rect -5066 18364 -4866 18410
rect -6384 18266 -6184 18312
rect -6004 18266 -5904 18312
rect -5346 18168 -5246 18214
rect -5066 18168 -4866 18214
rect -14518 17470 -8603 17646
rect -13115 16899 -5693 17005
rect -4604 16899 -4414 24189
rect -13115 16892 -4414 16899
rect -13115 16297 -13002 16892
rect -12736 16400 -12636 16446
rect -12126 16270 -11526 16316
rect -12736 16204 -12636 16250
rect -12967 16106 -12867 16152
rect -12736 16008 -12636 16054
rect -12967 15910 -12867 15956
rect -12736 15812 -12636 15858
rect -12126 15847 -11526 15893
rect -12126 15651 -11526 15697
rect -10806 16328 -10693 16892
rect -8115 16297 -8002 16892
rect -5806 16709 -4414 16892
rect -7736 16400 -7636 16446
rect -11214 16187 -10914 16233
rect -7126 16270 -6526 16316
rect -7736 16204 -7636 16250
rect -7967 16106 -7867 16152
rect -7736 16008 -7636 16054
rect -11214 15945 -10914 15991
rect -7967 15910 -7867 15956
rect -7736 15812 -7636 15858
rect -7126 15847 -6526 15893
rect -11214 15749 -10914 15795
rect -7126 15651 -6526 15697
rect -5806 16328 -5693 16709
rect -6214 16187 -5914 16233
rect -6214 15945 -5914 15991
rect -6214 15749 -5914 15795
rect -12937 15595 -12637 15641
rect -7937 15595 -7637 15641
rect -12937 15399 -12637 15445
rect -12038 15401 -11938 15447
rect -13474 15301 -13174 15347
rect -7937 15399 -7637 15445
rect -7038 15401 -6938 15447
rect -12937 15203 -12637 15249
rect -12038 15205 -11938 15251
rect -8474 15301 -8174 15347
rect -7937 15203 -7637 15249
rect -7038 15205 -6938 15251
rect -11807 15107 -11707 15153
rect -12038 15009 -11938 15055
rect -11807 14911 -11707 14957
rect -6807 15107 -6707 15153
rect -7038 15009 -6938 15055
rect -12966 14818 -12766 14864
rect -12038 14813 -11938 14859
rect -12966 14622 -12766 14668
rect -12037 14596 -11737 14642
rect -13296 14524 -13096 14570
rect -12966 14426 -12766 14472
rect -12037 14400 -11737 14446
rect -13296 14328 -13096 14374
rect -11500 14302 -11200 14348
rect -12966 14230 -12766 14276
rect -12037 14204 -11737 14250
rect -12434 13896 -12262 13961
rect -6807 14911 -6707 14957
rect -7966 14818 -7766 14864
rect -7038 14813 -6938 14859
rect -7966 14622 -7766 14668
rect -7037 14596 -6737 14642
rect -8296 14524 -8096 14570
rect -7966 14426 -7766 14472
rect -7037 14400 -6737 14446
rect -8296 14328 -8096 14374
rect -6500 14302 -6200 14348
rect -7966 14230 -7766 14276
rect -7037 14204 -6737 14250
rect -10498 13896 -10331 13922
rect -12434 13770 -10331 13896
rect -12434 13769 -12262 13770
rect -10498 13743 -10331 13770
rect -7789 13725 -7589 13771
rect -5874 13765 -5774 13811
rect -8497 13529 -8297 13575
rect -7789 13529 -7589 13575
rect -14060 12964 -13429 13140
rect -11700 13096 -11500 13142
rect -11208 12998 -10808 13044
rect -7789 12987 -7589 13033
rect -11700 12900 -11500 12946
rect -11208 12802 -10808 12848
rect -7789 12791 -7589 12837
rect -12650 12751 -12513 12768
rect -11542 12751 -11405 12774
rect -12650 12716 -11405 12751
rect -12650 12710 -12513 12716
rect -12573 12674 -12436 12675
rect -11370 12674 -11233 12697
rect -12573 12639 -11233 12674
rect -12573 12617 -12436 12639
rect -7789 12595 -7589 12641
rect -8496 12497 -8196 12543
rect -7789 12399 -7589 12445
rect -11699 12191 -11499 12237
rect -5874 13569 -5774 13615
rect -6105 13471 -6005 13517
rect -5874 13373 -5774 13419
rect -6105 13275 -6005 13321
rect -5874 13177 -5774 13223
rect -6075 12960 -5775 13006
rect -6075 12764 -5775 12810
rect -6612 12666 -6312 12712
rect -6075 12568 -5775 12614
rect -6278 12401 -6220 12491
rect -7100 12377 -6220 12401
rect -7104 12361 -6220 12377
rect -7104 12245 -7051 12361
rect -6278 12354 -6220 12361
rect -7013 12267 -6881 12282
rect -6171 12267 -6113 12396
rect -7013 12259 -6113 12267
rect -7100 12198 -7060 12245
rect -7013 12231 -6130 12259
rect -7013 12229 -6881 12231
rect -11207 12093 -10807 12139
rect -11699 11995 -11499 12041
rect -11207 11897 -10807 11943
rect -12494 11840 -12357 11854
rect -11540 11840 -11403 11856
rect -12494 11798 -11403 11840
rect -12494 11797 -11407 11798
rect -12494 11796 -12357 11797
rect -13896 11680 -13696 11726
rect -12415 11758 -12278 11761
rect -11369 11758 -11232 11781
rect -12415 11723 -11232 11758
rect -7783 11823 -7683 11869
rect -5853 11895 -5653 11941
rect -12415 11703 -12278 11723
rect -6561 11699 -6361 11745
rect -5853 11699 -5653 11745
rect -13289 11582 -12989 11628
rect -7783 11627 -7683 11673
rect -13896 11484 -13696 11530
rect -8014 11529 -7914 11575
rect -12815 11416 -12700 11425
rect -12288 11416 -12138 11459
rect -13896 11288 -13696 11334
rect -12815 11329 -12138 11416
rect -7783 11431 -7683 11477
rect -12815 11291 -12700 11329
rect -12288 11291 -12138 11329
rect -8014 11333 -7914 11379
rect -12815 11204 -12138 11291
rect -13896 11092 -13696 11138
rect -12815 11107 -12700 11204
rect -12288 11107 -12138 11204
rect -7783 11235 -7683 11281
rect -5853 11157 -5653 11203
rect -12815 11020 -12138 11107
rect -12815 10934 -12700 11020
rect -12288 10934 -12138 11020
rect -12042 10985 -11842 11031
rect -7984 11018 -7684 11064
rect -12815 10847 -12138 10934
rect -11478 10887 -10878 10933
rect -12815 10754 -12700 10847
rect -12288 10754 -12138 10847
rect -5853 10961 -5653 11007
rect -12042 10789 -11842 10835
rect -7984 10822 -7684 10868
rect -12815 10667 -12138 10754
rect -11478 10691 -10878 10737
rect -13896 10550 -13696 10596
rect -13188 10550 -12988 10596
rect -12815 10442 -12700 10667
rect -12288 10655 -12138 10667
rect -8521 10724 -8221 10770
rect -5853 10765 -5653 10811
rect -7984 10626 -7684 10672
rect -6560 10667 -6260 10713
rect -5853 10569 -5653 10615
rect -13896 10354 -13696 10400
rect -16157 10260 -16034 10306
rect -16157 10200 -7840 10260
rect -16157 10183 -16034 10200
rect -15790 10119 -15667 10155
rect -15790 10055 -8271 10119
rect -15790 10053 -15494 10055
rect -15790 10032 -15666 10053
rect -15485 10002 -15367 10003
rect -15485 9941 -6799 10002
rect -15485 9873 -15366 9941
rect -15400 9872 -15366 9873
rect -15205 9889 -15082 9890
rect -15205 9828 -6866 9889
rect -15205 9766 -15082 9828
rect -14948 9789 -14825 9796
rect -12005 9789 -11768 9790
rect -5939 9789 -5701 9790
rect -14948 9729 -5701 9789
rect -14948 9673 -14825 9729
rect -14715 9681 -14592 9690
rect -14715 9620 -5787 9681
rect -14715 9567 -14592 9620
rect -14516 9490 -14393 9499
rect -14516 9429 -5866 9490
rect -14516 9376 -14393 9429
rect -7268 9369 -7025 9382
rect -16414 9265 -16236 9325
rect -7311 9281 -7025 9369
rect -7311 9265 -7080 9281
rect -17836 9129 -7080 9265
rect -17836 565 -17700 9129
rect -16414 9112 -16236 9129
rect -16277 8494 -5438 8555
rect -16277 8032 -5433 8494
rect -6540 7273 -5433 8032
rect -12975 3566 -11404 6943
rect -3582 5554 -2367 39356
rect 16949 11350 17282 16839
rect 15933 10178 16018 10179
rect 15588 10127 15788 10173
rect 15933 10132 16218 10178
rect 16818 10132 17018 10178
rect 14785 9869 14985 9915
rect 15933 9663 15979 10132
rect 15933 9662 16018 9663
rect 15588 9611 15788 9657
rect 15933 9616 16218 9662
rect 16818 9616 17018 9662
rect 14785 9353 14985 9399
rect 15933 9146 15979 9616
rect 15588 9095 15788 9141
rect 15933 9100 16218 9146
rect 16818 9100 17018 9146
rect 3375 7565 4103 8200
rect 2866 4116 3250 4560
rect -13122 3329 -8953 3566
rect -13011 2361 -12663 3329
rect -11909 2361 -11561 3329
rect -11015 2361 -10667 3329
rect -10239 2361 -9891 3329
rect -9633 2361 -9285 3329
rect -13395 2124 -9226 2361
rect -13415 1504 -13369 1975
rect -13297 1575 -13251 1975
rect -13179 1504 -13133 1975
rect -13061 1575 -13015 1975
rect -12943 1504 -12897 1975
rect -12825 1575 -12779 1975
rect -12707 1504 -12661 1975
rect -12589 1575 -12543 1975
rect -12471 1504 -12425 1975
rect -12353 1575 -12307 1975
rect -12235 1504 -12189 1975
rect -12117 1575 -12071 1975
rect -11999 1504 -11953 1975
rect -11881 1575 -11835 1975
rect -11763 1504 -11717 1975
rect -11645 1575 -11599 1975
rect -11527 1504 -11481 1975
rect -11409 1575 -11363 1975
rect -11291 1504 -11245 1975
rect -11173 1575 -11127 1975
rect -11055 1504 -11009 1975
rect -10937 1575 -10891 1975
rect -10819 1504 -10773 1975
rect -10701 1575 -10655 1975
rect -10583 1504 -10537 1975
rect -10465 1575 -10419 1975
rect -10347 1504 -10301 1975
rect -10229 1575 -10183 1975
rect -10111 1504 -10065 1975
rect -9993 1575 -9947 1975
rect -9875 1504 -9829 1975
rect -9757 1575 -9711 1975
rect -9639 1504 -9593 1975
rect -9509 1575 -9463 1975
rect -9273 1575 -9227 1975
rect -9037 1575 -8991 1975
rect -8801 1575 -8755 1975
rect -8565 1575 -8519 1975
rect -8329 1575 -8283 1975
rect -8093 1575 -8047 1975
rect -7857 1575 -7811 1975
rect -7621 1575 -7575 1975
rect -7491 1575 -7445 1975
rect -7255 1575 -7209 1975
rect -7019 1575 -6973 1975
rect -6783 1575 -6737 1975
rect -6547 1575 -6501 1975
rect -6417 1575 -6371 1975
rect -6181 1575 -6135 1975
rect -5945 1575 -5899 1975
rect -3590 1837 -3544 2037
rect -3394 1837 -3348 2037
rect -3198 1837 -3152 2037
rect -2740 1837 -2694 2037
rect -2544 1837 -2498 2037
rect -2348 1837 -2302 2037
rect -13444 1430 -9567 1504
rect -9659 1314 -9613 1430
rect -9659 1268 -7961 1314
rect -9659 767 -9613 1268
rect -9423 767 -9377 1268
rect -9187 767 -9141 1268
rect -8951 767 -8905 1268
rect -8715 767 -8669 1268
rect -8479 767 -8433 1268
rect -8243 767 -8197 1268
rect -8007 767 -7961 1268
rect 3061 2508 3235 4116
rect 2809 2392 3235 2508
rect 2391 2356 3235 2392
rect 707 2001 753 2085
rect 1219 1990 1265 2110
rect 1509 1995 1555 2115
rect -2849 1278 -2047 1322
rect -5243 1178 -3681 1219
rect -2849 1178 -2805 1278
rect -5243 1134 -2805 1178
rect -5243 1073 -3681 1134
rect -2094 1108 -2048 1278
rect -18039 321 -17604 565
rect -5243 473 -5078 1073
rect -1898 1108 -1852 1308
rect -1702 1108 -1656 1308
rect -1506 1108 -1460 1308
rect -1310 1108 -1264 1308
rect -2740 762 -2694 962
rect -2544 762 -2498 962
rect -2348 762 -2302 962
rect -2094 762 -2048 962
rect -1898 762 -1852 962
rect -1702 762 -1656 962
rect -1506 762 -1460 962
rect -1310 762 -1264 962
rect -6599 389 -5077 473
rect -6600 308 -5077 389
rect 707 1653 753 1821
rect 1941 1970 1987 2122
rect 2177 1970 2223 2122
rect 2391 1970 2427 2356
rect 2809 2272 3235 2356
rect 2494 2001 2540 2085
rect 2803 1970 2849 2085
rect 1941 1934 2849 1970
rect 1043 1699 1089 1819
rect 1219 1699 1265 1819
rect 1395 1699 1441 1819
rect 1684 1639 1730 1819
rect 1830 1639 1876 1819
rect 2494 1653 2540 1821
rect 2803 1653 2849 1821
rect 707 1041 753 1209
rect 1043 1043 1089 1163
rect 1219 1043 1265 1163
rect 1395 1043 1441 1163
rect 1684 1043 1730 1223
rect 1830 1043 1876 1223
rect 707 777 753 861
rect 2494 1041 2540 1209
rect 2803 1041 2849 1209
rect 3061 1159 3235 2272
rect 3500 1279 3875 7565
rect 4509 2013 4555 2213
rect 4705 2013 4751 2213
rect 4901 2013 4947 2213
rect 5359 2013 5405 2213
rect 5555 2013 5601 2213
rect 5751 2013 5797 2213
rect 4509 1733 4555 1833
rect 4705 1733 4751 1833
rect 4901 1733 4947 1833
rect 5359 1733 5405 1833
rect 5555 1733 5601 1833
rect 5751 1733 5797 1833
rect 8138 6696 8184 7496
rect 9854 6696 9900 7496
rect 11570 6696 11616 7496
rect 11700 6696 11746 7496
rect 12616 6696 12662 7496
rect 8174 5643 8220 6443
rect 9890 5643 9936 6443
rect 11606 5643 11652 6443
rect 14484 7856 14591 7858
rect 14484 7749 14796 7856
rect 14484 7642 14795 7749
rect 14484 6213 14653 7642
rect 16043 9012 16101 9100
rect 17131 9012 17318 9181
rect 15726 8966 15886 9012
rect 16033 8966 17318 9012
rect 17202 8956 17318 8966
rect 14443 6016 14691 6213
rect 8174 4643 8220 5443
rect 9032 4643 9078 5443
rect 9890 4643 9936 5443
rect 10748 4643 10794 5443
rect 11606 4643 11652 5443
rect 15814 3722 16331 4171
rect 7612 1857 7658 2257
rect 7848 1857 7894 2257
rect 8084 1857 8130 2257
rect 8214 1857 8260 2257
rect 8450 1857 8496 2257
rect 8686 1857 8732 2257
rect 8922 1857 8968 2257
rect 9158 1857 9204 2257
rect 9288 1857 9334 2257
rect 9524 1857 9570 2257
rect 9760 1857 9806 2257
rect 9996 1857 10042 2257
rect 10232 1857 10278 2257
rect 10468 1857 10514 2257
rect 10704 1857 10750 2257
rect 10940 1857 10986 2257
rect 11176 1857 11222 2257
rect 11306 1786 11352 2257
rect 11424 1857 11470 2257
rect 11542 1786 11588 2257
rect 11660 1857 11706 2257
rect 11778 1786 11824 2257
rect 11896 1857 11942 2257
rect 12014 1786 12060 2257
rect 12132 1857 12178 2257
rect 12250 1786 12296 2257
rect 12368 1857 12414 2257
rect 12486 1786 12532 2257
rect 12604 1857 12650 2257
rect 12722 1786 12768 2257
rect 12840 1857 12886 2257
rect 12958 1786 13004 2257
rect 13076 1857 13122 2257
rect 13194 1786 13240 2257
rect 13312 1857 13358 2257
rect 13430 1786 13476 2257
rect 13548 1857 13594 2257
rect 13666 1786 13712 2257
rect 13784 1857 13830 2257
rect 13902 1786 13948 2257
rect 14020 1857 14066 2257
rect 14138 1786 14184 2257
rect 14256 1857 14302 2257
rect 14374 1786 14420 2257
rect 14492 1857 14538 2257
rect 14610 1786 14656 2257
rect 14728 1857 14774 2257
rect 14846 1786 14892 2257
rect 14964 1857 15010 2257
rect 15082 1786 15128 2257
rect 11280 1712 15157 1786
rect 4186 1385 4963 1519
rect 5250 1454 6052 1498
rect 4580 1384 4827 1385
rect 5250 1354 5294 1454
rect 4064 1310 5294 1354
rect 5359 1318 5405 1418
rect 5555 1318 5601 1418
rect 5751 1318 5797 1418
rect 3061 1101 3899 1159
rect 1219 752 1265 872
rect 1509 747 1555 867
rect 1941 892 2849 928
rect 1941 740 1987 892
rect 2177 740 2223 892
rect -6600 257 -5078 308
rect -6601 224 -5078 257
rect -31679 -62597 -30522 -8679
rect -29580 -46472 -28157 -10506
rect -6601 -11153 -6294 224
rect 2391 506 2427 892
rect 2494 777 2540 861
rect 2803 777 2849 892
rect 3061 589 3235 1101
rect 2794 506 3235 589
rect 2391 470 3235 506
rect 2794 439 3235 470
rect 2794 355 3099 439
rect -5058 -535 -5012 -335
rect -4862 -535 -4816 -335
rect -4666 -535 -4620 -335
rect -4208 -535 -4162 -335
rect -4012 -535 -3966 -335
rect -3816 -535 -3770 -335
rect -1581 -342 -1323 -85
rect -4208 -1610 -4162 -1410
rect -4012 -1610 -3966 -1410
rect -3816 -1610 -3770 -1410
rect -1517 -2369 -1361 -342
rect 3281 -911 3574 -645
rect -1585 -2584 -1283 -2369
rect 3313 -2539 3558 -911
rect 3841 -1011 3899 1101
rect 4064 265 4108 1310
rect 6005 1284 6051 1454
rect 4388 1066 4549 1243
rect 6201 1284 6247 1484
rect 6397 1284 6443 1484
rect 6593 1284 6639 1484
rect 6789 1284 6835 1484
rect 3985 76 4186 265
rect 4408 -15 4507 1066
rect 5359 938 5405 1138
rect 5555 938 5601 1138
rect 5751 938 5797 1138
rect 6005 938 6051 1138
rect 6201 938 6247 1138
rect 6397 938 6443 1138
rect 6593 938 6639 1138
rect 6789 938 6835 1138
rect 5730 686 6208 775
rect 5943 223 6135 686
rect 4383 -213 4585 -15
rect 5891 -122 6236 223
rect 4524 -677 4570 -477
rect 4720 -677 4766 -477
rect 4916 -677 4962 -477
rect 5374 -677 5420 -477
rect 5570 -677 5616 -477
rect 5766 -677 5812 -477
rect 4524 -957 4570 -857
rect 4720 -957 4766 -857
rect 4916 -957 4962 -857
rect 5374 -957 5420 -857
rect 5570 -957 5616 -857
rect 5766 -957 5812 -857
rect 3841 -1066 4999 -1011
rect 7904 1049 7950 1449
rect 11326 1596 11372 1712
rect 15522 1597 15742 1833
rect 8140 1049 8186 1449
rect 8376 1049 8422 1449
rect 8612 1049 8658 1449
rect 8848 1049 8894 1449
rect 9084 1049 9130 1449
rect 9320 1049 9366 1449
rect 9674 1550 11372 1596
rect 9556 1049 9602 1449
rect 9674 1049 9720 1550
rect 9792 1049 9838 1449
rect 9910 1049 9956 1550
rect 10028 1049 10074 1449
rect 10146 1049 10192 1550
rect 10264 1049 10310 1449
rect 10382 1049 10428 1550
rect 10500 1049 10546 1449
rect 10618 1049 10664 1550
rect 10736 1049 10782 1449
rect 10854 1049 10900 1550
rect 10972 1049 11018 1449
rect 11090 1049 11136 1550
rect 11208 1049 11254 1449
rect 11326 1049 11372 1550
rect 11444 1049 11490 1449
rect 11562 1049 11608 1449
rect 11680 1049 11726 1449
rect 11798 1049 11844 1449
rect 11916 1049 11962 1449
rect 12034 1049 12080 1449
rect 12152 1049 12198 1449
rect 12270 1049 12316 1449
rect 12388 1049 12434 1449
rect 12506 1049 12552 1449
rect 12624 1049 12670 1449
rect 12742 1049 12788 1449
rect 12860 1049 12906 1449
rect 12978 1049 13024 1449
rect 13096 1049 13142 1449
rect 13214 1049 13260 1449
rect 13332 1049 13378 1449
rect 13450 1049 13496 1449
rect 13568 1049 13614 1449
rect 13686 1049 13732 1449
rect 13804 1049 13850 1449
rect 13922 1049 13968 1449
rect 14040 1049 14086 1449
rect 14158 1049 14204 1449
rect 14276 1049 14322 1449
rect 14394 1049 14440 1449
rect 14512 1049 14558 1449
rect 14630 1049 14676 1449
rect 14748 1049 14794 1449
rect 14866 1049 14912 1449
rect 14984 1049 15030 1449
rect 7571 -899 7617 -499
rect 7807 -899 7853 -499
rect 8043 -899 8089 -499
rect 8173 -899 8219 -499
rect 8409 -899 8455 -499
rect 8645 -899 8691 -499
rect 8881 -899 8927 -499
rect 9117 -899 9163 -499
rect 9247 -899 9293 -499
rect 9483 -899 9529 -499
rect 9719 -899 9765 -499
rect 9955 -899 10001 -499
rect 10191 -899 10237 -499
rect 10427 -899 10473 -499
rect 10663 -899 10709 -499
rect 10899 -899 10945 -499
rect 11135 -899 11181 -499
rect 11265 -970 11311 -499
rect 11383 -899 11429 -499
rect 11501 -970 11547 -499
rect 11619 -899 11665 -499
rect 11737 -970 11783 -499
rect 11855 -899 11901 -499
rect 11973 -970 12019 -499
rect 12091 -899 12137 -499
rect 12209 -970 12255 -499
rect 12327 -899 12373 -499
rect 12445 -970 12491 -499
rect 12563 -899 12609 -499
rect 12681 -970 12727 -499
rect 12799 -899 12845 -499
rect 12917 -970 12963 -499
rect 13035 -899 13081 -499
rect 13153 -970 13199 -499
rect 13271 -899 13317 -499
rect 13389 -970 13435 -499
rect 13507 -899 13553 -499
rect 13625 -970 13671 -499
rect 13743 -899 13789 -499
rect 13861 -970 13907 -499
rect 13979 -899 14025 -499
rect 14097 -970 14143 -499
rect 14215 -899 14261 -499
rect 14333 -970 14379 -499
rect 14451 -899 14497 -499
rect 14569 -970 14615 -499
rect 14687 -899 14733 -499
rect 14805 -970 14851 -499
rect 14923 -899 14969 -499
rect 15041 -970 15087 -499
rect 3841 -1069 4601 -1066
rect 11239 -1044 15116 -970
rect 5265 -1236 6067 -1192
rect 5265 -1336 5309 -1236
rect 4333 -1380 5309 -1336
rect 5374 -1372 5420 -1272
rect 5570 -1372 5616 -1272
rect 5766 -1372 5812 -1272
rect 4353 -2171 4397 -1380
rect 6020 -1406 6066 -1236
rect 6216 -1406 6262 -1206
rect 6412 -1406 6458 -1206
rect 6608 -1406 6654 -1206
rect 6804 -1406 6850 -1206
rect 5374 -1752 5420 -1552
rect 5570 -1752 5616 -1552
rect 5766 -1752 5812 -1552
rect 6020 -1752 6066 -1552
rect 6216 -1752 6262 -1552
rect 6412 -1752 6458 -1552
rect 6608 -1752 6654 -1552
rect 6804 -1752 6850 -1552
rect 7863 -1707 7909 -1307
rect 11285 -1160 11331 -1044
rect 8099 -1707 8145 -1307
rect 8335 -1707 8381 -1307
rect 8571 -1707 8617 -1307
rect 8807 -1707 8853 -1307
rect 9043 -1707 9089 -1307
rect 9279 -1707 9325 -1307
rect 9633 -1206 11331 -1160
rect 9515 -1707 9561 -1307
rect 9633 -1707 9679 -1206
rect 9751 -1707 9797 -1307
rect 9869 -1707 9915 -1206
rect 9987 -1707 10033 -1307
rect 10105 -1707 10151 -1206
rect 10223 -1707 10269 -1307
rect 10341 -1707 10387 -1206
rect 10459 -1707 10505 -1307
rect 10577 -1707 10623 -1206
rect 10695 -1707 10741 -1307
rect 10813 -1707 10859 -1206
rect 10931 -1707 10977 -1307
rect 11049 -1707 11095 -1206
rect 11167 -1707 11213 -1307
rect 11285 -1707 11331 -1206
rect 11403 -1707 11449 -1307
rect 11521 -1707 11567 -1307
rect 11639 -1707 11685 -1307
rect 11757 -1707 11803 -1307
rect 11875 -1707 11921 -1307
rect 11993 -1707 12039 -1307
rect 12111 -1707 12157 -1307
rect 12229 -1707 12275 -1307
rect 12347 -1707 12393 -1307
rect 12465 -1707 12511 -1307
rect 12583 -1707 12629 -1307
rect 12701 -1707 12747 -1307
rect 12819 -1707 12865 -1307
rect 12937 -1707 12983 -1307
rect 13055 -1707 13101 -1307
rect 13173 -1707 13219 -1307
rect 13291 -1707 13337 -1307
rect 13409 -1707 13455 -1307
rect 13527 -1707 13573 -1307
rect 13645 -1707 13691 -1307
rect 13763 -1707 13809 -1307
rect 13881 -1707 13927 -1307
rect 13999 -1707 14045 -1307
rect 14117 -1707 14163 -1307
rect 14235 -1707 14281 -1307
rect 14353 -1707 14399 -1307
rect 14471 -1707 14517 -1307
rect 14589 -1707 14635 -1307
rect 14707 -1707 14753 -1307
rect 14825 -1707 14871 -1307
rect 14943 -1707 14989 -1307
rect 4310 -2309 4465 -2171
rect 3196 -2900 3624 -2539
rect 15547 -2842 15703 1597
rect 15814 -255 16329 3722
rect 16519 909 17132 8006
rect 26753 7623 38073 8844
rect 18137 3181 18324 3184
rect 18137 2985 18330 3181
rect 16519 296 17906 909
rect 16101 -1228 16445 -871
rect 15440 -3211 15853 -2842
rect 16133 -3292 16375 -1228
rect 16088 -3623 16483 -3292
rect 17293 -4848 17906 296
rect 18137 -4849 18324 2985
rect 17978 -5437 18468 -4849
rect 18621 -5532 18758 2557
rect 19788 3178 19834 3378
rect 19984 3178 20030 3378
rect 20180 3178 20226 3378
rect 20638 3178 20684 3378
rect 20834 3178 20880 3378
rect 21030 3178 21076 3378
rect 19788 2898 19834 2998
rect 19984 2898 20030 2998
rect 20180 2898 20226 2998
rect 19552 2862 19650 2892
rect 20638 2898 20684 2998
rect 20834 2898 20880 2998
rect 21030 2898 21076 2998
rect 19552 2858 19659 2862
rect 19552 2787 20314 2858
rect 20529 2619 21331 2663
rect 19341 2519 19481 2579
rect 20529 2519 20573 2619
rect 19341 2475 20573 2519
rect 20638 2483 20684 2583
rect 20834 2483 20880 2583
rect 21030 2483 21076 2583
rect 19341 2444 19481 2475
rect 21284 2449 21330 2619
rect 21480 2449 21526 2649
rect 21676 2449 21722 2649
rect 21872 2449 21918 2649
rect 22068 2449 22114 2649
rect 20638 2103 20684 2303
rect 20834 2103 20880 2303
rect 21030 2103 21076 2303
rect 21284 2103 21330 2303
rect 21480 2103 21526 2303
rect 21676 2103 21722 2303
rect 21872 2103 21918 2303
rect 22068 2103 22114 2303
rect 22436 1241 22925 1317
rect 19472 943 22925 1241
rect 19472 -496 19542 943
rect 22436 895 22925 943
rect 19960 -172 20006 28
rect 20156 -172 20202 28
rect 20352 -172 20398 28
rect 20810 -172 20856 28
rect 21006 -172 21052 28
rect 21202 -172 21248 28
rect 19960 -452 20006 -352
rect 20156 -452 20202 -352
rect 20352 -452 20398 -352
rect 20810 -452 20856 -352
rect 21006 -452 21052 -352
rect 21202 -452 21248 -352
rect 19472 -566 20517 -496
rect 26836 3886 28029 7623
rect 29111 3886 30304 7623
rect 31275 3886 32468 7623
rect 33884 3886 35077 7623
rect 36381 3886 37574 7623
rect 41672 4185 44640 4844
rect 26583 3483 38866 3886
rect 41865 3233 42195 4185
rect 42554 3233 42884 4185
rect 43243 3233 43573 4185
rect 43752 3233 44082 4185
rect 41827 3129 44196 3233
rect 26688 2653 26963 2876
rect 26762 646 26890 2653
rect 27715 1791 27761 1991
rect 27873 1791 27919 1991
rect 27715 1468 27761 1668
rect 27873 1468 27919 1668
rect 28261 1468 28307 2057
rect 28577 1468 28623 2057
rect 30324 2096 30370 2496
rect 30640 2096 30686 2496
rect 30956 2096 31002 2496
rect 31114 2096 31160 2496
rect 31272 2096 31318 2496
rect 31430 2096 31476 2496
rect 31588 2096 31634 2496
rect 35059 2118 35105 2518
rect 35375 2118 35421 2518
rect 35691 2118 35737 2518
rect 35849 2118 35895 2518
rect 36007 2118 36053 2518
rect 36165 2118 36211 2518
rect 36323 2118 36369 2518
rect 29023 1468 29069 2062
rect 29307 1800 29353 2062
rect 29465 1800 29511 2062
rect 29286 1763 29546 1800
rect 29286 1754 30129 1763
rect 29311 1467 29357 1754
rect 29469 1717 30129 1754
rect 29469 1467 29515 1717
rect 30083 1411 30129 1717
rect 30324 1411 30370 1840
rect 30640 1440 30686 1840
rect 30956 1440 31002 1840
rect 31272 1440 31318 1840
rect 30083 1365 30370 1411
rect 31588 1417 31634 1840
rect 32570 1784 32616 1984
rect 32728 1784 32774 1984
rect 32570 1417 32616 1661
rect 32728 1461 32774 1661
rect 31588 1371 32616 1417
rect 33116 1461 33162 2050
rect 33432 1461 33478 2050
rect 36780 2075 36826 2475
rect 37096 2075 37142 2475
rect 37412 2075 37458 2475
rect 37570 2075 37616 2475
rect 37728 2075 37774 2475
rect 37886 2075 37932 2475
rect 38044 2075 38090 2475
rect 33878 1461 33924 2055
rect 34162 1793 34208 2055
rect 34320 1793 34366 2055
rect 39180 2735 39226 2935
rect 39376 2735 39422 2935
rect 39572 2735 39618 2935
rect 40062 2735 40108 2935
rect 40258 2735 40304 2935
rect 40454 2735 40500 2935
rect 41805 2735 41851 2935
rect 42001 2735 42047 2935
rect 42197 2735 42243 2935
rect 39180 2455 39226 2555
rect 39376 2455 39422 2555
rect 39572 2455 39618 2555
rect 42762 2735 42808 2935
rect 42958 2735 43004 2935
rect 43154 2735 43200 2935
rect 44505 2735 44551 2935
rect 44701 2735 44747 2935
rect 44897 2735 44943 2935
rect 38805 2407 38941 2408
rect 38780 2288 38972 2407
rect 39453 2335 39590 2395
rect 39460 2288 39555 2335
rect 40062 2455 40108 2555
rect 40258 2455 40304 2555
rect 40454 2455 40500 2555
rect 41805 2455 41851 2555
rect 42001 2455 42047 2555
rect 42197 2455 42243 2555
rect 42080 2334 42217 2394
rect 38780 2193 39555 2288
rect 38780 2149 38972 2193
rect 39460 2126 39555 2193
rect 39440 2066 39572 2126
rect 34550 1793 34596 1841
rect 34141 1747 34596 1793
rect 34166 1460 34212 1747
rect 34324 1460 34370 1747
rect 26762 518 27180 646
rect 20701 -731 21503 -687
rect 19212 -831 19359 -829
rect 20701 -831 20745 -731
rect 19212 -875 20745 -831
rect 20810 -867 20856 -767
rect 21006 -867 21052 -767
rect 21202 -867 21248 -767
rect 18424 -6171 19081 -5532
rect 19212 -6293 19542 -875
rect 21456 -901 21502 -731
rect 21652 -901 21698 -701
rect 21848 -901 21894 -701
rect 22044 -901 22090 -701
rect 22240 -901 22286 -701
rect 27052 -38 27180 518
rect 27810 398 27856 1141
rect 27968 489 28014 1141
rect 27689 352 27856 398
rect 29116 937 29162 1137
rect 29274 937 29320 1137
rect 29115 489 29161 689
rect 27531 -23 27577 177
rect 27689 -23 27735 352
rect 29273 369 29319 689
rect 30324 440 30370 840
rect 30640 440 30686 840
rect 30956 440 31002 840
rect 31272 440 31318 840
rect 31588 440 31634 840
rect 32665 391 32711 1134
rect 32823 482 32869 1134
rect 29273 323 29546 369
rect 27961 -21 28007 179
rect 28277 -21 28323 179
rect 28593 -21 28639 179
rect 28909 -21 28955 179
rect 29225 -21 29271 179
rect 29500 -21 29546 323
rect 32544 345 32711 391
rect 33971 930 34017 1130
rect 34129 930 34175 1130
rect 34550 970 34596 1747
rect 35059 1462 35105 1862
rect 35375 1462 35421 1862
rect 35691 1462 35737 1862
rect 36007 1462 36053 1862
rect 36323 1462 36369 1862
rect 36780 1419 36826 1819
rect 37096 1419 37142 1819
rect 37412 1419 37458 1819
rect 37728 1419 37774 1819
rect 38044 1419 38090 1819
rect 41066 1797 41112 1897
rect 41262 1797 41308 1897
rect 41458 1797 41504 1897
rect 42104 2126 42199 2334
rect 42073 2066 42210 2126
rect 41903 1797 41949 1897
rect 42099 1797 42145 1897
rect 42295 1797 42341 1897
rect 50890 2634 50936 3034
rect 51126 2634 51172 3034
rect 51362 2634 51408 3034
rect 51492 2634 51538 3034
rect 51728 2634 51774 3034
rect 51964 2634 52010 3034
rect 52200 2634 52246 3034
rect 52436 2634 52482 3034
rect 52566 2634 52612 3034
rect 52802 2634 52848 3034
rect 53038 2634 53084 3034
rect 53274 2634 53320 3034
rect 53510 2634 53556 3034
rect 53746 2634 53792 3034
rect 53982 2634 54028 3034
rect 54218 2634 54264 3034
rect 54454 2634 54500 3034
rect 54584 2563 54630 3034
rect 54702 2634 54748 3034
rect 54820 2563 54866 3034
rect 54938 2634 54984 3034
rect 55056 2563 55102 3034
rect 55174 2634 55220 3034
rect 55292 2563 55338 3034
rect 55410 2634 55456 3034
rect 55528 2563 55574 3034
rect 55646 2634 55692 3034
rect 55764 2563 55810 3034
rect 55882 2634 55928 3034
rect 56000 2563 56046 3034
rect 56118 2634 56164 3034
rect 56236 2563 56282 3034
rect 56354 2634 56400 3034
rect 56472 2563 56518 3034
rect 56590 2634 56636 3034
rect 56708 2563 56754 3034
rect 56826 2634 56872 3034
rect 56944 2563 56990 3034
rect 57062 2634 57108 3034
rect 57180 2563 57226 3034
rect 57298 2634 57344 3034
rect 57416 2563 57462 3034
rect 57534 2634 57580 3034
rect 57652 2563 57698 3034
rect 57770 2634 57816 3034
rect 57888 2563 57934 3034
rect 58006 2634 58052 3034
rect 58124 2563 58170 3034
rect 58242 2634 58288 3034
rect 58360 2563 58406 3034
rect 42762 2455 42808 2555
rect 42958 2455 43004 2555
rect 43154 2455 43200 2555
rect 44505 2455 44551 2555
rect 44701 2455 44747 2555
rect 44897 2455 44943 2555
rect 54558 2489 58435 2563
rect 44684 2379 44816 2398
rect 45804 2379 45950 2441
rect 44684 2338 45950 2379
rect 44697 2335 45950 2338
rect 43766 1797 43812 1897
rect 43962 1797 44008 1897
rect 44158 1797 44204 1897
rect 44697 2120 44792 2335
rect 45804 2255 45950 2335
rect 44670 2060 44807 2120
rect 44603 1797 44649 1897
rect 44799 1797 44845 1897
rect 44995 1797 45041 1897
rect 45573 1887 45619 1987
rect 45769 1887 45815 1987
rect 45965 1887 46011 1987
rect 41066 1417 41112 1617
rect 41262 1417 41308 1617
rect 41458 1417 41504 1617
rect 41903 1417 41949 1617
rect 42099 1417 42145 1617
rect 42295 1417 42341 1617
rect 43766 1417 43812 1617
rect 43962 1417 44008 1617
rect 44158 1417 44204 1617
rect 44603 1417 44649 1617
rect 44799 1417 44845 1617
rect 44995 1417 45041 1617
rect 51182 1826 51228 2226
rect 54604 2373 54650 2489
rect 51418 1826 51464 2226
rect 51654 1826 51700 2226
rect 51890 1826 51936 2226
rect 52126 1826 52172 2226
rect 52362 1826 52408 2226
rect 52598 1826 52644 2226
rect 52952 2327 54650 2373
rect 52834 1826 52880 2226
rect 52952 1826 52998 2327
rect 53070 1826 53116 2226
rect 53188 1826 53234 2327
rect 53306 1826 53352 2226
rect 53424 1826 53470 2327
rect 53542 1826 53588 2226
rect 53660 1826 53706 2327
rect 53778 1826 53824 2226
rect 53896 1826 53942 2327
rect 54014 1826 54060 2226
rect 54132 1826 54178 2327
rect 54250 1826 54296 2226
rect 54368 1826 54414 2327
rect 54486 1826 54532 2226
rect 54604 1826 54650 2327
rect 58706 2260 59616 2704
rect 54722 1826 54768 2226
rect 54840 1826 54886 2226
rect 54958 1826 55004 2226
rect 55076 1826 55122 2226
rect 55194 1826 55240 2226
rect 55312 1826 55358 2226
rect 55430 1826 55476 2226
rect 55548 1826 55594 2226
rect 55666 1826 55712 2226
rect 55784 1826 55830 2226
rect 55902 1826 55948 2226
rect 56020 1826 56066 2226
rect 56138 1826 56184 2226
rect 56256 1826 56302 2226
rect 56374 1826 56420 2226
rect 56492 1826 56538 2226
rect 56610 1826 56656 2226
rect 56728 1826 56774 2226
rect 56846 1826 56892 2226
rect 56964 1826 57010 2226
rect 57082 1826 57128 2226
rect 57200 1826 57246 2226
rect 57318 1826 57364 2226
rect 57436 1826 57482 2226
rect 57554 1826 57600 2226
rect 57672 1826 57718 2226
rect 57790 1826 57836 2226
rect 57908 1826 57954 2226
rect 58026 1826 58072 2226
rect 58144 1826 58190 2226
rect 58262 1826 58308 2226
rect 45573 1507 45619 1707
rect 45769 1507 45815 1707
rect 45965 1507 46011 1707
rect 34550 924 35105 970
rect 33970 482 34016 682
rect 29658 -21 29704 179
rect 26988 -69 27304 -38
rect 26988 -149 27767 -69
rect 26988 -166 27304 -149
rect 27390 -306 27470 -149
rect 30324 -216 30370 184
rect 30640 -216 30686 184
rect 30956 -216 31002 184
rect 31114 -216 31160 184
rect 31272 -216 31318 184
rect 31430 -216 31476 184
rect 31588 -216 31634 184
rect 32386 -30 32432 170
rect 32544 -30 32590 345
rect 34128 362 34174 682
rect 35059 463 35105 924
rect 35375 463 35421 863
rect 35691 463 35737 863
rect 36007 463 36053 863
rect 36323 463 36369 863
rect 36780 506 36826 906
rect 37096 506 37142 906
rect 37412 506 37458 906
rect 37728 506 37774 906
rect 38044 506 38090 906
rect 34128 316 34401 362
rect 32816 -28 32862 172
rect 33132 -28 33178 172
rect 33448 -28 33494 172
rect 33764 -28 33810 172
rect 34080 -28 34126 172
rect 34355 -28 34401 316
rect 34513 -28 34559 172
rect 31866 -152 32623 -72
rect 31866 -306 31946 -152
rect 35059 -193 35105 207
rect 35375 -193 35421 207
rect 35691 -193 35737 207
rect 35849 -193 35895 207
rect 36007 -193 36053 207
rect 36165 -193 36211 207
rect 36323 -193 36369 207
rect 36780 -150 36826 250
rect 37096 -150 37142 250
rect 37412 -150 37458 250
rect 37570 -150 37616 250
rect 37728 -150 37774 250
rect 37886 -150 37932 250
rect 38044 -150 38090 250
rect 27390 -386 31946 -306
rect 19836 -1279 20093 -990
rect 20810 -1247 20856 -1047
rect 21006 -1247 21052 -1047
rect 21202 -1247 21248 -1047
rect 21456 -1247 21502 -1047
rect 21652 -1247 21698 -1047
rect 21848 -1247 21894 -1047
rect 22044 -1247 22090 -1047
rect 22240 -1247 22286 -1047
rect 18949 -6850 19611 -6293
rect 19868 -7025 20066 -1279
rect 46850 -4670 47412 -1960
rect 50687 -277 50733 123
rect 50923 -277 50969 123
rect 51159 -277 51205 123
rect 51289 -277 51335 123
rect 51525 -277 51571 123
rect 51761 -277 51807 123
rect 51997 -277 52043 123
rect 52233 -277 52279 123
rect 52363 -277 52409 123
rect 52599 -277 52645 123
rect 52835 -277 52881 123
rect 53071 -277 53117 123
rect 53307 -277 53353 123
rect 53543 -277 53589 123
rect 53779 -277 53825 123
rect 54015 -277 54061 123
rect 54251 -277 54297 123
rect 54381 -348 54427 123
rect 54499 -277 54545 123
rect 54617 -348 54663 123
rect 54735 -277 54781 123
rect 54853 -348 54899 123
rect 54971 -277 55017 123
rect 55089 -348 55135 123
rect 55207 -277 55253 123
rect 55325 -348 55371 123
rect 55443 -277 55489 123
rect 55561 -348 55607 123
rect 55679 -277 55725 123
rect 55797 -348 55843 123
rect 55915 -277 55961 123
rect 56033 -348 56079 123
rect 56151 -277 56197 123
rect 56269 -348 56315 123
rect 56387 -277 56433 123
rect 56505 -348 56551 123
rect 56623 -277 56669 123
rect 56741 -348 56787 123
rect 56859 -277 56905 123
rect 56977 -348 57023 123
rect 57095 -277 57141 123
rect 57213 -348 57259 123
rect 57331 -277 57377 123
rect 57449 -348 57495 123
rect 57567 -277 57613 123
rect 57685 -348 57731 123
rect 57803 -277 57849 123
rect 57921 -348 57967 123
rect 58039 -277 58085 123
rect 58157 -348 58203 123
rect 54355 -422 58232 -348
rect 50979 -1085 51025 -685
rect 54401 -538 54447 -422
rect 51215 -1085 51261 -685
rect 51451 -1085 51497 -685
rect 51687 -1085 51733 -685
rect 51923 -1085 51969 -685
rect 52159 -1085 52205 -685
rect 52395 -1085 52441 -685
rect 52749 -584 54447 -538
rect 52631 -1085 52677 -685
rect 52749 -1085 52795 -584
rect 52867 -1085 52913 -685
rect 52985 -1085 53031 -584
rect 53103 -1085 53149 -685
rect 53221 -1085 53267 -584
rect 53339 -1085 53385 -685
rect 53457 -1085 53503 -584
rect 53575 -1085 53621 -685
rect 53693 -1085 53739 -584
rect 53811 -1085 53857 -685
rect 53929 -1085 53975 -584
rect 54047 -1085 54093 -685
rect 54165 -1085 54211 -584
rect 54283 -1085 54329 -685
rect 54401 -1085 54447 -584
rect 54519 -1085 54565 -685
rect 54637 -1085 54683 -685
rect 54755 -1085 54801 -685
rect 54873 -1085 54919 -685
rect 54991 -1085 55037 -685
rect 55109 -1085 55155 -685
rect 55227 -1085 55273 -685
rect 55345 -1085 55391 -685
rect 55463 -1085 55509 -685
rect 55581 -1085 55627 -685
rect 55699 -1085 55745 -685
rect 55817 -1085 55863 -685
rect 55935 -1085 55981 -685
rect 56053 -1085 56099 -685
rect 56171 -1085 56217 -685
rect 56289 -1085 56335 -685
rect 56407 -1085 56453 -685
rect 56525 -1085 56571 -685
rect 56643 -1085 56689 -685
rect 56761 -1085 56807 -685
rect 56879 -1085 56925 -685
rect 56997 -1085 57043 -685
rect 57115 -1085 57161 -685
rect 57233 -1085 57279 -685
rect 57351 -1085 57397 -685
rect 57469 -1085 57515 -685
rect 57587 -1085 57633 -685
rect 57705 -1085 57751 -685
rect 57823 -1085 57869 -685
rect 57941 -1085 57987 -685
rect 58059 -1085 58105 -685
rect 50687 -3324 50733 -2924
rect 50923 -3324 50969 -2924
rect 51159 -3324 51205 -2924
rect 51289 -3324 51335 -2924
rect 51525 -3324 51571 -2924
rect 51761 -3324 51807 -2924
rect 51997 -3324 52043 -2924
rect 52233 -3324 52279 -2924
rect 52363 -3324 52409 -2924
rect 52599 -3324 52645 -2924
rect 52835 -3324 52881 -2924
rect 53071 -3324 53117 -2924
rect 53307 -3324 53353 -2924
rect 53543 -3324 53589 -2924
rect 53779 -3324 53825 -2924
rect 54015 -3324 54061 -2924
rect 54251 -3324 54297 -2924
rect 54499 -3324 54545 -2924
rect 54735 -3324 54781 -2924
rect 54971 -3324 55017 -2924
rect 55207 -3324 55253 -2924
rect 55443 -3324 55489 -2924
rect 55679 -3324 55725 -2924
rect 55915 -3324 55961 -2924
rect 56151 -3324 56197 -2924
rect 56387 -3324 56433 -2924
rect 56623 -3324 56669 -2924
rect 56859 -3324 56905 -2924
rect 57095 -3324 57141 -2924
rect 57331 -3324 57377 -2924
rect 57567 -3324 57613 -2924
rect 57803 -3324 57849 -2924
rect 58039 -3324 58085 -2924
rect 50979 -4132 51025 -3732
rect 51215 -4132 51261 -3732
rect 51451 -4132 51497 -3732
rect 51687 -4132 51733 -3732
rect 51923 -4132 51969 -3732
rect 52159 -4132 52205 -3732
rect 52395 -4132 52441 -3732
rect 52631 -4132 52677 -3732
rect 52867 -4132 52913 -3732
rect 53103 -4132 53149 -3732
rect 53339 -4132 53385 -3732
rect 53575 -4132 53621 -3732
rect 53811 -4132 53857 -3732
rect 54047 -4132 54093 -3732
rect 54283 -4132 54329 -3732
rect 54519 -4132 54565 -3732
rect 54637 -4132 54683 -3732
rect 54755 -4132 54801 -3732
rect 54873 -4132 54919 -3732
rect 54991 -4132 55037 -3732
rect 55109 -4132 55155 -3732
rect 55227 -4132 55273 -3732
rect 55345 -4132 55391 -3732
rect 55463 -4132 55509 -3732
rect 55581 -4132 55627 -3732
rect 55699 -4132 55745 -3732
rect 55817 -4132 55863 -3732
rect 55935 -4132 55981 -3732
rect 56053 -4132 56099 -3732
rect 56171 -4132 56217 -3732
rect 56289 -4132 56335 -3732
rect 56407 -4132 56453 -3732
rect 56525 -4132 56571 -3732
rect 56643 -4132 56689 -3732
rect 56761 -4132 56807 -3732
rect 56879 -4132 56925 -3732
rect 56997 -4132 57043 -3732
rect 57115 -4132 57161 -3732
rect 57233 -4132 57279 -3732
rect 57351 -4132 57397 -3732
rect 57469 -4132 57515 -3732
rect 57587 -4132 57633 -3732
rect 57705 -4132 57751 -3732
rect 57823 -4132 57869 -3732
rect 57941 -4132 57987 -3732
rect 58059 -4132 58105 -3732
rect 46778 -5304 47412 -4670
rect 19665 -7634 20295 -7025
rect 59172 -8831 59616 2260
rect 58913 -9909 59860 -8831
rect 60549 -9617 61159 -228
rect 62387 -3038 62433 -2838
rect 62583 -3038 62629 -2838
rect 62779 -3038 62825 -2838
rect 63237 -3038 63283 -2838
rect 63433 -3038 63479 -2838
rect 63629 -3038 63675 -2838
rect 61353 -3293 62176 -3228
rect 61353 -4779 61418 -3293
rect 62111 -3360 62176 -3293
rect 62387 -3318 62433 -3218
rect 62583 -3318 62629 -3218
rect 62779 -3318 62825 -3218
rect 63237 -3318 63283 -3218
rect 63433 -3318 63479 -3218
rect 63629 -3318 63675 -3218
rect 62111 -3425 62910 -3360
rect 62387 -3431 62910 -3425
rect 63128 -3597 63930 -3553
rect 63128 -3697 63172 -3597
rect 61655 -3741 63172 -3697
rect 63237 -3733 63283 -3633
rect 63433 -3733 63479 -3633
rect 63629 -3733 63675 -3633
rect 61261 -5041 61482 -4779
rect 60423 -10731 61454 -9617
rect 61655 -11116 62108 -3741
rect 63883 -3767 63929 -3597
rect 62432 -4139 62779 -3786
rect 64079 -3767 64125 -3567
rect 64275 -3767 64321 -3567
rect 64471 -3767 64517 -3567
rect 64667 -3767 64713 -3567
rect 63237 -4113 63283 -3913
rect 63433 -4113 63479 -3913
rect 63629 -4113 63675 -3913
rect 63883 -4113 63929 -3913
rect 64079 -4113 64125 -3913
rect 64275 -4113 64321 -3913
rect 64471 -4113 64517 -3913
rect 64667 -4113 64713 -3913
rect -6611 -11894 -5937 -11153
rect 61366 -11971 62272 -11116
rect 62465 -12441 62732 -4139
rect 62246 -13180 63072 -12441
rect -11299 -15829 -11253 -15328
rect -11063 -15829 -11017 -15328
rect -10827 -15829 -10781 -15328
rect -10591 -15829 -10545 -15328
rect -10355 -15829 -10309 -15328
rect -10119 -15829 -10073 -15328
rect -9883 -15829 -9837 -15328
rect -9647 -15829 -9601 -15328
rect -11299 -15875 -9601 -15829
rect -11299 -15991 -11253 -15875
rect -15084 -16065 -11207 -15991
rect -15055 -16536 -15009 -16065
rect -14937 -16536 -14891 -16136
rect -14819 -16536 -14773 -16065
rect -14701 -16536 -14655 -16136
rect -14583 -16536 -14537 -16065
rect -14465 -16536 -14419 -16136
rect -14347 -16536 -14301 -16065
rect -14229 -16536 -14183 -16136
rect -14111 -16536 -14065 -16065
rect -13993 -16536 -13947 -16136
rect -13875 -16536 -13829 -16065
rect -13757 -16536 -13711 -16136
rect -13639 -16536 -13593 -16065
rect -13521 -16536 -13475 -16136
rect -13403 -16536 -13357 -16065
rect -13285 -16536 -13239 -16136
rect -13167 -16536 -13121 -16065
rect -13049 -16536 -13003 -16136
rect -12931 -16536 -12885 -16065
rect -12813 -16536 -12767 -16136
rect -12695 -16536 -12649 -16065
rect -12577 -16536 -12531 -16136
rect -12459 -16536 -12413 -16065
rect -12341 -16536 -12295 -16136
rect -12223 -16536 -12177 -16065
rect -12105 -16536 -12059 -16136
rect -11987 -16536 -11941 -16065
rect -11869 -16536 -11823 -16136
rect -11751 -16536 -11705 -16065
rect -11633 -16536 -11587 -16136
rect -11515 -16536 -11469 -16065
rect -11397 -16536 -11351 -16136
rect -11279 -16536 -11233 -16065
rect -11149 -16536 -11103 -16136
rect -10913 -16536 -10867 -16136
rect -10677 -16536 -10631 -16136
rect -10441 -16536 -10395 -16136
rect -10205 -16536 -10159 -16136
rect -9969 -16536 -9923 -16136
rect -9733 -16536 -9687 -16136
rect -9497 -16536 -9451 -16136
rect -9261 -16536 -9215 -16136
rect -9131 -16536 -9085 -16136
rect -8895 -16536 -8849 -16136
rect -8659 -16536 -8613 -16136
rect -8423 -16536 -8377 -16136
rect -8187 -16536 -8141 -16136
rect -8057 -16536 -8011 -16136
rect -7821 -16536 -7775 -16136
rect -7585 -16536 -7539 -16136
rect -23884 -27924 -23823 -19397
rect -23937 -28047 -23814 -27924
rect -23693 -28123 -23632 -19318
rect -23584 -19470 -23523 -19232
rect -22744 -19384 -22698 -19184
rect -22548 -19384 -22502 -19184
rect -22352 -19384 -22306 -19184
rect -22156 -19384 -22110 -19184
rect -21614 -19384 -21568 -19184
rect -21418 -19384 -21372 -19184
rect -15145 -18597 -15099 -18397
rect -14949 -18597 -14903 -18397
rect -14753 -18597 -14707 -18397
rect -14308 -18597 -14262 -18397
rect -14112 -18597 -14066 -18397
rect -13916 -18597 -13870 -18397
rect -12445 -18597 -12399 -18397
rect -12249 -18597 -12203 -18397
rect -12053 -18597 -12007 -18397
rect -11608 -18597 -11562 -18397
rect -11412 -18597 -11366 -18397
rect -11216 -18597 -11170 -18397
rect -23584 -25299 -23524 -19470
rect -20745 -19606 -20699 -19306
rect -20549 -19606 -20503 -19306
rect -21054 -19661 -20917 -19644
rect -21082 -19702 -20917 -19661
rect -23584 -25536 -23523 -25299
rect -23746 -28246 -23623 -28123
rect -23584 -28356 -23524 -25536
rect -23640 -28479 -23517 -28356
rect -23485 -28613 -23424 -20397
rect -23547 -28736 -23423 -28613
rect -23372 -28897 -23311 -20330
rect -23441 -28898 -23311 -28897
rect -23441 -28931 -23310 -28898
rect -23440 -29016 -23310 -28931
rect -23258 -29025 -23194 -21802
rect -23260 -29197 -23194 -29025
rect -23281 -29198 -23194 -29197
rect -23281 -29321 -23158 -29198
rect -23113 -29565 -23053 -21371
rect -22687 -21515 -22641 -21215
rect -22491 -21515 -22445 -21215
rect -22295 -21515 -22249 -21215
rect -22078 -21314 -22032 -21214
rect -21882 -21314 -21836 -21214
rect -21686 -21314 -21640 -21214
rect -21490 -21314 -21444 -21214
rect -21082 -20412 -21046 -19702
rect -20959 -19809 -20822 -19751
rect -21084 -20544 -21031 -20412
rect -20952 -20582 -20912 -19809
rect -20353 -19606 -20307 -19306
rect -20136 -19405 -20090 -19305
rect -19940 -19405 -19894 -19305
rect -19744 -19405 -19698 -19305
rect -19548 -19405 -19502 -19305
rect -21068 -20591 -20912 -20582
rect -21115 -20631 -20912 -20591
rect -21068 -20635 -20936 -20631
rect -20914 -21320 -20868 -21120
rect -20718 -21320 -20672 -21120
rect -20522 -21320 -20476 -21120
rect -20326 -21320 -20280 -21120
rect -19784 -21320 -19738 -21120
rect -19588 -21320 -19542 -21120
rect -19109 -20568 -19063 -20268
rect -18913 -20568 -18867 -20268
rect -18717 -20568 -18671 -20268
rect -18500 -20569 -18454 -20469
rect -18304 -20569 -18258 -20469
rect -18108 -20569 -18062 -20469
rect -17912 -20569 -17866 -20469
rect -17662 -20657 -17616 -20057
rect -17466 -20657 -17420 -20057
rect -17043 -20657 -16997 -20057
rect -19083 -21497 -19037 -21297
rect -18887 -21497 -18841 -21297
rect -18691 -21497 -18645 -21297
rect -18495 -21497 -18449 -21297
rect -18110 -21468 -18064 -21168
rect -17914 -21468 -17868 -21168
rect -17718 -21468 -17672 -21168
rect -17501 -21267 -17455 -21167
rect -17305 -21267 -17259 -21167
rect -17109 -21267 -17063 -21167
rect -16913 -21267 -16867 -21167
rect -8783 -19007 -8737 -18407
rect -8360 -19007 -8314 -18407
rect -8164 -19007 -8118 -18407
rect -6675 -18803 -6629 -18603
rect -6479 -18803 -6433 -18603
rect -6283 -18803 -6237 -18603
rect -6169 -18803 -6123 -18603
rect -5973 -18803 -5927 -18603
rect -5860 -18803 -5814 -18603
rect -5664 -18803 -5618 -18603
rect -4175 -18803 -4129 -18603
rect -3979 -18803 -3933 -18603
rect -3783 -18803 -3737 -18603
rect -3669 -18803 -3623 -18603
rect -3473 -18803 -3427 -18603
rect -3360 -18803 -3314 -18603
rect -3164 -18803 -3118 -18603
rect -1675 -18803 -1629 -18603
rect -1479 -18803 -1433 -18603
rect -1283 -18803 -1237 -18603
rect -1169 -18803 -1123 -18603
rect -973 -18803 -927 -18603
rect -860 -18803 -814 -18603
rect -664 -18803 -618 -18603
rect 825 -18803 871 -18603
rect 1021 -18803 1067 -18603
rect 1217 -18803 1263 -18603
rect 1331 -18803 1377 -18603
rect 1527 -18803 1573 -18603
rect 1640 -18803 1686 -18603
rect 1836 -18803 1882 -18603
rect 3325 -18803 3371 -18603
rect 3521 -18803 3567 -18603
rect 3717 -18803 3763 -18603
rect 3831 -18803 3877 -18603
rect 4027 -18803 4073 -18603
rect 4140 -18803 4186 -18603
rect 4336 -18803 4382 -18603
rect 6325 -18803 6371 -18603
rect 6521 -18803 6567 -18603
rect 6717 -18803 6763 -18603
rect 6831 -18803 6877 -18603
rect 7027 -18803 7073 -18603
rect 7140 -18803 7186 -18603
rect 7336 -18803 7382 -18603
rect -15047 -19915 -15001 -19715
rect -14851 -19915 -14805 -19715
rect -14655 -19915 -14609 -19715
rect -13304 -19915 -13258 -19715
rect -13108 -19915 -13062 -19715
rect -12912 -19915 -12866 -19715
rect -12347 -19915 -12301 -19715
rect -12151 -19915 -12105 -19715
rect -11955 -19915 -11909 -19715
rect -10604 -19915 -10558 -19715
rect -10408 -19915 -10362 -19715
rect -10212 -19915 -10166 -19715
rect -9722 -19915 -9676 -19715
rect -9526 -19915 -9480 -19715
rect -9330 -19915 -9284 -19715
rect -14375 -21103 -14178 -21049
rect -19570 -24029 -19391 -23862
rect -22622 -25009 -22576 -24409
rect -22426 -25009 -22380 -24409
rect -21416 -24738 -21370 -24338
rect -21220 -24738 -21174 -24338
rect -20511 -24739 -20465 -24339
rect -20315 -24739 -20269 -24339
rect -21590 -24900 -21532 -24763
rect -21590 -25809 -21555 -24900
rect -20674 -24901 -20616 -24764
rect -21515 -24938 -21457 -24934
rect -21516 -25071 -21457 -24938
rect -21610 -25946 -21552 -25809
rect -21516 -25888 -21473 -25071
rect -21517 -26025 -21459 -25888
rect -20674 -25967 -20639 -24901
rect -20597 -25073 -20539 -24936
rect -20696 -26104 -20638 -25967
rect -20597 -26044 -20562 -25073
rect -20603 -26181 -20545 -26044
rect -22959 -27427 -22913 -27227
rect -22763 -27427 -22717 -27227
rect -22221 -27427 -22175 -27227
rect -22025 -27427 -21979 -27227
rect -21829 -27427 -21783 -27227
rect -21633 -27427 -21587 -27227
rect -20349 -27591 -20173 -26960
rect -19543 -25793 -19417 -24029
rect -14232 -22134 -14178 -21103
rect -14120 -21544 -14074 -21244
rect -13924 -21544 -13878 -21244
rect -13728 -21544 -13682 -21244
rect -13511 -21545 -13465 -21445
rect -13315 -21545 -13269 -21445
rect -13119 -21545 -13073 -21445
rect -12923 -21545 -12877 -21445
rect -12673 -21633 -12627 -21033
rect -12477 -21633 -12431 -21033
rect -12054 -21633 -12008 -21033
rect -15843 -22310 -14178 -22134
rect -19544 -25965 -19352 -25793
rect -19109 -25568 -19063 -25268
rect -18913 -25568 -18867 -25268
rect -18717 -25568 -18671 -25268
rect -18500 -25569 -18454 -25469
rect -18304 -25569 -18258 -25469
rect -18108 -25569 -18062 -25469
rect -17912 -25569 -17866 -25469
rect -17662 -25657 -17616 -25057
rect -17466 -25657 -17420 -25057
rect -17043 -25657 -16997 -25057
rect -19083 -26497 -19037 -26297
rect -18887 -26497 -18841 -26297
rect -18691 -26497 -18645 -26297
rect -18495 -26497 -18449 -26297
rect -18110 -26468 -18064 -26168
rect -17914 -26468 -17868 -26168
rect -17718 -26468 -17672 -26168
rect -17501 -26267 -17455 -26167
rect -17305 -26267 -17259 -26167
rect -17109 -26267 -17063 -26167
rect -16913 -26267 -16867 -26167
rect -15843 -28049 -15667 -22310
rect -14232 -22507 -14178 -22310
rect -14094 -22473 -14048 -22273
rect -14282 -22657 -14152 -22507
rect -13898 -22473 -13852 -22273
rect -13702 -22473 -13656 -22273
rect -13506 -22473 -13460 -22273
rect -13121 -22444 -13075 -22144
rect -12925 -22444 -12879 -22144
rect -12729 -22444 -12683 -22144
rect -12512 -22243 -12466 -22143
rect -12316 -22243 -12270 -22143
rect -12120 -22243 -12074 -22143
rect -11924 -22243 -11878 -22143
rect -15145 -23524 -15099 -23324
rect -14949 -23524 -14903 -23324
rect -14753 -23524 -14707 -23324
rect -14308 -23524 -14262 -23324
rect -14112 -23524 -14066 -23324
rect -13916 -23524 -13870 -23324
rect -12445 -23524 -12399 -23324
rect -12249 -23524 -12203 -23324
rect -12053 -23524 -12007 -23324
rect -11608 -23524 -11562 -23324
rect -11412 -23524 -11366 -23324
rect -11216 -23524 -11170 -23324
rect -15047 -24842 -15001 -24642
rect -14851 -24842 -14805 -24642
rect -14655 -24842 -14609 -24642
rect -13304 -24842 -13258 -24642
rect -13108 -24842 -13062 -24642
rect -12912 -24842 -12866 -24642
rect -12347 -24842 -12301 -24642
rect -12151 -24842 -12105 -24642
rect -11955 -24842 -11909 -24642
rect -10604 -24842 -10558 -24642
rect -10408 -24842 -10362 -24642
rect -10212 -24842 -10166 -24642
rect -9722 -24842 -9676 -24642
rect -9526 -24842 -9480 -24642
rect -9330 -24842 -9284 -24642
rect -8756 -23941 -8710 -23341
rect -8333 -23941 -8287 -23341
rect -8137 -23941 -8091 -23341
rect -7140 -19864 -7004 -19790
rect -7140 -20246 -7089 -19864
rect -7014 -20132 -6968 -19932
rect -6818 -20132 -6772 -19932
rect -6622 -20132 -6576 -19932
rect -4564 -19070 -4425 -19061
rect -3486 -19068 -3347 -19067
rect -3486 -19070 -2898 -19068
rect -4564 -19096 -2898 -19070
rect -4564 -19098 -3347 -19096
rect -4564 -19115 -4425 -19098
rect -3486 -19121 -3347 -19098
rect -5347 -19361 -5224 -19225
rect -5343 -19992 -5229 -19361
rect -5348 -20128 -5225 -19992
rect -2926 -20100 -2898 -19096
rect -2064 -19070 -1925 -19061
rect -986 -19068 -847 -19067
rect -986 -19070 -414 -19068
rect -2064 -19096 -414 -19070
rect -2064 -19098 -847 -19096
rect -2064 -19115 -1925 -19098
rect -986 -19121 -847 -19098
rect -2780 -19396 -2657 -19260
rect -2776 -19848 -2662 -19396
rect -2781 -19984 -2658 -19848
rect -442 -19961 -414 -19096
rect 436 -19070 575 -19061
rect 1514 -19068 1653 -19067
rect 1514 -19070 2052 -19068
rect 436 -19096 2052 -19070
rect 436 -19098 1653 -19096
rect 436 -19115 575 -19098
rect 1514 -19121 1653 -19098
rect -297 -19396 -174 -19260
rect -293 -19813 -179 -19396
rect -298 -19814 -175 -19813
rect -298 -19876 8 -19814
rect 2024 -19841 2052 -19096
rect 2936 -19070 3075 -19061
rect 4014 -19068 4153 -19067
rect 4014 -19070 5373 -19068
rect 2936 -19096 5373 -19070
rect 2936 -19098 4153 -19096
rect 2936 -19115 3075 -19098
rect 4014 -19121 4153 -19098
rect 5345 -19694 5373 -19096
rect 5936 -19070 6075 -19061
rect 7014 -19068 7153 -19067
rect 6912 -19070 9523 -19068
rect 5936 -19096 9523 -19070
rect 5936 -19098 7153 -19096
rect 5936 -19115 6075 -19098
rect 7014 -19121 7153 -19098
rect 5345 -19722 9372 -19694
rect 2024 -19869 9213 -19841
rect -442 -19989 9051 -19961
rect -2926 -20136 8892 -20100
rect -7140 -20297 8725 -20246
rect 3367 -20655 3490 -20646
rect 3768 -20655 3891 -20644
rect -1522 -20670 -1399 -20658
rect -1228 -20670 -1105 -20657
rect -1522 -20785 -1105 -20670
rect -1522 -20794 -1399 -20785
rect -1228 -20793 -1105 -20785
rect 1750 -20685 1873 -20670
rect 2139 -20685 2262 -20669
rect 1750 -20792 2262 -20685
rect 3367 -20762 3891 -20655
rect 3367 -20782 3490 -20762
rect 3768 -20780 3891 -20762
rect 5124 -20662 5247 -20649
rect 6340 -20662 6463 -20650
rect 5124 -20767 6463 -20662
rect 5124 -20785 5247 -20767
rect 6340 -20786 6463 -20767
rect 1750 -20806 1873 -20792
rect 2139 -20805 2262 -20792
rect -7173 -21035 -7127 -20835
rect -6977 -21035 -6931 -20835
rect -6781 -21035 -6735 -20835
rect -5430 -21035 -5384 -20835
rect -5234 -21035 -5188 -20835
rect -5038 -21035 -4992 -20835
rect -4473 -21035 -4427 -20835
rect -4277 -21035 -4231 -20835
rect -4081 -21035 -4035 -20835
rect -2730 -21035 -2684 -20835
rect -2534 -21035 -2488 -20835
rect -2338 -21035 -2292 -20835
rect -1848 -21035 -1802 -20835
rect -1652 -21035 -1606 -20835
rect -1456 -21035 -1410 -20835
rect -1114 -21052 -1068 -20852
rect -918 -21052 -872 -20852
rect -376 -21052 -330 -20852
rect -180 -21052 -134 -20852
rect 16 -21052 62 -20852
rect 212 -21052 258 -20852
rect 619 -20965 665 -20865
rect 815 -20965 861 -20865
rect 1011 -20965 1057 -20865
rect 1207 -20965 1253 -20865
rect -7271 -22353 -7225 -22153
rect -7075 -22353 -7029 -22153
rect -6879 -22353 -6833 -22153
rect 1424 -21166 1470 -20866
rect 1620 -21166 1666 -20866
rect 1816 -21166 1862 -20866
rect 2224 -20967 2270 -20867
rect 2420 -20967 2466 -20867
rect 2616 -20967 2662 -20867
rect 2812 -20967 2858 -20867
rect 3029 -21168 3075 -20868
rect 3225 -21168 3271 -20868
rect 3421 -21168 3467 -20868
rect 3848 -21043 3894 -20843
rect 4044 -21043 4090 -20843
rect 4586 -21043 4632 -20843
rect 4782 -21043 4828 -20843
rect 4978 -21043 5024 -20843
rect 5174 -21043 5220 -20843
rect 6335 -21054 6381 -20854
rect 6531 -21054 6577 -20854
rect 6727 -21054 6773 -20854
rect 6841 -21054 6887 -20854
rect 7037 -21054 7083 -20854
rect 7150 -21054 7196 -20854
rect 7346 -21054 7392 -20854
rect 5946 -21321 6085 -21312
rect 7024 -21319 7163 -21318
rect 8354 -21319 8405 -21311
rect 7024 -21321 8405 -21319
rect 5946 -21347 8405 -21321
rect 5946 -21349 7163 -21347
rect 5946 -21366 6085 -21349
rect 7024 -21372 7163 -21349
rect 8354 -21362 8405 -21347
rect -6434 -22353 -6388 -22153
rect -6238 -22353 -6192 -22153
rect -6042 -22353 -5996 -22153
rect -4571 -22353 -4525 -22153
rect -4375 -22353 -4329 -22153
rect -4179 -22353 -4133 -22153
rect -3734 -22353 -3688 -22153
rect -3538 -22353 -3492 -22153
rect -3342 -22353 -3296 -22153
rect -7271 -23791 -7225 -23591
rect -7075 -23791 -7029 -23591
rect -6879 -23791 -6833 -23591
rect -6434 -23791 -6388 -23591
rect -6238 -23791 -6192 -23591
rect -6042 -23791 -5996 -23591
rect -4571 -23791 -4525 -23591
rect -4375 -23791 -4329 -23591
rect -4179 -23791 -4133 -23591
rect -3734 -23791 -3688 -23591
rect -3538 -23791 -3492 -23591
rect -3342 -23791 -3296 -23591
rect -7173 -25109 -7127 -24909
rect -6977 -25109 -6931 -24909
rect -6781 -25109 -6735 -24909
rect -5430 -25109 -5384 -24909
rect -5234 -25109 -5188 -24909
rect -5038 -25109 -4992 -24909
rect -4473 -25109 -4427 -24909
rect -4277 -25109 -4231 -24909
rect -4081 -25109 -4035 -24909
rect -2730 -25109 -2684 -24909
rect -2534 -25109 -2488 -24909
rect -2338 -25109 -2292 -24909
rect -1848 -25109 -1802 -24909
rect -1652 -25109 -1606 -24909
rect -1456 -25109 -1410 -24909
rect -1114 -25092 -1068 -24892
rect -918 -25092 -872 -24892
rect -376 -25092 -330 -24892
rect -180 -25092 -134 -24892
rect 16 -25092 62 -24892
rect 212 -25092 258 -24892
rect 619 -25079 665 -24979
rect 815 -25079 861 -24979
rect 1011 -25079 1057 -24979
rect 1207 -25079 1253 -24979
rect 1424 -25078 1470 -24778
rect 1620 -25078 1666 -24778
rect 1816 -25078 1862 -24778
rect 2224 -25077 2270 -24977
rect 2420 -25077 2466 -24977
rect 2616 -25077 2662 -24977
rect 2812 -25077 2858 -24977
rect 3029 -25076 3075 -24776
rect 5946 -24595 6085 -24578
rect 7024 -24595 7163 -24572
rect 5946 -24597 7163 -24595
rect 8135 -24597 8280 -24502
rect 8367 -24597 8395 -21362
rect 5946 -24623 8397 -24597
rect 5946 -24632 6085 -24623
rect 7024 -24625 8397 -24623
rect 7024 -24626 7163 -24625
rect 8135 -24637 8280 -24625
rect 3225 -25076 3271 -24776
rect 3421 -25076 3467 -24776
rect 3848 -25101 3894 -24901
rect 4044 -25101 4090 -24901
rect 4586 -25101 4632 -24901
rect 4782 -25101 4828 -24901
rect 4978 -25101 5024 -24901
rect 5174 -25101 5220 -24901
rect 6335 -25090 6381 -24890
rect 6531 -25090 6577 -24890
rect 6727 -25090 6773 -24890
rect 6841 -25090 6887 -24890
rect 7037 -25090 7083 -24890
rect 7150 -25090 7196 -24890
rect 7346 -25090 7392 -24890
rect -1522 -25159 -1399 -25150
rect -1228 -25159 -1105 -25151
rect -1522 -25274 -1105 -25159
rect 1750 -25152 1873 -25138
rect 2139 -25152 2262 -25139
rect 1750 -25259 2262 -25152
rect 1750 -25274 1873 -25259
rect -1522 -25286 -1399 -25274
rect -1228 -25287 -1105 -25274
rect 2139 -25275 2262 -25259
rect 3367 -25182 3490 -25162
rect 3768 -25182 3891 -25164
rect 3367 -25289 3891 -25182
rect 3367 -25298 3490 -25289
rect 3768 -25300 3891 -25289
rect 5124 -25177 5247 -25159
rect 6340 -25177 6463 -25158
rect 5124 -25282 6463 -25177
rect 5124 -25295 5247 -25282
rect 6340 -25294 6463 -25282
rect 8674 -25647 8725 -20297
rect -5483 -25698 8725 -25647
rect -7064 -26846 -6925 -26829
rect -5986 -26846 -5847 -26823
rect -7064 -26848 -5847 -26846
rect -5483 -26848 -5455 -25698
rect -7064 -26874 -5455 -26848
rect -7064 -26883 -6925 -26874
rect -5986 -26876 -5455 -26874
rect -5986 -26877 -5847 -26876
rect 8585 -25808 8733 -25800
rect 8856 -25808 8892 -20136
rect -5348 -25952 -5225 -25816
rect -2926 -25844 8892 -25808
rect -5343 -26583 -5229 -25952
rect -5347 -26719 -5224 -26583
rect -4564 -26846 -4425 -26829
rect -3486 -26846 -3347 -26823
rect -4564 -26848 -3347 -26846
rect -2926 -26848 -2898 -25844
rect 8585 -25848 8733 -25844
rect -4564 -26874 -2898 -26848
rect -4564 -26883 -4425 -26874
rect -3486 -26876 -2898 -26874
rect -3486 -26877 -3347 -26876
rect 8425 -25955 8568 -25937
rect 9023 -25955 9051 -19989
rect -2781 -26096 -2658 -25960
rect -442 -25983 9051 -25955
rect -2776 -26548 -2662 -26096
rect -2780 -26684 -2657 -26548
rect -2064 -26846 -1925 -26829
rect -986 -26846 -847 -26823
rect -2064 -26848 -847 -26846
rect -442 -26848 -414 -25983
rect 8425 -25984 8568 -25983
rect -2064 -26874 -414 -26848
rect -2064 -26883 -1925 -26874
rect -986 -26876 -414 -26874
rect -986 -26877 -847 -26876
rect -298 -26130 8 -26068
rect 8299 -26075 8443 -26068
rect 9185 -26075 9213 -19869
rect 2024 -26103 9213 -26075
rect -298 -26131 -175 -26130
rect -293 -26548 -179 -26131
rect -297 -26684 -174 -26548
rect 436 -26846 575 -26829
rect 1514 -26846 1653 -26823
rect 436 -26848 1653 -26846
rect 2024 -26848 2052 -26103
rect 8299 -26115 8443 -26103
rect 436 -26874 2052 -26848
rect 436 -26883 575 -26874
rect 1514 -26876 2052 -26874
rect 1514 -26877 1653 -26876
rect 7986 -26222 8125 -26207
rect 9344 -26222 9372 -19722
rect 5345 -26250 9372 -26222
rect 2936 -26846 3075 -26829
rect 4014 -26846 4153 -26823
rect 2936 -26848 4153 -26846
rect 5345 -26848 5373 -26250
rect 7986 -26254 8125 -26250
rect 2936 -26874 5373 -26848
rect 2936 -26883 3075 -26874
rect 4014 -26876 5373 -26874
rect 4014 -26877 4153 -26876
rect 5936 -26846 6075 -26829
rect 7014 -26846 7153 -26823
rect 5936 -26848 7153 -26846
rect 7951 -26848 8016 -26744
rect 9495 -26848 9523 -19096
rect 5936 -26874 9523 -26848
rect 5936 -26883 6075 -26874
rect 6912 -26876 9523 -26874
rect 7014 -26877 7153 -26876
rect 7951 -26881 8016 -26876
rect -6675 -27341 -6629 -27141
rect -6479 -27341 -6433 -27141
rect -6283 -27341 -6237 -27141
rect -6169 -27341 -6123 -27141
rect -5973 -27341 -5927 -27141
rect -5860 -27341 -5814 -27141
rect -5664 -27341 -5618 -27141
rect -4175 -27341 -4129 -27141
rect -3979 -27341 -3933 -27141
rect -3783 -27341 -3737 -27141
rect -3669 -27341 -3623 -27141
rect -3473 -27341 -3427 -27141
rect -3360 -27341 -3314 -27141
rect -3164 -27341 -3118 -27141
rect -1675 -27341 -1629 -27141
rect -1479 -27341 -1433 -27141
rect -1283 -27341 -1237 -27141
rect -1169 -27341 -1123 -27141
rect -973 -27341 -927 -27141
rect -860 -27341 -814 -27141
rect -664 -27341 -618 -27141
rect 825 -27341 871 -27141
rect 1021 -27341 1067 -27141
rect 1217 -27341 1263 -27141
rect 1331 -27341 1377 -27141
rect 1527 -27341 1573 -27141
rect 1640 -27341 1686 -27141
rect 1836 -27341 1882 -27141
rect 3325 -27341 3371 -27141
rect 3521 -27341 3567 -27141
rect 3717 -27341 3763 -27141
rect 3831 -27341 3877 -27141
rect 4027 -27341 4073 -27141
rect 4140 -27341 4186 -27141
rect 4336 -27341 4382 -27141
rect 6325 -27341 6371 -27141
rect 6521 -27341 6567 -27141
rect 6717 -27341 6763 -27141
rect 6831 -27341 6877 -27141
rect 7027 -27341 7073 -27141
rect 7140 -27341 7186 -27141
rect 7336 -27341 7382 -27141
rect -23130 -29688 -23007 -29565
rect 7946 -28118 8007 -27514
rect 8064 -27518 8108 -27515
rect 7893 -28241 8016 -28118
rect 8055 -28351 8115 -27518
rect 7999 -28474 8122 -28351
rect 8154 -28608 8215 -27661
rect 8092 -28731 8216 -28608
rect 8267 -28892 8328 -27515
rect 8198 -28893 8328 -28892
rect 8198 -28926 8329 -28893
rect 8199 -29011 8329 -28926
rect 8381 -29020 8445 -27511
rect 8379 -29192 8445 -29020
rect 8358 -29193 8445 -29192
rect 8358 -29316 8481 -29193
rect 8526 -29560 8586 -27475
rect 8509 -29683 8632 -29560
rect 20580 -21304 20626 -21104
rect 20776 -21304 20822 -21104
rect 20972 -21304 21018 -21104
rect 21417 -21304 21463 -21104
rect 21613 -21304 21659 -21104
rect 21809 -21304 21855 -21104
rect 23280 -21304 23326 -21104
rect 23476 -21304 23522 -21104
rect 23672 -21304 23718 -21104
rect 24117 -21304 24163 -21104
rect 24313 -21304 24359 -21104
rect 24509 -21304 24555 -21104
rect 17373 -22502 17419 -21902
rect 17569 -22502 17615 -21902
rect 18694 -22622 18740 -22422
rect 18890 -22622 18936 -22422
rect 19086 -22622 19132 -22422
rect 19576 -22622 19622 -22422
rect 19772 -22622 19818 -22422
rect 19968 -22622 20014 -22422
rect 21319 -22622 21365 -22422
rect 21515 -22622 21561 -22422
rect 21711 -22622 21757 -22422
rect 22276 -22622 22322 -22422
rect 22472 -22622 22518 -22422
rect 22668 -22622 22714 -22422
rect 24019 -22622 24065 -22422
rect 24215 -22622 24261 -22422
rect 24411 -22622 24457 -22422
rect 17368 -24848 17414 -24448
rect 17564 -24848 17610 -24448
rect 18314 -24848 18360 -24448
rect 18510 -24848 18556 -24448
rect 21139 -23574 21185 -23174
rect 21335 -23574 21381 -23174
rect 21531 -23574 21577 -23174
rect 19230 -24882 19276 -24682
rect 19426 -24882 19472 -24682
rect 19622 -24882 19668 -24682
rect 19818 -24882 19864 -24682
rect 20360 -24882 20406 -24682
rect 20556 -24882 20602 -24682
rect 21089 -24875 21135 -24675
rect 21285 -24875 21331 -24675
rect 21481 -24875 21527 -24675
rect 21969 -24804 22015 -24104
rect 22165 -24804 22211 -24104
rect 22369 -24804 22415 -24104
rect 22565 -24804 22611 -24104
rect 22969 -24804 23015 -24104
rect 23165 -24804 23211 -24104
rect 23369 -24804 23415 -24104
rect 23565 -24804 23611 -24104
rect 23969 -24804 24015 -24104
rect 24165 -24804 24211 -24104
rect 24369 -24804 24415 -24104
rect 24565 -24804 24611 -24104
rect 10566 -25860 10612 -25660
rect 10762 -25860 10808 -25660
rect 10958 -25860 11004 -25660
rect 11448 -25860 11494 -25660
rect 11644 -25860 11690 -25660
rect 11840 -25860 11886 -25660
rect 13191 -25860 13237 -25660
rect 13387 -25860 13433 -25660
rect 13583 -25860 13629 -25660
rect 14148 -25860 14194 -25660
rect 14344 -25860 14390 -25660
rect 14540 -25860 14586 -25660
rect 15891 -25860 15937 -25660
rect 16087 -25860 16133 -25660
rect 16283 -25860 16329 -25660
rect 12452 -27178 12498 -26978
rect 12648 -27178 12694 -26978
rect 12844 -27178 12890 -26978
rect 13289 -27178 13335 -26978
rect 13485 -27178 13531 -26978
rect 13681 -27178 13727 -26978
rect 15152 -27178 15198 -26978
rect 15348 -27178 15394 -26978
rect 15544 -27178 15590 -26978
rect 15989 -27178 16035 -26978
rect 16185 -27178 16231 -26978
rect 16381 -27178 16427 -26978
rect 26952 -20951 26998 -20751
rect 27148 -20951 27194 -20751
rect 27344 -20951 27390 -20751
rect 27540 -20951 27586 -20751
rect 27925 -21080 27971 -20780
rect 28121 -21080 28167 -20780
rect 28317 -21080 28363 -20780
rect 28534 -21081 28580 -20981
rect 28730 -21081 28776 -20981
rect 28926 -21081 28972 -20981
rect 29122 -21081 29168 -20981
rect 29204 -21396 29278 -21380
rect 29432 -21396 29542 -21360
rect 29204 -21492 29542 -21396
rect 29204 -21498 29278 -21492
rect 29432 -21510 29542 -21492
rect 26926 -21980 26972 -21680
rect 27122 -21980 27168 -21680
rect 27318 -21980 27364 -21680
rect 27535 -21779 27581 -21679
rect 27731 -21779 27777 -21679
rect 27927 -21779 27973 -21679
rect 28123 -21779 28169 -21679
rect 28373 -22191 28419 -21591
rect 28569 -22191 28615 -21591
rect 28992 -22191 29038 -21591
rect 30365 -21949 30411 -21449
rect 30561 -21949 30607 -21449
rect 31156 -21949 31202 -21449
rect 31286 -21949 31332 -21449
rect 31514 -21749 31560 -21449
rect 31710 -21749 31756 -21449
rect 26944 -24404 26990 -24204
rect 27140 -24404 27186 -24204
rect 27336 -24404 27382 -24204
rect 27532 -24404 27578 -24204
rect 27917 -24533 27963 -24233
rect 28113 -24533 28159 -24233
rect 28309 -24533 28355 -24233
rect 28526 -24534 28572 -24434
rect 28722 -24534 28768 -24434
rect 28918 -24534 28964 -24434
rect 29114 -24534 29160 -24434
rect 28119 -24808 28302 -24767
rect 29422 -24808 29518 -24779
rect 28119 -24890 29518 -24808
rect 28119 -24897 28302 -24890
rect 29422 -24916 29518 -24890
rect 26918 -25433 26964 -25133
rect 27114 -25433 27160 -25133
rect 27310 -25433 27356 -25133
rect 27527 -25232 27573 -25132
rect 27723 -25232 27769 -25132
rect 27919 -25232 27965 -25132
rect 28115 -25232 28161 -25132
rect 28365 -25644 28411 -25044
rect 28561 -25644 28607 -25044
rect 28984 -25644 29030 -25044
rect 30612 -24435 30658 -24235
rect 30808 -24435 30854 -24235
rect 31004 -24435 31050 -24235
rect 31200 -24435 31246 -24235
rect 31585 -24564 31631 -24264
rect 31781 -24564 31827 -24264
rect 31977 -24564 32023 -24264
rect 32194 -24565 32240 -24465
rect 32390 -24565 32436 -24465
rect 32586 -24565 32632 -24465
rect 32782 -24565 32828 -24465
rect 32842 -24830 32933 -24818
rect 33092 -24830 33243 -24803
rect 32842 -24969 33243 -24830
rect 32842 -24981 32933 -24969
rect 33092 -24994 33243 -24969
rect 30586 -25464 30632 -25164
rect 30782 -25464 30828 -25164
rect 30978 -25464 31024 -25164
rect 31195 -25263 31241 -25163
rect 31391 -25263 31437 -25163
rect 31587 -25263 31633 -25163
rect 31783 -25263 31829 -25163
rect 32033 -25675 32079 -25075
rect 32229 -25675 32275 -25075
rect 32652 -25675 32698 -25075
rect 35392 -20962 35438 -20762
rect 35588 -20962 35634 -20762
rect 35784 -20962 35830 -20762
rect 35980 -20962 36026 -20762
rect 36365 -21091 36411 -20791
rect 36561 -21091 36607 -20791
rect 36757 -21091 36803 -20791
rect 36974 -21092 37020 -20992
rect 37170 -21092 37216 -20992
rect 37366 -21092 37412 -20992
rect 37562 -21092 37608 -20992
rect 37644 -21407 37718 -21391
rect 37872 -21407 37982 -21371
rect 37644 -21503 37982 -21407
rect 37644 -21509 37718 -21503
rect 37872 -21521 37982 -21503
rect 35366 -21991 35412 -21691
rect 35562 -21991 35608 -21691
rect 35758 -21991 35804 -21691
rect 35975 -21790 36021 -21690
rect 36171 -21790 36217 -21690
rect 36367 -21790 36413 -21690
rect 36563 -21790 36609 -21690
rect 36813 -22202 36859 -21602
rect 37009 -22202 37055 -21602
rect 37432 -22202 37478 -21602
rect 38805 -21960 38851 -21460
rect 39001 -21960 39047 -21460
rect 39596 -21960 39642 -21460
rect 39726 -21960 39772 -21460
rect 39954 -21760 40000 -21460
rect 40150 -21760 40196 -21460
rect 35384 -24415 35430 -24215
rect 35580 -24415 35626 -24215
rect 35776 -24415 35822 -24215
rect 35972 -24415 36018 -24215
rect 36357 -24544 36403 -24244
rect 36553 -24544 36599 -24244
rect 36749 -24544 36795 -24244
rect 36966 -24545 37012 -24445
rect 37162 -24545 37208 -24445
rect 37358 -24545 37404 -24445
rect 37554 -24545 37600 -24445
rect 36559 -24819 36742 -24778
rect 37862 -24819 37958 -24790
rect 36559 -24901 37958 -24819
rect 36559 -24908 36742 -24901
rect 37862 -24927 37958 -24901
rect 35358 -25444 35404 -25144
rect 35554 -25444 35600 -25144
rect 35750 -25444 35796 -25144
rect 35967 -25243 36013 -25143
rect 36163 -25243 36209 -25143
rect 36359 -25243 36405 -25143
rect 36555 -25243 36601 -25143
rect 36805 -25655 36851 -25055
rect 37001 -25655 37047 -25055
rect 37424 -25655 37470 -25055
rect 39052 -24446 39098 -24246
rect 39248 -24446 39294 -24246
rect 39444 -24446 39490 -24246
rect 39640 -24446 39686 -24246
rect 40025 -24575 40071 -24275
rect 40221 -24575 40267 -24275
rect 40417 -24575 40463 -24275
rect 40634 -24576 40680 -24476
rect 40830 -24576 40876 -24476
rect 41026 -24576 41072 -24476
rect 41222 -24576 41268 -24476
rect 41282 -24841 41373 -24829
rect 41532 -24841 41683 -24814
rect 41282 -24980 41683 -24841
rect 41282 -24992 41373 -24980
rect 41532 -25005 41683 -24980
rect 39026 -25475 39072 -25175
rect 39222 -25475 39268 -25175
rect 39418 -25475 39464 -25175
rect 39635 -25274 39681 -25174
rect 39831 -25274 39877 -25174
rect 40027 -25274 40073 -25174
rect 40223 -25274 40269 -25174
rect 40473 -25686 40519 -25086
rect 40669 -25686 40715 -25086
rect 41092 -25686 41138 -25086
rect 44255 -21001 44301 -20801
rect 44451 -21001 44497 -20801
rect 44647 -21001 44693 -20801
rect 44843 -21001 44889 -20801
rect 45228 -21130 45274 -20830
rect 45424 -21130 45470 -20830
rect 45620 -21130 45666 -20830
rect 45837 -21131 45883 -21031
rect 46033 -21131 46079 -21031
rect 46229 -21131 46275 -21031
rect 46425 -21131 46471 -21031
rect 46507 -21446 46581 -21430
rect 46735 -21446 46845 -21410
rect 46507 -21542 46845 -21446
rect 46507 -21548 46581 -21542
rect 46735 -21560 46845 -21542
rect 44229 -22030 44275 -21730
rect 44425 -22030 44471 -21730
rect 44621 -22030 44667 -21730
rect 44838 -21829 44884 -21729
rect 45034 -21829 45080 -21729
rect 45230 -21829 45276 -21729
rect 45426 -21829 45472 -21729
rect 45676 -22241 45722 -21641
rect 45872 -22241 45918 -21641
rect 46295 -22241 46341 -21641
rect 47668 -21999 47714 -21499
rect 47864 -21999 47910 -21499
rect 48459 -21999 48505 -21499
rect 48589 -21999 48635 -21499
rect 48817 -21799 48863 -21499
rect 49013 -21799 49059 -21499
rect 44247 -24454 44293 -24254
rect 44443 -24454 44489 -24254
rect 44639 -24454 44685 -24254
rect 44835 -24454 44881 -24254
rect 45220 -24583 45266 -24283
rect 45416 -24583 45462 -24283
rect 45612 -24583 45658 -24283
rect 45829 -24584 45875 -24484
rect 46025 -24584 46071 -24484
rect 46221 -24584 46267 -24484
rect 46417 -24584 46463 -24484
rect 45422 -24858 45605 -24817
rect 46725 -24858 46821 -24829
rect 45422 -24940 46821 -24858
rect 45422 -24947 45605 -24940
rect 46725 -24966 46821 -24940
rect 44221 -25483 44267 -25183
rect 44417 -25483 44463 -25183
rect 44613 -25483 44659 -25183
rect 44830 -25282 44876 -25182
rect 45026 -25282 45072 -25182
rect 45222 -25282 45268 -25182
rect 45418 -25282 45464 -25182
rect 45668 -25694 45714 -25094
rect 45864 -25694 45910 -25094
rect 46287 -25694 46333 -25094
rect 47915 -24485 47961 -24285
rect 48111 -24485 48157 -24285
rect 48307 -24485 48353 -24285
rect 48503 -24485 48549 -24285
rect 48888 -24614 48934 -24314
rect 49084 -24614 49130 -24314
rect 49280 -24614 49326 -24314
rect 49497 -24615 49543 -24515
rect 49693 -24615 49739 -24515
rect 49889 -24615 49935 -24515
rect 50085 -24615 50131 -24515
rect 50145 -24880 50236 -24868
rect 50395 -24880 50546 -24853
rect 50145 -25019 50546 -24880
rect 50145 -25031 50236 -25019
rect 50395 -25044 50546 -25019
rect 47889 -25514 47935 -25214
rect 48085 -25514 48131 -25214
rect 48281 -25514 48327 -25214
rect 48498 -25313 48544 -25213
rect 48694 -25313 48740 -25213
rect 48890 -25313 48936 -25213
rect 49086 -25313 49132 -25213
rect 49336 -25725 49382 -25125
rect 49532 -25725 49578 -25125
rect 49955 -25725 50001 -25125
rect 53453 -20967 53499 -20767
rect 53649 -20967 53695 -20767
rect 53845 -20967 53891 -20767
rect 54041 -20967 54087 -20767
rect 54426 -21096 54472 -20796
rect 54622 -21096 54668 -20796
rect 54818 -21096 54864 -20796
rect 55035 -21097 55081 -20997
rect 55231 -21097 55277 -20997
rect 55427 -21097 55473 -20997
rect 55623 -21097 55669 -20997
rect 55705 -21412 55779 -21396
rect 55933 -21412 56043 -21376
rect 55705 -21508 56043 -21412
rect 55705 -21514 55779 -21508
rect 55933 -21526 56043 -21508
rect 53427 -21996 53473 -21696
rect 53623 -21996 53669 -21696
rect 53819 -21996 53865 -21696
rect 54036 -21795 54082 -21695
rect 54232 -21795 54278 -21695
rect 54428 -21795 54474 -21695
rect 54624 -21795 54670 -21695
rect 54874 -22207 54920 -21607
rect 55070 -22207 55116 -21607
rect 55493 -22207 55539 -21607
rect 56866 -21965 56912 -21465
rect 57062 -21965 57108 -21465
rect 57657 -21965 57703 -21465
rect 57787 -21965 57833 -21465
rect 58015 -21765 58061 -21465
rect 58211 -21765 58257 -21465
rect 53445 -24420 53491 -24220
rect 53641 -24420 53687 -24220
rect 53837 -24420 53883 -24220
rect 54033 -24420 54079 -24220
rect 54418 -24549 54464 -24249
rect 54614 -24549 54660 -24249
rect 54810 -24549 54856 -24249
rect 55027 -24550 55073 -24450
rect 55223 -24550 55269 -24450
rect 55419 -24550 55465 -24450
rect 55615 -24550 55661 -24450
rect 54620 -24824 54803 -24783
rect 55923 -24824 56019 -24795
rect 54620 -24906 56019 -24824
rect 54620 -24913 54803 -24906
rect 55923 -24932 56019 -24906
rect 53419 -25449 53465 -25149
rect 53615 -25449 53661 -25149
rect 53811 -25449 53857 -25149
rect 54028 -25248 54074 -25148
rect 54224 -25248 54270 -25148
rect 54420 -25248 54466 -25148
rect 54616 -25248 54662 -25148
rect 54866 -25660 54912 -25060
rect 55062 -25660 55108 -25060
rect 55485 -25660 55531 -25060
rect 57113 -24451 57159 -24251
rect 57309 -24451 57355 -24251
rect 57505 -24451 57551 -24251
rect 57701 -24451 57747 -24251
rect 58086 -24580 58132 -24280
rect 58282 -24580 58328 -24280
rect 58478 -24580 58524 -24280
rect 58695 -24581 58741 -24481
rect 58891 -24581 58937 -24481
rect 59087 -24581 59133 -24481
rect 59283 -24581 59329 -24481
rect 59343 -24846 59434 -24834
rect 59593 -24846 59744 -24819
rect 59343 -24985 59744 -24846
rect 59343 -24997 59434 -24985
rect 59593 -25010 59744 -24985
rect 57087 -25480 57133 -25180
rect 57283 -25480 57329 -25180
rect 57479 -25480 57525 -25180
rect 57696 -25279 57742 -25179
rect 57892 -25279 57938 -25179
rect 58088 -25279 58134 -25179
rect 58284 -25279 58330 -25179
rect 58534 -25691 58580 -25091
rect 58730 -25691 58776 -25091
rect 59153 -25691 59199 -25091
rect 62207 -20901 62253 -20701
rect 62403 -20901 62449 -20701
rect 62599 -20901 62645 -20701
rect 62795 -20901 62841 -20701
rect 63180 -21030 63226 -20730
rect 63376 -21030 63422 -20730
rect 63572 -21030 63618 -20730
rect 63789 -21031 63835 -20931
rect 63985 -21031 64031 -20931
rect 64181 -21031 64227 -20931
rect 64377 -21031 64423 -20931
rect 64459 -21346 64533 -21330
rect 64687 -21346 64797 -21310
rect 64459 -21442 64797 -21346
rect 64459 -21448 64533 -21442
rect 64687 -21460 64797 -21442
rect 62181 -21930 62227 -21630
rect 62377 -21930 62423 -21630
rect 62573 -21930 62619 -21630
rect 62790 -21729 62836 -21629
rect 62986 -21729 63032 -21629
rect 63182 -21729 63228 -21629
rect 63378 -21729 63424 -21629
rect 63628 -22141 63674 -21541
rect 63824 -22141 63870 -21541
rect 64247 -22141 64293 -21541
rect 65620 -21899 65666 -21399
rect 65816 -21899 65862 -21399
rect 66411 -21899 66457 -21399
rect 66541 -21899 66587 -21399
rect 66769 -21699 66815 -21399
rect 66965 -21699 67011 -21399
rect 62199 -24354 62245 -24154
rect 62395 -24354 62441 -24154
rect 62591 -24354 62637 -24154
rect 62787 -24354 62833 -24154
rect 63172 -24483 63218 -24183
rect 63368 -24483 63414 -24183
rect 63564 -24483 63610 -24183
rect 63781 -24484 63827 -24384
rect 63977 -24484 64023 -24384
rect 64173 -24484 64219 -24384
rect 64369 -24484 64415 -24384
rect 63374 -24758 63557 -24717
rect 64677 -24758 64773 -24729
rect 63374 -24840 64773 -24758
rect 63374 -24847 63557 -24840
rect 64677 -24866 64773 -24840
rect 62173 -25383 62219 -25083
rect 62369 -25383 62415 -25083
rect 62565 -25383 62611 -25083
rect 62782 -25182 62828 -25082
rect 62978 -25182 63024 -25082
rect 63174 -25182 63220 -25082
rect 63370 -25182 63416 -25082
rect 63620 -25594 63666 -24994
rect 63816 -25594 63862 -24994
rect 64239 -25594 64285 -24994
rect 65867 -24385 65913 -24185
rect 66063 -24385 66109 -24185
rect 66259 -24385 66305 -24185
rect 66455 -24385 66501 -24185
rect 66840 -24514 66886 -24214
rect 67036 -24514 67082 -24214
rect 67232 -24514 67278 -24214
rect 67449 -24515 67495 -24415
rect 67645 -24515 67691 -24415
rect 67841 -24515 67887 -24415
rect 68037 -24515 68083 -24415
rect 68097 -24780 68188 -24768
rect 68347 -24780 68498 -24753
rect 68097 -24919 68498 -24780
rect 68097 -24931 68188 -24919
rect 68347 -24944 68498 -24919
rect 65841 -25414 65887 -25114
rect 66037 -25414 66083 -25114
rect 66233 -25414 66279 -25114
rect 66450 -25213 66496 -25113
rect 66646 -25213 66692 -25113
rect 66842 -25213 66888 -25113
rect 67038 -25213 67084 -25113
rect 67288 -25625 67334 -25025
rect 67484 -25625 67530 -25025
rect 67907 -25625 67953 -25025
rect 71360 -20884 71406 -20684
rect 71556 -20884 71602 -20684
rect 71752 -20884 71798 -20684
rect 71948 -20884 71994 -20684
rect 72333 -21013 72379 -20713
rect 72529 -21013 72575 -20713
rect 72725 -21013 72771 -20713
rect 72942 -21014 72988 -20914
rect 73138 -21014 73184 -20914
rect 73334 -21014 73380 -20914
rect 73530 -21014 73576 -20914
rect 73612 -21329 73686 -21313
rect 73840 -21329 73950 -21293
rect 73612 -21425 73950 -21329
rect 73612 -21431 73686 -21425
rect 73840 -21443 73950 -21425
rect 71334 -21913 71380 -21613
rect 71530 -21913 71576 -21613
rect 71726 -21913 71772 -21613
rect 71943 -21712 71989 -21612
rect 72139 -21712 72185 -21612
rect 72335 -21712 72381 -21612
rect 72531 -21712 72577 -21612
rect 72781 -22124 72827 -21524
rect 72977 -22124 73023 -21524
rect 73400 -22124 73446 -21524
rect 74773 -21882 74819 -21382
rect 74969 -21882 75015 -21382
rect 75564 -21882 75610 -21382
rect 75694 -21882 75740 -21382
rect 75922 -21682 75968 -21382
rect 76118 -21682 76164 -21382
rect 71352 -24337 71398 -24137
rect 71548 -24337 71594 -24137
rect 71744 -24337 71790 -24137
rect 71940 -24337 71986 -24137
rect 72325 -24466 72371 -24166
rect 72521 -24466 72567 -24166
rect 72717 -24466 72763 -24166
rect 72934 -24467 72980 -24367
rect 73130 -24467 73176 -24367
rect 73326 -24467 73372 -24367
rect 73522 -24467 73568 -24367
rect 72527 -24741 72710 -24700
rect 73830 -24741 73926 -24712
rect 72527 -24823 73926 -24741
rect 72527 -24830 72710 -24823
rect 73830 -24849 73926 -24823
rect 71326 -25366 71372 -25066
rect 71522 -25366 71568 -25066
rect 71718 -25366 71764 -25066
rect 71935 -25165 71981 -25065
rect 72131 -25165 72177 -25065
rect 72327 -25165 72373 -25065
rect 72523 -25165 72569 -25065
rect 72773 -25577 72819 -24977
rect 72969 -25577 73015 -24977
rect 73392 -25577 73438 -24977
rect 75020 -24368 75066 -24168
rect 75216 -24368 75262 -24168
rect 75412 -24368 75458 -24168
rect 75608 -24368 75654 -24168
rect 75993 -24497 76039 -24197
rect 76189 -24497 76235 -24197
rect 76385 -24497 76431 -24197
rect 76602 -24498 76648 -24398
rect 76798 -24498 76844 -24398
rect 76994 -24498 77040 -24398
rect 77190 -24498 77236 -24398
rect 77250 -24763 77341 -24751
rect 77500 -24763 77651 -24736
rect 77250 -24902 77651 -24763
rect 77250 -24914 77341 -24902
rect 77500 -24927 77651 -24902
rect 74994 -25397 75040 -25097
rect 75190 -25397 75236 -25097
rect 75386 -25397 75432 -25097
rect 75603 -25196 75649 -25096
rect 75799 -25196 75845 -25096
rect 75995 -25196 76041 -25096
rect 76191 -25196 76237 -25096
rect 76441 -25608 76487 -25008
rect 76637 -25608 76683 -25008
rect 77060 -25608 77106 -25008
rect 80724 -20846 80770 -20646
rect 80920 -20846 80966 -20646
rect 81116 -20846 81162 -20646
rect 81312 -20846 81358 -20646
rect 81697 -20975 81743 -20675
rect 81893 -20975 81939 -20675
rect 82089 -20975 82135 -20675
rect 82306 -20976 82352 -20876
rect 82502 -20976 82548 -20876
rect 82698 -20976 82744 -20876
rect 82894 -20976 82940 -20876
rect 82976 -21291 83050 -21275
rect 83204 -21291 83314 -21255
rect 82976 -21387 83314 -21291
rect 82976 -21393 83050 -21387
rect 83204 -21405 83314 -21387
rect 80698 -21875 80744 -21575
rect 80894 -21875 80940 -21575
rect 81090 -21875 81136 -21575
rect 81307 -21674 81353 -21574
rect 81503 -21674 81549 -21574
rect 81699 -21674 81745 -21574
rect 81895 -21674 81941 -21574
rect 82145 -22086 82191 -21486
rect 82341 -22086 82387 -21486
rect 82764 -22086 82810 -21486
rect 84137 -21844 84183 -21344
rect 84333 -21844 84379 -21344
rect 84928 -21844 84974 -21344
rect 85058 -21844 85104 -21344
rect 85286 -21644 85332 -21344
rect 85482 -21644 85528 -21344
rect 80716 -24299 80762 -24099
rect 80912 -24299 80958 -24099
rect 81108 -24299 81154 -24099
rect 81304 -24299 81350 -24099
rect 81689 -24428 81735 -24128
rect 81885 -24428 81931 -24128
rect 82081 -24428 82127 -24128
rect 82298 -24429 82344 -24329
rect 82494 -24429 82540 -24329
rect 82690 -24429 82736 -24329
rect 82886 -24429 82932 -24329
rect 81891 -24703 82074 -24662
rect 83194 -24703 83290 -24674
rect 81891 -24785 83290 -24703
rect 81891 -24792 82074 -24785
rect 83194 -24811 83290 -24785
rect 80690 -25328 80736 -25028
rect 80886 -25328 80932 -25028
rect 81082 -25328 81128 -25028
rect 81299 -25127 81345 -25027
rect 81495 -25127 81541 -25027
rect 81691 -25127 81737 -25027
rect 81887 -25127 81933 -25027
rect 82137 -25539 82183 -24939
rect 82333 -25539 82379 -24939
rect 82756 -25539 82802 -24939
rect 84384 -24330 84430 -24130
rect 84580 -24330 84626 -24130
rect 84776 -24330 84822 -24130
rect 84972 -24330 85018 -24130
rect 85357 -24459 85403 -24159
rect 85553 -24459 85599 -24159
rect 85749 -24459 85795 -24159
rect 85966 -24460 86012 -24360
rect 86162 -24460 86208 -24360
rect 86358 -24460 86404 -24360
rect 86554 -24460 86600 -24360
rect 86614 -24725 86705 -24713
rect 86864 -24725 87015 -24698
rect 86614 -24864 87015 -24725
rect 86614 -24876 86705 -24864
rect 86864 -24889 87015 -24864
rect 84358 -25359 84404 -25059
rect 84554 -25359 84600 -25059
rect 84750 -25359 84796 -25059
rect 84967 -25158 85013 -25058
rect 85163 -25158 85209 -25058
rect 85359 -25158 85405 -25058
rect 85555 -25158 85601 -25058
rect 85805 -25570 85851 -24970
rect 86001 -25570 86047 -24970
rect 86424 -25570 86470 -24970
rect 89990 -7667 92959 -4698
rect -26157 -34013 -26083 -33984
rect -26157 -34059 -25612 -34013
rect -26157 -34249 -26083 -34059
rect -26012 -34177 -25612 -34131
rect -26157 -34295 -25612 -34249
rect -26157 -34485 -26083 -34295
rect -26012 -34413 -25612 -34367
rect -26157 -34531 -25612 -34485
rect -26157 -34721 -26083 -34531
rect -26012 -34649 -25612 -34603
rect -26157 -34767 -25612 -34721
rect -26157 -34957 -26083 -34767
rect -26012 -34885 -25612 -34839
rect -26157 -35003 -25612 -34957
rect -26157 -35193 -26083 -35003
rect -26012 -35121 -25612 -35075
rect -26157 -35239 -25612 -35193
rect -26157 -35429 -26083 -35239
rect -26012 -35357 -25612 -35311
rect -26157 -35475 -25612 -35429
rect -26157 -35665 -26083 -35475
rect -26012 -35593 -25612 -35547
rect -26157 -35711 -25612 -35665
rect -26157 -35901 -26083 -35711
rect -26012 -35829 -25612 -35783
rect -26157 -35947 -25612 -35901
rect -26157 -36137 -26083 -35947
rect -26012 -36065 -25612 -36019
rect -26157 -36183 -25612 -36137
rect -26157 -36373 -26083 -36183
rect -26012 -36301 -25612 -36255
rect -26157 -36419 -25612 -36373
rect -26157 -36609 -26083 -36419
rect -26012 -36537 -25612 -36491
rect -26157 -36655 -25612 -36609
rect -26157 -36845 -26083 -36655
rect -26012 -36773 -25612 -36727
rect -26157 -36891 -25612 -36845
rect -26157 -37081 -26083 -36891
rect -26012 -37009 -25612 -36963
rect -26157 -37127 -25612 -37081
rect -26157 -37317 -26083 -37127
rect -26012 -37245 -25612 -37199
rect -23334 -37202 -23233 -37147
rect -26157 -37363 -25612 -37317
rect -26157 -37553 -26083 -37363
rect -23486 -37390 -23233 -37202
rect -23486 -37433 -23246 -37390
rect -26012 -37481 -25612 -37435
rect -26157 -37599 -25612 -37553
rect -26157 -37769 -26083 -37599
rect -26012 -37717 -25612 -37671
rect -26820 -37789 -26083 -37769
rect -26820 -37815 -25612 -37789
rect -26319 -38005 -26273 -37815
rect -26157 -37835 -25612 -37815
rect -26157 -37861 -26083 -37835
rect -26820 -38051 -26273 -38005
rect -26319 -38241 -26273 -38051
rect -26820 -38287 -26273 -38241
rect -26319 -38477 -26273 -38287
rect -26820 -38523 -26273 -38477
rect -26319 -38713 -26273 -38523
rect -26820 -38759 -26273 -38713
rect -26319 -38949 -26273 -38759
rect -26820 -38995 -26273 -38949
rect -26319 -39185 -26273 -38995
rect -26820 -39231 -26273 -39185
rect -26319 -39421 -26273 -39231
rect -26820 -39467 -26273 -39421
rect -26012 -37965 -25612 -37919
rect -26012 -38201 -25612 -38155
rect -26012 -38437 -25612 -38391
rect -26012 -38673 -25612 -38627
rect -26012 -38909 -25612 -38863
rect -26012 -39145 -25612 -39099
rect -26012 -39381 -25612 -39335
rect -26012 -39617 -25612 -39571
rect -26012 -39853 -25612 -39807
rect -26012 -39983 -25612 -39937
rect -26012 -40219 -25612 -40173
rect -26012 -40455 -25612 -40409
rect -26012 -40691 -25612 -40645
rect -26012 -40927 -25612 -40881
rect -26012 -41057 -25612 -41011
rect -26012 -41293 -25612 -41247
rect -26012 -41529 -25612 -41483
rect -23486 -46358 -23350 -37433
rect -23186 -44515 -23125 -35988
rect -23239 -44638 -23116 -44515
rect -22995 -44714 -22934 -35909
rect -22886 -36061 -22825 -35823
rect -22046 -35975 -22000 -35775
rect -21850 -35975 -21804 -35775
rect -21654 -35975 -21608 -35775
rect -21458 -35975 -21412 -35775
rect -20916 -35975 -20870 -35775
rect -20720 -35975 -20674 -35775
rect -14447 -35188 -14401 -34988
rect -14251 -35188 -14205 -34988
rect -14055 -35188 -14009 -34988
rect -13610 -35188 -13564 -34988
rect -13414 -35188 -13368 -34988
rect -13218 -35188 -13172 -34988
rect -11747 -35188 -11701 -34988
rect -11551 -35188 -11505 -34988
rect -11355 -35188 -11309 -34988
rect -10910 -35188 -10864 -34988
rect -10714 -35188 -10668 -34988
rect -10518 -35188 -10472 -34988
rect -22886 -41890 -22826 -36061
rect -20047 -36197 -20001 -35897
rect -19851 -36197 -19805 -35897
rect -22886 -42127 -22825 -41890
rect -23048 -44837 -22925 -44714
rect -22886 -44947 -22826 -42127
rect -22942 -45070 -22819 -44947
rect -22787 -45204 -22726 -36988
rect -22849 -45327 -22725 -45204
rect -21989 -38106 -21943 -37806
rect -21793 -38106 -21747 -37806
rect -21597 -38106 -21551 -37806
rect -21380 -37905 -21334 -37805
rect -21184 -37905 -21138 -37805
rect -20988 -37905 -20942 -37805
rect -20792 -37905 -20746 -37805
rect -20261 -36400 -20124 -36342
rect -20254 -37173 -20214 -36400
rect -19655 -36197 -19609 -35897
rect -19438 -35996 -19392 -35896
rect -19242 -35996 -19196 -35896
rect -19046 -35996 -19000 -35896
rect -18850 -35996 -18804 -35896
rect -20370 -37182 -20214 -37173
rect -20417 -37222 -20214 -37182
rect -20370 -37226 -20238 -37222
rect -20216 -37911 -20170 -37711
rect -20020 -37911 -19974 -37711
rect -19824 -37911 -19778 -37711
rect -19628 -37911 -19582 -37711
rect -19086 -37911 -19040 -37711
rect -18890 -37911 -18844 -37711
rect -18411 -37159 -18365 -36859
rect -18215 -37159 -18169 -36859
rect -18019 -37159 -17973 -36859
rect -17802 -37160 -17756 -37060
rect -17606 -37160 -17560 -37060
rect -17410 -37160 -17364 -37060
rect -17214 -37160 -17168 -37060
rect -16964 -37248 -16918 -36648
rect -16768 -37248 -16722 -36648
rect -16345 -37248 -16299 -36648
rect -18385 -38088 -18339 -37888
rect -18189 -38088 -18143 -37888
rect -17993 -38088 -17947 -37888
rect -17797 -38088 -17751 -37888
rect -17412 -38059 -17366 -37759
rect -17216 -38059 -17170 -37759
rect -17020 -38059 -16974 -37759
rect -16803 -37858 -16757 -37758
rect -16607 -37858 -16561 -37758
rect -16411 -37858 -16365 -37758
rect -16215 -37858 -16169 -37758
rect -8085 -35598 -8039 -34998
rect -7662 -35598 -7616 -34998
rect -7466 -35598 -7420 -34998
rect -5977 -35394 -5931 -35194
rect -5781 -35394 -5735 -35194
rect -5585 -35394 -5539 -35194
rect -5471 -35394 -5425 -35194
rect -5275 -35394 -5229 -35194
rect -5162 -35394 -5116 -35194
rect -4966 -35394 -4920 -35194
rect -3477 -35394 -3431 -35194
rect -3281 -35394 -3235 -35194
rect -3085 -35394 -3039 -35194
rect -2971 -35394 -2925 -35194
rect -2775 -35394 -2729 -35194
rect -2662 -35394 -2616 -35194
rect -2466 -35394 -2420 -35194
rect -977 -35394 -931 -35194
rect -781 -35394 -735 -35194
rect -585 -35394 -539 -35194
rect -471 -35394 -425 -35194
rect -275 -35394 -229 -35194
rect -162 -35394 -116 -35194
rect 34 -35394 80 -35194
rect 1523 -35394 1569 -35194
rect 1719 -35394 1765 -35194
rect 1915 -35394 1961 -35194
rect 2029 -35394 2075 -35194
rect 2225 -35394 2271 -35194
rect 2338 -35394 2384 -35194
rect 2534 -35394 2580 -35194
rect 4023 -35394 4069 -35194
rect 4219 -35394 4265 -35194
rect 4415 -35394 4461 -35194
rect 4529 -35394 4575 -35194
rect 4725 -35394 4771 -35194
rect 4838 -35394 4884 -35194
rect 5034 -35394 5080 -35194
rect 7023 -35394 7069 -35194
rect 7219 -35394 7265 -35194
rect 7415 -35394 7461 -35194
rect 7529 -35394 7575 -35194
rect 7725 -35394 7771 -35194
rect 7838 -35394 7884 -35194
rect 8034 -35394 8080 -35194
rect -14349 -36506 -14303 -36306
rect -14153 -36506 -14107 -36306
rect -13957 -36506 -13911 -36306
rect -12606 -36506 -12560 -36306
rect -12410 -36506 -12364 -36306
rect -12214 -36506 -12168 -36306
rect -11649 -36506 -11603 -36306
rect -11453 -36506 -11407 -36306
rect -11257 -36506 -11211 -36306
rect -9906 -36506 -9860 -36306
rect -9710 -36506 -9664 -36306
rect -9514 -36506 -9468 -36306
rect -9024 -36506 -8978 -36306
rect -8828 -36506 -8782 -36306
rect -8632 -36506 -8586 -36306
rect -13677 -37694 -13480 -37640
rect -18872 -40620 -18693 -40453
rect -21924 -41600 -21878 -41000
rect -21728 -41600 -21682 -41000
rect -20718 -41329 -20672 -40929
rect -20522 -41329 -20476 -40929
rect -19813 -41330 -19767 -40930
rect -19617 -41330 -19571 -40930
rect -20892 -41491 -20834 -41354
rect -20892 -42400 -20857 -41491
rect -20912 -42537 -20854 -42400
rect -22261 -44018 -22215 -43818
rect -22065 -44018 -22019 -43818
rect -21523 -44018 -21477 -43818
rect -21327 -44018 -21281 -43818
rect -21131 -44018 -21085 -43818
rect -20935 -44018 -20889 -43818
rect -19651 -44182 -19475 -43551
rect -18845 -42384 -18719 -40620
rect -13534 -38725 -13480 -37694
rect -13422 -38135 -13376 -37835
rect -13226 -38135 -13180 -37835
rect -13030 -38135 -12984 -37835
rect -12813 -38136 -12767 -38036
rect -12617 -38136 -12571 -38036
rect -12421 -38136 -12375 -38036
rect -12225 -38136 -12179 -38036
rect -11975 -38224 -11929 -37624
rect -11779 -38224 -11733 -37624
rect -11356 -38224 -11310 -37624
rect -15145 -38901 -13480 -38725
rect -18846 -42556 -18654 -42384
rect -18411 -42159 -18365 -41859
rect -18215 -42159 -18169 -41859
rect -18019 -42159 -17973 -41859
rect -17802 -42160 -17756 -42060
rect -17606 -42160 -17560 -42060
rect -17410 -42160 -17364 -42060
rect -17214 -42160 -17168 -42060
rect -16964 -42248 -16918 -41648
rect -16768 -42248 -16722 -41648
rect -16345 -42248 -16299 -41648
rect -18385 -43088 -18339 -42888
rect -18189 -43088 -18143 -42888
rect -17993 -43088 -17947 -42888
rect -17797 -43088 -17751 -42888
rect -17412 -43059 -17366 -42759
rect -17216 -43059 -17170 -42759
rect -17020 -43059 -16974 -42759
rect -16803 -42858 -16757 -42758
rect -16607 -42858 -16561 -42758
rect -16411 -42858 -16365 -42758
rect -16215 -42858 -16169 -42758
rect -15145 -44640 -14969 -38901
rect -13534 -39098 -13480 -38901
rect -13396 -39064 -13350 -38864
rect -13584 -39248 -13454 -39098
rect -13200 -39064 -13154 -38864
rect -13004 -39064 -12958 -38864
rect -12808 -39064 -12762 -38864
rect -12423 -39035 -12377 -38735
rect -12227 -39035 -12181 -38735
rect -12031 -39035 -11985 -38735
rect -11814 -38834 -11768 -38734
rect -11618 -38834 -11572 -38734
rect -11422 -38834 -11376 -38734
rect -11226 -38834 -11180 -38734
rect -14447 -40115 -14401 -39915
rect -14251 -40115 -14205 -39915
rect -14055 -40115 -14009 -39915
rect -13610 -40115 -13564 -39915
rect -13414 -40115 -13368 -39915
rect -13218 -40115 -13172 -39915
rect -11747 -40115 -11701 -39915
rect -11551 -40115 -11505 -39915
rect -11355 -40115 -11309 -39915
rect -10910 -40115 -10864 -39915
rect -10714 -40115 -10668 -39915
rect -10518 -40115 -10472 -39915
rect -14349 -41433 -14303 -41233
rect -14153 -41433 -14107 -41233
rect -13957 -41433 -13911 -41233
rect -12606 -41433 -12560 -41233
rect -12410 -41433 -12364 -41233
rect -12214 -41433 -12168 -41233
rect -11649 -41433 -11603 -41233
rect -11453 -41433 -11407 -41233
rect -11257 -41433 -11211 -41233
rect -9906 -41433 -9860 -41233
rect -9710 -41433 -9664 -41233
rect -9514 -41433 -9468 -41233
rect -9024 -41433 -8978 -41233
rect -8828 -41433 -8782 -41233
rect -8632 -41433 -8586 -41233
rect -8058 -40532 -8012 -39932
rect -7635 -40532 -7589 -39932
rect -7439 -40532 -7393 -39932
rect -6442 -36455 -6306 -36381
rect -6442 -36837 -6391 -36455
rect -6316 -36723 -6270 -36523
rect -6120 -36723 -6074 -36523
rect -5924 -36723 -5878 -36523
rect -4649 -35952 -4526 -35816
rect -4645 -36583 -4531 -35952
rect -4650 -36719 -4527 -36583
rect -2082 -35987 -1959 -35851
rect -2078 -36439 -1964 -35987
rect -2083 -36575 -1960 -36439
rect 401 -35987 524 -35851
rect 405 -36404 519 -35987
rect 400 -36405 523 -36404
rect 400 -36467 706 -36405
rect 3634 -35661 3773 -35652
rect 4712 -35659 4851 -35658
rect 4712 -35661 6071 -35659
rect 3634 -35687 6071 -35661
rect 3634 -35689 4851 -35687
rect 3634 -35706 3773 -35689
rect 4712 -35712 4851 -35689
rect 6043 -36285 6071 -35687
rect 6634 -35661 6773 -35652
rect 7712 -35659 7851 -35658
rect 7610 -35661 10221 -35659
rect 6634 -35687 10221 -35661
rect 6634 -35689 7851 -35687
rect 6634 -35706 6773 -35689
rect 7712 -35712 7851 -35689
rect 6043 -36313 10070 -36285
rect -6442 -36888 9423 -36837
rect -665 -37145 9298 -37094
rect 4065 -37246 4188 -37237
rect 4466 -37246 4589 -37235
rect -824 -37261 -701 -37249
rect -530 -37261 -407 -37248
rect -824 -37376 -407 -37261
rect -824 -37385 -701 -37376
rect -530 -37384 -407 -37376
rect 2448 -37276 2571 -37261
rect 2837 -37276 2960 -37260
rect 2448 -37383 2960 -37276
rect 4065 -37353 4589 -37246
rect 4065 -37373 4188 -37353
rect 4466 -37371 4589 -37353
rect 5822 -37253 5945 -37240
rect 7038 -37253 7161 -37241
rect 5822 -37358 7161 -37253
rect 5822 -37376 5945 -37358
rect 7038 -37377 7161 -37358
rect 2448 -37397 2571 -37383
rect 2837 -37396 2960 -37383
rect -6475 -37626 -6429 -37426
rect -6279 -37626 -6233 -37426
rect -6083 -37626 -6037 -37426
rect -4732 -37626 -4686 -37426
rect -4536 -37626 -4490 -37426
rect -4340 -37626 -4294 -37426
rect -3775 -37626 -3729 -37426
rect -3579 -37626 -3533 -37426
rect -3383 -37626 -3337 -37426
rect -2032 -37626 -1986 -37426
rect -1836 -37626 -1790 -37426
rect -1640 -37626 -1594 -37426
rect -1150 -37626 -1104 -37426
rect -954 -37626 -908 -37426
rect -758 -37626 -712 -37426
rect -416 -37643 -370 -37443
rect -220 -37643 -174 -37443
rect 322 -37643 368 -37443
rect 518 -37643 564 -37443
rect 714 -37643 760 -37443
rect 910 -37643 956 -37443
rect 1317 -37556 1363 -37456
rect -5950 -38123 -5818 -38063
rect -5914 -38590 -5854 -38123
rect 1513 -37556 1559 -37456
rect 1709 -37556 1755 -37456
rect 1905 -37556 1951 -37456
rect -6573 -38944 -6527 -38744
rect -6377 -38944 -6331 -38744
rect -6181 -38944 -6135 -38744
rect 2122 -37757 2168 -37457
rect 2318 -37757 2364 -37457
rect 2514 -37757 2560 -37457
rect 2922 -37558 2968 -37458
rect 3118 -37558 3164 -37458
rect 3314 -37558 3360 -37458
rect 3510 -37558 3556 -37458
rect 3727 -37759 3773 -37459
rect 3923 -37759 3969 -37459
rect 4119 -37759 4165 -37459
rect 4546 -37634 4592 -37434
rect 4742 -37634 4788 -37434
rect 5284 -37634 5330 -37434
rect 5480 -37634 5526 -37434
rect 5676 -37634 5722 -37434
rect 5872 -37634 5918 -37434
rect 7033 -37645 7079 -37445
rect 7229 -37645 7275 -37445
rect 7425 -37645 7471 -37445
rect 7539 -37645 7585 -37445
rect 7735 -37645 7781 -37445
rect 7848 -37645 7894 -37445
rect 8044 -37645 8090 -37445
rect 6644 -37912 6783 -37903
rect 7722 -37910 7861 -37909
rect 9052 -37910 9103 -37902
rect 7722 -37912 9103 -37910
rect 6644 -37938 9103 -37912
rect 6644 -37940 7861 -37938
rect 6644 -37957 6783 -37940
rect 7722 -37963 7861 -37940
rect 9052 -37953 9103 -37938
rect -5736 -38944 -5690 -38744
rect -5540 -38944 -5494 -38744
rect -5344 -38944 -5298 -38744
rect -3873 -38944 -3827 -38744
rect -3677 -38944 -3631 -38744
rect -3481 -38944 -3435 -38744
rect -3036 -38944 -2990 -38744
rect -2840 -38944 -2794 -38744
rect -2644 -38944 -2598 -38744
rect -6573 -40382 -6527 -40182
rect -6377 -40382 -6331 -40182
rect -6181 -40382 -6135 -40182
rect -5736 -40382 -5690 -40182
rect -5540 -40382 -5494 -40182
rect -5344 -40382 -5298 -40182
rect -3873 -40382 -3827 -40182
rect -3677 -40382 -3631 -40182
rect -3481 -40382 -3435 -40182
rect -3036 -40382 -2990 -40182
rect -2840 -40382 -2794 -40182
rect -2644 -40382 -2598 -40182
rect -4177 -40974 -4040 -40914
rect -4128 -41422 -4068 -40974
rect -3202 -40915 -3142 -40551
rect -3231 -40975 -3099 -40915
rect -6475 -41700 -6429 -41500
rect -6279 -41700 -6233 -41500
rect -6083 -41700 -6037 -41500
rect -4732 -41700 -4686 -41500
rect -4536 -41700 -4490 -41500
rect -4340 -41700 -4294 -41500
rect -3775 -41700 -3729 -41500
rect -3579 -41700 -3533 -41500
rect -3383 -41700 -3337 -41500
rect -2032 -41700 -1986 -41500
rect -1836 -41700 -1790 -41500
rect -1640 -41700 -1594 -41500
rect -1150 -41700 -1104 -41500
rect -954 -41700 -908 -41500
rect -758 -41700 -712 -41500
rect -416 -41683 -370 -41483
rect -220 -41683 -174 -41483
rect 322 -41683 368 -41483
rect 518 -41683 564 -41483
rect 714 -41683 760 -41483
rect 910 -41683 956 -41483
rect 1317 -41670 1363 -41570
rect 1513 -41670 1559 -41570
rect 1709 -41670 1755 -41570
rect 1905 -41670 1951 -41570
rect 2122 -41669 2168 -41369
rect 2318 -41669 2364 -41369
rect 2514 -41669 2560 -41369
rect 2922 -41668 2968 -41568
rect 3118 -41668 3164 -41568
rect 3314 -41668 3360 -41568
rect 3510 -41668 3556 -41568
rect 3727 -41667 3773 -41367
rect 6644 -41186 6783 -41169
rect 7722 -41186 7861 -41163
rect 6644 -41188 7861 -41186
rect 8833 -41188 8978 -41093
rect 9065 -41188 9093 -37953
rect 6644 -41214 9095 -41188
rect 6644 -41223 6783 -41214
rect 7722 -41216 9095 -41214
rect 7722 -41217 7861 -41216
rect 8833 -41228 8978 -41216
rect 3923 -41667 3969 -41367
rect 4119 -41667 4165 -41367
rect 4546 -41692 4592 -41492
rect 4742 -41692 4788 -41492
rect 5284 -41692 5330 -41492
rect 5480 -41692 5526 -41492
rect 5676 -41692 5722 -41492
rect 5872 -41692 5918 -41492
rect 7033 -41681 7079 -41481
rect 7229 -41681 7275 -41481
rect 7425 -41681 7471 -41481
rect 7539 -41681 7585 -41481
rect 7735 -41681 7781 -41481
rect 7848 -41681 7894 -41481
rect 8044 -41681 8090 -41481
rect -824 -41750 -701 -41741
rect -530 -41750 -407 -41742
rect -824 -41865 -407 -41750
rect 2448 -41743 2571 -41729
rect 2837 -41743 2960 -41730
rect 2448 -41850 2960 -41743
rect 2448 -41865 2571 -41850
rect -824 -41877 -701 -41865
rect -530 -41878 -407 -41865
rect 2837 -41866 2960 -41850
rect 4065 -41773 4188 -41753
rect 4466 -41773 4589 -41755
rect 4065 -41880 4589 -41773
rect 4065 -41889 4188 -41880
rect 4466 -41891 4589 -41880
rect 5822 -41768 5945 -41750
rect 7038 -41768 7161 -41749
rect 5822 -41873 7161 -41768
rect 5822 -41886 5945 -41873
rect 7038 -41885 7161 -41873
rect 9247 -41981 9298 -37145
rect -665 -42032 9298 -41981
rect 9247 -42103 9298 -42032
rect 9127 -42210 9318 -42103
rect 9372 -42238 9423 -36888
rect -4785 -42289 9423 -42238
rect -6366 -43437 -6227 -43420
rect -5288 -43437 -5149 -43414
rect -6366 -43439 -5149 -43437
rect -4785 -43439 -4757 -42289
rect -6366 -43465 -4757 -43439
rect -6366 -43474 -6227 -43465
rect -5288 -43467 -4757 -43465
rect -5288 -43468 -5149 -43467
rect -4650 -42543 -4527 -42407
rect -4645 -43174 -4531 -42543
rect -4649 -43310 -4526 -43174
rect -2083 -42687 -1960 -42551
rect -2078 -43139 -1964 -42687
rect -2082 -43275 -1959 -43139
rect 400 -42721 706 -42659
rect 400 -42722 523 -42721
rect 405 -43139 519 -42722
rect 401 -43275 524 -43139
rect 8684 -42813 8823 -42798
rect 10042 -42813 10070 -36313
rect 6043 -42841 10070 -42813
rect 3634 -43437 3773 -43420
rect 4712 -43437 4851 -43414
rect 3634 -43439 4851 -43437
rect 6043 -43439 6071 -42841
rect 8684 -42845 8823 -42841
rect 3634 -43465 6071 -43439
rect 3634 -43474 3773 -43465
rect 4712 -43467 6071 -43465
rect 4712 -43468 4851 -43467
rect 6634 -43437 6773 -43420
rect 7712 -43437 7851 -43414
rect 6634 -43439 7851 -43437
rect 8649 -43439 8714 -43335
rect 10193 -43439 10221 -35687
rect 6634 -43465 10221 -43439
rect 6634 -43474 6773 -43465
rect 7610 -43467 10221 -43465
rect 7712 -43468 7851 -43467
rect 8649 -43472 8714 -43467
rect -5977 -43932 -5931 -43732
rect -5781 -43932 -5735 -43732
rect -5585 -43932 -5539 -43732
rect -5471 -43932 -5425 -43732
rect -5275 -43932 -5229 -43732
rect -5162 -43932 -5116 -43732
rect -4966 -43932 -4920 -43732
rect -3477 -43932 -3431 -43732
rect -3281 -43932 -3235 -43732
rect -3085 -43932 -3039 -43732
rect -2971 -43932 -2925 -43732
rect -2775 -43932 -2729 -43732
rect -2662 -43932 -2616 -43732
rect -2466 -43932 -2420 -43732
rect -977 -43932 -931 -43732
rect -781 -43932 -735 -43732
rect -585 -43932 -539 -43732
rect -471 -43932 -425 -43732
rect -275 -43932 -229 -43732
rect -162 -43932 -116 -43732
rect 34 -43932 80 -43732
rect 1523 -43932 1569 -43732
rect 1719 -43932 1765 -43732
rect 1915 -43932 1961 -43732
rect 2029 -43932 2075 -43732
rect 2225 -43932 2271 -43732
rect 2338 -43932 2384 -43732
rect 2534 -43932 2580 -43732
rect 4023 -43932 4069 -43732
rect 4219 -43932 4265 -43732
rect 4415 -43932 4461 -43732
rect 4529 -43932 4575 -43732
rect 4725 -43932 4771 -43732
rect 4838 -43932 4884 -43732
rect 5034 -43932 5080 -43732
rect 7023 -43932 7069 -43732
rect 7219 -43932 7265 -43732
rect 7415 -43932 7461 -43732
rect 7529 -43932 7575 -43732
rect 7725 -43932 7771 -43732
rect 7838 -43932 7884 -43732
rect 8034 -43932 8080 -43732
rect 10557 -43995 10852 -36705
rect -23503 -46536 -23290 -46358
rect 8644 -44709 8705 -44105
rect 8762 -44109 8806 -44106
rect 8591 -44832 8714 -44709
rect 8753 -44942 8813 -44109
rect 8697 -45065 8820 -44942
rect 8852 -45199 8913 -44252
rect 8790 -45322 8914 -45199
rect 9505 -44264 10852 -43995
rect 10557 -46526 10852 -44264
rect 15894 -36662 26127 -36622
rect 15894 -36956 26307 -36662
rect 15894 -36974 26272 -36956
rect 17738 -37818 17917 -37742
rect 17738 -37893 19408 -37818
rect 17738 -37931 17917 -37893
rect 19333 -37968 19408 -37893
rect 21278 -37895 21324 -37695
rect 21474 -37895 21520 -37695
rect 21670 -37895 21716 -37695
rect 22115 -37895 22161 -37695
rect 22311 -37895 22357 -37695
rect 22507 -37895 22553 -37695
rect 23978 -37895 24024 -37695
rect 24174 -37895 24220 -37695
rect 24370 -37895 24416 -37695
rect 19306 -38103 19438 -37968
rect 24815 -37895 24861 -37695
rect 25011 -37895 25057 -37695
rect 25207 -37895 25253 -37695
rect 18071 -39093 18117 -38493
rect 18267 -39093 18313 -38493
rect 21822 -38428 21882 -38064
rect 21779 -38488 21911 -38428
rect 22720 -38487 22857 -38427
rect 22748 -38935 22808 -38487
rect 19392 -39213 19438 -39013
rect 19588 -39213 19634 -39013
rect 19784 -39213 19830 -39013
rect 20274 -39213 20320 -39013
rect 20470 -39213 20516 -39013
rect 20666 -39213 20712 -39013
rect 22017 -39213 22063 -39013
rect 22213 -39213 22259 -39013
rect 22409 -39213 22455 -39013
rect 22974 -39213 23020 -39013
rect 23170 -39213 23216 -39013
rect 23366 -39213 23412 -39013
rect 24717 -39213 24763 -39013
rect 24913 -39213 24959 -39013
rect 25109 -39213 25155 -39013
rect 18066 -41439 18112 -41039
rect 18262 -41439 18308 -41039
rect 19012 -41439 19058 -41039
rect 19208 -41439 19254 -41039
rect 21837 -40165 21883 -39765
rect 22033 -40165 22079 -39765
rect 22229 -40165 22275 -39765
rect 19928 -41473 19974 -41273
rect 20124 -41473 20170 -41273
rect 20320 -41473 20366 -41273
rect 20516 -41473 20562 -41273
rect 21058 -41473 21104 -41273
rect 21254 -41473 21300 -41273
rect 21787 -41466 21833 -41266
rect 21983 -41466 22029 -41266
rect 22179 -41466 22225 -41266
rect 22667 -41395 22713 -40695
rect 22863 -41395 22909 -40695
rect 23067 -41395 23113 -40695
rect 23263 -41395 23309 -40695
rect 23667 -41395 23713 -40695
rect 23863 -41395 23909 -40695
rect 24067 -41395 24113 -40695
rect 24263 -41395 24309 -40695
rect 24667 -41395 24713 -40695
rect 24863 -41395 24909 -40695
rect 25067 -41395 25113 -40695
rect 25263 -41395 25309 -40695
rect 11264 -42451 11310 -42251
rect 11460 -42451 11506 -42251
rect 11656 -42451 11702 -42251
rect 12146 -42451 12192 -42251
rect 12342 -42451 12388 -42251
rect 12538 -42451 12584 -42251
rect 13889 -42451 13935 -42251
rect 14085 -42451 14131 -42251
rect 14281 -42451 14327 -42251
rect 14846 -42451 14892 -42251
rect 15042 -42451 15088 -42251
rect 15238 -42451 15284 -42251
rect 16589 -42451 16635 -42251
rect 16785 -42451 16831 -42251
rect 16981 -42451 17027 -42251
rect 13651 -43036 13783 -42976
rect 13694 -43400 13754 -43036
rect 14620 -42977 14680 -42529
rect 14592 -43037 14729 -42977
rect 13150 -43769 13196 -43569
rect 13346 -43769 13392 -43569
rect 13542 -43769 13588 -43569
rect 13987 -43769 14033 -43569
rect 14183 -43769 14229 -43569
rect 14379 -43769 14425 -43569
rect 15850 -43769 15896 -43569
rect 16046 -43769 16092 -43569
rect 16242 -43769 16288 -43569
rect 16687 -43769 16733 -43569
rect 16883 -43769 16929 -43569
rect 17079 -43769 17125 -43569
rect 26027 -44073 26272 -36974
rect 26895 -36814 27108 -36775
rect 26895 -36868 28333 -36814
rect 26895 -36908 27108 -36868
rect 28279 -37158 28333 -36868
rect 28279 -37212 28607 -37158
rect 28553 -37267 28607 -37212
rect 26896 -38735 27155 -38472
rect 27650 -37542 27696 -37342
rect 27846 -37542 27892 -37342
rect 28042 -37542 28088 -37342
rect 28527 -37325 28686 -37267
rect 28238 -37542 28284 -37342
rect 28623 -37671 28669 -37371
rect 28819 -37671 28865 -37371
rect 29015 -37671 29061 -37371
rect 29232 -37672 29278 -37572
rect 29428 -37672 29474 -37572
rect 29624 -37672 29670 -37572
rect 29820 -37672 29866 -37572
rect 29902 -37987 29976 -37971
rect 30130 -37987 30240 -37951
rect 29902 -38083 30240 -37987
rect 29902 -38089 29976 -38083
rect 30130 -38101 30240 -38083
rect 27624 -38571 27670 -38271
rect 27820 -38571 27866 -38271
rect 28016 -38571 28062 -38271
rect 28233 -38370 28279 -38270
rect 28429 -38370 28475 -38270
rect 28625 -38370 28671 -38270
rect 28821 -38370 28867 -38270
rect 29071 -38782 29117 -38182
rect 29267 -38782 29313 -38182
rect 29690 -38782 29736 -38182
rect 31063 -38540 31109 -38040
rect 31259 -38540 31305 -38040
rect 31854 -38540 31900 -38040
rect 31984 -38540 32030 -38040
rect 32212 -38340 32258 -38040
rect 32408 -38340 32454 -38040
rect 27642 -40995 27688 -40795
rect 27838 -40995 27884 -40795
rect 28034 -40995 28080 -40795
rect 28230 -40995 28276 -40795
rect 28615 -41124 28661 -40824
rect 28811 -41124 28857 -40824
rect 29007 -41124 29053 -40824
rect 29224 -41125 29270 -41025
rect 29420 -41125 29466 -41025
rect 29616 -41125 29662 -41025
rect 29812 -41125 29858 -41025
rect 28817 -41399 29000 -41358
rect 30120 -41399 30216 -41370
rect 28817 -41481 30216 -41399
rect 28817 -41488 29000 -41481
rect 30120 -41507 30216 -41481
rect 27616 -42024 27662 -41724
rect 27812 -42024 27858 -41724
rect 28008 -42024 28054 -41724
rect 28225 -41823 28271 -41723
rect 28421 -41823 28467 -41723
rect 28617 -41823 28663 -41723
rect 28813 -41823 28859 -41723
rect 29063 -42235 29109 -41635
rect 29259 -42235 29305 -41635
rect 29682 -42235 29728 -41635
rect 31310 -41026 31356 -40826
rect 31506 -41026 31552 -40826
rect 31702 -41026 31748 -40826
rect 31898 -41026 31944 -40826
rect 32283 -41155 32329 -40855
rect 32479 -41155 32525 -40855
rect 32675 -41155 32721 -40855
rect 32892 -41156 32938 -41056
rect 33088 -41156 33134 -41056
rect 33284 -41156 33330 -41056
rect 33480 -41156 33526 -41056
rect 33540 -41421 33631 -41409
rect 33790 -41421 33941 -41394
rect 33540 -41560 33941 -41421
rect 33540 -41572 33631 -41560
rect 33790 -41585 33941 -41560
rect 31284 -42055 31330 -41755
rect 31480 -42055 31526 -41755
rect 31676 -42055 31722 -41755
rect 31893 -41854 31939 -41754
rect 32089 -41854 32135 -41754
rect 32285 -41854 32331 -41754
rect 32481 -41854 32527 -41754
rect 32731 -42266 32777 -41666
rect 32927 -42266 32973 -41666
rect 33350 -42266 33396 -41666
rect 36090 -37553 36136 -37353
rect 36286 -37553 36332 -37353
rect 36482 -37553 36528 -37353
rect 36678 -37553 36724 -37353
rect 37063 -37682 37109 -37382
rect 37259 -37682 37305 -37382
rect 37455 -37682 37501 -37382
rect 37672 -37683 37718 -37583
rect 37868 -37683 37914 -37583
rect 38064 -37683 38110 -37583
rect 38260 -37683 38306 -37583
rect 38342 -37998 38416 -37982
rect 38570 -37998 38680 -37962
rect 38342 -38094 38680 -37998
rect 38342 -38100 38416 -38094
rect 38570 -38112 38680 -38094
rect 36064 -38582 36110 -38282
rect 36260 -38582 36306 -38282
rect 36456 -38582 36502 -38282
rect 36673 -38381 36719 -38281
rect 36869 -38381 36915 -38281
rect 37065 -38381 37111 -38281
rect 37261 -38381 37307 -38281
rect 37511 -38793 37557 -38193
rect 37707 -38793 37753 -38193
rect 38130 -38793 38176 -38193
rect 39503 -38551 39549 -38051
rect 39699 -38551 39745 -38051
rect 40294 -38551 40340 -38051
rect 40424 -38551 40470 -38051
rect 40652 -38351 40698 -38051
rect 40848 -38351 40894 -38051
rect 36082 -41006 36128 -40806
rect 36278 -41006 36324 -40806
rect 36474 -41006 36520 -40806
rect 36670 -41006 36716 -40806
rect 37055 -41135 37101 -40835
rect 37251 -41135 37297 -40835
rect 37447 -41135 37493 -40835
rect 37664 -41136 37710 -41036
rect 37860 -41136 37906 -41036
rect 38056 -41136 38102 -41036
rect 38252 -41136 38298 -41036
rect 37257 -41410 37440 -41369
rect 38560 -41410 38656 -41381
rect 37257 -41492 38656 -41410
rect 37257 -41499 37440 -41492
rect 38560 -41518 38656 -41492
rect 36056 -42035 36102 -41735
rect 36252 -42035 36298 -41735
rect 36448 -42035 36494 -41735
rect 36665 -41834 36711 -41734
rect 36861 -41834 36907 -41734
rect 37057 -41834 37103 -41734
rect 37253 -41834 37299 -41734
rect 37503 -42246 37549 -41646
rect 37699 -42246 37745 -41646
rect 38122 -42246 38168 -41646
rect 39750 -41037 39796 -40837
rect 39946 -41037 39992 -40837
rect 40142 -41037 40188 -40837
rect 40338 -41037 40384 -40837
rect 40723 -41166 40769 -40866
rect 40919 -41166 40965 -40866
rect 41115 -41166 41161 -40866
rect 41332 -41167 41378 -41067
rect 41528 -41167 41574 -41067
rect 41724 -41167 41770 -41067
rect 41920 -41167 41966 -41067
rect 41980 -41432 42071 -41420
rect 42230 -41432 42381 -41405
rect 41980 -41571 42381 -41432
rect 41980 -41583 42071 -41571
rect 42230 -41596 42381 -41571
rect 39724 -42066 39770 -41766
rect 39920 -42066 39966 -41766
rect 40116 -42066 40162 -41766
rect 40333 -41865 40379 -41765
rect 40529 -41865 40575 -41765
rect 40725 -41865 40771 -41765
rect 40921 -41865 40967 -41765
rect 41171 -42277 41217 -41677
rect 41367 -42277 41413 -41677
rect 41790 -42277 41836 -41677
rect 44953 -37592 44999 -37392
rect 45149 -37592 45195 -37392
rect 45345 -37592 45391 -37392
rect 45541 -37592 45587 -37392
rect 45926 -37721 45972 -37421
rect 46122 -37721 46168 -37421
rect 46318 -37721 46364 -37421
rect 46535 -37722 46581 -37622
rect 46731 -37722 46777 -37622
rect 46927 -37722 46973 -37622
rect 47123 -37722 47169 -37622
rect 47205 -38037 47279 -38021
rect 47433 -38037 47543 -38001
rect 47205 -38133 47543 -38037
rect 47205 -38139 47279 -38133
rect 47433 -38151 47543 -38133
rect 44927 -38621 44973 -38321
rect 45123 -38621 45169 -38321
rect 45319 -38621 45365 -38321
rect 45536 -38420 45582 -38320
rect 45732 -38420 45778 -38320
rect 45928 -38420 45974 -38320
rect 46124 -38420 46170 -38320
rect 46374 -38832 46420 -38232
rect 46570 -38832 46616 -38232
rect 46993 -38832 47039 -38232
rect 48366 -38590 48412 -38090
rect 48562 -38590 48608 -38090
rect 49157 -38590 49203 -38090
rect 49287 -38590 49333 -38090
rect 49515 -38390 49561 -38090
rect 49711 -38390 49757 -38090
rect 44945 -41045 44991 -40845
rect 45141 -41045 45187 -40845
rect 45337 -41045 45383 -40845
rect 45533 -41045 45579 -40845
rect 45918 -41174 45964 -40874
rect 46114 -41174 46160 -40874
rect 46310 -41174 46356 -40874
rect 46527 -41175 46573 -41075
rect 46723 -41175 46769 -41075
rect 46919 -41175 46965 -41075
rect 47115 -41175 47161 -41075
rect 46120 -41449 46303 -41408
rect 47423 -41449 47519 -41420
rect 46120 -41531 47519 -41449
rect 46120 -41538 46303 -41531
rect 47423 -41557 47519 -41531
rect 44919 -42074 44965 -41774
rect 45115 -42074 45161 -41774
rect 45311 -42074 45357 -41774
rect 45528 -41873 45574 -41773
rect 45724 -41873 45770 -41773
rect 45920 -41873 45966 -41773
rect 46116 -41873 46162 -41773
rect 46366 -42285 46412 -41685
rect 46562 -42285 46608 -41685
rect 46985 -42285 47031 -41685
rect 48613 -41076 48659 -40876
rect 48809 -41076 48855 -40876
rect 49005 -41076 49051 -40876
rect 49201 -41076 49247 -40876
rect 49586 -41205 49632 -40905
rect 49782 -41205 49828 -40905
rect 49978 -41205 50024 -40905
rect 50195 -41206 50241 -41106
rect 50391 -41206 50437 -41106
rect 50587 -41206 50633 -41106
rect 50783 -41206 50829 -41106
rect 50843 -41471 50934 -41459
rect 51093 -41471 51244 -41444
rect 50843 -41610 51244 -41471
rect 50843 -41622 50934 -41610
rect 51093 -41635 51244 -41610
rect 48587 -42105 48633 -41805
rect 48783 -42105 48829 -41805
rect 48979 -42105 49025 -41805
rect 49196 -41904 49242 -41804
rect 49392 -41904 49438 -41804
rect 49588 -41904 49634 -41804
rect 49784 -41904 49830 -41804
rect 50034 -42316 50080 -41716
rect 50230 -42316 50276 -41716
rect 50653 -42316 50699 -41716
rect 54151 -37558 54197 -37358
rect 54347 -37558 54393 -37358
rect 54543 -37558 54589 -37358
rect 54739 -37558 54785 -37358
rect 55124 -37687 55170 -37387
rect 55320 -37687 55366 -37387
rect 55516 -37687 55562 -37387
rect 55733 -37688 55779 -37588
rect 55929 -37688 55975 -37588
rect 56125 -37688 56171 -37588
rect 56321 -37688 56367 -37588
rect 56403 -38003 56477 -37987
rect 56631 -38003 56741 -37967
rect 56403 -38099 56741 -38003
rect 56403 -38105 56477 -38099
rect 56631 -38117 56741 -38099
rect 54125 -38587 54171 -38287
rect 54321 -38587 54367 -38287
rect 54517 -38587 54563 -38287
rect 54734 -38386 54780 -38286
rect 54930 -38386 54976 -38286
rect 55126 -38386 55172 -38286
rect 55322 -38386 55368 -38286
rect 55572 -38798 55618 -38198
rect 55768 -38798 55814 -38198
rect 56191 -38798 56237 -38198
rect 57564 -38556 57610 -38056
rect 57760 -38556 57806 -38056
rect 58355 -38556 58401 -38056
rect 58485 -38556 58531 -38056
rect 58713 -38356 58759 -38056
rect 58909 -38356 58955 -38056
rect 54143 -41011 54189 -40811
rect 54339 -41011 54385 -40811
rect 54535 -41011 54581 -40811
rect 54731 -41011 54777 -40811
rect 55116 -41140 55162 -40840
rect 55312 -41140 55358 -40840
rect 55508 -41140 55554 -40840
rect 55725 -41141 55771 -41041
rect 55921 -41141 55967 -41041
rect 56117 -41141 56163 -41041
rect 56313 -41141 56359 -41041
rect 55318 -41415 55501 -41374
rect 56621 -41415 56717 -41386
rect 55318 -41497 56717 -41415
rect 55318 -41504 55501 -41497
rect 56621 -41523 56717 -41497
rect 54117 -42040 54163 -41740
rect 54313 -42040 54359 -41740
rect 54509 -42040 54555 -41740
rect 54726 -41839 54772 -41739
rect 54922 -41839 54968 -41739
rect 55118 -41839 55164 -41739
rect 55314 -41839 55360 -41739
rect 55564 -42251 55610 -41651
rect 55760 -42251 55806 -41651
rect 56183 -42251 56229 -41651
rect 57811 -41042 57857 -40842
rect 58007 -41042 58053 -40842
rect 58203 -41042 58249 -40842
rect 58399 -41042 58445 -40842
rect 58784 -41171 58830 -40871
rect 58980 -41171 59026 -40871
rect 59176 -41171 59222 -40871
rect 59393 -41172 59439 -41072
rect 59589 -41172 59635 -41072
rect 59785 -41172 59831 -41072
rect 59981 -41172 60027 -41072
rect 60041 -41437 60132 -41425
rect 60291 -41437 60442 -41410
rect 60041 -41576 60442 -41437
rect 60041 -41588 60132 -41576
rect 60291 -41601 60442 -41576
rect 57785 -42071 57831 -41771
rect 57981 -42071 58027 -41771
rect 58177 -42071 58223 -41771
rect 58394 -41870 58440 -41770
rect 58590 -41870 58636 -41770
rect 58786 -41870 58832 -41770
rect 58982 -41870 59028 -41770
rect 59232 -42282 59278 -41682
rect 59428 -42282 59474 -41682
rect 59851 -42282 59897 -41682
rect 62905 -37492 62951 -37292
rect 63101 -37492 63147 -37292
rect 63297 -37492 63343 -37292
rect 63493 -37492 63539 -37292
rect 63878 -37621 63924 -37321
rect 64074 -37621 64120 -37321
rect 64270 -37621 64316 -37321
rect 64487 -37622 64533 -37522
rect 64683 -37622 64729 -37522
rect 64879 -37622 64925 -37522
rect 65075 -37622 65121 -37522
rect 65157 -37937 65231 -37921
rect 65385 -37937 65495 -37901
rect 65157 -38033 65495 -37937
rect 65157 -38039 65231 -38033
rect 65385 -38051 65495 -38033
rect 62879 -38521 62925 -38221
rect 63075 -38521 63121 -38221
rect 63271 -38521 63317 -38221
rect 63488 -38320 63534 -38220
rect 63684 -38320 63730 -38220
rect 63880 -38320 63926 -38220
rect 64076 -38320 64122 -38220
rect 64326 -38732 64372 -38132
rect 64522 -38732 64568 -38132
rect 64945 -38732 64991 -38132
rect 66318 -38490 66364 -37990
rect 66514 -38490 66560 -37990
rect 67109 -38490 67155 -37990
rect 67239 -38490 67285 -37990
rect 67467 -38290 67513 -37990
rect 67663 -38290 67709 -37990
rect 62897 -40945 62943 -40745
rect 63093 -40945 63139 -40745
rect 63289 -40945 63335 -40745
rect 63485 -40945 63531 -40745
rect 63870 -41074 63916 -40774
rect 64066 -41074 64112 -40774
rect 64262 -41074 64308 -40774
rect 64479 -41075 64525 -40975
rect 64675 -41075 64721 -40975
rect 64871 -41075 64917 -40975
rect 65067 -41075 65113 -40975
rect 64072 -41349 64255 -41308
rect 65375 -41349 65471 -41320
rect 64072 -41431 65471 -41349
rect 64072 -41438 64255 -41431
rect 65375 -41457 65471 -41431
rect 62871 -41974 62917 -41674
rect 63067 -41974 63113 -41674
rect 63263 -41974 63309 -41674
rect 63480 -41773 63526 -41673
rect 63676 -41773 63722 -41673
rect 63872 -41773 63918 -41673
rect 64068 -41773 64114 -41673
rect 64318 -42185 64364 -41585
rect 64514 -42185 64560 -41585
rect 64937 -42185 64983 -41585
rect 66565 -40976 66611 -40776
rect 66761 -40976 66807 -40776
rect 66957 -40976 67003 -40776
rect 67153 -40976 67199 -40776
rect 67538 -41105 67584 -40805
rect 67734 -41105 67780 -40805
rect 67930 -41105 67976 -40805
rect 68147 -41106 68193 -41006
rect 68343 -41106 68389 -41006
rect 68539 -41106 68585 -41006
rect 68735 -41106 68781 -41006
rect 68795 -41371 68886 -41359
rect 69045 -41371 69196 -41344
rect 68795 -41510 69196 -41371
rect 68795 -41522 68886 -41510
rect 69045 -41535 69196 -41510
rect 66539 -42005 66585 -41705
rect 66735 -42005 66781 -41705
rect 66931 -42005 66977 -41705
rect 67148 -41804 67194 -41704
rect 67344 -41804 67390 -41704
rect 67540 -41804 67586 -41704
rect 67736 -41804 67782 -41704
rect 67986 -42216 68032 -41616
rect 68182 -42216 68228 -41616
rect 68605 -42216 68651 -41616
rect 72058 -37475 72104 -37275
rect 72254 -37475 72300 -37275
rect 72450 -37475 72496 -37275
rect 72646 -37475 72692 -37275
rect 73031 -37604 73077 -37304
rect 73227 -37604 73273 -37304
rect 73423 -37604 73469 -37304
rect 73640 -37605 73686 -37505
rect 73836 -37605 73882 -37505
rect 74032 -37605 74078 -37505
rect 74228 -37605 74274 -37505
rect 74310 -37920 74384 -37904
rect 74538 -37920 74648 -37884
rect 74310 -38016 74648 -37920
rect 74310 -38022 74384 -38016
rect 74538 -38034 74648 -38016
rect 72032 -38504 72078 -38204
rect 72228 -38504 72274 -38204
rect 72424 -38504 72470 -38204
rect 72641 -38303 72687 -38203
rect 72837 -38303 72883 -38203
rect 73033 -38303 73079 -38203
rect 73229 -38303 73275 -38203
rect 73479 -38715 73525 -38115
rect 73675 -38715 73721 -38115
rect 74098 -38715 74144 -38115
rect 75471 -38473 75517 -37973
rect 75667 -38473 75713 -37973
rect 76262 -38473 76308 -37973
rect 76392 -38473 76438 -37973
rect 76620 -38273 76666 -37973
rect 76816 -38273 76862 -37973
rect 72050 -40928 72096 -40728
rect 72246 -40928 72292 -40728
rect 72442 -40928 72488 -40728
rect 72638 -40928 72684 -40728
rect 73023 -41057 73069 -40757
rect 73219 -41057 73265 -40757
rect 73415 -41057 73461 -40757
rect 73632 -41058 73678 -40958
rect 73828 -41058 73874 -40958
rect 74024 -41058 74070 -40958
rect 74220 -41058 74266 -40958
rect 73225 -41332 73408 -41291
rect 74528 -41332 74624 -41303
rect 73225 -41414 74624 -41332
rect 73225 -41421 73408 -41414
rect 74528 -41440 74624 -41414
rect 72024 -41957 72070 -41657
rect 72220 -41957 72266 -41657
rect 72416 -41957 72462 -41657
rect 72633 -41756 72679 -41656
rect 72829 -41756 72875 -41656
rect 73025 -41756 73071 -41656
rect 73221 -41756 73267 -41656
rect 73471 -42168 73517 -41568
rect 73667 -42168 73713 -41568
rect 74090 -42168 74136 -41568
rect 75718 -40959 75764 -40759
rect 75914 -40959 75960 -40759
rect 76110 -40959 76156 -40759
rect 76306 -40959 76352 -40759
rect 76691 -41088 76737 -40788
rect 76887 -41088 76933 -40788
rect 77083 -41088 77129 -40788
rect 77300 -41089 77346 -40989
rect 77496 -41089 77542 -40989
rect 77692 -41089 77738 -40989
rect 77888 -41089 77934 -40989
rect 77948 -41354 78039 -41342
rect 78198 -41354 78349 -41327
rect 77948 -41493 78349 -41354
rect 77948 -41505 78039 -41493
rect 78198 -41518 78349 -41493
rect 75692 -41988 75738 -41688
rect 75888 -41988 75934 -41688
rect 76084 -41988 76130 -41688
rect 76301 -41787 76347 -41687
rect 76497 -41787 76543 -41687
rect 76693 -41787 76739 -41687
rect 76889 -41787 76935 -41687
rect 77139 -42199 77185 -41599
rect 77335 -42199 77381 -41599
rect 77758 -42199 77804 -41599
rect 81422 -37437 81468 -37237
rect 81618 -37437 81664 -37237
rect 81814 -37437 81860 -37237
rect 82010 -37437 82056 -37237
rect 82395 -37566 82441 -37266
rect 82591 -37566 82637 -37266
rect 82787 -37566 82833 -37266
rect 83004 -37567 83050 -37467
rect 83200 -37567 83246 -37467
rect 83396 -37567 83442 -37467
rect 83592 -37567 83638 -37467
rect 83674 -37882 83748 -37866
rect 83902 -37882 84012 -37846
rect 83674 -37978 84012 -37882
rect 83674 -37984 83748 -37978
rect 83902 -37996 84012 -37978
rect 81396 -38466 81442 -38166
rect 81592 -38466 81638 -38166
rect 81788 -38466 81834 -38166
rect 82005 -38265 82051 -38165
rect 82201 -38265 82247 -38165
rect 82397 -38265 82443 -38165
rect 82593 -38265 82639 -38165
rect 82843 -38677 82889 -38077
rect 83039 -38677 83085 -38077
rect 83462 -38677 83508 -38077
rect 84835 -38435 84881 -37935
rect 85031 -38435 85077 -37935
rect 85626 -38435 85672 -37935
rect 85756 -38435 85802 -37935
rect 85984 -38235 86030 -37935
rect 86180 -38235 86226 -37935
rect 81414 -40890 81460 -40690
rect 81610 -40890 81656 -40690
rect 81806 -40890 81852 -40690
rect 82002 -40890 82048 -40690
rect 82387 -41019 82433 -40719
rect 82583 -41019 82629 -40719
rect 82779 -41019 82825 -40719
rect 82996 -41020 83042 -40920
rect 83192 -41020 83238 -40920
rect 83388 -41020 83434 -40920
rect 83584 -41020 83630 -40920
rect 82589 -41294 82772 -41253
rect 83892 -41294 83988 -41265
rect 82589 -41376 83988 -41294
rect 82589 -41383 82772 -41376
rect 83892 -41402 83988 -41376
rect 81388 -41919 81434 -41619
rect 81584 -41919 81630 -41619
rect 81780 -41919 81826 -41619
rect 81997 -41718 82043 -41618
rect 82193 -41718 82239 -41618
rect 82389 -41718 82435 -41618
rect 82585 -41718 82631 -41618
rect 82835 -42130 82881 -41530
rect 83031 -42130 83077 -41530
rect 83454 -42130 83500 -41530
rect 85082 -40921 85128 -40721
rect 85278 -40921 85324 -40721
rect 85474 -40921 85520 -40721
rect 85670 -40921 85716 -40721
rect 86055 -41050 86101 -40750
rect 86251 -41050 86297 -40750
rect 86447 -41050 86493 -40750
rect 86664 -41051 86710 -40951
rect 86860 -41051 86906 -40951
rect 87056 -41051 87102 -40951
rect 87252 -41051 87298 -40951
rect 87312 -41316 87403 -41304
rect 87562 -41316 87713 -41289
rect 87312 -41455 87713 -41316
rect 87312 -41467 87403 -41455
rect 87562 -41480 87713 -41455
rect 85056 -41950 85102 -41650
rect 85252 -41950 85298 -41650
rect 85448 -41950 85494 -41650
rect 85665 -41749 85711 -41649
rect 85861 -41749 85907 -41649
rect 86057 -41749 86103 -41649
rect 86253 -41749 86299 -41649
rect 86503 -42161 86549 -41561
rect 86699 -42161 86745 -41561
rect 87122 -42161 87168 -41561
rect 26027 -44318 82025 -44073
rect -27977 -52158 -27903 -52129
rect -27977 -52204 -27432 -52158
rect -27977 -52394 -27903 -52204
rect -27832 -52322 -27432 -52276
rect -27977 -52440 -27432 -52394
rect -27977 -52630 -27903 -52440
rect -27832 -52558 -27432 -52512
rect -27977 -52676 -27432 -52630
rect -27977 -52866 -27903 -52676
rect -27832 -52794 -27432 -52748
rect -27977 -52912 -27432 -52866
rect -27977 -53102 -27903 -52912
rect -27832 -53030 -27432 -52984
rect -27977 -53148 -27432 -53102
rect -27977 -53338 -27903 -53148
rect -27832 -53266 -27432 -53220
rect -27977 -53384 -27432 -53338
rect -27977 -53574 -27903 -53384
rect -27832 -53502 -27432 -53456
rect -27977 -53620 -27432 -53574
rect -27977 -53810 -27903 -53620
rect -27832 -53738 -27432 -53692
rect -27977 -53856 -27432 -53810
rect -27977 -54046 -27903 -53856
rect -27832 -53974 -27432 -53928
rect -27977 -54092 -27432 -54046
rect -27977 -54282 -27903 -54092
rect -27832 -54210 -27432 -54164
rect -27977 -54328 -27432 -54282
rect -27977 -54518 -27903 -54328
rect -27832 -54446 -27432 -54400
rect -27977 -54564 -27432 -54518
rect -27977 -54754 -27903 -54564
rect -27832 -54682 -27432 -54636
rect -27977 -54800 -27432 -54754
rect -27977 -54990 -27903 -54800
rect -27832 -54918 -27432 -54872
rect -27977 -55036 -27432 -54990
rect -27977 -55226 -27903 -55036
rect -27832 -55154 -27432 -55108
rect -27977 -55272 -27432 -55226
rect -27977 -55462 -27903 -55272
rect -22631 -55313 -22530 -55258
rect -27832 -55390 -27432 -55344
rect -27977 -55508 -27432 -55462
rect -22783 -55501 -22530 -55313
rect -27977 -55698 -27903 -55508
rect -22783 -55544 -22543 -55501
rect -27832 -55626 -27432 -55580
rect -27977 -55744 -27432 -55698
rect -27977 -55914 -27903 -55744
rect -27832 -55862 -27432 -55816
rect -28640 -55934 -27903 -55914
rect -28640 -55960 -27432 -55934
rect -28139 -56150 -28093 -55960
rect -27977 -55980 -27432 -55960
rect -27977 -56006 -27903 -55980
rect -28640 -56196 -28093 -56150
rect -28139 -56386 -28093 -56196
rect -28640 -56432 -28093 -56386
rect -28139 -56622 -28093 -56432
rect -28640 -56668 -28093 -56622
rect -28139 -56858 -28093 -56668
rect -28640 -56904 -28093 -56858
rect -28139 -57094 -28093 -56904
rect -28640 -57140 -28093 -57094
rect -28139 -57330 -28093 -57140
rect -28640 -57376 -28093 -57330
rect -28139 -57566 -28093 -57376
rect -28640 -57612 -28093 -57566
rect -27832 -56110 -27432 -56064
rect -27832 -56346 -27432 -56300
rect -27832 -56582 -27432 -56536
rect -27832 -56818 -27432 -56772
rect -27832 -57054 -27432 -57008
rect -27832 -57290 -27432 -57244
rect -27832 -57526 -27432 -57480
rect -27832 -57762 -27432 -57716
rect -27832 -57998 -27432 -57952
rect -27832 -58128 -27432 -58082
rect -27832 -58364 -27432 -58318
rect -27832 -58600 -27432 -58554
rect -27832 -58836 -27432 -58790
rect -27832 -59072 -27432 -59026
rect -27832 -59202 -27432 -59156
rect -27832 -59438 -27432 -59392
rect -27832 -59674 -27432 -59628
rect -31679 -63836 -30520 -62597
rect -31679 -64865 -30522 -63836
rect -22783 -64469 -22647 -55544
rect -22483 -62626 -22422 -54099
rect -22536 -62749 -22413 -62626
rect -22292 -62825 -22231 -54020
rect -22183 -54172 -22122 -53934
rect -21343 -54086 -21297 -53886
rect -21147 -54086 -21101 -53886
rect -20951 -54086 -20905 -53886
rect -20755 -54086 -20709 -53886
rect -20213 -54086 -20167 -53886
rect -20017 -54086 -19971 -53886
rect -13744 -53299 -13698 -53099
rect -13548 -53299 -13502 -53099
rect -13352 -53299 -13306 -53099
rect -12907 -53299 -12861 -53099
rect -12711 -53299 -12665 -53099
rect -12515 -53299 -12469 -53099
rect -11044 -53299 -10998 -53099
rect -10848 -53299 -10802 -53099
rect -10652 -53299 -10606 -53099
rect -10207 -53299 -10161 -53099
rect -10011 -53299 -9965 -53099
rect -9815 -53299 -9769 -53099
rect -22183 -60001 -22123 -54172
rect -19344 -54308 -19298 -54008
rect -19148 -54308 -19102 -54008
rect -22183 -60238 -22122 -60001
rect -22345 -62948 -22222 -62825
rect -22183 -63058 -22123 -60238
rect -22239 -63181 -22116 -63058
rect -22084 -63315 -22023 -55099
rect -22146 -63438 -22022 -63315
rect -21286 -56217 -21240 -55917
rect -21090 -56217 -21044 -55917
rect -20894 -56217 -20848 -55917
rect -20677 -56016 -20631 -55916
rect -20481 -56016 -20435 -55916
rect -20285 -56016 -20239 -55916
rect -20089 -56016 -20043 -55916
rect -19558 -54511 -19421 -54453
rect -19551 -55284 -19511 -54511
rect -18952 -54308 -18906 -54008
rect -18735 -54107 -18689 -54007
rect -18539 -54107 -18493 -54007
rect -18343 -54107 -18297 -54007
rect -18147 -54107 -18101 -54007
rect -19667 -55293 -19511 -55284
rect -19714 -55333 -19511 -55293
rect -19667 -55337 -19535 -55333
rect -19513 -56022 -19467 -55822
rect -19317 -56022 -19271 -55822
rect -19121 -56022 -19075 -55822
rect -18925 -56022 -18879 -55822
rect -18383 -56022 -18337 -55822
rect -18187 -56022 -18141 -55822
rect -17708 -55270 -17662 -54970
rect -17512 -55270 -17466 -54970
rect -17316 -55270 -17270 -54970
rect -17099 -55271 -17053 -55171
rect -16903 -55271 -16857 -55171
rect -16707 -55271 -16661 -55171
rect -16511 -55271 -16465 -55171
rect -16261 -55359 -16215 -54759
rect -16065 -55359 -16019 -54759
rect -15642 -55359 -15596 -54759
rect -17682 -56199 -17636 -55999
rect -17486 -56199 -17440 -55999
rect -17290 -56199 -17244 -55999
rect -17094 -56199 -17048 -55999
rect -16709 -56170 -16663 -55870
rect -16513 -56170 -16467 -55870
rect -16317 -56170 -16271 -55870
rect -16100 -55969 -16054 -55869
rect -15904 -55969 -15858 -55869
rect -15708 -55969 -15662 -55869
rect -15512 -55969 -15466 -55869
rect -7382 -53709 -7336 -53109
rect -6959 -53709 -6913 -53109
rect -6763 -53709 -6717 -53109
rect -5274 -53505 -5228 -53305
rect -5078 -53505 -5032 -53305
rect -4882 -53505 -4836 -53305
rect -4768 -53505 -4722 -53305
rect -4572 -53505 -4526 -53305
rect -4459 -53505 -4413 -53305
rect -4263 -53505 -4217 -53305
rect -2774 -53505 -2728 -53305
rect -2578 -53505 -2532 -53305
rect -2382 -53505 -2336 -53305
rect -2268 -53505 -2222 -53305
rect -2072 -53505 -2026 -53305
rect -1959 -53505 -1913 -53305
rect -1763 -53505 -1717 -53305
rect -274 -53505 -228 -53305
rect -78 -53505 -32 -53305
rect 118 -53505 164 -53305
rect 232 -53505 278 -53305
rect 428 -53505 474 -53305
rect 541 -53505 587 -53305
rect 737 -53505 783 -53305
rect 2226 -53505 2272 -53305
rect 2422 -53505 2468 -53305
rect 2618 -53505 2664 -53305
rect 2732 -53505 2778 -53305
rect 2928 -53505 2974 -53305
rect 3041 -53505 3087 -53305
rect 3237 -53505 3283 -53305
rect 4726 -53505 4772 -53305
rect 4922 -53505 4968 -53305
rect 5118 -53505 5164 -53305
rect 5232 -53505 5278 -53305
rect 5428 -53505 5474 -53305
rect 5541 -53505 5587 -53305
rect 5737 -53505 5783 -53305
rect 7726 -53505 7772 -53305
rect 7922 -53505 7968 -53305
rect 8118 -53505 8164 -53305
rect 8232 -53505 8278 -53305
rect 8428 -53505 8474 -53305
rect 8541 -53505 8587 -53305
rect 8737 -53505 8783 -53305
rect -13646 -54617 -13600 -54417
rect -13450 -54617 -13404 -54417
rect -13254 -54617 -13208 -54417
rect -11903 -54617 -11857 -54417
rect -11707 -54617 -11661 -54417
rect -11511 -54617 -11465 -54417
rect -10946 -54617 -10900 -54417
rect -10750 -54617 -10704 -54417
rect -10554 -54617 -10508 -54417
rect -9203 -54617 -9157 -54417
rect -9007 -54617 -8961 -54417
rect -8811 -54617 -8765 -54417
rect -8321 -54617 -8275 -54417
rect -8125 -54617 -8079 -54417
rect -7929 -54617 -7883 -54417
rect -12974 -55805 -12777 -55751
rect -18169 -58731 -17990 -58564
rect -21221 -59711 -21175 -59111
rect -21025 -59711 -20979 -59111
rect -20015 -59440 -19969 -59040
rect -19819 -59440 -19773 -59040
rect -19110 -59441 -19064 -59041
rect -18914 -59441 -18868 -59041
rect -20189 -59602 -20131 -59465
rect -20189 -60511 -20154 -59602
rect -20209 -60648 -20151 -60511
rect -21558 -62129 -21512 -61929
rect -21362 -62129 -21316 -61929
rect -20820 -62129 -20774 -61929
rect -20624 -62129 -20578 -61929
rect -20428 -62129 -20382 -61929
rect -20232 -62129 -20186 -61929
rect -18948 -62293 -18772 -61662
rect -18142 -60495 -18016 -58731
rect -12831 -56836 -12777 -55805
rect -12719 -56246 -12673 -55946
rect -12523 -56246 -12477 -55946
rect -12327 -56246 -12281 -55946
rect -12110 -56247 -12064 -56147
rect -11914 -56247 -11868 -56147
rect -11718 -56247 -11672 -56147
rect -11522 -56247 -11476 -56147
rect -11272 -56335 -11226 -55735
rect -11076 -56335 -11030 -55735
rect -10653 -56335 -10607 -55735
rect -14442 -57012 -12777 -56836
rect -18143 -60667 -17951 -60495
rect -17708 -60270 -17662 -59970
rect -17512 -60270 -17466 -59970
rect -17316 -60270 -17270 -59970
rect -17099 -60271 -17053 -60171
rect -16903 -60271 -16857 -60171
rect -16707 -60271 -16661 -60171
rect -16511 -60271 -16465 -60171
rect -16261 -60359 -16215 -59759
rect -16065 -60359 -16019 -59759
rect -15642 -60359 -15596 -59759
rect -17682 -61199 -17636 -60999
rect -17486 -61199 -17440 -60999
rect -17290 -61199 -17244 -60999
rect -17094 -61199 -17048 -60999
rect -16709 -61170 -16663 -60870
rect -16513 -61170 -16467 -60870
rect -16317 -61170 -16271 -60870
rect -16100 -60969 -16054 -60869
rect -15904 -60969 -15858 -60869
rect -15708 -60969 -15662 -60869
rect -15512 -60969 -15466 -60869
rect -14442 -62751 -14266 -57012
rect -12831 -57209 -12777 -57012
rect -12693 -57175 -12647 -56975
rect -12881 -57359 -12751 -57209
rect -12497 -57175 -12451 -56975
rect -12301 -57175 -12255 -56975
rect -12105 -57175 -12059 -56975
rect -11720 -57146 -11674 -56846
rect -11524 -57146 -11478 -56846
rect -11328 -57146 -11282 -56846
rect -11111 -56945 -11065 -56845
rect -10915 -56945 -10869 -56845
rect -10719 -56945 -10673 -56845
rect -10523 -56945 -10477 -56845
rect -13744 -58226 -13698 -58026
rect -13548 -58226 -13502 -58026
rect -13352 -58226 -13306 -58026
rect -12907 -58226 -12861 -58026
rect -12711 -58226 -12665 -58026
rect -12515 -58226 -12469 -58026
rect -11044 -58226 -10998 -58026
rect -10848 -58226 -10802 -58026
rect -10652 -58226 -10606 -58026
rect -10207 -58226 -10161 -58026
rect -10011 -58226 -9965 -58026
rect -9815 -58226 -9769 -58026
rect -13646 -59544 -13600 -59344
rect -13450 -59544 -13404 -59344
rect -13254 -59544 -13208 -59344
rect -11903 -59544 -11857 -59344
rect -11707 -59544 -11661 -59344
rect -11511 -59544 -11465 -59344
rect -10946 -59544 -10900 -59344
rect -10750 -59544 -10704 -59344
rect -10554 -59544 -10508 -59344
rect -9203 -59544 -9157 -59344
rect -9007 -59544 -8961 -59344
rect -8811 -59544 -8765 -59344
rect -8321 -59544 -8275 -59344
rect -8125 -59544 -8079 -59344
rect -7929 -59544 -7883 -59344
rect -7355 -58643 -7309 -58043
rect -6932 -58643 -6886 -58043
rect -6736 -58643 -6690 -58043
rect -5739 -54566 -5603 -54492
rect -5739 -54948 -5688 -54566
rect -5613 -54834 -5567 -54634
rect -5417 -54834 -5371 -54634
rect -5221 -54834 -5175 -54634
rect -3946 -54063 -3823 -53927
rect -3942 -54694 -3828 -54063
rect -3947 -54830 -3824 -54694
rect -1379 -54098 -1256 -53962
rect -1375 -54550 -1261 -54098
rect -1380 -54686 -1257 -54550
rect 1104 -54098 1227 -53962
rect 1108 -54515 1222 -54098
rect 1103 -54516 1226 -54515
rect 1103 -54578 1409 -54516
rect 4337 -53772 4476 -53763
rect 5415 -53770 5554 -53769
rect 5415 -53772 6774 -53770
rect 4337 -53798 6774 -53772
rect 4337 -53800 5554 -53798
rect 4337 -53817 4476 -53800
rect 5415 -53823 5554 -53800
rect 6746 -54396 6774 -53798
rect 7337 -53772 7476 -53763
rect 8415 -53770 8554 -53769
rect 8313 -53772 10924 -53770
rect 7337 -53798 10924 -53772
rect 7337 -53800 8554 -53798
rect 7337 -53817 7476 -53800
rect 8415 -53823 8554 -53800
rect 6746 -54424 10773 -54396
rect -5739 -54999 10126 -54948
rect 38 -55256 10001 -55205
rect 4768 -55357 4891 -55348
rect 5169 -55357 5292 -55346
rect -121 -55372 2 -55360
rect 173 -55372 296 -55359
rect -121 -55487 296 -55372
rect -121 -55496 2 -55487
rect 173 -55495 296 -55487
rect 3151 -55387 3274 -55372
rect 3540 -55387 3663 -55371
rect 3151 -55494 3663 -55387
rect 4768 -55464 5292 -55357
rect 4768 -55484 4891 -55464
rect 5169 -55482 5292 -55464
rect 6525 -55364 6648 -55351
rect 7741 -55364 7864 -55352
rect 6525 -55469 7864 -55364
rect 6525 -55487 6648 -55469
rect 7741 -55488 7864 -55469
rect 3151 -55508 3274 -55494
rect 3540 -55507 3663 -55494
rect -5772 -55737 -5726 -55537
rect -5576 -55737 -5530 -55537
rect -5380 -55737 -5334 -55537
rect -4029 -55737 -3983 -55537
rect -3833 -55737 -3787 -55537
rect -3637 -55737 -3591 -55537
rect -3072 -55737 -3026 -55537
rect -2876 -55737 -2830 -55537
rect -2680 -55737 -2634 -55537
rect -1329 -55737 -1283 -55537
rect -1133 -55737 -1087 -55537
rect -937 -55737 -891 -55537
rect -447 -55737 -401 -55537
rect -251 -55737 -205 -55537
rect -55 -55737 -9 -55537
rect 287 -55754 333 -55554
rect 483 -55754 529 -55554
rect 1025 -55754 1071 -55554
rect 1221 -55754 1267 -55554
rect 1417 -55754 1463 -55554
rect 1613 -55754 1659 -55554
rect 2020 -55667 2066 -55567
rect -5247 -56234 -5115 -56174
rect -5211 -56701 -5151 -56234
rect 2216 -55667 2262 -55567
rect 2412 -55667 2458 -55567
rect 2608 -55667 2654 -55567
rect -5870 -57055 -5824 -56855
rect -5674 -57055 -5628 -56855
rect -5478 -57055 -5432 -56855
rect 2825 -55868 2871 -55568
rect 3021 -55868 3067 -55568
rect 3217 -55868 3263 -55568
rect 3625 -55669 3671 -55569
rect 3821 -55669 3867 -55569
rect 4017 -55669 4063 -55569
rect 4213 -55669 4259 -55569
rect 4430 -55870 4476 -55570
rect 4626 -55870 4672 -55570
rect 4822 -55870 4868 -55570
rect 5249 -55745 5295 -55545
rect 5445 -55745 5491 -55545
rect 5987 -55745 6033 -55545
rect 6183 -55745 6229 -55545
rect 6379 -55745 6425 -55545
rect 6575 -55745 6621 -55545
rect 7736 -55756 7782 -55556
rect 7932 -55756 7978 -55556
rect 8128 -55756 8174 -55556
rect 8242 -55756 8288 -55556
rect 8438 -55756 8484 -55556
rect 8551 -55756 8597 -55556
rect 8747 -55756 8793 -55556
rect 7347 -56023 7486 -56014
rect 8425 -56021 8564 -56020
rect 9755 -56021 9806 -56013
rect 8425 -56023 9806 -56021
rect 7347 -56049 9806 -56023
rect 7347 -56051 8564 -56049
rect 7347 -56068 7486 -56051
rect 8425 -56074 8564 -56051
rect 9755 -56064 9806 -56049
rect -5033 -57055 -4987 -56855
rect -4837 -57055 -4791 -56855
rect -4641 -57055 -4595 -56855
rect -3170 -57055 -3124 -56855
rect -2974 -57055 -2928 -56855
rect -2778 -57055 -2732 -56855
rect -2333 -57055 -2287 -56855
rect -2137 -57055 -2091 -56855
rect -1941 -57055 -1895 -56855
rect -5870 -58493 -5824 -58293
rect -5674 -58493 -5628 -58293
rect -5478 -58493 -5432 -58293
rect -5033 -58493 -4987 -58293
rect -4837 -58493 -4791 -58293
rect -4641 -58493 -4595 -58293
rect -3170 -58493 -3124 -58293
rect -2974 -58493 -2928 -58293
rect -2778 -58493 -2732 -58293
rect -2333 -58493 -2287 -58293
rect -2137 -58493 -2091 -58293
rect -1941 -58493 -1895 -58293
rect -3474 -59085 -3337 -59025
rect -3425 -59533 -3365 -59085
rect -2499 -59026 -2439 -58662
rect -2528 -59086 -2396 -59026
rect -5772 -59811 -5726 -59611
rect -5576 -59811 -5530 -59611
rect -5380 -59811 -5334 -59611
rect -4029 -59811 -3983 -59611
rect -3833 -59811 -3787 -59611
rect -3637 -59811 -3591 -59611
rect -3072 -59811 -3026 -59611
rect -2876 -59811 -2830 -59611
rect -2680 -59811 -2634 -59611
rect -1329 -59811 -1283 -59611
rect -1133 -59811 -1087 -59611
rect -937 -59811 -891 -59611
rect -447 -59811 -401 -59611
rect -251 -59811 -205 -59611
rect -55 -59811 -9 -59611
rect 287 -59794 333 -59594
rect 483 -59794 529 -59594
rect 1025 -59794 1071 -59594
rect 1221 -59794 1267 -59594
rect 1417 -59794 1463 -59594
rect 1613 -59794 1659 -59594
rect 2020 -59781 2066 -59681
rect 2216 -59781 2262 -59681
rect 2412 -59781 2458 -59681
rect 2608 -59781 2654 -59681
rect 2825 -59780 2871 -59480
rect 3021 -59780 3067 -59480
rect 3217 -59780 3263 -59480
rect 3625 -59779 3671 -59679
rect 3821 -59779 3867 -59679
rect 4017 -59779 4063 -59679
rect 4213 -59779 4259 -59679
rect 4430 -59778 4476 -59478
rect 7347 -59297 7486 -59280
rect 8425 -59297 8564 -59274
rect 7347 -59299 8564 -59297
rect 9536 -59299 9681 -59204
rect 9768 -59299 9796 -56064
rect 7347 -59325 9798 -59299
rect 7347 -59334 7486 -59325
rect 8425 -59327 9798 -59325
rect 8425 -59328 8564 -59327
rect 9536 -59339 9681 -59327
rect 4626 -59778 4672 -59478
rect 4822 -59778 4868 -59478
rect 5249 -59803 5295 -59603
rect 5445 -59803 5491 -59603
rect 5987 -59803 6033 -59603
rect 6183 -59803 6229 -59603
rect 6379 -59803 6425 -59603
rect 6575 -59803 6621 -59603
rect 7736 -59792 7782 -59592
rect 7932 -59792 7978 -59592
rect 8128 -59792 8174 -59592
rect 8242 -59792 8288 -59592
rect 8438 -59792 8484 -59592
rect 8551 -59792 8597 -59592
rect 8747 -59792 8793 -59592
rect -121 -59861 2 -59852
rect 173 -59861 296 -59853
rect -121 -59976 296 -59861
rect 3151 -59854 3274 -59840
rect 3540 -59854 3663 -59841
rect 3151 -59961 3663 -59854
rect 3151 -59976 3274 -59961
rect -121 -59988 2 -59976
rect 173 -59989 296 -59976
rect 3540 -59977 3663 -59961
rect 4768 -59884 4891 -59864
rect 5169 -59884 5292 -59866
rect 4768 -59991 5292 -59884
rect 4768 -60000 4891 -59991
rect 5169 -60002 5292 -59991
rect 6525 -59879 6648 -59861
rect 7741 -59879 7864 -59860
rect 6525 -59984 7864 -59879
rect 6525 -59997 6648 -59984
rect 7741 -59996 7864 -59984
rect 9950 -60092 10001 -55256
rect 38 -60143 10001 -60092
rect 9950 -60214 10001 -60143
rect 9830 -60321 10021 -60214
rect 10075 -60349 10126 -54999
rect -4082 -60400 10126 -60349
rect -5663 -61548 -5524 -61531
rect -4585 -61548 -4446 -61525
rect -5663 -61550 -4446 -61548
rect -4082 -61550 -4054 -60400
rect -5663 -61576 -4054 -61550
rect -5663 -61585 -5524 -61576
rect -4585 -61578 -4054 -61576
rect -4585 -61579 -4446 -61578
rect -3947 -60654 -3824 -60518
rect -3942 -61285 -3828 -60654
rect -3946 -61421 -3823 -61285
rect -1380 -60798 -1257 -60662
rect -1375 -61250 -1261 -60798
rect -1379 -61386 -1256 -61250
rect 1103 -60832 1409 -60770
rect 1103 -60833 1226 -60832
rect 1108 -61250 1222 -60833
rect 1104 -61386 1227 -61250
rect 9387 -60924 9526 -60909
rect 10745 -60924 10773 -54424
rect 6746 -60952 10773 -60924
rect 4337 -61548 4476 -61531
rect 5415 -61548 5554 -61525
rect 4337 -61550 5554 -61548
rect 6746 -61550 6774 -60952
rect 9387 -60956 9526 -60952
rect 4337 -61576 6774 -61550
rect 4337 -61585 4476 -61576
rect 5415 -61578 6774 -61576
rect 5415 -61579 5554 -61578
rect 7337 -61548 7476 -61531
rect 8415 -61548 8554 -61525
rect 7337 -61550 8554 -61548
rect 9352 -61550 9417 -61446
rect 10896 -61550 10924 -53798
rect 7337 -61576 10924 -61550
rect 7337 -61585 7476 -61576
rect 8313 -61578 10924 -61576
rect 8415 -61579 8554 -61578
rect 9352 -61583 9417 -61578
rect -5274 -62043 -5228 -61843
rect -5078 -62043 -5032 -61843
rect -4882 -62043 -4836 -61843
rect -4768 -62043 -4722 -61843
rect -4572 -62043 -4526 -61843
rect -4459 -62043 -4413 -61843
rect -4263 -62043 -4217 -61843
rect -2774 -62043 -2728 -61843
rect -2578 -62043 -2532 -61843
rect -2382 -62043 -2336 -61843
rect -2268 -62043 -2222 -61843
rect -2072 -62043 -2026 -61843
rect -1959 -62043 -1913 -61843
rect -1763 -62043 -1717 -61843
rect -274 -62043 -228 -61843
rect -78 -62043 -32 -61843
rect 118 -62043 164 -61843
rect 232 -62043 278 -61843
rect 428 -62043 474 -61843
rect 541 -62043 587 -61843
rect 737 -62043 783 -61843
rect 2226 -62043 2272 -61843
rect 2422 -62043 2468 -61843
rect 2618 -62043 2664 -61843
rect 2732 -62043 2778 -61843
rect 2928 -62043 2974 -61843
rect 3041 -62043 3087 -61843
rect 3237 -62043 3283 -61843
rect 4726 -62043 4772 -61843
rect 4922 -62043 4968 -61843
rect 5118 -62043 5164 -61843
rect 5232 -62043 5278 -61843
rect 5428 -62043 5474 -61843
rect 5541 -62043 5587 -61843
rect 5737 -62043 5783 -61843
rect 7726 -62043 7772 -61843
rect 7922 -62043 7968 -61843
rect 8118 -62043 8164 -61843
rect 8232 -62043 8278 -61843
rect 8428 -62043 8474 -61843
rect 8541 -62043 8587 -61843
rect 8737 -62043 8783 -61843
rect 11260 -62106 11555 -54816
rect -22800 -64647 -22587 -64469
rect 9347 -62820 9408 -62216
rect 9465 -62220 9509 -62217
rect 9294 -62943 9417 -62820
rect 9456 -63053 9516 -62220
rect 9400 -63176 9523 -63053
rect 9555 -63310 9616 -62363
rect 9493 -63433 9617 -63310
rect 10208 -62375 11555 -62106
rect 11260 -64637 11555 -62375
rect 16597 -54773 26830 -54733
rect 16597 -55067 27010 -54773
rect 16597 -55085 26975 -55067
rect 18441 -55929 18620 -55853
rect 18441 -56004 20111 -55929
rect 18441 -56042 18620 -56004
rect 20036 -56079 20111 -56004
rect 21981 -56006 22027 -55806
rect 22177 -56006 22223 -55806
rect 22373 -56006 22419 -55806
rect 22818 -56006 22864 -55806
rect 23014 -56006 23060 -55806
rect 23210 -56006 23256 -55806
rect 24681 -56006 24727 -55806
rect 24877 -56006 24923 -55806
rect 25073 -56006 25119 -55806
rect 20009 -56214 20141 -56079
rect 25518 -56006 25564 -55806
rect 25714 -56006 25760 -55806
rect 25910 -56006 25956 -55806
rect 18774 -57204 18820 -56604
rect 18970 -57204 19016 -56604
rect 22525 -56539 22585 -56175
rect 22482 -56599 22614 -56539
rect 23423 -56598 23560 -56538
rect 23451 -57046 23511 -56598
rect 20095 -57324 20141 -57124
rect 20291 -57324 20337 -57124
rect 20487 -57324 20533 -57124
rect 20977 -57324 21023 -57124
rect 21173 -57324 21219 -57124
rect 21369 -57324 21415 -57124
rect 22720 -57324 22766 -57124
rect 22916 -57324 22962 -57124
rect 23112 -57324 23158 -57124
rect 23677 -57324 23723 -57124
rect 23873 -57324 23919 -57124
rect 24069 -57324 24115 -57124
rect 25420 -57324 25466 -57124
rect 25616 -57324 25662 -57124
rect 25812 -57324 25858 -57124
rect 18769 -59550 18815 -59150
rect 18965 -59550 19011 -59150
rect 19715 -59550 19761 -59150
rect 19911 -59550 19957 -59150
rect 22540 -58276 22586 -57876
rect 22736 -58276 22782 -57876
rect 22932 -58276 22978 -57876
rect 20631 -59584 20677 -59384
rect 20827 -59584 20873 -59384
rect 21023 -59584 21069 -59384
rect 21219 -59584 21265 -59384
rect 21761 -59584 21807 -59384
rect 21957 -59584 22003 -59384
rect 22490 -59577 22536 -59377
rect 22686 -59577 22732 -59377
rect 22882 -59577 22928 -59377
rect 23370 -59506 23416 -58806
rect 23566 -59506 23612 -58806
rect 23770 -59506 23816 -58806
rect 23966 -59506 24012 -58806
rect 24370 -59506 24416 -58806
rect 24566 -59506 24612 -58806
rect 24770 -59506 24816 -58806
rect 24966 -59506 25012 -58806
rect 25370 -59506 25416 -58806
rect 25566 -59506 25612 -58806
rect 25770 -59506 25816 -58806
rect 25966 -59506 26012 -58806
rect 11967 -60562 12013 -60362
rect 12163 -60562 12209 -60362
rect 12359 -60562 12405 -60362
rect 12849 -60562 12895 -60362
rect 13045 -60562 13091 -60362
rect 13241 -60562 13287 -60362
rect 14592 -60562 14638 -60362
rect 14788 -60562 14834 -60362
rect 14984 -60562 15030 -60362
rect 15549 -60562 15595 -60362
rect 15745 -60562 15791 -60362
rect 15941 -60562 15987 -60362
rect 17292 -60562 17338 -60362
rect 17488 -60562 17534 -60362
rect 17684 -60562 17730 -60362
rect 14354 -61147 14486 -61087
rect 14397 -61511 14457 -61147
rect 15323 -61088 15383 -60640
rect 15295 -61148 15432 -61088
rect 13853 -61880 13899 -61680
rect 14049 -61880 14095 -61680
rect 14245 -61880 14291 -61680
rect 14690 -61880 14736 -61680
rect 14886 -61880 14932 -61680
rect 15082 -61880 15128 -61680
rect 16553 -61880 16599 -61680
rect 16749 -61880 16795 -61680
rect 16945 -61880 16991 -61680
rect 17390 -61880 17436 -61680
rect 17586 -61880 17632 -61680
rect 17782 -61880 17828 -61680
rect 26730 -62184 26975 -55085
rect 27598 -54925 27811 -54886
rect 27598 -54979 29036 -54925
rect 27598 -55019 27811 -54979
rect 28982 -55269 29036 -54979
rect 28982 -55323 29310 -55269
rect 29256 -55378 29310 -55323
rect 27599 -56846 27858 -56583
rect 28353 -55653 28399 -55453
rect 28549 -55653 28595 -55453
rect 28745 -55653 28791 -55453
rect 29230 -55436 29389 -55378
rect 28941 -55653 28987 -55453
rect 29326 -55782 29372 -55482
rect 29522 -55782 29568 -55482
rect 29718 -55782 29764 -55482
rect 29935 -55783 29981 -55683
rect 30131 -55783 30177 -55683
rect 30327 -55783 30373 -55683
rect 30523 -55783 30569 -55683
rect 30605 -56098 30679 -56082
rect 30833 -56098 30943 -56062
rect 30605 -56194 30943 -56098
rect 30605 -56200 30679 -56194
rect 30833 -56212 30943 -56194
rect 28327 -56682 28373 -56382
rect 28523 -56682 28569 -56382
rect 28719 -56682 28765 -56382
rect 28936 -56481 28982 -56381
rect 29132 -56481 29178 -56381
rect 29328 -56481 29374 -56381
rect 29524 -56481 29570 -56381
rect 29774 -56893 29820 -56293
rect 29970 -56893 30016 -56293
rect 30393 -56893 30439 -56293
rect 31766 -56651 31812 -56151
rect 31962 -56651 32008 -56151
rect 32557 -56651 32603 -56151
rect 32687 -56651 32733 -56151
rect 32915 -56451 32961 -56151
rect 33111 -56451 33157 -56151
rect 28345 -59106 28391 -58906
rect 28541 -59106 28587 -58906
rect 28737 -59106 28783 -58906
rect 28933 -59106 28979 -58906
rect 29318 -59235 29364 -58935
rect 29514 -59235 29560 -58935
rect 29710 -59235 29756 -58935
rect 29927 -59236 29973 -59136
rect 30123 -59236 30169 -59136
rect 30319 -59236 30365 -59136
rect 30515 -59236 30561 -59136
rect 29520 -59510 29703 -59469
rect 30823 -59510 30919 -59481
rect 29520 -59592 30919 -59510
rect 29520 -59599 29703 -59592
rect 30823 -59618 30919 -59592
rect 28319 -60135 28365 -59835
rect 28515 -60135 28561 -59835
rect 28711 -60135 28757 -59835
rect 28928 -59934 28974 -59834
rect 29124 -59934 29170 -59834
rect 29320 -59934 29366 -59834
rect 29516 -59934 29562 -59834
rect 29766 -60346 29812 -59746
rect 29962 -60346 30008 -59746
rect 30385 -60346 30431 -59746
rect 32013 -59137 32059 -58937
rect 32209 -59137 32255 -58937
rect 32405 -59137 32451 -58937
rect 32601 -59137 32647 -58937
rect 32986 -59266 33032 -58966
rect 33182 -59266 33228 -58966
rect 33378 -59266 33424 -58966
rect 33595 -59267 33641 -59167
rect 33791 -59267 33837 -59167
rect 33987 -59267 34033 -59167
rect 34183 -59267 34229 -59167
rect 34243 -59532 34334 -59520
rect 34493 -59532 34644 -59505
rect 34243 -59671 34644 -59532
rect 34243 -59683 34334 -59671
rect 34493 -59696 34644 -59671
rect 31987 -60166 32033 -59866
rect 32183 -60166 32229 -59866
rect 32379 -60166 32425 -59866
rect 32596 -59965 32642 -59865
rect 32792 -59965 32838 -59865
rect 32988 -59965 33034 -59865
rect 33184 -59965 33230 -59865
rect 33434 -60377 33480 -59777
rect 33630 -60377 33676 -59777
rect 34053 -60377 34099 -59777
rect 36793 -55664 36839 -55464
rect 36989 -55664 37035 -55464
rect 37185 -55664 37231 -55464
rect 37381 -55664 37427 -55464
rect 37766 -55793 37812 -55493
rect 37962 -55793 38008 -55493
rect 38158 -55793 38204 -55493
rect 38375 -55794 38421 -55694
rect 38571 -55794 38617 -55694
rect 38767 -55794 38813 -55694
rect 38963 -55794 39009 -55694
rect 39045 -56109 39119 -56093
rect 39273 -56109 39383 -56073
rect 39045 -56205 39383 -56109
rect 39045 -56211 39119 -56205
rect 39273 -56223 39383 -56205
rect 36767 -56693 36813 -56393
rect 36963 -56693 37009 -56393
rect 37159 -56693 37205 -56393
rect 37376 -56492 37422 -56392
rect 37572 -56492 37618 -56392
rect 37768 -56492 37814 -56392
rect 37964 -56492 38010 -56392
rect 38214 -56904 38260 -56304
rect 38410 -56904 38456 -56304
rect 38833 -56904 38879 -56304
rect 40206 -56662 40252 -56162
rect 40402 -56662 40448 -56162
rect 40997 -56662 41043 -56162
rect 41127 -56662 41173 -56162
rect 41355 -56462 41401 -56162
rect 41551 -56462 41597 -56162
rect 36785 -59117 36831 -58917
rect 36981 -59117 37027 -58917
rect 37177 -59117 37223 -58917
rect 37373 -59117 37419 -58917
rect 37758 -59246 37804 -58946
rect 37954 -59246 38000 -58946
rect 38150 -59246 38196 -58946
rect 38367 -59247 38413 -59147
rect 38563 -59247 38609 -59147
rect 38759 -59247 38805 -59147
rect 38955 -59247 39001 -59147
rect 37960 -59521 38143 -59480
rect 39263 -59521 39359 -59492
rect 37960 -59603 39359 -59521
rect 37960 -59610 38143 -59603
rect 39263 -59629 39359 -59603
rect 36759 -60146 36805 -59846
rect 36955 -60146 37001 -59846
rect 37151 -60146 37197 -59846
rect 37368 -59945 37414 -59845
rect 37564 -59945 37610 -59845
rect 37760 -59945 37806 -59845
rect 37956 -59945 38002 -59845
rect 38206 -60357 38252 -59757
rect 38402 -60357 38448 -59757
rect 38825 -60357 38871 -59757
rect 40453 -59148 40499 -58948
rect 40649 -59148 40695 -58948
rect 40845 -59148 40891 -58948
rect 41041 -59148 41087 -58948
rect 41426 -59277 41472 -58977
rect 41622 -59277 41668 -58977
rect 41818 -59277 41864 -58977
rect 42035 -59278 42081 -59178
rect 42231 -59278 42277 -59178
rect 42427 -59278 42473 -59178
rect 42623 -59278 42669 -59178
rect 42683 -59543 42774 -59531
rect 42933 -59543 43084 -59516
rect 42683 -59682 43084 -59543
rect 42683 -59694 42774 -59682
rect 42933 -59707 43084 -59682
rect 40427 -60177 40473 -59877
rect 40623 -60177 40669 -59877
rect 40819 -60177 40865 -59877
rect 41036 -59976 41082 -59876
rect 41232 -59976 41278 -59876
rect 41428 -59976 41474 -59876
rect 41624 -59976 41670 -59876
rect 41874 -60388 41920 -59788
rect 42070 -60388 42116 -59788
rect 42493 -60388 42539 -59788
rect 45656 -55703 45702 -55503
rect 45852 -55703 45898 -55503
rect 46048 -55703 46094 -55503
rect 46244 -55703 46290 -55503
rect 46629 -55832 46675 -55532
rect 46825 -55832 46871 -55532
rect 47021 -55832 47067 -55532
rect 47238 -55833 47284 -55733
rect 47434 -55833 47480 -55733
rect 47630 -55833 47676 -55733
rect 47826 -55833 47872 -55733
rect 47908 -56148 47982 -56132
rect 48136 -56148 48246 -56112
rect 47908 -56244 48246 -56148
rect 47908 -56250 47982 -56244
rect 48136 -56262 48246 -56244
rect 45630 -56732 45676 -56432
rect 45826 -56732 45872 -56432
rect 46022 -56732 46068 -56432
rect 46239 -56531 46285 -56431
rect 46435 -56531 46481 -56431
rect 46631 -56531 46677 -56431
rect 46827 -56531 46873 -56431
rect 47077 -56943 47123 -56343
rect 47273 -56943 47319 -56343
rect 47696 -56943 47742 -56343
rect 49069 -56701 49115 -56201
rect 49265 -56701 49311 -56201
rect 49860 -56701 49906 -56201
rect 49990 -56701 50036 -56201
rect 50218 -56501 50264 -56201
rect 50414 -56501 50460 -56201
rect 45648 -59156 45694 -58956
rect 45844 -59156 45890 -58956
rect 46040 -59156 46086 -58956
rect 46236 -59156 46282 -58956
rect 46621 -59285 46667 -58985
rect 46817 -59285 46863 -58985
rect 47013 -59285 47059 -58985
rect 47230 -59286 47276 -59186
rect 47426 -59286 47472 -59186
rect 47622 -59286 47668 -59186
rect 47818 -59286 47864 -59186
rect 46823 -59560 47006 -59519
rect 48126 -59560 48222 -59531
rect 46823 -59642 48222 -59560
rect 46823 -59649 47006 -59642
rect 48126 -59668 48222 -59642
rect 45622 -60185 45668 -59885
rect 45818 -60185 45864 -59885
rect 46014 -60185 46060 -59885
rect 46231 -59984 46277 -59884
rect 46427 -59984 46473 -59884
rect 46623 -59984 46669 -59884
rect 46819 -59984 46865 -59884
rect 47069 -60396 47115 -59796
rect 47265 -60396 47311 -59796
rect 47688 -60396 47734 -59796
rect 49316 -59187 49362 -58987
rect 49512 -59187 49558 -58987
rect 49708 -59187 49754 -58987
rect 49904 -59187 49950 -58987
rect 50289 -59316 50335 -59016
rect 50485 -59316 50531 -59016
rect 50681 -59316 50727 -59016
rect 50898 -59317 50944 -59217
rect 51094 -59317 51140 -59217
rect 51290 -59317 51336 -59217
rect 51486 -59317 51532 -59217
rect 51546 -59582 51637 -59570
rect 51796 -59582 51947 -59555
rect 51546 -59721 51947 -59582
rect 51546 -59733 51637 -59721
rect 51796 -59746 51947 -59721
rect 49290 -60216 49336 -59916
rect 49486 -60216 49532 -59916
rect 49682 -60216 49728 -59916
rect 49899 -60015 49945 -59915
rect 50095 -60015 50141 -59915
rect 50291 -60015 50337 -59915
rect 50487 -60015 50533 -59915
rect 50737 -60427 50783 -59827
rect 50933 -60427 50979 -59827
rect 51356 -60427 51402 -59827
rect 54854 -55669 54900 -55469
rect 55050 -55669 55096 -55469
rect 55246 -55669 55292 -55469
rect 55442 -55669 55488 -55469
rect 55827 -55798 55873 -55498
rect 56023 -55798 56069 -55498
rect 56219 -55798 56265 -55498
rect 56436 -55799 56482 -55699
rect 56632 -55799 56678 -55699
rect 56828 -55799 56874 -55699
rect 57024 -55799 57070 -55699
rect 57106 -56114 57180 -56098
rect 57334 -56114 57444 -56078
rect 57106 -56210 57444 -56114
rect 57106 -56216 57180 -56210
rect 57334 -56228 57444 -56210
rect 54828 -56698 54874 -56398
rect 55024 -56698 55070 -56398
rect 55220 -56698 55266 -56398
rect 55437 -56497 55483 -56397
rect 55633 -56497 55679 -56397
rect 55829 -56497 55875 -56397
rect 56025 -56497 56071 -56397
rect 56275 -56909 56321 -56309
rect 56471 -56909 56517 -56309
rect 56894 -56909 56940 -56309
rect 58267 -56667 58313 -56167
rect 58463 -56667 58509 -56167
rect 59058 -56667 59104 -56167
rect 59188 -56667 59234 -56167
rect 59416 -56467 59462 -56167
rect 59612 -56467 59658 -56167
rect 54846 -59122 54892 -58922
rect 55042 -59122 55088 -58922
rect 55238 -59122 55284 -58922
rect 55434 -59122 55480 -58922
rect 55819 -59251 55865 -58951
rect 56015 -59251 56061 -58951
rect 56211 -59251 56257 -58951
rect 56428 -59252 56474 -59152
rect 56624 -59252 56670 -59152
rect 56820 -59252 56866 -59152
rect 57016 -59252 57062 -59152
rect 56021 -59526 56204 -59485
rect 57324 -59526 57420 -59497
rect 56021 -59608 57420 -59526
rect 56021 -59615 56204 -59608
rect 57324 -59634 57420 -59608
rect 54820 -60151 54866 -59851
rect 55016 -60151 55062 -59851
rect 55212 -60151 55258 -59851
rect 55429 -59950 55475 -59850
rect 55625 -59950 55671 -59850
rect 55821 -59950 55867 -59850
rect 56017 -59950 56063 -59850
rect 56267 -60362 56313 -59762
rect 56463 -60362 56509 -59762
rect 56886 -60362 56932 -59762
rect 58514 -59153 58560 -58953
rect 58710 -59153 58756 -58953
rect 58906 -59153 58952 -58953
rect 59102 -59153 59148 -58953
rect 59487 -59282 59533 -58982
rect 59683 -59282 59729 -58982
rect 59879 -59282 59925 -58982
rect 60096 -59283 60142 -59183
rect 60292 -59283 60338 -59183
rect 60488 -59283 60534 -59183
rect 60684 -59283 60730 -59183
rect 60744 -59548 60835 -59536
rect 60994 -59548 61145 -59521
rect 60744 -59687 61145 -59548
rect 60744 -59699 60835 -59687
rect 60994 -59712 61145 -59687
rect 58488 -60182 58534 -59882
rect 58684 -60182 58730 -59882
rect 58880 -60182 58926 -59882
rect 59097 -59981 59143 -59881
rect 59293 -59981 59339 -59881
rect 59489 -59981 59535 -59881
rect 59685 -59981 59731 -59881
rect 59935 -60393 59981 -59793
rect 60131 -60393 60177 -59793
rect 60554 -60393 60600 -59793
rect 63608 -55603 63654 -55403
rect 63804 -55603 63850 -55403
rect 64000 -55603 64046 -55403
rect 64196 -55603 64242 -55403
rect 64581 -55732 64627 -55432
rect 64777 -55732 64823 -55432
rect 64973 -55732 65019 -55432
rect 65190 -55733 65236 -55633
rect 65386 -55733 65432 -55633
rect 65582 -55733 65628 -55633
rect 65778 -55733 65824 -55633
rect 65860 -56048 65934 -56032
rect 66088 -56048 66198 -56012
rect 65860 -56144 66198 -56048
rect 65860 -56150 65934 -56144
rect 66088 -56162 66198 -56144
rect 63582 -56632 63628 -56332
rect 63778 -56632 63824 -56332
rect 63974 -56632 64020 -56332
rect 64191 -56431 64237 -56331
rect 64387 -56431 64433 -56331
rect 64583 -56431 64629 -56331
rect 64779 -56431 64825 -56331
rect 65029 -56843 65075 -56243
rect 65225 -56843 65271 -56243
rect 65648 -56843 65694 -56243
rect 67021 -56601 67067 -56101
rect 67217 -56601 67263 -56101
rect 67812 -56601 67858 -56101
rect 67942 -56601 67988 -56101
rect 68170 -56401 68216 -56101
rect 68366 -56401 68412 -56101
rect 63600 -59056 63646 -58856
rect 63796 -59056 63842 -58856
rect 63992 -59056 64038 -58856
rect 64188 -59056 64234 -58856
rect 64573 -59185 64619 -58885
rect 64769 -59185 64815 -58885
rect 64965 -59185 65011 -58885
rect 65182 -59186 65228 -59086
rect 65378 -59186 65424 -59086
rect 65574 -59186 65620 -59086
rect 65770 -59186 65816 -59086
rect 64775 -59460 64958 -59419
rect 66078 -59460 66174 -59431
rect 64775 -59542 66174 -59460
rect 64775 -59549 64958 -59542
rect 66078 -59568 66174 -59542
rect 63574 -60085 63620 -59785
rect 63770 -60085 63816 -59785
rect 63966 -60085 64012 -59785
rect 64183 -59884 64229 -59784
rect 64379 -59884 64425 -59784
rect 64575 -59884 64621 -59784
rect 64771 -59884 64817 -59784
rect 65021 -60296 65067 -59696
rect 65217 -60296 65263 -59696
rect 65640 -60296 65686 -59696
rect 67268 -59087 67314 -58887
rect 67464 -59087 67510 -58887
rect 67660 -59087 67706 -58887
rect 67856 -59087 67902 -58887
rect 68241 -59216 68287 -58916
rect 68437 -59216 68483 -58916
rect 68633 -59216 68679 -58916
rect 68850 -59217 68896 -59117
rect 69046 -59217 69092 -59117
rect 69242 -59217 69288 -59117
rect 69438 -59217 69484 -59117
rect 69498 -59482 69589 -59470
rect 69748 -59482 69899 -59455
rect 69498 -59621 69899 -59482
rect 69498 -59633 69589 -59621
rect 69748 -59646 69899 -59621
rect 67242 -60116 67288 -59816
rect 67438 -60116 67484 -59816
rect 67634 -60116 67680 -59816
rect 67851 -59915 67897 -59815
rect 68047 -59915 68093 -59815
rect 68243 -59915 68289 -59815
rect 68439 -59915 68485 -59815
rect 68689 -60327 68735 -59727
rect 68885 -60327 68931 -59727
rect 69308 -60327 69354 -59727
rect 72761 -55586 72807 -55386
rect 72957 -55586 73003 -55386
rect 73153 -55586 73199 -55386
rect 73349 -55586 73395 -55386
rect 73734 -55715 73780 -55415
rect 73930 -55715 73976 -55415
rect 74126 -55715 74172 -55415
rect 74343 -55716 74389 -55616
rect 74539 -55716 74585 -55616
rect 74735 -55716 74781 -55616
rect 74931 -55716 74977 -55616
rect 75013 -56031 75087 -56015
rect 75241 -56031 75351 -55995
rect 75013 -56127 75351 -56031
rect 75013 -56133 75087 -56127
rect 75241 -56145 75351 -56127
rect 72735 -56615 72781 -56315
rect 72931 -56615 72977 -56315
rect 73127 -56615 73173 -56315
rect 73344 -56414 73390 -56314
rect 73540 -56414 73586 -56314
rect 73736 -56414 73782 -56314
rect 73932 -56414 73978 -56314
rect 74182 -56826 74228 -56226
rect 74378 -56826 74424 -56226
rect 74801 -56826 74847 -56226
rect 76174 -56584 76220 -56084
rect 76370 -56584 76416 -56084
rect 76965 -56584 77011 -56084
rect 77095 -56584 77141 -56084
rect 77323 -56384 77369 -56084
rect 77519 -56384 77565 -56084
rect 72753 -59039 72799 -58839
rect 72949 -59039 72995 -58839
rect 73145 -59039 73191 -58839
rect 73341 -59039 73387 -58839
rect 73726 -59168 73772 -58868
rect 73922 -59168 73968 -58868
rect 74118 -59168 74164 -58868
rect 74335 -59169 74381 -59069
rect 74531 -59169 74577 -59069
rect 74727 -59169 74773 -59069
rect 74923 -59169 74969 -59069
rect 73928 -59443 74111 -59402
rect 75231 -59443 75327 -59414
rect 73928 -59525 75327 -59443
rect 73928 -59532 74111 -59525
rect 75231 -59551 75327 -59525
rect 72727 -60068 72773 -59768
rect 72923 -60068 72969 -59768
rect 73119 -60068 73165 -59768
rect 73336 -59867 73382 -59767
rect 73532 -59867 73578 -59767
rect 73728 -59867 73774 -59767
rect 73924 -59867 73970 -59767
rect 74174 -60279 74220 -59679
rect 74370 -60279 74416 -59679
rect 74793 -60279 74839 -59679
rect 76421 -59070 76467 -58870
rect 76617 -59070 76663 -58870
rect 76813 -59070 76859 -58870
rect 77009 -59070 77055 -58870
rect 77394 -59199 77440 -58899
rect 77590 -59199 77636 -58899
rect 77786 -59199 77832 -58899
rect 78003 -59200 78049 -59100
rect 78199 -59200 78245 -59100
rect 78395 -59200 78441 -59100
rect 78591 -59200 78637 -59100
rect 78651 -59465 78742 -59453
rect 78901 -59465 79052 -59438
rect 78651 -59604 79052 -59465
rect 78651 -59616 78742 -59604
rect 78901 -59629 79052 -59604
rect 76395 -60099 76441 -59799
rect 76591 -60099 76637 -59799
rect 76787 -60099 76833 -59799
rect 77004 -59898 77050 -59798
rect 77200 -59898 77246 -59798
rect 77396 -59898 77442 -59798
rect 77592 -59898 77638 -59798
rect 77842 -60310 77888 -59710
rect 78038 -60310 78084 -59710
rect 78461 -60310 78507 -59710
rect 82125 -55548 82171 -55348
rect 82321 -55548 82367 -55348
rect 82517 -55548 82563 -55348
rect 82713 -55548 82759 -55348
rect 83098 -55677 83144 -55377
rect 83294 -55677 83340 -55377
rect 83490 -55677 83536 -55377
rect 83707 -55678 83753 -55578
rect 83903 -55678 83949 -55578
rect 84099 -55678 84145 -55578
rect 84295 -55678 84341 -55578
rect 84377 -55993 84451 -55977
rect 84605 -55993 84715 -55957
rect 84377 -56089 84715 -55993
rect 84377 -56095 84451 -56089
rect 84605 -56107 84715 -56089
rect 82099 -56577 82145 -56277
rect 82295 -56577 82341 -56277
rect 82491 -56577 82537 -56277
rect 82708 -56376 82754 -56276
rect 82904 -56376 82950 -56276
rect 83100 -56376 83146 -56276
rect 83296 -56376 83342 -56276
rect 83546 -56788 83592 -56188
rect 83742 -56788 83788 -56188
rect 84165 -56788 84211 -56188
rect 85538 -56546 85584 -56046
rect 85734 -56546 85780 -56046
rect 86329 -56546 86375 -56046
rect 86459 -56546 86505 -56046
rect 86687 -56346 86733 -56046
rect 86883 -56346 86929 -56046
rect 82117 -59001 82163 -58801
rect 82313 -59001 82359 -58801
rect 82509 -59001 82555 -58801
rect 82705 -59001 82751 -58801
rect 83090 -59130 83136 -58830
rect 83286 -59130 83332 -58830
rect 83482 -59130 83528 -58830
rect 83699 -59131 83745 -59031
rect 83895 -59131 83941 -59031
rect 84091 -59131 84137 -59031
rect 84287 -59131 84333 -59031
rect 83292 -59405 83475 -59364
rect 84595 -59405 84691 -59376
rect 83292 -59487 84691 -59405
rect 83292 -59494 83475 -59487
rect 84595 -59513 84691 -59487
rect 82091 -60030 82137 -59730
rect 82287 -60030 82333 -59730
rect 82483 -60030 82529 -59730
rect 82700 -59829 82746 -59729
rect 82896 -59829 82942 -59729
rect 83092 -59829 83138 -59729
rect 83288 -59829 83334 -59729
rect 83538 -60241 83584 -59641
rect 83734 -60241 83780 -59641
rect 84157 -60241 84203 -59641
rect 85785 -59032 85831 -58832
rect 85981 -59032 86027 -58832
rect 86177 -59032 86223 -58832
rect 86373 -59032 86419 -58832
rect 86758 -59161 86804 -58861
rect 86954 -59161 87000 -58861
rect 87150 -59161 87196 -58861
rect 87367 -59162 87413 -59062
rect 87563 -59162 87609 -59062
rect 87759 -59162 87805 -59062
rect 87955 -59162 88001 -59062
rect 88015 -59427 88106 -59415
rect 88265 -59427 88416 -59400
rect 88015 -59566 88416 -59427
rect 88015 -59578 88106 -59566
rect 88265 -59591 88416 -59566
rect 85759 -60061 85805 -59761
rect 85955 -60061 86001 -59761
rect 86151 -60061 86197 -59761
rect 86368 -59860 86414 -59760
rect 86564 -59860 86610 -59760
rect 86760 -59860 86806 -59760
rect 86956 -59860 87002 -59760
rect 87206 -60272 87252 -59672
rect 87402 -60272 87448 -59672
rect 87825 -60272 87871 -59672
rect 90119 -54278 92731 -7667
rect 26730 -62429 82728 -62184
<< obsm1 >>
rect -12466 121009 -12123 121054
rect -12466 120725 -1630 121009
rect -12466 120695 -12123 120725
rect -12170 120137 -12098 120171
rect -12318 120072 -12098 120137
rect -12651 119752 -12351 119798
rect -12651 119314 -12351 119360
rect -12318 119117 -12253 120072
rect -12170 120066 -12098 120072
rect -12039 119835 -11439 119881
rect -10773 119815 -10727 120014
rect -10929 119769 -10727 119815
rect -10773 119717 -10727 119769
rect -8615 120289 -8553 120302
rect -8615 120070 -6144 120289
rect -10775 119671 -10598 119717
rect -12039 119623 -11439 119669
rect -10775 119619 -10727 119671
rect -10929 119573 -10727 119619
rect -12039 119525 -11439 119571
rect -10775 119521 -10727 119573
rect -10775 119475 -10598 119521
rect -12039 119427 -11439 119473
rect -10773 119423 -10727 119475
rect -10929 119377 -10727 119423
rect -12039 119216 -11439 119262
rect -10391 119062 -10008 119108
rect -11729 118816 -11683 119015
rect -10928 118964 -10091 119010
rect -10055 118912 -10008 119062
rect -10391 118866 -10008 118912
rect -11729 118770 -11527 118816
rect -11729 118718 -11683 118770
rect -10928 118768 -10628 118814
rect -11858 118672 -11681 118718
rect -11729 118620 -11681 118672
rect -10582 118654 -10524 118733
rect -10055 118716 -10008 118866
rect -9109 118795 -8809 118841
rect -8615 118746 -8553 120070
rect -10391 118670 -10008 118716
rect -8624 118680 -8541 118746
rect -8113 118697 -7813 118743
rect -10092 118669 -10008 118670
rect -11729 118574 -11527 118620
rect -10582 118600 -10415 118654
rect -10582 118574 -10524 118600
rect -11729 118522 -11681 118574
rect -11858 118476 -11681 118522
rect -11729 118424 -11683 118476
rect -11729 118378 -11527 118424
rect -10543 118233 -10497 118432
rect -10469 118380 -10415 118600
rect -9109 118567 -8609 118613
rect -9109 118469 -8609 118515
rect -8538 118508 -8400 118562
rect -10469 118326 -10071 118380
rect -10799 118187 -10497 118233
rect -10543 118135 -10497 118187
rect -12448 118063 -12065 118109
rect -10545 118089 -10269 118135
rect -12448 117913 -12401 118063
rect -10545 118037 -10497 118089
rect -12365 117965 -11528 118011
rect -10799 117991 -10497 118037
rect -10545 117939 -10497 117991
rect -12448 117867 -12065 117913
rect -10545 117893 -10269 117939
rect -12448 117717 -12401 117867
rect -10543 117841 -10497 117893
rect -11828 117769 -11528 117815
rect -10799 117795 -10497 117841
rect -12448 117671 -12065 117717
rect -12448 117670 -12364 117671
rect -10565 117613 -10415 117639
rect -12023 117559 -10415 117613
rect -12023 117416 -11969 117559
rect -10565 117509 -10415 117559
rect -10125 117368 -10071 118326
rect -8517 118261 -8473 118508
rect -8313 118469 -7813 118515
rect -9109 118143 -8609 118189
rect -8523 118123 -8469 118261
rect -8313 118143 -7813 118189
rect -9109 118018 -8609 118064
rect -9109 117920 -8609 117966
rect -9109 117548 -8809 117594
rect -8517 117455 -8473 118123
rect -8313 118013 -7813 118059
rect -8313 117915 -7813 117961
rect -8313 117817 -7813 117863
rect -8313 117548 -7813 117594
rect -10131 117271 -10065 117368
rect -8523 117317 -8469 117455
rect -8860 117247 -8769 117259
rect -9572 117168 -8769 117247
rect -12139 116469 -12067 116503
rect -12287 116404 -12067 116469
rect -12620 116084 -12320 116130
rect -12620 115646 -12320 115692
rect -12287 115449 -12222 116404
rect -12139 116398 -12067 116404
rect -12008 116167 -11408 116213
rect -12008 115955 -11408 116001
rect -12008 115857 -11408 115903
rect -12008 115759 -11408 115805
rect -12008 115548 -11408 115594
rect -10024 116747 -9927 116758
rect -9572 116747 -9493 117168
rect -8860 117156 -8769 117168
rect -10024 116668 -9493 116747
rect -10024 116642 -9927 116668
rect -8686 116477 -8614 116511
rect -10742 116147 -10696 116346
rect -10898 116101 -10696 116147
rect -10742 116049 -10696 116101
rect -8834 116412 -8614 116477
rect -9167 116092 -8867 116138
rect -10744 116003 -10567 116049
rect -10744 115951 -10696 116003
rect -10898 115905 -10696 115951
rect -10744 115853 -10696 115905
rect -10744 115807 -10567 115853
rect -10742 115755 -10696 115807
rect -10898 115709 -10696 115755
rect -9167 115654 -8867 115700
rect -8834 115457 -8769 116412
rect -8686 116406 -8614 116412
rect -8555 116175 -7955 116221
rect -7289 116155 -7243 116354
rect -7445 116109 -7243 116155
rect -7289 116057 -7243 116109
rect -7291 116011 -7114 116057
rect -8555 115963 -7955 116009
rect -7291 115959 -7243 116011
rect -7445 115913 -7243 115959
rect -8555 115865 -7955 115911
rect -7291 115861 -7243 115913
rect -7291 115815 -7114 115861
rect -8555 115767 -7955 115813
rect -7289 115763 -7243 115815
rect -7445 115717 -7243 115763
rect -8555 115556 -7955 115602
rect -10360 115394 -9977 115440
rect -6907 115402 -6524 115448
rect -11698 115148 -11652 115347
rect -10897 115296 -10060 115342
rect -10024 115244 -9977 115394
rect -10360 115198 -9977 115244
rect -11698 115102 -11496 115148
rect -11698 115050 -11652 115102
rect -10897 115100 -10597 115146
rect -11827 115004 -11650 115050
rect -11698 114952 -11650 115004
rect -10551 114986 -10493 115065
rect -10024 115048 -9977 115198
rect -8245 115156 -8199 115355
rect -7444 115304 -6607 115350
rect -6571 115252 -6524 115402
rect -6907 115206 -6524 115252
rect -8245 115110 -8043 115156
rect -8245 115058 -8199 115110
rect -7444 115108 -7144 115154
rect -10360 115002 -9977 115048
rect -8374 115012 -8197 115058
rect -10061 115001 -9977 115002
rect -11698 114906 -11496 114952
rect -10551 114932 -10384 114986
rect -8245 114960 -8197 115012
rect -7098 114994 -7040 115073
rect -6571 115056 -6524 115206
rect -6907 115010 -6524 115056
rect -6608 115009 -6524 115010
rect -10551 114906 -10493 114932
rect -11698 114854 -11650 114906
rect -11827 114808 -11650 114854
rect -11698 114756 -11652 114808
rect -11698 114710 -11496 114756
rect -14622 76452 -14337 114640
rect -17317 76167 -14337 76452
rect -17317 57173 -17032 76167
rect -14701 75156 -14324 75216
rect -16789 74856 -14324 75156
rect -16789 58539 -16489 74856
rect -14701 74847 -14324 74856
rect -13782 75207 -13601 114640
rect -10512 114565 -10466 114764
rect -10438 114712 -10384 114932
rect -8245 114914 -8043 114960
rect -7098 114940 -6931 114994
rect -7098 114914 -7040 114940
rect -8245 114862 -8197 114914
rect -8374 114816 -8197 114862
rect -8245 114764 -8199 114816
rect -8245 114718 -8043 114764
rect -10438 114658 -10040 114712
rect -10768 114519 -10466 114565
rect -10512 114467 -10466 114519
rect -12417 114395 -12034 114441
rect -10514 114421 -10238 114467
rect -12417 114245 -12370 114395
rect -10514 114369 -10466 114421
rect -12334 114297 -11497 114343
rect -10768 114323 -10466 114369
rect -10514 114271 -10466 114323
rect -12417 114199 -12034 114245
rect -10514 114225 -10238 114271
rect -12417 114049 -12370 114199
rect -10512 114173 -10466 114225
rect -11797 114101 -11497 114147
rect -10768 114127 -10466 114173
rect -12417 114003 -12034 114049
rect -12417 114002 -12333 114003
rect -10534 113945 -10384 113971
rect -11992 113891 -10384 113945
rect -11992 113748 -11938 113891
rect -10534 113841 -10384 113891
rect -10094 113549 -10040 114658
rect -7059 114573 -7013 114772
rect -6985 114720 -6931 114940
rect -6985 114666 -6587 114720
rect -7315 114527 -7013 114573
rect -7059 114475 -7013 114527
rect -8964 114403 -8581 114449
rect -7061 114429 -6785 114475
rect -8964 114253 -8917 114403
rect -7061 114377 -7013 114429
rect -8881 114305 -8044 114351
rect -7315 114331 -7013 114377
rect -7061 114279 -7013 114331
rect -8964 114207 -8581 114253
rect -7061 114233 -6785 114279
rect -8964 114057 -8917 114207
rect -7059 114181 -7013 114233
rect -8344 114109 -8044 114155
rect -7315 114135 -7013 114181
rect -8964 114011 -8581 114057
rect -8964 114010 -8880 114011
rect -7081 113953 -6931 113979
rect -8539 113899 -6931 113953
rect -8539 113756 -8485 113899
rect -7081 113849 -6931 113899
rect -10220 111989 -10001 113549
rect -6641 113518 -6587 114666
rect -6745 113223 -6472 113518
rect -6363 111989 -6144 120070
rect -10220 111770 -6144 111989
rect -12491 111194 -2536 111505
rect -12208 110773 -12136 110807
rect -12356 110708 -12136 110773
rect -12689 110388 -12389 110434
rect -12689 109950 -12389 109996
rect -12356 109753 -12291 110708
rect -12208 110702 -12136 110708
rect -12077 110471 -11477 110517
rect -10811 110451 -10765 110650
rect -10967 110405 -10765 110451
rect -10811 110353 -10765 110405
rect -8653 110933 -8591 110938
rect -8653 110626 -6145 110933
rect -10813 110307 -10636 110353
rect -12077 110259 -11477 110305
rect -10813 110255 -10765 110307
rect -10967 110209 -10765 110255
rect -12077 110161 -11477 110207
rect -10813 110157 -10765 110209
rect -10813 110111 -10636 110157
rect -12077 110063 -11477 110109
rect -10811 110059 -10765 110111
rect -10967 110013 -10765 110059
rect -12077 109852 -11477 109898
rect -10429 109698 -10046 109744
rect -11767 109452 -11721 109651
rect -10966 109600 -10129 109646
rect -10093 109548 -10046 109698
rect -10429 109502 -10046 109548
rect -11767 109406 -11565 109452
rect -11767 109354 -11721 109406
rect -10966 109404 -10666 109450
rect -11896 109308 -11719 109354
rect -11767 109256 -11719 109308
rect -10620 109290 -10562 109369
rect -10093 109352 -10046 109502
rect -9147 109431 -8847 109477
rect -8653 109382 -8591 110626
rect -10429 109306 -10046 109352
rect -8662 109316 -8579 109382
rect -8151 109333 -7851 109379
rect -10130 109305 -10046 109306
rect -11767 109210 -11565 109256
rect -10620 109236 -10453 109290
rect -10620 109210 -10562 109236
rect -11767 109158 -11719 109210
rect -11896 109112 -11719 109158
rect -11767 109060 -11721 109112
rect -11767 109014 -11565 109060
rect -10581 108869 -10535 109068
rect -10507 109016 -10453 109236
rect -9147 109203 -8647 109249
rect -9147 109105 -8647 109151
rect -8576 109144 -8438 109198
rect -10507 108962 -10109 109016
rect -10837 108823 -10535 108869
rect -10581 108771 -10535 108823
rect -12486 108699 -12103 108745
rect -10583 108725 -10307 108771
rect -12486 108549 -12439 108699
rect -10583 108673 -10535 108725
rect -12403 108601 -11566 108647
rect -10837 108627 -10535 108673
rect -10583 108575 -10535 108627
rect -12486 108503 -12103 108549
rect -10583 108529 -10307 108575
rect -12486 108353 -12439 108503
rect -10581 108477 -10535 108529
rect -11866 108405 -11566 108451
rect -10837 108431 -10535 108477
rect -12486 108307 -12103 108353
rect -12486 108306 -12402 108307
rect -10603 108249 -10453 108275
rect -12061 108195 -10453 108249
rect -12061 108052 -12007 108195
rect -10603 108145 -10453 108195
rect -10163 108004 -10109 108962
rect -8555 108897 -8511 109144
rect -8351 109105 -7851 109151
rect -9147 108779 -8647 108825
rect -8561 108759 -8507 108897
rect -8351 108779 -7851 108825
rect -9147 108654 -8647 108700
rect -9147 108556 -8647 108602
rect -9147 108184 -8847 108230
rect -8555 108091 -8511 108759
rect -8351 108649 -7851 108695
rect -8351 108551 -7851 108597
rect -8351 108453 -7851 108499
rect -8351 108184 -7851 108230
rect -10169 107907 -10103 108004
rect -8561 107953 -8507 108091
rect -8898 107883 -8807 107895
rect -9610 107804 -8807 107883
rect -12177 107105 -12105 107139
rect -12325 107040 -12105 107105
rect -12658 106720 -12358 106766
rect -12658 106282 -12358 106328
rect -12325 106085 -12260 107040
rect -12177 107034 -12105 107040
rect -12046 106803 -11446 106849
rect -12046 106591 -11446 106637
rect -12046 106493 -11446 106539
rect -12046 106395 -11446 106441
rect -12046 106184 -11446 106230
rect -10062 107383 -9965 107394
rect -9610 107383 -9531 107804
rect -8898 107792 -8807 107804
rect -10062 107304 -9531 107383
rect -10062 107278 -9965 107304
rect -8724 107113 -8652 107147
rect -10780 106783 -10734 106982
rect -10936 106737 -10734 106783
rect -10780 106685 -10734 106737
rect -8872 107048 -8652 107113
rect -9205 106728 -8905 106774
rect -10782 106639 -10605 106685
rect -10782 106587 -10734 106639
rect -10936 106541 -10734 106587
rect -10782 106489 -10734 106541
rect -10782 106443 -10605 106489
rect -10780 106391 -10734 106443
rect -10936 106345 -10734 106391
rect -9205 106290 -8905 106336
rect -8872 106093 -8807 107048
rect -8724 107042 -8652 107048
rect -8593 106811 -7993 106857
rect -7327 106791 -7281 106990
rect -7483 106745 -7281 106791
rect -7327 106693 -7281 106745
rect -7329 106647 -7152 106693
rect -8593 106599 -7993 106645
rect -7329 106595 -7281 106647
rect -7483 106549 -7281 106595
rect -8593 106501 -7993 106547
rect -7329 106497 -7281 106549
rect -7329 106451 -7152 106497
rect -8593 106403 -7993 106449
rect -7327 106399 -7281 106451
rect -7483 106353 -7281 106399
rect -8593 106192 -7993 106238
rect -10398 106030 -10015 106076
rect -6945 106038 -6562 106084
rect -11736 105784 -11690 105983
rect -10935 105932 -10098 105978
rect -10062 105880 -10015 106030
rect -10398 105834 -10015 105880
rect -11736 105738 -11534 105784
rect -11736 105686 -11690 105738
rect -10935 105736 -10635 105782
rect -11865 105640 -11688 105686
rect -11736 105588 -11688 105640
rect -10589 105622 -10531 105701
rect -10062 105684 -10015 105834
rect -8283 105792 -8237 105991
rect -7482 105940 -6645 105986
rect -6609 105888 -6562 106038
rect -6945 105842 -6562 105888
rect -8283 105746 -8081 105792
rect -8283 105694 -8237 105746
rect -7482 105744 -7182 105790
rect -10398 105638 -10015 105684
rect -8412 105648 -8235 105694
rect -10099 105637 -10015 105638
rect -11736 105542 -11534 105588
rect -10589 105568 -10422 105622
rect -8283 105596 -8235 105648
rect -7136 105630 -7078 105709
rect -6609 105692 -6562 105842
rect -6945 105646 -6562 105692
rect -6646 105645 -6562 105646
rect -10589 105542 -10531 105568
rect -11736 105490 -11688 105542
rect -11865 105444 -11688 105490
rect -11736 105392 -11690 105444
rect -11736 105346 -11534 105392
rect -10550 105201 -10504 105400
rect -10476 105348 -10422 105568
rect -8283 105550 -8081 105596
rect -7136 105576 -6969 105630
rect -7136 105550 -7078 105576
rect -8283 105498 -8235 105550
rect -8412 105452 -8235 105498
rect -8283 105400 -8237 105452
rect -8283 105354 -8081 105400
rect -10476 105294 -10078 105348
rect -10806 105155 -10504 105201
rect -10550 105103 -10504 105155
rect -12455 105031 -12072 105077
rect -10552 105057 -10276 105103
rect -12455 104881 -12408 105031
rect -10552 105005 -10504 105057
rect -12372 104933 -11535 104979
rect -10806 104959 -10504 105005
rect -10552 104907 -10504 104959
rect -12455 104835 -12072 104881
rect -10552 104861 -10276 104907
rect -12455 104685 -12408 104835
rect -10550 104809 -10504 104861
rect -11835 104737 -11535 104783
rect -10806 104763 -10504 104809
rect -12455 104639 -12072 104685
rect -12455 104638 -12371 104639
rect -10572 104581 -10422 104607
rect -12030 104527 -10422 104581
rect -12030 104384 -11976 104527
rect -10572 104477 -10422 104527
rect -10132 104035 -10078 105294
rect -7097 105209 -7051 105408
rect -7023 105356 -6969 105576
rect -7023 105302 -6625 105356
rect -7353 105163 -7051 105209
rect -7097 105111 -7051 105163
rect -9002 105039 -8619 105085
rect -7099 105065 -6823 105111
rect -9002 104889 -8955 105039
rect -7099 105013 -7051 105065
rect -8919 104941 -8082 104987
rect -7353 104967 -7051 105013
rect -7099 104915 -7051 104967
rect -9002 104843 -8619 104889
rect -7099 104869 -6823 104915
rect -9002 104693 -8955 104843
rect -7097 104817 -7051 104869
rect -8382 104745 -8082 104791
rect -7353 104771 -7051 104817
rect -9002 104647 -8619 104693
rect -9002 104646 -8918 104647
rect -7119 104589 -6969 104615
rect -8577 104535 -6969 104589
rect -8577 104392 -8523 104535
rect -7119 104485 -6969 104535
rect -6679 104236 -6625 105302
rect -10195 102845 -9895 104035
rect -6774 103968 -6534 104236
rect -6445 102845 -6145 110626
rect -10195 102545 -6145 102845
rect -12471 102237 -12167 102279
rect -6770 102237 -6479 102318
rect -12471 102060 -3120 102237
rect -12471 102018 -12167 102060
rect -6770 101980 -6479 102060
rect -12225 101620 -12153 101654
rect -12373 101555 -12153 101620
rect -12706 101235 -12406 101281
rect -12706 100797 -12406 100843
rect -12373 100600 -12308 101555
rect -12225 101549 -12153 101555
rect -12094 101318 -11494 101364
rect -10828 101298 -10782 101497
rect -10984 101252 -10782 101298
rect -10828 101200 -10782 101252
rect -8670 101743 -8608 101785
rect -8670 101505 -6199 101743
rect -10830 101154 -10653 101200
rect -12094 101106 -11494 101152
rect -10830 101102 -10782 101154
rect -10984 101056 -10782 101102
rect -12094 101008 -11494 101054
rect -10830 101004 -10782 101056
rect -10830 100958 -10653 101004
rect -12094 100910 -11494 100956
rect -10828 100906 -10782 100958
rect -10984 100860 -10782 100906
rect -12094 100699 -11494 100745
rect -10446 100545 -10063 100591
rect -11784 100299 -11738 100498
rect -10983 100447 -10146 100493
rect -10110 100395 -10063 100545
rect -10446 100349 -10063 100395
rect -11784 100253 -11582 100299
rect -11784 100201 -11738 100253
rect -10983 100251 -10683 100297
rect -11913 100155 -11736 100201
rect -11784 100103 -11736 100155
rect -10637 100137 -10579 100216
rect -10110 100199 -10063 100349
rect -9164 100278 -8864 100324
rect -8670 100229 -8608 101505
rect -10446 100153 -10063 100199
rect -8679 100163 -8596 100229
rect -8168 100180 -7868 100226
rect -10147 100152 -10063 100153
rect -11784 100057 -11582 100103
rect -10637 100083 -10470 100137
rect -10637 100057 -10579 100083
rect -11784 100005 -11736 100057
rect -11913 99959 -11736 100005
rect -11784 99907 -11738 99959
rect -11784 99861 -11582 99907
rect -10598 99716 -10552 99915
rect -10524 99863 -10470 100083
rect -9164 100050 -8664 100096
rect -9164 99952 -8664 99998
rect -8593 99991 -8455 100045
rect -10524 99809 -10126 99863
rect -10854 99670 -10552 99716
rect -10598 99618 -10552 99670
rect -12503 99546 -12120 99592
rect -10600 99572 -10324 99618
rect -12503 99396 -12456 99546
rect -10600 99520 -10552 99572
rect -12420 99448 -11583 99494
rect -10854 99474 -10552 99520
rect -10600 99422 -10552 99474
rect -12503 99350 -12120 99396
rect -10600 99376 -10324 99422
rect -12503 99200 -12456 99350
rect -10598 99324 -10552 99376
rect -11883 99252 -11583 99298
rect -10854 99278 -10552 99324
rect -12503 99154 -12120 99200
rect -12503 99153 -12419 99154
rect -10620 99096 -10470 99122
rect -12078 99042 -10470 99096
rect -12078 98899 -12024 99042
rect -10620 98992 -10470 99042
rect -10180 98851 -10126 99809
rect -8572 99744 -8528 99991
rect -8368 99952 -7868 99998
rect -9164 99626 -8664 99672
rect -8578 99606 -8524 99744
rect -8368 99626 -7868 99672
rect -9164 99501 -8664 99547
rect -9164 99403 -8664 99449
rect -9164 99031 -8864 99077
rect -8572 98938 -8528 99606
rect -8368 99496 -7868 99542
rect -8368 99398 -7868 99444
rect -8368 99300 -7868 99346
rect -8368 99031 -7868 99077
rect -10186 98754 -10120 98851
rect -8578 98800 -8524 98938
rect -8915 98730 -8824 98742
rect -9627 98651 -8824 98730
rect -12194 97952 -12122 97986
rect -12342 97887 -12122 97952
rect -12675 97567 -12375 97613
rect -12675 97129 -12375 97175
rect -12342 96932 -12277 97887
rect -12194 97881 -12122 97887
rect -12063 97650 -11463 97696
rect -12063 97438 -11463 97484
rect -12063 97340 -11463 97386
rect -12063 97242 -11463 97288
rect -12063 97031 -11463 97077
rect -10079 98230 -9982 98241
rect -9627 98230 -9548 98651
rect -8915 98639 -8824 98651
rect -10079 98151 -9548 98230
rect -10079 98125 -9982 98151
rect -8741 97960 -8669 97994
rect -10797 97630 -10751 97829
rect -10953 97584 -10751 97630
rect -10797 97532 -10751 97584
rect -8889 97895 -8669 97960
rect -9222 97575 -8922 97621
rect -10799 97486 -10622 97532
rect -10799 97434 -10751 97486
rect -10953 97388 -10751 97434
rect -10799 97336 -10751 97388
rect -10799 97290 -10622 97336
rect -10797 97238 -10751 97290
rect -10953 97192 -10751 97238
rect -9222 97137 -8922 97183
rect -8889 96940 -8824 97895
rect -8741 97889 -8669 97895
rect -8610 97658 -8010 97704
rect -7344 97638 -7298 97837
rect -7500 97592 -7298 97638
rect -7344 97540 -7298 97592
rect -7346 97494 -7169 97540
rect -8610 97446 -8010 97492
rect -7346 97442 -7298 97494
rect -7500 97396 -7298 97442
rect -8610 97348 -8010 97394
rect -7346 97344 -7298 97396
rect -7346 97298 -7169 97344
rect -8610 97250 -8010 97296
rect -7344 97246 -7298 97298
rect -7500 97200 -7298 97246
rect -8610 97039 -8010 97085
rect -10415 96877 -10032 96923
rect -6962 96885 -6579 96931
rect -11753 96631 -11707 96830
rect -10952 96779 -10115 96825
rect -10079 96727 -10032 96877
rect -10415 96681 -10032 96727
rect -11753 96585 -11551 96631
rect -11753 96533 -11707 96585
rect -10952 96583 -10652 96629
rect -11882 96487 -11705 96533
rect -11753 96435 -11705 96487
rect -10606 96469 -10548 96548
rect -10079 96531 -10032 96681
rect -8300 96639 -8254 96838
rect -7499 96787 -6662 96833
rect -6626 96735 -6579 96885
rect -6962 96689 -6579 96735
rect -8300 96593 -8098 96639
rect -8300 96541 -8254 96593
rect -7499 96591 -7199 96637
rect -10415 96485 -10032 96531
rect -8429 96495 -8252 96541
rect -10116 96484 -10032 96485
rect -11753 96389 -11551 96435
rect -10606 96415 -10439 96469
rect -8300 96443 -8252 96495
rect -7153 96477 -7095 96556
rect -6626 96539 -6579 96689
rect -6962 96493 -6579 96539
rect -6663 96492 -6579 96493
rect -10606 96389 -10548 96415
rect -11753 96337 -11705 96389
rect -11882 96291 -11705 96337
rect -11753 96239 -11707 96291
rect -11753 96193 -11551 96239
rect -10567 96048 -10521 96247
rect -10493 96195 -10439 96415
rect -8300 96397 -8098 96443
rect -7153 96423 -6986 96477
rect -7153 96397 -7095 96423
rect -8300 96345 -8252 96397
rect -8429 96299 -8252 96345
rect -8300 96247 -8254 96299
rect -8300 96201 -8098 96247
rect -10493 96141 -10095 96195
rect -10823 96002 -10521 96048
rect -10567 95950 -10521 96002
rect -12472 95878 -12089 95924
rect -10569 95904 -10293 95950
rect -12472 95728 -12425 95878
rect -10569 95852 -10521 95904
rect -12389 95780 -11552 95826
rect -10823 95806 -10521 95852
rect -10569 95754 -10521 95806
rect -12472 95682 -12089 95728
rect -10569 95708 -10293 95754
rect -12472 95532 -12425 95682
rect -10567 95656 -10521 95708
rect -11852 95584 -11552 95630
rect -10823 95610 -10521 95656
rect -12472 95486 -12089 95532
rect -12472 95485 -12388 95486
rect -10589 95428 -10439 95454
rect -12047 95374 -10439 95428
rect -12047 95231 -11993 95374
rect -10589 95324 -10439 95374
rect -10149 94895 -10095 96141
rect -7114 96056 -7068 96255
rect -7040 96203 -6986 96423
rect -7040 96149 -6642 96203
rect -7370 96010 -7068 96056
rect -7114 95958 -7068 96010
rect -9019 95886 -8636 95932
rect -7116 95912 -6840 95958
rect -9019 95736 -8972 95886
rect -7116 95860 -7068 95912
rect -8936 95788 -8099 95834
rect -7370 95814 -7068 95860
rect -7116 95762 -7068 95814
rect -9019 95690 -8636 95736
rect -7116 95716 -6840 95762
rect -9019 95540 -8972 95690
rect -7114 95664 -7068 95716
rect -8399 95592 -8099 95638
rect -7370 95618 -7068 95664
rect -9019 95494 -8636 95540
rect -9019 95493 -8935 95494
rect -7136 95436 -6986 95462
rect -8594 95382 -6986 95436
rect -8594 95239 -8540 95382
rect -7136 95332 -6986 95382
rect -6696 95055 -6642 96149
rect -10199 93997 -9961 94895
rect -6771 94805 -6542 95055
rect -6437 93997 -6199 101505
rect -10199 93759 -6199 93997
rect -12524 93528 -12225 93545
rect -6788 93528 -6474 93580
rect -12524 93307 -3635 93528
rect -12524 93253 -12225 93307
rect -6788 93204 -6474 93307
rect -12291 92866 -12219 92900
rect -12439 92801 -12219 92866
rect -12772 92481 -12472 92527
rect -12772 92043 -12472 92089
rect -12439 91846 -12374 92801
rect -12291 92795 -12219 92801
rect -12160 92564 -11560 92610
rect -10894 92544 -10848 92743
rect -11050 92498 -10848 92544
rect -10894 92446 -10848 92498
rect -8736 92956 -8674 93031
rect -8736 92697 -6158 92956
rect -10896 92400 -10719 92446
rect -12160 92352 -11560 92398
rect -10896 92348 -10848 92400
rect -11050 92302 -10848 92348
rect -12160 92254 -11560 92300
rect -10896 92250 -10848 92302
rect -10896 92204 -10719 92250
rect -12160 92156 -11560 92202
rect -10894 92152 -10848 92204
rect -11050 92106 -10848 92152
rect -12160 91945 -11560 91991
rect -10512 91791 -10129 91837
rect -11850 91545 -11804 91744
rect -11049 91693 -10212 91739
rect -10176 91641 -10129 91791
rect -10512 91595 -10129 91641
rect -11850 91499 -11648 91545
rect -11850 91447 -11804 91499
rect -11049 91497 -10749 91543
rect -11979 91401 -11802 91447
rect -11850 91349 -11802 91401
rect -10703 91383 -10645 91462
rect -10176 91445 -10129 91595
rect -9230 91524 -8930 91570
rect -8736 91475 -8674 92697
rect -10512 91399 -10129 91445
rect -8745 91409 -8662 91475
rect -8234 91426 -7934 91472
rect -10213 91398 -10129 91399
rect -11850 91303 -11648 91349
rect -10703 91329 -10536 91383
rect -10703 91303 -10645 91329
rect -11850 91251 -11802 91303
rect -11979 91205 -11802 91251
rect -11850 91153 -11804 91205
rect -11850 91107 -11648 91153
rect -10664 90962 -10618 91161
rect -10590 91109 -10536 91329
rect -9230 91296 -8730 91342
rect -9230 91198 -8730 91244
rect -8659 91237 -8521 91291
rect -10590 91055 -10192 91109
rect -10920 90916 -10618 90962
rect -10664 90864 -10618 90916
rect -12569 90792 -12186 90838
rect -10666 90818 -10390 90864
rect -12569 90642 -12522 90792
rect -10666 90766 -10618 90818
rect -12486 90694 -11649 90740
rect -10920 90720 -10618 90766
rect -10666 90668 -10618 90720
rect -12569 90596 -12186 90642
rect -10666 90622 -10390 90668
rect -12569 90446 -12522 90596
rect -10664 90570 -10618 90622
rect -11949 90498 -11649 90544
rect -10920 90524 -10618 90570
rect -12569 90400 -12186 90446
rect -12569 90399 -12485 90400
rect -10686 90342 -10536 90368
rect -12144 90288 -10536 90342
rect -12144 90145 -12090 90288
rect -10686 90238 -10536 90288
rect -10246 90097 -10192 91055
rect -8638 90990 -8594 91237
rect -8434 91198 -7934 91244
rect -9230 90872 -8730 90918
rect -8644 90852 -8590 90990
rect -8434 90872 -7934 90918
rect -9230 90747 -8730 90793
rect -9230 90649 -8730 90695
rect -9230 90277 -8930 90323
rect -8638 90184 -8594 90852
rect -8434 90742 -7934 90788
rect -8434 90644 -7934 90690
rect -8434 90546 -7934 90592
rect -8434 90277 -7934 90323
rect -10252 90000 -10186 90097
rect -8644 90046 -8590 90184
rect -8981 89976 -8890 89988
rect -9693 89897 -8890 89976
rect -12260 89198 -12188 89232
rect -12408 89133 -12188 89198
rect -12741 88813 -12441 88859
rect -12741 88375 -12441 88421
rect -12408 88178 -12343 89133
rect -12260 89127 -12188 89133
rect -12129 88896 -11529 88942
rect -12129 88684 -11529 88730
rect -12129 88586 -11529 88632
rect -12129 88488 -11529 88534
rect -12129 88277 -11529 88323
rect -10145 89476 -10048 89487
rect -9693 89476 -9614 89897
rect -8981 89885 -8890 89897
rect -10145 89397 -9614 89476
rect -10145 89371 -10048 89397
rect -8807 89206 -8735 89240
rect -10863 88876 -10817 89075
rect -11019 88830 -10817 88876
rect -10863 88778 -10817 88830
rect -8955 89141 -8735 89206
rect -9288 88821 -8988 88867
rect -10865 88732 -10688 88778
rect -10865 88680 -10817 88732
rect -11019 88634 -10817 88680
rect -10865 88582 -10817 88634
rect -10865 88536 -10688 88582
rect -10863 88484 -10817 88536
rect -11019 88438 -10817 88484
rect -9288 88383 -8988 88429
rect -8955 88186 -8890 89141
rect -8807 89135 -8735 89141
rect -8676 88904 -8076 88950
rect -7410 88884 -7364 89083
rect -7566 88838 -7364 88884
rect -7410 88786 -7364 88838
rect -7412 88740 -7235 88786
rect -8676 88692 -8076 88738
rect -7412 88688 -7364 88740
rect -7566 88642 -7364 88688
rect -8676 88594 -8076 88640
rect -7412 88590 -7364 88642
rect -7412 88544 -7235 88590
rect -8676 88496 -8076 88542
rect -7410 88492 -7364 88544
rect -7566 88446 -7364 88492
rect -8676 88285 -8076 88331
rect -10481 88123 -10098 88169
rect -7028 88131 -6645 88177
rect -11819 87877 -11773 88076
rect -11018 88025 -10181 88071
rect -10145 87973 -10098 88123
rect -10481 87927 -10098 87973
rect -11819 87831 -11617 87877
rect -11819 87779 -11773 87831
rect -11018 87829 -10718 87875
rect -11948 87733 -11771 87779
rect -11819 87681 -11771 87733
rect -10672 87715 -10614 87794
rect -10145 87777 -10098 87927
rect -8366 87885 -8320 88084
rect -7565 88033 -6728 88079
rect -6692 87981 -6645 88131
rect -7028 87935 -6645 87981
rect -8366 87839 -8164 87885
rect -8366 87787 -8320 87839
rect -7565 87837 -7265 87883
rect -10481 87731 -10098 87777
rect -8495 87741 -8318 87787
rect -10182 87730 -10098 87731
rect -11819 87635 -11617 87681
rect -10672 87661 -10505 87715
rect -8366 87689 -8318 87741
rect -7219 87723 -7161 87802
rect -6692 87785 -6645 87935
rect -7028 87739 -6645 87785
rect -6729 87738 -6645 87739
rect -10672 87635 -10614 87661
rect -11819 87583 -11771 87635
rect -11948 87537 -11771 87583
rect -11819 87485 -11773 87537
rect -11819 87439 -11617 87485
rect -10633 87294 -10587 87493
rect -10559 87441 -10505 87661
rect -8366 87643 -8164 87689
rect -7219 87669 -7052 87723
rect -7219 87643 -7161 87669
rect -8366 87591 -8318 87643
rect -8495 87545 -8318 87591
rect -8366 87493 -8320 87545
rect -8366 87447 -8164 87493
rect -10559 87387 -10161 87441
rect -10889 87248 -10587 87294
rect -10633 87196 -10587 87248
rect -12538 87124 -12155 87170
rect -10635 87150 -10359 87196
rect -12538 86974 -12491 87124
rect -10635 87098 -10587 87150
rect -12455 87026 -11618 87072
rect -10889 87052 -10587 87098
rect -10635 87000 -10587 87052
rect -12538 86928 -12155 86974
rect -10635 86954 -10359 87000
rect -12538 86778 -12491 86928
rect -10633 86902 -10587 86954
rect -11918 86830 -11618 86876
rect -10889 86856 -10587 86902
rect -12538 86732 -12155 86778
rect -12538 86731 -12454 86732
rect -10655 86674 -10505 86700
rect -12113 86620 -10505 86674
rect -12113 86477 -12059 86620
rect -10655 86570 -10505 86620
rect -10215 86178 -10161 87387
rect -7180 87302 -7134 87501
rect -7106 87449 -7052 87669
rect -7106 87395 -6708 87449
rect -7436 87256 -7134 87302
rect -7180 87204 -7134 87256
rect -9085 87132 -8702 87178
rect -7182 87158 -6906 87204
rect -9085 86982 -9038 87132
rect -7182 87106 -7134 87158
rect -9002 87034 -8165 87080
rect -7436 87060 -7134 87106
rect -7182 87008 -7134 87060
rect -9085 86936 -8702 86982
rect -7182 86962 -6906 87008
rect -9085 86786 -9038 86936
rect -7180 86910 -7134 86962
rect -8465 86838 -8165 86884
rect -7436 86864 -7134 86910
rect -9085 86740 -8702 86786
rect -9085 86739 -9001 86740
rect -7202 86682 -7052 86708
rect -8660 86628 -7052 86682
rect -8660 86485 -8606 86628
rect -7202 86578 -7052 86628
rect -10280 85229 -10021 86178
rect -6762 86012 -6708 87395
rect -6832 85766 -6612 86012
rect -6417 85229 -6158 92697
rect -10280 84970 -6158 85229
rect -12587 84339 -12087 84389
rect -12587 84113 -4187 84339
rect -12587 84091 -12087 84113
rect -12325 83668 -12253 83702
rect -12473 83603 -12253 83668
rect -12806 83283 -12506 83329
rect -12806 82845 -12506 82891
rect -12473 82648 -12408 83603
rect -12325 83597 -12253 83603
rect -12194 83366 -11594 83412
rect -10928 83346 -10882 83545
rect -11084 83300 -10882 83346
rect -10928 83248 -10882 83300
rect -8770 83652 -8708 83833
rect -8770 83450 -6150 83652
rect -10930 83202 -10753 83248
rect -12194 83154 -11594 83200
rect -10930 83150 -10882 83202
rect -11084 83104 -10882 83150
rect -12194 83056 -11594 83102
rect -10930 83052 -10882 83104
rect -10930 83006 -10753 83052
rect -12194 82958 -11594 83004
rect -10928 82954 -10882 83006
rect -11084 82908 -10882 82954
rect -12194 82747 -11594 82793
rect -10546 82593 -10163 82639
rect -11884 82347 -11838 82546
rect -11083 82495 -10246 82541
rect -10210 82443 -10163 82593
rect -10546 82397 -10163 82443
rect -11884 82301 -11682 82347
rect -11884 82249 -11838 82301
rect -11083 82299 -10783 82345
rect -12013 82203 -11836 82249
rect -11884 82151 -11836 82203
rect -10737 82185 -10679 82264
rect -10210 82247 -10163 82397
rect -9264 82326 -8964 82372
rect -8770 82277 -8708 83450
rect -10546 82201 -10163 82247
rect -8779 82211 -8696 82277
rect -8268 82228 -7968 82274
rect -10247 82200 -10163 82201
rect -11884 82105 -11682 82151
rect -10737 82131 -10570 82185
rect -10737 82105 -10679 82131
rect -11884 82053 -11836 82105
rect -12013 82007 -11836 82053
rect -11884 81955 -11838 82007
rect -11884 81909 -11682 81955
rect -10698 81764 -10652 81963
rect -10624 81911 -10570 82131
rect -9264 82098 -8764 82144
rect -9264 82000 -8764 82046
rect -8693 82039 -8555 82093
rect -10624 81857 -10226 81911
rect -10954 81718 -10652 81764
rect -10698 81666 -10652 81718
rect -12603 81594 -12220 81640
rect -10700 81620 -10424 81666
rect -12603 81444 -12556 81594
rect -10700 81568 -10652 81620
rect -12520 81496 -11683 81542
rect -10954 81522 -10652 81568
rect -10700 81470 -10652 81522
rect -12603 81398 -12220 81444
rect -10700 81424 -10424 81470
rect -12603 81248 -12556 81398
rect -10698 81372 -10652 81424
rect -11983 81300 -11683 81346
rect -10954 81326 -10652 81372
rect -12603 81202 -12220 81248
rect -12603 81201 -12519 81202
rect -10720 81144 -10570 81170
rect -12178 81090 -10570 81144
rect -12178 80947 -12124 81090
rect -10720 81040 -10570 81090
rect -10280 80899 -10226 81857
rect -8672 81792 -8628 82039
rect -8468 82000 -7968 82046
rect -9264 81674 -8764 81720
rect -8678 81654 -8624 81792
rect -8468 81674 -7968 81720
rect -9264 81549 -8764 81595
rect -9264 81451 -8764 81497
rect -9264 81079 -8964 81125
rect -8672 80986 -8628 81654
rect -8468 81544 -7968 81590
rect -8468 81446 -7968 81492
rect -8468 81348 -7968 81394
rect -8468 81079 -7968 81125
rect -10286 80802 -10220 80899
rect -8678 80848 -8624 80986
rect -9015 80778 -8924 80790
rect -9727 80699 -8924 80778
rect -12294 80000 -12222 80034
rect -12442 79935 -12222 80000
rect -12775 79615 -12475 79661
rect -12775 79177 -12475 79223
rect -12442 78980 -12377 79935
rect -12294 79929 -12222 79935
rect -12163 79698 -11563 79744
rect -12163 79486 -11563 79532
rect -12163 79388 -11563 79434
rect -12163 79290 -11563 79336
rect -12163 79079 -11563 79125
rect -10179 80278 -10082 80289
rect -9727 80278 -9648 80699
rect -9015 80687 -8924 80699
rect -10179 80199 -9648 80278
rect -10179 80173 -10082 80199
rect -8841 80008 -8769 80042
rect -10897 79678 -10851 79877
rect -11053 79632 -10851 79678
rect -10897 79580 -10851 79632
rect -8989 79943 -8769 80008
rect -9322 79623 -9022 79669
rect -10899 79534 -10722 79580
rect -10899 79482 -10851 79534
rect -11053 79436 -10851 79482
rect -10899 79384 -10851 79436
rect -10899 79338 -10722 79384
rect -10897 79286 -10851 79338
rect -11053 79240 -10851 79286
rect -9322 79185 -9022 79231
rect -8989 78988 -8924 79943
rect -8841 79937 -8769 79943
rect -8710 79706 -8110 79752
rect -7444 79686 -7398 79885
rect -7600 79640 -7398 79686
rect -7444 79588 -7398 79640
rect -7446 79542 -7269 79588
rect -8710 79494 -8110 79540
rect -7446 79490 -7398 79542
rect -7600 79444 -7398 79490
rect -8710 79396 -8110 79442
rect -7446 79392 -7398 79444
rect -7446 79346 -7269 79392
rect -8710 79298 -8110 79344
rect -7444 79294 -7398 79346
rect -7600 79248 -7398 79294
rect -8710 79087 -8110 79133
rect -10515 78925 -10132 78971
rect -7062 78933 -6679 78979
rect -11853 78679 -11807 78878
rect -11052 78827 -10215 78873
rect -10179 78775 -10132 78925
rect -10515 78729 -10132 78775
rect -11853 78633 -11651 78679
rect -11853 78581 -11807 78633
rect -11052 78631 -10752 78677
rect -11982 78535 -11805 78581
rect -11853 78483 -11805 78535
rect -10706 78517 -10648 78596
rect -10179 78579 -10132 78729
rect -8400 78687 -8354 78886
rect -7599 78835 -6762 78881
rect -6726 78783 -6679 78933
rect -7062 78737 -6679 78783
rect -8400 78641 -8198 78687
rect -8400 78589 -8354 78641
rect -7599 78639 -7299 78685
rect -10515 78533 -10132 78579
rect -8529 78543 -8352 78589
rect -10216 78532 -10132 78533
rect -11853 78437 -11651 78483
rect -10706 78463 -10539 78517
rect -8400 78491 -8352 78543
rect -7253 78525 -7195 78604
rect -6726 78587 -6679 78737
rect -7062 78541 -6679 78587
rect -6763 78540 -6679 78541
rect -10706 78437 -10648 78463
rect -11853 78385 -11805 78437
rect -11982 78339 -11805 78385
rect -11853 78287 -11807 78339
rect -11853 78241 -11651 78287
rect -10667 78096 -10621 78295
rect -10593 78243 -10539 78463
rect -8400 78445 -8198 78491
rect -7253 78471 -7086 78525
rect -7253 78445 -7195 78471
rect -8400 78393 -8352 78445
rect -8529 78347 -8352 78393
rect -8400 78295 -8354 78347
rect -8400 78249 -8198 78295
rect -10593 78189 -10195 78243
rect -10923 78050 -10621 78096
rect -10667 77998 -10621 78050
rect -12572 77926 -12189 77972
rect -10669 77952 -10393 77998
rect -12572 77776 -12525 77926
rect -10669 77900 -10621 77952
rect -12489 77828 -11652 77874
rect -10923 77854 -10621 77900
rect -10669 77802 -10621 77854
rect -12572 77730 -12189 77776
rect -10669 77756 -10393 77802
rect -12572 77580 -12525 77730
rect -10667 77704 -10621 77756
rect -11952 77632 -11652 77678
rect -10923 77658 -10621 77704
rect -12572 77534 -12189 77580
rect -12572 77533 -12488 77534
rect -10689 77476 -10539 77502
rect -12147 77422 -10539 77476
rect -12147 77279 -12093 77422
rect -10689 77372 -10539 77422
rect -10249 77021 -10195 78189
rect -7214 78104 -7168 78303
rect -7140 78251 -7086 78471
rect -7140 78197 -6742 78251
rect -7470 78058 -7168 78104
rect -7214 78006 -7168 78058
rect -9119 77934 -8736 77980
rect -7216 77960 -6940 78006
rect -9119 77784 -9072 77934
rect -7216 77908 -7168 77960
rect -9036 77836 -8199 77882
rect -7470 77862 -7168 77908
rect -7216 77810 -7168 77862
rect -9119 77738 -8736 77784
rect -7216 77764 -6940 77810
rect -9119 77588 -9072 77738
rect -7214 77712 -7168 77764
rect -8499 77640 -8199 77686
rect -7470 77666 -7168 77712
rect -9119 77542 -8736 77588
rect -9119 77541 -9035 77542
rect -7236 77484 -7086 77510
rect -8694 77430 -7086 77484
rect -8694 77287 -8640 77430
rect -7236 77380 -7086 77430
rect -6796 77072 -6742 78197
rect -10344 75893 -10142 77021
rect -6878 76775 -6656 77072
rect -6352 75893 -6150 83450
rect -10344 75691 -6150 75893
rect -12557 75514 -12226 75586
rect -12557 75249 -4628 75514
rect -13809 74890 -13518 75207
rect -12286 74805 -12214 74839
rect -12434 74740 -12214 74805
rect -12767 74420 -12467 74466
rect -12767 73982 -12467 74028
rect -12434 73785 -12369 74740
rect -12286 74734 -12214 74740
rect -12155 74503 -11555 74549
rect -10889 74483 -10843 74682
rect -11045 74437 -10843 74483
rect -10889 74385 -10843 74437
rect -10891 74339 -10714 74385
rect -12155 74291 -11555 74337
rect -10891 74287 -10843 74339
rect -11045 74241 -10843 74287
rect -8731 74277 -8669 74970
rect -12155 74193 -11555 74239
rect -10891 74189 -10843 74241
rect -10891 74143 -10714 74189
rect -12155 74095 -11555 74141
rect -10889 74091 -10843 74143
rect -11045 74045 -10843 74091
rect -8731 74061 -6168 74277
rect -12155 73884 -11555 73930
rect -10507 73730 -10124 73776
rect -11845 73484 -11799 73683
rect -11044 73632 -10207 73678
rect -10171 73580 -10124 73730
rect -10507 73534 -10124 73580
rect -11845 73438 -11643 73484
rect -11845 73386 -11799 73438
rect -11044 73436 -10744 73482
rect -11974 73340 -11797 73386
rect -11845 73288 -11797 73340
rect -10698 73322 -10640 73401
rect -10171 73384 -10124 73534
rect -9225 73463 -8925 73509
rect -8731 73414 -8669 74061
rect -10507 73338 -10124 73384
rect -8740 73348 -8657 73414
rect -8229 73365 -7929 73411
rect -10208 73337 -10124 73338
rect -11845 73242 -11643 73288
rect -10698 73268 -10531 73322
rect -10698 73242 -10640 73268
rect -11845 73190 -11797 73242
rect -11974 73144 -11797 73190
rect -11845 73092 -11799 73144
rect -11845 73046 -11643 73092
rect -10659 72901 -10613 73100
rect -10585 73048 -10531 73268
rect -9225 73235 -8725 73281
rect -9225 73137 -8725 73183
rect -8654 73176 -8516 73230
rect -10585 72994 -10187 73048
rect -10915 72855 -10613 72901
rect -10659 72803 -10613 72855
rect -12564 72731 -12181 72777
rect -10661 72757 -10385 72803
rect -12564 72581 -12517 72731
rect -10661 72705 -10613 72757
rect -12481 72633 -11644 72679
rect -10915 72659 -10613 72705
rect -10661 72607 -10613 72659
rect -12564 72535 -12181 72581
rect -10661 72561 -10385 72607
rect -12564 72385 -12517 72535
rect -10659 72509 -10613 72561
rect -11944 72437 -11644 72483
rect -10915 72463 -10613 72509
rect -12564 72339 -12181 72385
rect -12564 72338 -12480 72339
rect -10681 72281 -10531 72307
rect -12139 72227 -10531 72281
rect -12139 72084 -12085 72227
rect -10681 72177 -10531 72227
rect -10241 72036 -10187 72994
rect -8633 72929 -8589 73176
rect -8429 73137 -7929 73183
rect -9225 72811 -8725 72857
rect -8639 72791 -8585 72929
rect -8429 72811 -7929 72857
rect -9225 72686 -8725 72732
rect -9225 72588 -8725 72634
rect -9225 72216 -8925 72262
rect -8633 72123 -8589 72791
rect -8429 72681 -7929 72727
rect -8429 72583 -7929 72629
rect -8429 72485 -7929 72531
rect -8429 72216 -7929 72262
rect -10247 71939 -10181 72036
rect -8639 71985 -8585 72123
rect -8976 71915 -8885 71927
rect -9688 71836 -8885 71915
rect -12255 71137 -12183 71171
rect -12403 71072 -12183 71137
rect -12736 70752 -12436 70798
rect -12736 70314 -12436 70360
rect -12403 70117 -12338 71072
rect -12255 71066 -12183 71072
rect -12124 70835 -11524 70881
rect -12124 70623 -11524 70669
rect -12124 70525 -11524 70571
rect -12124 70427 -11524 70473
rect -12124 70216 -11524 70262
rect -10140 71415 -10043 71426
rect -9688 71415 -9609 71836
rect -8976 71824 -8885 71836
rect -10140 71336 -9609 71415
rect -10140 71310 -10043 71336
rect -8802 71145 -8730 71179
rect -10858 70815 -10812 71014
rect -11014 70769 -10812 70815
rect -10858 70717 -10812 70769
rect -8950 71080 -8730 71145
rect -9283 70760 -8983 70806
rect -10860 70671 -10683 70717
rect -10860 70619 -10812 70671
rect -11014 70573 -10812 70619
rect -10860 70521 -10812 70573
rect -10860 70475 -10683 70521
rect -10858 70423 -10812 70475
rect -11014 70377 -10812 70423
rect -9283 70322 -8983 70368
rect -8950 70125 -8885 71080
rect -8802 71074 -8730 71080
rect -8671 70843 -8071 70889
rect -7405 70823 -7359 71022
rect -7561 70777 -7359 70823
rect -7405 70725 -7359 70777
rect -7407 70679 -7230 70725
rect -8671 70631 -8071 70677
rect -7407 70627 -7359 70679
rect -7561 70581 -7359 70627
rect -8671 70533 -8071 70579
rect -7407 70529 -7359 70581
rect -7407 70483 -7230 70529
rect -8671 70435 -8071 70481
rect -7405 70431 -7359 70483
rect -7561 70385 -7359 70431
rect -8671 70224 -8071 70270
rect -10476 70062 -10093 70108
rect -7023 70070 -6640 70116
rect -11814 69816 -11768 70015
rect -11013 69964 -10176 70010
rect -10140 69912 -10093 70062
rect -10476 69866 -10093 69912
rect -11814 69770 -11612 69816
rect -11814 69718 -11768 69770
rect -11013 69768 -10713 69814
rect -11943 69672 -11766 69718
rect -11814 69620 -11766 69672
rect -10667 69654 -10609 69733
rect -10140 69716 -10093 69866
rect -8361 69824 -8315 70023
rect -7560 69972 -6723 70018
rect -6687 69920 -6640 70070
rect -7023 69874 -6640 69920
rect -8361 69778 -8159 69824
rect -8361 69726 -8315 69778
rect -7560 69776 -7260 69822
rect -10476 69670 -10093 69716
rect -8490 69680 -8313 69726
rect -10177 69669 -10093 69670
rect -11814 69574 -11612 69620
rect -10667 69600 -10500 69654
rect -8361 69628 -8313 69680
rect -7214 69662 -7156 69741
rect -6687 69724 -6640 69874
rect -7023 69678 -6640 69724
rect -6724 69677 -6640 69678
rect -10667 69574 -10609 69600
rect -11814 69522 -11766 69574
rect -11943 69476 -11766 69522
rect -11814 69424 -11768 69476
rect -11814 69378 -11612 69424
rect -10628 69233 -10582 69432
rect -10554 69380 -10500 69600
rect -8361 69582 -8159 69628
rect -7214 69608 -7047 69662
rect -7214 69582 -7156 69608
rect -8361 69530 -8313 69582
rect -8490 69484 -8313 69530
rect -8361 69432 -8315 69484
rect -8361 69386 -8159 69432
rect -10554 69326 -10156 69380
rect -10884 69187 -10582 69233
rect -10628 69135 -10582 69187
rect -12533 69063 -12150 69109
rect -10630 69089 -10354 69135
rect -12533 68913 -12486 69063
rect -10630 69037 -10582 69089
rect -12450 68965 -11613 69011
rect -10884 68991 -10582 69037
rect -10630 68939 -10582 68991
rect -12533 68867 -12150 68913
rect -10630 68893 -10354 68939
rect -12533 68717 -12486 68867
rect -10628 68841 -10582 68893
rect -11913 68769 -11613 68815
rect -10884 68795 -10582 68841
rect -12533 68671 -12150 68717
rect -12533 68670 -12449 68671
rect -10650 68613 -10500 68639
rect -12108 68559 -10500 68613
rect -12108 68416 -12054 68559
rect -10650 68509 -10500 68559
rect -10210 68045 -10156 69326
rect -7175 69241 -7129 69440
rect -7101 69388 -7047 69608
rect -7101 69334 -6703 69388
rect -7431 69195 -7129 69241
rect -7175 69143 -7129 69195
rect -9080 69071 -8697 69117
rect -7177 69097 -6901 69143
rect -9080 68921 -9033 69071
rect -7177 69045 -7129 69097
rect -8997 68973 -8160 69019
rect -7431 68999 -7129 69045
rect -7177 68947 -7129 68999
rect -9080 68875 -8697 68921
rect -7177 68901 -6901 68947
rect -9080 68725 -9033 68875
rect -7175 68849 -7129 68901
rect -8460 68777 -8160 68823
rect -7431 68803 -7129 68849
rect -9080 68679 -8697 68725
rect -9080 68678 -8996 68679
rect -7197 68621 -7047 68647
rect -8655 68567 -7047 68621
rect -8655 68424 -8601 68567
rect -7197 68517 -7047 68567
rect -6757 68228 -6703 69334
rect -13782 59190 -13601 67990
rect -10264 67386 -10073 68045
rect -6834 67871 -6567 68228
rect -6359 67386 -6168 74061
rect -10264 67195 -6168 67386
rect -6723 67050 -6669 67056
rect -6800 67033 -6533 67050
rect -12289 67023 -5050 67033
rect -12458 66800 -5050 67023
rect -12289 66784 -5050 66800
rect -6800 66693 -6533 66784
rect -12275 66365 -12203 66399
rect -12423 66300 -12203 66365
rect -12756 65980 -12456 66026
rect -12756 65542 -12456 65588
rect -12423 65345 -12358 66300
rect -12275 66294 -12203 66300
rect -12144 66063 -11544 66109
rect -10878 66043 -10832 66242
rect -11034 65997 -10832 66043
rect -10878 65945 -10832 65997
rect -10880 65899 -10703 65945
rect -12144 65851 -11544 65897
rect -10880 65847 -10832 65899
rect -11034 65801 -10832 65847
rect -12144 65753 -11544 65799
rect -10880 65749 -10832 65801
rect -10880 65703 -10703 65749
rect -12144 65655 -11544 65701
rect -10878 65651 -10832 65703
rect -8720 65677 -8658 66530
rect -11034 65605 -10832 65651
rect -8720 65508 -6242 65677
rect -12144 65444 -11544 65490
rect -10496 65290 -10113 65336
rect -11834 65044 -11788 65243
rect -11033 65192 -10196 65238
rect -10160 65140 -10113 65290
rect -10496 65094 -10113 65140
rect -11834 64998 -11632 65044
rect -11834 64946 -11788 64998
rect -11033 64996 -10733 65042
rect -11963 64900 -11786 64946
rect -11834 64848 -11786 64900
rect -10687 64882 -10629 64961
rect -10160 64944 -10113 65094
rect -9214 65023 -8914 65069
rect -8720 64974 -8658 65508
rect -10496 64898 -10113 64944
rect -8729 64908 -8646 64974
rect -8218 64925 -7918 64971
rect -10197 64897 -10113 64898
rect -11834 64802 -11632 64848
rect -10687 64828 -10520 64882
rect -10687 64802 -10629 64828
rect -11834 64750 -11786 64802
rect -11963 64704 -11786 64750
rect -11834 64652 -11788 64704
rect -11834 64606 -11632 64652
rect -10648 64461 -10602 64660
rect -10574 64608 -10520 64828
rect -9214 64795 -8714 64841
rect -9214 64697 -8714 64743
rect -8643 64736 -8505 64790
rect -10574 64554 -10176 64608
rect -10904 64415 -10602 64461
rect -10648 64363 -10602 64415
rect -12553 64291 -12170 64337
rect -10650 64317 -10374 64363
rect -12553 64141 -12506 64291
rect -10650 64265 -10602 64317
rect -12470 64193 -11633 64239
rect -10904 64219 -10602 64265
rect -10650 64167 -10602 64219
rect -12553 64095 -12170 64141
rect -10650 64121 -10374 64167
rect -12553 63945 -12506 64095
rect -10648 64069 -10602 64121
rect -11933 63997 -11633 64043
rect -10904 64023 -10602 64069
rect -12553 63899 -12170 63945
rect -12553 63898 -12469 63899
rect -10670 63841 -10520 63867
rect -12128 63787 -10520 63841
rect -12128 63644 -12074 63787
rect -10670 63737 -10520 63787
rect -10230 63596 -10176 64554
rect -8622 64489 -8578 64736
rect -8418 64697 -7918 64743
rect -9214 64371 -8714 64417
rect -8628 64351 -8574 64489
rect -8418 64371 -7918 64417
rect -9214 64246 -8714 64292
rect -9214 64148 -8714 64194
rect -9214 63776 -8914 63822
rect -8622 63683 -8578 64351
rect -8418 64241 -7918 64287
rect -8418 64143 -7918 64189
rect -8418 64045 -7918 64091
rect -8418 63776 -7918 63822
rect -10236 63499 -10170 63596
rect -8628 63545 -8574 63683
rect -8965 63475 -8874 63487
rect -9677 63396 -8874 63475
rect -12244 62697 -12172 62731
rect -12392 62632 -12172 62697
rect -12725 62312 -12425 62358
rect -12725 61874 -12425 61920
rect -12392 61677 -12327 62632
rect -12244 62626 -12172 62632
rect -12113 62395 -11513 62441
rect -12113 62183 -11513 62229
rect -12113 62085 -11513 62131
rect -12113 61987 -11513 62033
rect -12113 61776 -11513 61822
rect -10129 62975 -10032 62986
rect -9677 62975 -9598 63396
rect -8965 63384 -8874 63396
rect -10129 62896 -9598 62975
rect -10129 62870 -10032 62896
rect -8791 62705 -8719 62739
rect -10847 62375 -10801 62574
rect -11003 62329 -10801 62375
rect -10847 62277 -10801 62329
rect -8939 62640 -8719 62705
rect -9272 62320 -8972 62366
rect -10849 62231 -10672 62277
rect -10849 62179 -10801 62231
rect -11003 62133 -10801 62179
rect -10849 62081 -10801 62133
rect -10849 62035 -10672 62081
rect -10847 61983 -10801 62035
rect -11003 61937 -10801 61983
rect -9272 61882 -8972 61928
rect -8939 61685 -8874 62640
rect -8791 62634 -8719 62640
rect -8660 62403 -8060 62449
rect -7394 62383 -7348 62582
rect -7550 62337 -7348 62383
rect -7394 62285 -7348 62337
rect -7396 62239 -7219 62285
rect -8660 62191 -8060 62237
rect -7396 62187 -7348 62239
rect -7550 62141 -7348 62187
rect -8660 62093 -8060 62139
rect -7396 62089 -7348 62141
rect -7396 62043 -7219 62089
rect -8660 61995 -8060 62041
rect -7394 61991 -7348 62043
rect -7550 61945 -7348 61991
rect -8660 61784 -8060 61830
rect -10465 61622 -10082 61668
rect -7012 61630 -6629 61676
rect -11803 61376 -11757 61575
rect -11002 61524 -10165 61570
rect -10129 61472 -10082 61622
rect -10465 61426 -10082 61472
rect -11803 61330 -11601 61376
rect -11803 61278 -11757 61330
rect -11002 61328 -10702 61374
rect -11932 61232 -11755 61278
rect -11803 61180 -11755 61232
rect -10656 61214 -10598 61293
rect -10129 61276 -10082 61426
rect -8350 61384 -8304 61583
rect -7549 61532 -6712 61578
rect -6676 61480 -6629 61630
rect -7012 61434 -6629 61480
rect -8350 61338 -8148 61384
rect -8350 61286 -8304 61338
rect -7549 61336 -7249 61382
rect -10465 61230 -10082 61276
rect -8479 61240 -8302 61286
rect -10166 61229 -10082 61230
rect -11803 61134 -11601 61180
rect -10656 61160 -10489 61214
rect -8350 61188 -8302 61240
rect -6676 61284 -6629 61434
rect -7012 61238 -6629 61284
rect -6713 61237 -6629 61238
rect -10656 61134 -10598 61160
rect -11803 61082 -11755 61134
rect -11932 61036 -11755 61082
rect -11803 60984 -11757 61036
rect -11803 60938 -11601 60984
rect -10617 60793 -10571 60992
rect -10543 60940 -10489 61160
rect -8350 61142 -8148 61188
rect -8350 61090 -8302 61142
rect -8479 61044 -8302 61090
rect -8350 60992 -8304 61044
rect -8350 60946 -8148 60992
rect -10543 60886 -10145 60940
rect -10873 60747 -10571 60793
rect -10617 60695 -10571 60747
rect -12522 60623 -12139 60669
rect -10619 60649 -10343 60695
rect -12522 60473 -12475 60623
rect -10619 60597 -10571 60649
rect -12439 60525 -11602 60571
rect -10873 60551 -10571 60597
rect -10619 60499 -10571 60551
rect -12522 60427 -12139 60473
rect -10619 60453 -10343 60499
rect -12522 60277 -12475 60427
rect -10617 60401 -10571 60453
rect -11902 60329 -11602 60375
rect -10873 60355 -10571 60401
rect -12522 60231 -12139 60277
rect -12522 60230 -12438 60231
rect -10639 60173 -10489 60199
rect -12097 60119 -10489 60173
rect -12097 59976 -12043 60119
rect -10639 60069 -10489 60119
rect -10199 59562 -10145 60886
rect -7164 60801 -7118 61000
rect -7420 60755 -7118 60801
rect -7164 60703 -7118 60755
rect -9069 60631 -8686 60677
rect -7166 60657 -6890 60703
rect -9069 60481 -9022 60631
rect -7166 60605 -7118 60657
rect -8986 60533 -8149 60579
rect -7420 60559 -7118 60605
rect -7166 60507 -7118 60559
rect -9069 60435 -8686 60481
rect -7166 60461 -6890 60507
rect -9069 60285 -9022 60435
rect -7164 60409 -7118 60461
rect -8449 60337 -8149 60383
rect -7420 60363 -7118 60409
rect -9069 60239 -8686 60285
rect -9069 60238 -8985 60239
rect -7186 60181 -7036 60207
rect -8644 60127 -7036 60181
rect -8644 59984 -8590 60127
rect -7186 60077 -7036 60127
rect -10228 59381 -10059 59562
rect -6411 59381 -6242 65508
rect -10228 59212 -6242 59381
rect -16789 58418 -10422 58539
rect -16789 57378 -16489 58418
rect -14248 58285 -11470 58311
rect -14248 58251 -11308 58285
rect -14248 58190 -11470 58251
rect -17212 57031 -17091 57173
rect -14248 57031 -14127 58190
rect -13798 57694 -13578 57876
rect -11407 57694 -11373 58197
rect -13798 57624 -11373 57694
rect -13798 57505 -13578 57624
rect -17212 56910 -14127 57031
rect -11407 56101 -11373 57624
rect -11342 57011 -11308 58251
rect -10490 57985 -10445 58418
rect -9655 58253 -7041 58408
rect -10499 57867 -10441 57985
rect -11273 57780 -10573 57826
rect -10388 57780 -9688 57826
rect -11273 57380 -10573 57426
rect -10388 57380 -9688 57426
rect -9655 57226 -9585 58253
rect -8398 58068 -8334 58191
rect -10386 57156 -9585 57226
rect -10511 57011 -10453 57089
rect -11342 56977 -10453 57011
rect -10511 56971 -10453 56977
rect -11273 56780 -10573 56826
rect -10388 56780 -9688 56826
rect -11273 56380 -10573 56426
rect -10388 56380 -9688 56426
rect -9655 56235 -9585 57156
rect -10385 56165 -9585 56235
rect -11407 56067 -10438 56101
rect -10472 56012 -10438 56067
rect -10484 55894 -10426 56012
rect -11273 55780 -10573 55826
rect -10388 55780 -9688 55826
rect -11273 55380 -10573 55426
rect -10388 55380 -9688 55426
rect -9655 55191 -9585 56165
rect -9834 55121 -9585 55191
rect -9358 57982 -8334 58068
rect -9358 57978 -8287 57982
rect -11344 54892 -11144 54938
rect -10964 54892 -10864 54938
rect -10230 54925 -9517 54982
rect -10230 54896 -10096 54925
rect -10497 54760 -10297 54806
rect -10043 54746 -9643 54792
rect -11344 54696 -11144 54742
rect -10964 54696 -10864 54742
rect -10497 54662 -10297 54708
rect -10497 54550 -10297 54596
rect -10043 54550 -9643 54596
rect -11344 54500 -11144 54546
rect -10964 54500 -10864 54546
rect -11062 54161 -11002 54428
rect -10247 54442 -10189 54443
rect -10248 54161 -10188 54442
rect -9764 54161 -9632 54193
rect -11062 54101 -9632 54161
rect -10892 54022 -10832 54054
rect -10147 54022 -10087 54062
rect -9764 54033 -9632 54101
rect -10892 53962 -10087 54022
rect -10892 53923 -10832 53962
rect -10147 53930 -10087 53962
rect -11351 53771 -11151 53817
rect -10643 53771 -10443 53817
rect -10743 53358 -10443 53404
rect -10743 53260 -10443 53306
rect -10743 53162 -10443 53208
rect -11351 53033 -11151 53079
rect -10743 53049 -10443 53095
rect -10743 52951 -10443 52997
rect -11351 52837 -11151 52883
rect -10743 52853 -10443 52899
rect -10744 52739 -10444 52785
rect -11351 52641 -11151 52687
rect -10744 52543 -10444 52589
rect -11195 52390 -11063 52400
rect -11195 52348 -10139 52390
rect -11195 52340 -11063 52348
rect -10945 52225 -10813 52285
rect -11317 52132 -10917 52178
rect -11317 52034 -10917 52080
rect -11317 51936 -10917 51982
rect -11317 51725 -10917 51771
rect -10885 51318 -10843 52225
rect -10804 51860 -10744 51992
rect -10797 51473 -10755 51860
rect -10625 51823 -10425 51869
rect -10724 51637 -10664 51769
rect -10181 51662 -10139 52348
rect -9574 51767 -9517 54925
rect -9358 54196 -9268 57978
rect -8424 57922 -8287 57978
rect -9091 57822 -8891 57868
rect -8711 57822 -8611 57868
rect -8053 57724 -7953 57770
rect -7773 57724 -7573 57770
rect -9091 57626 -8891 57672
rect -8711 57626 -8611 57672
rect -8053 57528 -7953 57574
rect -7773 57528 -7573 57574
rect -9091 57430 -8891 57476
rect -8711 57430 -8611 57476
rect -8053 57332 -7953 57378
rect -7773 57332 -7573 57378
rect -8454 57209 -8394 57245
rect -8454 57149 -7927 57209
rect -8454 57113 -8394 57149
rect -7883 57091 -7591 57148
rect -8616 57030 -8414 57032
rect -9076 56984 -8976 57030
rect -8661 56984 -8414 57030
rect -9076 56886 -8976 56932
rect -8661 56886 -8561 56932
rect -8462 56840 -8414 56984
rect -8053 56887 -7953 56933
rect -8580 56834 -8414 56840
rect -9076 56788 -8976 56834
rect -8661 56788 -8414 56834
rect -8580 56779 -8414 56788
rect -9076 56690 -8976 56736
rect -8661 56690 -8561 56736
rect -8462 56644 -8414 56779
rect -8053 56691 -7953 56737
rect -8582 56638 -8414 56644
rect -9076 56592 -8976 56638
rect -8661 56592 -8414 56638
rect -8582 56583 -8414 56592
rect -9076 56494 -8976 56540
rect -8661 56494 -8561 56540
rect -9076 56396 -8976 56442
rect -9076 56298 -8976 56344
rect -8848 56301 -8774 56470
rect -8462 56453 -8414 56583
rect -8053 56495 -7953 56541
rect -8580 56442 -8414 56453
rect -8661 56396 -8414 56442
rect -8580 56392 -8414 56396
rect -9091 56079 -8891 56125
rect -9091 55883 -8891 55929
rect -9091 55687 -8891 55733
rect -8838 55529 -8781 56301
rect -8661 56298 -8561 56344
rect -8711 56079 -8611 56125
rect -8711 55883 -8611 55929
rect -8711 55687 -8611 55733
rect -9073 55472 -8781 55529
rect -8462 55542 -8414 56392
rect -8103 56276 -8003 56322
rect -7883 56319 -7826 57091
rect -7773 56887 -7573 56933
rect -7773 56691 -7573 56737
rect -7773 56495 -7573 56541
rect -8103 56178 -8003 56224
rect -7890 56150 -7816 56319
rect -7688 56276 -7588 56322
rect -7688 56178 -7588 56224
rect -8103 56080 -8003 56126
rect -7688 56080 -7588 56126
rect -8103 55982 -8003 56028
rect -7688 55982 -7588 56028
rect -8103 55884 -8003 55930
rect -7688 55884 -7588 55930
rect -8103 55786 -8003 55832
rect -7688 55786 -7588 55832
rect -8103 55688 -8003 55734
rect -7688 55688 -7588 55734
rect -8103 55590 -8003 55636
rect -7929 55542 -7869 55637
rect -7688 55590 -7588 55636
rect -8462 55501 -7868 55542
rect -7929 55500 -7869 55501
rect -8788 55307 -8656 55308
rect -8788 55248 -7842 55307
rect -8701 55247 -7842 55248
rect -9091 55122 -8891 55168
rect -8711 55122 -8611 55168
rect -7908 55164 -7848 55247
rect -9091 54926 -8891 54972
rect -8711 54926 -8611 54972
rect -8053 55024 -7953 55070
rect -7773 55024 -7573 55070
rect -8053 54828 -7953 54874
rect -7773 54828 -7573 54874
rect -9091 54730 -8891 54776
rect -8711 54730 -8611 54776
rect -8053 54632 -7953 54678
rect -7773 54632 -7573 54678
rect -7883 54391 -7591 54448
rect -9076 54284 -8976 54330
rect -8661 54327 -8561 54330
rect -8661 54281 -8418 54327
rect -9449 54036 -9268 54196
rect -9076 54186 -8976 54232
rect -8661 54186 -8561 54232
rect -9076 54088 -8976 54134
rect -8661 54132 -8561 54134
rect -8464 54132 -8418 54281
rect -8053 54187 -7953 54233
rect -8661 54090 -8418 54132
rect -8661 54088 -8561 54090
rect -9076 53990 -8976 54036
rect -8661 53990 -8561 54036
rect -9076 53892 -8976 53938
rect -8661 53937 -8561 53938
rect -8464 53937 -8418 54090
rect -8053 53991 -7953 54037
rect -8661 53895 -8418 53937
rect -8661 53892 -8561 53895
rect -9076 53794 -8976 53840
rect -8661 53794 -8561 53840
rect -9076 53696 -8976 53742
rect -9076 53598 -8976 53644
rect -8848 53601 -8774 53770
rect -8661 53741 -8561 53742
rect -8464 53741 -8418 53895
rect -8053 53795 -7953 53841
rect -8661 53699 -8418 53741
rect -8661 53696 -8561 53699
rect -9091 53379 -8891 53425
rect -9091 53183 -8891 53229
rect -9091 52987 -8891 53033
rect -8838 52829 -8781 53601
rect -8661 53598 -8561 53644
rect -8464 53613 -8418 53699
rect -8464 53567 -8206 53613
rect -8103 53576 -8003 53622
rect -7883 53619 -7826 54391
rect -7773 54187 -7573 54233
rect -7773 53991 -7573 54037
rect -7773 53795 -7573 53841
rect -8711 53379 -8611 53425
rect -8711 53183 -8611 53229
rect -8711 52987 -8611 53033
rect -8252 52840 -8206 53567
rect -8103 53478 -8003 53524
rect -7890 53450 -7816 53619
rect -7688 53576 -7588 53622
rect -7688 53478 -7588 53524
rect -8103 53380 -8003 53426
rect -7688 53380 -7588 53426
rect -8103 53282 -8003 53328
rect -7688 53282 -7588 53328
rect -8103 53184 -8003 53230
rect -7688 53184 -7588 53230
rect -8103 53086 -8003 53132
rect -7688 53086 -7588 53132
rect -8103 52988 -8003 53034
rect -7688 52988 -7588 53034
rect -8103 52890 -8003 52936
rect -7931 52840 -7871 52948
rect -7688 52890 -7588 52936
rect -9073 52772 -8287 52829
rect -8252 52802 -7871 52840
rect -8251 52794 -7871 52802
rect -8812 52689 -8680 52691
rect -8452 52689 -8392 52722
rect -8812 52631 -8392 52689
rect -8452 52590 -8392 52631
rect -8344 52620 -8287 52772
rect -8344 52563 -8109 52620
rect -9091 52497 -8891 52543
rect -8711 52497 -8611 52543
rect -9091 52301 -8891 52347
rect -8711 52301 -8611 52347
rect -9091 52105 -8891 52151
rect -8711 52105 -8611 52151
rect -8166 51767 -8109 52563
rect -9574 51710 -8109 51767
rect -8105 51662 -8045 51670
rect -10713 51563 -10671 51637
rect -10181 51620 -8041 51662
rect -10713 51521 -10068 51563
rect -10797 51431 -10142 51473
rect -10730 51318 -10670 51321
rect -10885 51276 -10670 51318
rect -11317 51186 -10917 51232
rect -10730 51189 -10670 51276
rect -11317 51088 -10917 51134
rect -11317 50990 -10917 51036
rect -10625 50877 -10425 50923
rect -11317 50779 -10917 50825
rect -16664 50122 -12822 50250
rect -16664 50117 -16528 50122
rect -12886 49854 -12822 50122
rect -10184 50062 -10142 51431
rect -10110 50731 -10068 51521
rect -8971 51501 -8371 51547
rect -8105 51538 -8045 51620
rect -8971 51403 -8371 51449
rect -8971 51305 -8371 51351
rect -8971 51192 -8371 51238
rect -8971 51094 -8371 51140
rect -8007 51078 -7807 51124
rect -8971 50996 -8371 51042
rect -8007 50882 -7807 50928
rect -8971 50784 -8371 50830
rect -10110 50729 -9914 50731
rect -10110 50533 -9712 50729
rect -10110 50526 -10068 50533
rect -12933 49794 -12796 49854
rect -12609 49694 -12509 49740
rect -12329 49694 -12129 49740
rect -13647 49596 -13447 49642
rect -13267 49596 -13167 49642
rect -12609 49498 -12509 49544
rect -12329 49498 -12129 49544
rect -13647 49400 -13447 49446
rect -13267 49400 -13167 49446
rect -12609 49302 -12509 49348
rect -12329 49302 -12129 49348
rect -13647 49204 -13447 49250
rect -13267 49204 -13167 49250
rect -12826 49081 -12766 49117
rect -13293 49021 -12766 49081
rect -13629 48963 -13337 49020
rect -12826 48985 -12766 49021
rect -13647 48759 -13447 48805
rect -13647 48563 -13447 48609
rect -13647 48367 -13447 48413
rect -13632 48148 -13532 48194
rect -13394 48191 -13337 48963
rect -12806 48902 -12604 48904
rect -12806 48856 -12559 48902
rect -12244 48856 -12144 48902
rect -13267 48759 -13167 48805
rect -12806 48712 -12758 48856
rect -12659 48758 -12559 48804
rect -12244 48758 -12144 48804
rect -12806 48706 -12640 48712
rect -12806 48660 -12559 48706
rect -12244 48660 -12144 48706
rect -12806 48651 -12640 48660
rect -13267 48563 -13167 48609
rect -12806 48516 -12758 48651
rect -12659 48562 -12559 48608
rect -12244 48562 -12144 48608
rect -12806 48510 -12638 48516
rect -12806 48464 -12559 48510
rect -12244 48464 -12144 48510
rect -12806 48455 -12638 48464
rect -13267 48367 -13167 48413
rect -12806 48325 -12758 48455
rect -12659 48366 -12559 48412
rect -12244 48366 -12144 48412
rect -12806 48314 -12640 48325
rect -12806 48268 -12559 48314
rect -12806 48264 -12640 48268
rect -13632 48050 -13532 48096
rect -13404 48022 -13330 48191
rect -13217 48148 -13117 48194
rect -13217 48050 -13117 48096
rect -13632 47952 -13532 47998
rect -13217 47952 -13117 47998
rect -13632 47854 -13532 47900
rect -13217 47854 -13117 47900
rect -13632 47756 -13532 47802
rect -13217 47756 -13117 47802
rect -13632 47658 -13532 47704
rect -13217 47658 -13117 47704
rect -13632 47560 -13532 47606
rect -13217 47560 -13117 47606
rect -13632 47462 -13532 47508
rect -13351 47414 -13291 47509
rect -13217 47462 -13117 47508
rect -12806 47414 -12758 48264
rect -12659 48170 -12559 48216
rect -12446 48173 -12372 48342
rect -12244 48268 -12144 48314
rect -12609 47951 -12509 47997
rect -12609 47755 -12509 47801
rect -12609 47559 -12509 47605
rect -13352 47373 -12758 47414
rect -12439 47401 -12382 48173
rect -12244 48170 -12144 48216
rect -10219 48169 -10129 50062
rect -9908 48619 -9712 50533
rect -7705 48757 -7554 49584
rect -7196 48761 -7041 58253
rect -7261 48494 -6963 48761
rect -6119 48812 -5978 49377
rect -6119 48527 -5979 48812
rect -5299 48786 -5050 66784
rect -4893 49068 -4628 75249
rect -4413 49460 -4187 84113
rect -7964 48169 -7800 48173
rect -3856 48169 -3635 93307
rect -10219 48079 -3635 48169
rect -7964 48075 -7800 48079
rect -12329 47951 -12129 47997
rect -12329 47755 -12129 47801
rect -12329 47559 -12129 47605
rect -13351 47372 -13291 47373
rect -12439 47344 -12147 47401
rect -10005 47298 -9580 47377
rect -3297 47298 -3120 102060
rect -12564 47179 -12432 47180
rect -13378 47120 -12432 47179
rect -13378 47119 -12519 47120
rect -13372 47036 -13312 47119
rect -12609 46994 -12509 47040
rect -12329 46994 -12129 47040
rect -10005 46967 -3120 47298
rect -13647 46896 -13447 46942
rect -13267 46896 -13167 46942
rect -10005 46863 -9580 46967
rect -12609 46798 -12509 46844
rect -12329 46798 -12129 46844
rect -13647 46700 -13447 46746
rect -13267 46700 -13167 46746
rect -12609 46602 -12509 46648
rect -12329 46602 -12129 46648
rect -11060 46631 -10830 46652
rect -2847 46631 -2536 111194
rect -13647 46504 -13447 46550
rect -13267 46504 -13167 46550
rect -13629 46263 -13337 46320
rect -11060 46380 -2536 46631
rect -11060 46364 -10830 46380
rect -13647 46059 -13447 46105
rect -13647 45863 -13447 45909
rect -13647 45667 -13447 45713
rect -13632 45448 -13532 45494
rect -13394 45491 -13337 46263
rect -12659 46199 -12559 46202
rect -12802 46153 -12559 46199
rect -12244 46156 -12144 46202
rect -13267 46059 -13167 46105
rect -12802 46004 -12756 46153
rect -12659 46058 -12559 46104
rect -12244 46058 -12144 46104
rect -12659 46004 -12559 46006
rect -12802 45962 -12559 46004
rect -13267 45863 -13167 45909
rect -12802 45809 -12756 45962
rect -12659 45960 -12559 45962
rect -12244 45960 -12144 46006
rect -12659 45862 -12559 45908
rect -12244 45862 -12144 45908
rect -12659 45809 -12559 45810
rect -12802 45767 -12559 45809
rect -13267 45667 -13167 45713
rect -12802 45613 -12756 45767
rect -12659 45764 -12559 45767
rect -12244 45764 -12144 45810
rect -12659 45666 -12559 45712
rect -12244 45666 -12144 45712
rect -10881 45657 -10540 45713
rect -1914 45657 -1630 120725
rect -12659 45613 -12559 45614
rect -12802 45571 -12559 45613
rect -13632 45350 -13532 45396
rect -13404 45322 -13330 45491
rect -13217 45448 -13117 45494
rect -12802 45485 -12756 45571
rect -12659 45568 -12559 45571
rect -13014 45439 -12756 45485
rect -12659 45470 -12559 45516
rect -12446 45473 -12372 45642
rect -12244 45568 -12144 45614
rect -13217 45350 -13117 45396
rect -13632 45252 -13532 45298
rect -13217 45252 -13117 45298
rect -13632 45154 -13532 45200
rect -13217 45154 -13117 45200
rect -13632 45056 -13532 45102
rect -13217 45056 -13117 45102
rect -13632 44958 -13532 45004
rect -13217 44958 -13117 45004
rect -13632 44860 -13532 44906
rect -13217 44860 -13117 44906
rect -13632 44762 -13532 44808
rect -13349 44712 -13289 44820
rect -13217 44762 -13117 44808
rect -13014 44712 -12968 45439
rect -12609 45251 -12509 45297
rect -12609 45055 -12509 45101
rect -12609 44859 -12509 44905
rect -13349 44674 -12968 44712
rect -12439 44701 -12382 45473
rect -12244 45470 -12144 45516
rect -10881 45388 -1630 45657
rect -10881 45327 -10540 45388
rect -12329 45251 -12129 45297
rect -12329 45055 -12129 45101
rect -12329 44859 -12129 44905
rect -13349 44666 -12969 44674
rect -12933 44644 -12147 44701
rect -12933 44492 -12876 44644
rect -13111 44435 -12876 44492
rect -12828 44561 -12768 44594
rect -12540 44561 -12408 44563
rect -12828 44503 -12408 44561
rect -12828 44462 -12768 44503
rect -13111 43724 -13054 44435
rect -12609 44369 -12509 44415
rect -12329 44369 -12129 44415
rect -12609 44173 -12509 44219
rect -12329 44173 -12129 44219
rect -12609 43977 -12509 44023
rect -12329 43977 -12129 44023
rect -16901 43524 -6998 43724
rect -13482 42882 -5400 42910
rect -13482 40779 -13454 42882
rect -12779 42745 -6103 42754
rect -12779 42726 -5986 42745
rect -13494 40640 -13440 40779
rect -13810 40551 -13610 40597
rect -13810 40242 -13610 40288
rect -13482 40164 -13454 40640
rect -13426 40453 -13380 40589
rect -13204 40551 -13004 40597
rect -13500 40025 -13446 40164
rect -13810 39932 -13610 39978
rect -13810 39736 -13610 39782
rect -13417 39755 -13389 40453
rect -13426 39616 -13372 39755
rect -13810 39374 -13610 39420
rect -13282 40147 -13236 40278
rect -13204 40242 -13004 40288
rect -13810 39276 -13610 39322
rect -13810 39178 -13610 39224
rect -13270 39221 -13242 40147
rect -13204 40030 -13004 40076
rect -13204 39932 -13004 39978
rect -13204 39736 -13004 39782
rect -13204 39638 -13004 39684
rect -13204 39374 -13004 39420
rect -13443 39193 -13242 39221
rect -13810 39058 -13610 39104
rect -13443 39006 -13415 39193
rect -13810 38960 -13610 39006
rect -13810 38862 -13610 38908
rect -13456 38867 -13402 39006
rect -13204 38960 -13004 39006
rect -12779 38753 -12751 42726
rect -7941 42601 -7808 42613
rect -12646 42563 -6236 42601
rect -12646 41798 -12608 42563
rect -13482 38725 -12751 38753
rect -13482 37779 -13454 38725
rect -12646 41118 -12618 41798
rect -10163 42449 -10045 42465
rect -12509 42421 -6373 42449
rect -13494 37640 -13440 37779
rect -13810 37551 -13610 37597
rect -13810 37242 -13610 37288
rect -13482 37164 -13454 37640
rect -13426 37453 -13380 37589
rect -13169 38589 -13033 38590
rect -12737 38589 -12691 38628
rect -13169 38545 -12691 38589
rect -13169 38544 -13033 38545
rect -12737 38492 -12691 38545
rect -13204 37551 -13004 37597
rect -13500 37025 -13446 37164
rect -13810 36932 -13610 36978
rect -13810 36736 -13610 36782
rect -13417 36755 -13389 37453
rect -13426 36616 -13372 36755
rect -13810 36374 -13610 36420
rect -13282 37147 -13236 37278
rect -13204 37242 -13004 37288
rect -13810 36276 -13610 36322
rect -13810 36178 -13610 36224
rect -13270 36221 -13242 37147
rect -13204 37030 -13004 37076
rect -13204 36932 -13004 36978
rect -13204 36736 -13004 36782
rect -13204 36638 -13004 36684
rect -13204 36374 -13004 36420
rect -13443 36193 -13242 36221
rect -13810 36058 -13610 36104
rect -13443 36006 -13415 36193
rect -13810 35960 -13610 36006
rect -13810 35862 -13610 35908
rect -13456 35867 -13402 36006
rect -13204 35960 -13004 36006
rect -13169 35684 -13033 35685
rect -12721 35684 -12675 35723
rect -13169 35640 -12675 35684
rect -13169 35639 -13033 35640
rect -12721 35587 -12675 35640
rect -12646 35448 -12608 41118
rect -13482 35420 -12608 35448
rect -13482 35279 -13454 35420
rect -13494 35140 -13440 35279
rect -13810 35051 -13610 35097
rect -13810 34742 -13610 34788
rect -13482 34664 -13454 35140
rect -13426 34953 -13380 35089
rect -13204 35051 -13004 35097
rect -13500 34525 -13446 34664
rect -13810 34432 -13610 34478
rect -13810 34236 -13610 34282
rect -13417 34255 -13389 34953
rect -13426 34116 -13372 34255
rect -13810 33874 -13610 33920
rect -13282 34647 -13236 34778
rect -13204 34742 -13004 34788
rect -13810 33776 -13610 33822
rect -13810 33678 -13610 33724
rect -13270 33721 -13242 34647
rect -13204 34530 -13004 34576
rect -13204 34432 -13004 34478
rect -13204 34236 -13004 34282
rect -13204 34138 -13004 34184
rect -13204 33874 -13004 33920
rect -13443 33693 -13242 33721
rect -13810 33558 -13610 33604
rect -13443 33506 -13415 33693
rect -13810 33460 -13610 33506
rect -13810 33362 -13610 33408
rect -13456 33367 -13402 33506
rect -13204 33460 -13004 33506
rect -12784 33404 -12738 33540
rect -13169 33267 -13033 33268
rect -12783 33267 -12739 33404
rect -13169 33223 -12739 33267
rect -13169 33222 -13033 33223
rect -12509 32973 -12481 42421
rect -10163 42401 -10045 42421
rect -11296 42290 -11157 42302
rect -12383 42239 -6486 42290
rect -12383 41903 -12345 42239
rect -11296 42233 -11157 42239
rect -10460 42134 -10365 42139
rect -12241 42083 -6636 42134
rect -13482 32945 -12481 32973
rect -13482 32779 -13454 32945
rect -12376 41710 -12345 41903
rect -13494 32640 -13440 32779
rect -13810 32551 -13610 32597
rect -13810 32242 -13610 32288
rect -13482 32164 -13454 32640
rect -13426 32453 -13380 32589
rect -13204 32551 -13004 32597
rect -13500 32025 -13446 32164
rect -13810 31932 -13610 31978
rect -13810 31736 -13610 31782
rect -13417 31755 -13389 32453
rect -13426 31616 -13372 31755
rect -13810 31374 -13610 31420
rect -13282 32147 -13236 32278
rect -13204 32242 -13004 32288
rect -13810 31276 -13610 31322
rect -13810 31178 -13610 31224
rect -13270 31221 -13242 32147
rect -13204 32030 -13004 32076
rect -13204 31932 -13004 31978
rect -13204 31736 -13004 31782
rect -13204 31638 -13004 31684
rect -13204 31374 -13004 31420
rect -13443 31193 -13242 31221
rect -13810 31058 -13610 31104
rect -13443 31006 -13415 31193
rect -13810 30960 -13610 31006
rect -13810 30862 -13610 30908
rect -13456 30867 -13402 31006
rect -13204 30960 -13004 31006
rect -12797 30907 -12751 31043
rect -13169 30787 -13033 30788
rect -12796 30787 -12752 30907
rect -13169 30743 -12752 30787
rect -13169 30742 -13033 30743
rect -12796 30742 -12752 30743
rect -12396 30501 -12345 41710
rect -13482 30473 -12345 30501
rect -13482 30279 -13454 30473
rect -12241 41710 -12195 42083
rect -10460 42080 -10365 42083
rect -13494 30140 -13440 30279
rect -13810 30051 -13610 30097
rect -13810 29742 -13610 29788
rect -13482 29664 -13454 30140
rect -13426 29953 -13380 30089
rect -13204 30051 -13004 30097
rect -13500 29525 -13446 29664
rect -13810 29432 -13610 29478
rect -13810 29236 -13610 29282
rect -13417 29255 -13389 29953
rect -13426 29116 -13372 29255
rect -13810 28874 -13610 28920
rect -13282 29647 -13236 29778
rect -13204 29742 -13004 29788
rect -13810 28776 -13610 28822
rect -13810 28678 -13610 28724
rect -13270 28721 -13242 29647
rect -13204 29530 -13004 29576
rect -13204 29432 -13004 29478
rect -13204 29236 -13004 29282
rect -13204 29138 -13004 29184
rect -13204 28874 -13004 28920
rect -13443 28693 -13242 28721
rect -13810 28558 -13610 28604
rect -13443 28506 -13415 28693
rect -13810 28460 -13610 28506
rect -13810 28362 -13610 28408
rect -13456 28367 -13402 28506
rect -13204 28460 -13004 28506
rect -13173 28239 -13037 28240
rect -12467 28239 -12331 28240
rect -13173 28195 -12331 28239
rect -13173 28194 -13037 28195
rect -12467 28194 -12331 28195
rect -12246 27930 -12195 41710
rect -13482 27902 -12195 27930
rect -13482 27779 -13454 27902
rect -12080 35246 -12034 35382
rect -12076 28333 -12034 35246
rect -11996 35142 -11950 35297
rect -12078 28197 -12032 28333
rect -13494 27640 -13440 27779
rect -13810 27551 -13610 27597
rect -13810 27242 -13610 27288
rect -13482 27164 -13454 27640
rect -13426 27453 -13380 27589
rect -13204 27551 -13004 27597
rect -13500 27025 -13446 27164
rect -13810 26932 -13610 26978
rect -13810 26736 -13610 26782
rect -13417 26755 -13389 27453
rect -13426 26616 -13372 26755
rect -13810 26374 -13610 26420
rect -13282 27147 -13236 27278
rect -13204 27242 -13004 27288
rect -13810 26276 -13610 26322
rect -13810 26178 -13610 26224
rect -13270 26221 -13242 27147
rect -13204 27030 -13004 27076
rect -13204 26932 -13004 26978
rect -13204 26736 -13004 26782
rect -13204 26638 -13004 26684
rect -13204 26374 -13004 26420
rect -13443 26193 -13242 26221
rect -13810 26058 -13610 26104
rect -13443 26006 -13415 26193
rect -13810 25960 -13610 26006
rect -13810 25862 -13610 25908
rect -13456 25867 -13402 26006
rect -13204 25960 -13004 26006
rect -11994 25853 -11952 35142
rect -7674 41776 -7585 41799
rect -11238 41748 -7585 41776
rect -11238 40890 -11210 41748
rect -11238 40789 -11203 40890
rect -11243 40650 -11189 40789
rect -11559 40561 -11359 40607
rect -11559 40252 -11359 40298
rect -11231 40174 -11203 40650
rect -11175 40463 -11129 40599
rect -10953 40561 -10753 40607
rect -8129 40561 -7929 40607
rect -7674 41581 -7585 41748
rect -7672 40890 -7644 41581
rect -7679 40789 -7644 40890
rect -7693 40650 -7639 40789
rect -11249 40035 -11195 40174
rect -11559 39942 -11359 39988
rect -11559 39746 -11359 39792
rect -11166 39765 -11138 40463
rect -7753 40463 -7707 40599
rect -11175 39626 -11121 39765
rect -11559 39384 -11359 39430
rect -11031 40157 -10985 40288
rect -10953 40252 -10753 40298
rect -8129 40252 -7929 40298
rect -7897 40157 -7851 40288
rect -11559 39286 -11359 39332
rect -11559 39188 -11359 39234
rect -11019 39231 -10991 40157
rect -10953 40040 -10753 40086
rect -8129 40040 -7929 40086
rect -10953 39942 -10753 39988
rect -8129 39942 -7929 39988
rect -10953 39746 -10753 39792
rect -8129 39746 -7929 39792
rect -10953 39648 -10753 39694
rect -8129 39648 -7929 39694
rect -10953 39384 -10753 39430
rect -8129 39384 -7929 39430
rect -11192 39203 -10991 39231
rect -7891 39231 -7863 40157
rect -7744 39765 -7716 40463
rect -7679 40174 -7651 40650
rect -7523 40561 -7323 40607
rect -7523 40252 -7323 40298
rect -7687 40035 -7633 40174
rect -7523 39942 -7323 39988
rect -7761 39626 -7707 39765
rect -7523 39746 -7323 39792
rect -7523 39384 -7323 39430
rect -7523 39286 -7323 39332
rect -7891 39203 -7690 39231
rect -11559 39068 -11359 39114
rect -11192 39016 -11164 39203
rect -7718 39016 -7690 39203
rect -7523 39188 -7323 39234
rect -7523 39068 -7323 39114
rect -11559 38970 -11282 39016
rect -11559 38872 -11359 38918
rect -11328 38604 -11282 38970
rect -11205 38877 -11151 39016
rect -10953 38970 -10753 39016
rect -8129 38970 -7929 39016
rect -7731 38877 -7677 39016
rect -7600 38970 -7323 39016
rect -7600 38604 -7554 38970
rect -7523 38872 -7323 38918
rect -11328 38468 -11273 38604
rect -10963 38487 -10663 38533
rect -8219 38487 -7919 38533
rect -7609 38468 -7554 38604
rect -11328 38464 -11282 38468
rect -7600 38464 -7554 38468
rect -11570 38389 -11370 38435
rect -7512 38389 -7312 38435
rect -10963 38291 -10663 38337
rect -8219 38291 -7919 38337
rect -11570 38193 -11370 38239
rect -10962 38177 -10662 38223
rect -8220 38177 -7920 38223
rect -7512 38193 -7312 38239
rect -10962 38079 -10662 38125
rect -8220 38079 -7920 38125
rect -11570 37997 -11370 38043
rect -10962 37981 -10662 38027
rect -8220 37981 -7920 38027
rect -7512 37997 -7312 38043
rect -10962 37868 -10662 37914
rect -8220 37868 -7920 37914
rect -10962 37770 -10662 37816
rect -8220 37770 -7920 37816
rect -10962 37672 -10662 37718
rect -8220 37672 -7920 37718
rect -11570 37259 -11370 37305
rect -10862 37259 -10662 37305
rect -8220 37259 -8020 37305
rect -7512 37259 -7312 37305
rect -10709 36780 -10625 36781
rect -11008 36734 -10625 36780
rect -11545 36636 -11245 36682
rect -10672 36584 -10625 36734
rect -11008 36538 -10625 36584
rect -11545 36440 -10708 36486
rect -10672 36388 -10625 36538
rect -11008 36342 -10625 36388
rect -11546 36027 -11344 36073
rect -11390 35975 -11344 36027
rect -11392 35929 -11215 35975
rect -11392 35877 -11344 35929
rect -11546 35831 -11344 35877
rect -11392 35779 -11344 35831
rect -11392 35733 -11215 35779
rect -11390 35681 -11344 35733
rect -11546 35635 -11344 35681
rect -11390 35610 -11344 35635
rect -10711 35175 -10627 35176
rect -11010 35129 -10627 35175
rect -11547 35031 -11247 35077
rect -10674 34979 -10627 35129
rect -11010 34933 -10627 34979
rect -11547 34835 -10710 34881
rect -10674 34783 -10627 34933
rect -11010 34737 -10627 34783
rect -11548 34422 -11346 34468
rect -11392 34370 -11346 34422
rect -11394 34324 -11217 34370
rect -11394 34272 -11346 34324
rect -11548 34226 -11346 34272
rect -11394 34174 -11346 34226
rect -11394 34128 -11217 34174
rect -11392 34076 -11346 34128
rect -11548 34030 -11346 34076
rect -11392 34005 -11346 34030
rect -11228 33844 -11182 33870
rect -10573 33844 -10527 35547
rect -11228 33798 -10527 33844
rect -11228 33734 -11182 33798
rect -11402 33691 -11266 33699
rect -10461 33691 -10415 37115
rect -11402 33653 -10415 33691
rect -11400 33645 -10415 33653
rect -8467 33691 -8421 37115
rect -8257 36780 -8173 36781
rect -8257 36734 -7874 36780
rect -8257 36584 -8210 36734
rect -7637 36636 -7337 36682
rect -8257 36538 -7874 36584
rect -8257 36388 -8210 36538
rect -8174 36440 -7337 36486
rect -8257 36342 -7874 36388
rect -7538 36027 -7336 36073
rect -7538 35975 -7492 36027
rect -7667 35929 -7490 35975
rect -7538 35877 -7490 35929
rect -7538 35831 -7336 35877
rect -7538 35779 -7490 35831
rect -7667 35733 -7490 35779
rect -7538 35681 -7492 35733
rect -7538 35635 -7336 35681
rect -7538 35610 -7492 35635
rect -8355 33844 -8309 35547
rect -8255 35175 -8171 35176
rect -8255 35129 -7872 35175
rect -8255 34979 -8208 35129
rect -7635 35031 -7335 35077
rect -8255 34933 -7872 34979
rect -8255 34783 -8208 34933
rect -8172 34835 -7335 34881
rect -8255 34737 -7872 34783
rect -7536 34422 -7334 34468
rect -7536 34370 -7490 34422
rect -7665 34324 -7488 34370
rect -7536 34272 -7488 34324
rect -7536 34226 -7334 34272
rect -7536 34174 -7488 34226
rect -7665 34128 -7488 34174
rect -7536 34076 -7490 34128
rect -7536 34030 -7334 34076
rect -7536 34005 -7490 34030
rect -7700 33844 -7654 33870
rect -8355 33798 -7654 33844
rect -7700 33734 -7654 33798
rect -7616 33691 -7480 33699
rect -8467 33653 -7480 33691
rect -8467 33645 -7482 33653
rect -10954 33525 -10654 33571
rect -8228 33525 -7928 33571
rect -11561 33427 -11361 33473
rect -7521 33427 -7321 33473
rect -10954 33329 -10654 33375
rect -8228 33329 -7928 33375
rect -11561 33231 -11361 33277
rect -10953 33215 -10653 33261
rect -8229 33215 -7929 33261
rect -7521 33231 -7321 33277
rect -10953 33117 -10653 33163
rect -8229 33117 -7929 33163
rect -11561 33035 -11361 33081
rect -10953 33019 -10653 33065
rect -8229 33019 -7929 33065
rect -7521 33035 -7321 33081
rect -10953 32906 -10653 32952
rect -8229 32906 -7929 32952
rect -10953 32808 -10653 32854
rect -8229 32808 -7929 32854
rect -10953 32710 -10653 32756
rect -8229 32710 -7929 32756
rect -11561 32297 -11361 32343
rect -10853 32297 -10653 32343
rect -8229 32297 -8029 32343
rect -7521 32297 -7321 32343
rect -11155 32209 -11102 32293
rect -7780 32209 -7727 32293
rect -11155 32152 -10596 32209
rect -11578 31759 -11378 31805
rect -11198 31759 -11098 31805
rect -11578 31563 -11378 31609
rect -11198 31563 -11098 31609
rect -11578 31367 -11378 31413
rect -11198 31367 -11098 31413
rect -10653 31347 -10596 32152
rect -10939 31279 -10879 31320
rect -11299 31221 -10879 31279
rect -11299 31219 -11167 31221
rect -10939 31188 -10879 31221
rect -10831 31290 -10596 31347
rect -8286 32152 -7727 32209
rect -8286 31347 -8229 32152
rect -6932 35142 -6886 35297
rect -6848 35246 -6802 35382
rect -7784 31759 -7684 31805
rect -7504 31759 -7304 31805
rect -7784 31563 -7684 31609
rect -7504 31563 -7304 31609
rect -8090 31460 -8030 31530
rect -8090 31402 -7943 31460
rect -8090 31398 -8030 31402
rect -8286 31290 -8051 31347
rect -10831 31138 -10774 31290
rect -11560 31081 -10774 31138
rect -8108 31138 -8051 31290
rect -8001 31279 -7943 31402
rect -7784 31367 -7684 31413
rect -7504 31367 -7304 31413
rect -8001 31221 -7583 31279
rect -7715 31219 -7583 31221
rect -10738 31108 -10358 31116
rect -11578 30877 -11378 30923
rect -11578 30681 -11378 30727
rect -11578 30485 -11378 30531
rect -11563 30266 -11463 30312
rect -11325 30309 -11268 31081
rect -10739 31070 -10358 31108
rect -11198 30877 -11098 30923
rect -11198 30681 -11098 30727
rect -11198 30485 -11098 30531
rect -10739 30343 -10693 31070
rect -10590 30974 -10490 31020
rect -10418 30962 -10358 31070
rect -8524 31108 -8144 31116
rect -8524 31070 -8143 31108
rect -8108 31081 -7322 31138
rect -10175 30974 -10075 31020
rect -8807 30974 -8707 31020
rect -8524 30962 -8464 31070
rect -8392 30974 -8292 31020
rect -10590 30876 -10490 30922
rect -10175 30876 -10075 30922
rect -8807 30876 -8707 30922
rect -8392 30876 -8292 30922
rect -10590 30778 -10490 30824
rect -10175 30778 -10075 30824
rect -8807 30778 -8707 30824
rect -8392 30778 -8292 30824
rect -10590 30680 -10490 30726
rect -10175 30680 -10075 30726
rect -8807 30680 -8707 30726
rect -8392 30680 -8292 30726
rect -10590 30582 -10490 30628
rect -10175 30582 -10075 30628
rect -8807 30582 -8707 30628
rect -8392 30582 -8292 30628
rect -10590 30484 -10490 30530
rect -10175 30484 -10075 30530
rect -8807 30484 -8707 30530
rect -8392 30484 -8292 30530
rect -10590 30386 -10490 30432
rect -11563 30168 -11463 30214
rect -11335 30140 -11261 30309
rect -11148 30266 -11048 30312
rect -10951 30297 -10693 30343
rect -11148 30211 -11048 30214
rect -10951 30211 -10905 30297
rect -10590 30288 -10490 30334
rect -10377 30291 -10303 30460
rect -10175 30386 -10075 30432
rect -8807 30386 -8707 30432
rect -11148 30169 -10905 30211
rect -11148 30168 -11048 30169
rect -11563 30070 -11463 30116
rect -11148 30070 -11048 30116
rect -11563 29972 -11463 30018
rect -11148 30015 -11048 30018
rect -10951 30015 -10905 30169
rect -10540 30069 -10440 30115
rect -11148 29973 -10905 30015
rect -11148 29972 -11048 29973
rect -11563 29874 -11463 29920
rect -11148 29874 -11048 29920
rect -11563 29776 -11463 29822
rect -11148 29820 -11048 29822
rect -10951 29820 -10905 29973
rect -10540 29873 -10440 29919
rect -11148 29778 -10905 29820
rect -11148 29776 -11048 29778
rect -11563 29678 -11463 29724
rect -11148 29678 -11048 29724
rect -10951 29629 -10905 29778
rect -10540 29677 -10440 29723
rect -11563 29580 -11463 29626
rect -11148 29583 -10905 29629
rect -11148 29580 -11048 29583
rect -10370 29519 -10313 30291
rect -10175 30288 -10075 30334
rect -8807 30288 -8707 30334
rect -8579 30291 -8505 30460
rect -8392 30386 -8292 30432
rect -8189 30343 -8143 31070
rect -7784 30877 -7684 30923
rect -7784 30681 -7684 30727
rect -7784 30485 -7684 30531
rect -10260 30069 -10060 30115
rect -8822 30069 -8622 30115
rect -10260 29873 -10060 29919
rect -8822 29873 -8622 29919
rect -10260 29677 -10060 29723
rect -8822 29677 -8622 29723
rect -8569 29519 -8512 30291
rect -8392 30288 -8292 30334
rect -8189 30297 -7931 30343
rect -7977 30211 -7931 30297
rect -7834 30266 -7734 30312
rect -7614 30309 -7557 31081
rect -7504 30877 -7304 30923
rect -7504 30681 -7304 30727
rect -7504 30485 -7304 30531
rect -7834 30211 -7734 30214
rect -7977 30169 -7734 30211
rect -8442 30069 -8342 30115
rect -7977 30015 -7931 30169
rect -7834 30168 -7734 30169
rect -7621 30140 -7547 30309
rect -7419 30266 -7319 30312
rect -7419 30168 -7319 30214
rect -7834 30070 -7734 30116
rect -7419 30070 -7319 30116
rect -7834 30015 -7734 30018
rect -7977 29973 -7734 30015
rect -8442 29873 -8342 29919
rect -7977 29820 -7931 29973
rect -7834 29972 -7734 29973
rect -7419 29972 -7319 30018
rect -7834 29874 -7734 29920
rect -7419 29874 -7319 29920
rect -7834 29820 -7734 29822
rect -7977 29778 -7734 29820
rect -8442 29677 -8342 29723
rect -7977 29629 -7931 29778
rect -7834 29776 -7734 29778
rect -7419 29776 -7319 29822
rect -7834 29678 -7734 29724
rect -7419 29678 -7319 29724
rect -7977 29583 -7734 29629
rect -7834 29580 -7734 29583
rect -7419 29580 -7319 29626
rect -10370 29462 -10078 29519
rect -8804 29462 -8512 29519
rect -8089 29473 -8029 29516
rect -8453 29413 -8029 29473
rect -8089 29384 -8029 29413
rect -10540 29232 -10440 29278
rect -10260 29232 -10060 29278
rect -8822 29232 -8622 29278
rect -8442 29232 -8342 29278
rect -11578 29134 -11378 29180
rect -11198 29134 -11098 29180
rect -7784 29134 -7684 29180
rect -7504 29134 -7304 29180
rect -10540 29036 -10440 29082
rect -10260 29036 -10060 29082
rect -8822 29036 -8622 29082
rect -8442 29036 -8342 29082
rect -11578 28938 -11378 28984
rect -11198 28938 -11098 28984
rect -10540 28840 -10440 28886
rect -10260 28840 -10060 28886
rect -8822 28840 -8622 28886
rect -8442 28840 -8342 28886
rect -7784 28938 -7684 28984
rect -7504 28938 -7304 28984
rect -11578 28742 -11378 28788
rect -11198 28742 -11098 28788
rect -10395 28663 -10335 28746
rect -8547 28663 -8487 28746
rect -7784 28742 -7684 28788
rect -7504 28742 -7304 28788
rect -11188 28662 -10329 28663
rect -11275 28603 -10329 28662
rect -8553 28662 -7694 28663
rect -8553 28603 -7607 28662
rect -11275 28602 -11143 28603
rect -7739 28602 -7607 28603
rect -8090 28547 -8030 28575
rect -8090 28487 -7582 28547
rect -8090 28438 -8030 28487
rect -11560 28381 -11268 28438
rect -10416 28409 -10356 28410
rect -8526 28409 -8466 28410
rect -11578 28177 -11378 28223
rect -11578 27981 -11378 28027
rect -11578 27785 -11378 27831
rect -11563 27566 -11463 27612
rect -11325 27609 -11268 28381
rect -10949 28368 -10355 28409
rect -8527 28368 -7933 28409
rect -11198 28177 -11098 28223
rect -11198 27981 -11098 28027
rect -11198 27785 -11098 27831
rect -11563 27468 -11463 27514
rect -11335 27440 -11261 27609
rect -11148 27566 -11048 27612
rect -10949 27518 -10901 28368
rect -10590 28274 -10490 28320
rect -10416 28273 -10356 28368
rect -10175 28274 -10075 28320
rect -8807 28274 -8707 28320
rect -8526 28273 -8466 28368
rect -8392 28274 -8292 28320
rect -10590 28176 -10490 28222
rect -10175 28176 -10075 28222
rect -8807 28176 -8707 28222
rect -8392 28176 -8292 28222
rect -10590 28078 -10490 28124
rect -10175 28078 -10075 28124
rect -8807 28078 -8707 28124
rect -8392 28078 -8292 28124
rect -10590 27980 -10490 28026
rect -10175 27980 -10075 28026
rect -8807 27980 -8707 28026
rect -8392 27980 -8292 28026
rect -10590 27882 -10490 27928
rect -10175 27882 -10075 27928
rect -8807 27882 -8707 27928
rect -8392 27882 -8292 27928
rect -10590 27784 -10490 27830
rect -10175 27784 -10075 27830
rect -8807 27784 -8707 27830
rect -8392 27784 -8292 27830
rect -10590 27686 -10490 27732
rect -10590 27588 -10490 27634
rect -10377 27591 -10303 27760
rect -10175 27686 -10075 27732
rect -8807 27686 -8707 27732
rect -11067 27514 -10901 27518
rect -11148 27468 -10901 27514
rect -11067 27457 -10901 27468
rect -11563 27370 -11463 27416
rect -11148 27370 -11048 27416
rect -10949 27327 -10901 27457
rect -10540 27369 -10440 27415
rect -11069 27318 -10901 27327
rect -11563 27272 -11463 27318
rect -11148 27272 -10901 27318
rect -11069 27266 -10901 27272
rect -11563 27174 -11463 27220
rect -11148 27174 -11048 27220
rect -10949 27131 -10901 27266
rect -10540 27173 -10440 27219
rect -11067 27122 -10901 27131
rect -11563 27076 -11463 27122
rect -11148 27076 -10901 27122
rect -11067 27070 -10901 27076
rect -11563 26978 -11463 27024
rect -11148 26978 -11048 27024
rect -10949 26926 -10901 27070
rect -10540 26977 -10440 27023
rect -11563 26880 -11463 26926
rect -11148 26880 -10901 26926
rect -11103 26878 -10901 26880
rect -10370 26819 -10313 27591
rect -10175 27588 -10075 27634
rect -8807 27588 -8707 27634
rect -8579 27591 -8505 27760
rect -8392 27686 -8292 27732
rect -10260 27369 -10060 27415
rect -8822 27369 -8622 27415
rect -10260 27173 -10060 27219
rect -8822 27173 -8622 27219
rect -10260 26977 -10060 27023
rect -8822 26977 -8622 27023
rect -8569 26819 -8512 27591
rect -8392 27588 -8292 27634
rect -7981 27518 -7933 28368
rect -7614 28381 -7322 28438
rect -7784 28177 -7684 28223
rect -7784 27981 -7684 28027
rect -7784 27785 -7684 27831
rect -7834 27566 -7734 27612
rect -7614 27609 -7557 28381
rect -7504 28177 -7304 28223
rect -7504 27981 -7304 28027
rect -7504 27785 -7304 27831
rect -7981 27514 -7815 27518
rect -7981 27468 -7734 27514
rect -7981 27457 -7815 27468
rect -8442 27369 -8342 27415
rect -7981 27327 -7933 27457
rect -7621 27440 -7547 27609
rect -7419 27566 -7319 27612
rect -7419 27468 -7319 27514
rect -7834 27370 -7734 27416
rect -7419 27370 -7319 27416
rect -7981 27318 -7813 27327
rect -7981 27272 -7734 27318
rect -7419 27272 -7319 27318
rect -7981 27266 -7813 27272
rect -8442 27173 -8342 27219
rect -7981 27131 -7933 27266
rect -7834 27174 -7734 27220
rect -7419 27174 -7319 27220
rect -7981 27122 -7815 27131
rect -7981 27076 -7734 27122
rect -7419 27076 -7319 27122
rect -7981 27070 -7815 27076
rect -8442 26977 -8342 27023
rect -7981 26926 -7933 27070
rect -7834 26978 -7734 27024
rect -7419 26978 -7319 27024
rect -7981 26880 -7734 26926
rect -7419 26880 -7319 26926
rect -7981 26878 -7779 26880
rect -10941 26761 -10881 26797
rect -10370 26762 -10078 26819
rect -8804 26762 -8512 26819
rect -10941 26701 -10414 26761
rect -10941 26665 -10881 26701
rect -10540 26532 -10440 26578
rect -10260 26532 -10060 26578
rect -8822 26532 -8622 26578
rect -8442 26532 -8342 26578
rect -11578 26434 -11378 26480
rect -11198 26434 -11098 26480
rect -7784 26434 -7684 26480
rect -7504 26434 -7304 26480
rect -10540 26336 -10440 26382
rect -10260 26336 -10060 26382
rect -8822 26336 -8622 26382
rect -8442 26336 -8342 26382
rect -11578 26238 -11378 26284
rect -11198 26238 -11098 26284
rect -11578 26042 -11378 26088
rect -11198 26042 -11098 26088
rect -7784 26238 -7684 26284
rect -7504 26238 -7304 26284
rect -10540 26140 -10440 26186
rect -10260 26140 -10060 26186
rect -8822 26140 -8622 26186
rect -8442 26140 -8342 26186
rect -7784 26042 -7684 26088
rect -7504 26042 -7304 26088
rect -10911 25928 -10774 25988
rect -8108 25928 -7971 25988
rect -12005 25841 -11952 25853
rect -12005 25717 -11959 25841
rect -10885 25757 -10821 25928
rect -10916 25582 -10602 25757
rect -8061 25590 -7997 25928
rect -6930 25853 -6888 35142
rect -6848 28333 -6806 35246
rect -6850 28197 -6804 28333
rect -6687 27930 -6636 42083
rect -6537 30501 -6486 42239
rect -6401 32973 -6373 42421
rect -6274 35448 -6236 42563
rect -6131 41553 -5986 42726
rect -6131 38753 -6103 41553
rect -5878 40551 -5678 40597
rect -5428 41541 -5400 42882
rect -5428 41341 -5048 41541
rect -5428 40779 -5400 41341
rect -5442 40640 -5388 40779
rect -5502 40453 -5456 40589
rect -5878 40242 -5678 40288
rect -5646 40147 -5600 40278
rect -5878 40030 -5678 40076
rect -5878 39932 -5678 39978
rect -5878 39736 -5678 39782
rect -5878 39638 -5678 39684
rect -5878 39374 -5678 39420
rect -5640 39221 -5612 40147
rect -5493 39755 -5465 40453
rect -5428 40164 -5400 40640
rect -5272 40551 -5072 40597
rect -5272 40242 -5072 40288
rect -5436 40025 -5382 40164
rect -5272 39932 -5072 39978
rect -5510 39616 -5456 39755
rect -5272 39736 -5072 39782
rect -5272 39374 -5072 39420
rect -5272 39276 -5072 39322
rect -5640 39193 -5439 39221
rect -5467 39006 -5439 39193
rect -5272 39178 -5072 39224
rect -5272 39058 -5072 39104
rect -5878 38960 -5678 39006
rect -5480 38867 -5426 39006
rect -5272 38960 -5072 39006
rect -5272 38862 -5072 38908
rect -6131 38725 -5400 38753
rect -6191 38589 -6145 38628
rect -5849 38589 -5713 38590
rect -6191 38545 -5713 38589
rect -6191 38492 -6145 38545
rect -5849 38544 -5713 38545
rect -5878 37551 -5678 37597
rect -5428 37779 -5400 38725
rect -5442 37640 -5388 37779
rect -5502 37453 -5456 37589
rect -5878 37242 -5678 37288
rect -5646 37147 -5600 37278
rect -5878 37030 -5678 37076
rect -5878 36932 -5678 36978
rect -5878 36736 -5678 36782
rect -5878 36638 -5678 36684
rect -5878 36374 -5678 36420
rect -5640 36221 -5612 37147
rect -5493 36755 -5465 37453
rect -5428 37164 -5400 37640
rect -5272 37551 -5072 37597
rect -5272 37242 -5072 37288
rect -5436 37025 -5382 37164
rect -5272 36932 -5072 36978
rect -5510 36616 -5456 36755
rect -5272 36736 -5072 36782
rect -5272 36374 -5072 36420
rect -5272 36276 -5072 36322
rect -5640 36193 -5439 36221
rect -5467 36006 -5439 36193
rect -5272 36178 -5072 36224
rect -5272 36058 -5072 36104
rect -5878 35960 -5678 36006
rect -5480 35867 -5426 36006
rect -5272 35960 -5072 36006
rect -5272 35862 -5072 35908
rect -6207 35684 -6161 35723
rect -5849 35684 -5713 35685
rect -6207 35640 -5713 35684
rect -6207 35587 -6161 35640
rect -5849 35639 -5713 35640
rect -6274 35420 -5400 35448
rect -5878 35051 -5678 35097
rect -5428 35279 -5400 35420
rect -5442 35140 -5388 35279
rect -5502 34953 -5456 35089
rect -5878 34742 -5678 34788
rect -5646 34647 -5600 34778
rect -5878 34530 -5678 34576
rect -5878 34432 -5678 34478
rect -5878 34236 -5678 34282
rect -5878 34138 -5678 34184
rect -5878 33874 -5678 33920
rect -5640 33721 -5612 34647
rect -5493 34255 -5465 34953
rect -5428 34664 -5400 35140
rect -5272 35051 -5072 35097
rect -5272 34742 -5072 34788
rect -5436 34525 -5382 34664
rect -5272 34432 -5072 34478
rect -5510 34116 -5456 34255
rect -5272 34236 -5072 34282
rect -5272 33874 -5072 33920
rect -5272 33776 -5072 33822
rect -5640 33693 -5439 33721
rect -6144 33404 -6098 33540
rect -5467 33506 -5439 33693
rect -5272 33678 -5072 33724
rect -5272 33558 -5072 33604
rect -5878 33460 -5678 33506
rect -6143 33267 -6099 33404
rect -5480 33367 -5426 33506
rect -5272 33460 -5072 33506
rect -5272 33362 -5072 33408
rect -5849 33267 -5713 33268
rect -6143 33223 -5713 33267
rect -5849 33222 -5713 33223
rect -6401 32945 -5400 32973
rect -5878 32551 -5678 32597
rect -5428 32779 -5400 32945
rect -5442 32640 -5388 32779
rect -5502 32453 -5456 32589
rect -5878 32242 -5678 32288
rect -5646 32147 -5600 32278
rect -5878 32030 -5678 32076
rect -5878 31932 -5678 31978
rect -5878 31736 -5678 31782
rect -5878 31638 -5678 31684
rect -5878 31374 -5678 31420
rect -5640 31221 -5612 32147
rect -5493 31755 -5465 32453
rect -5428 32164 -5400 32640
rect -5272 32551 -5072 32597
rect -5272 32242 -5072 32288
rect -5436 32025 -5382 32164
rect -5272 31932 -5072 31978
rect -5510 31616 -5456 31755
rect -5272 31736 -5072 31782
rect -5272 31374 -5072 31420
rect -5272 31276 -5072 31322
rect -5640 31193 -5439 31221
rect -6131 30907 -6085 31043
rect -5467 31006 -5439 31193
rect -5272 31178 -5072 31224
rect -5272 31058 -5072 31104
rect -5878 30960 -5678 31006
rect -6130 30787 -6086 30907
rect -5480 30867 -5426 31006
rect -5272 30960 -5072 31006
rect -5272 30862 -5072 30908
rect -5849 30787 -5713 30788
rect -6130 30743 -5713 30787
rect -6130 30742 -6086 30743
rect -5849 30742 -5713 30743
rect -6537 30473 -5400 30501
rect -5878 30051 -5678 30097
rect -5428 30279 -5400 30473
rect -5442 30140 -5388 30279
rect -5502 29953 -5456 30089
rect -5878 29742 -5678 29788
rect -5646 29647 -5600 29778
rect -5878 29530 -5678 29576
rect -5878 29432 -5678 29478
rect -5878 29236 -5678 29282
rect -5878 29138 -5678 29184
rect -5878 28874 -5678 28920
rect -5640 28721 -5612 29647
rect -5493 29255 -5465 29953
rect -5428 29664 -5400 30140
rect -5272 30051 -5072 30097
rect -5272 29742 -5072 29788
rect -5436 29525 -5382 29664
rect -5272 29432 -5072 29478
rect -5510 29116 -5456 29255
rect -5272 29236 -5072 29282
rect -5272 28874 -5072 28920
rect -5272 28776 -5072 28822
rect -5640 28693 -5439 28721
rect -5467 28506 -5439 28693
rect -5272 28678 -5072 28724
rect -5272 28558 -5072 28604
rect -5878 28460 -5678 28506
rect -5480 28367 -5426 28506
rect -5272 28460 -5072 28506
rect -5272 28362 -5072 28408
rect -6551 28239 -6415 28240
rect -5845 28239 -5709 28240
rect -6551 28195 -5709 28239
rect -6551 28194 -6415 28195
rect -5845 28194 -5709 28195
rect -6687 27902 -5400 27930
rect -6340 27830 -5537 27858
rect -6340 27812 -6204 27830
rect -5878 27551 -5678 27597
rect -5565 27466 -5537 27830
rect -5428 27779 -5400 27902
rect -5442 27640 -5388 27779
rect -5590 27327 -5536 27466
rect -5502 27453 -5456 27589
rect -5878 27242 -5678 27288
rect -5646 27147 -5600 27278
rect -5878 27030 -5678 27076
rect -5878 26932 -5678 26978
rect -6601 26789 -6401 26835
rect -6221 26789 -6121 26835
rect -5878 26736 -5678 26782
rect -6601 26593 -6401 26639
rect -6221 26593 -6121 26639
rect -5878 26638 -5678 26684
rect -6601 26397 -6401 26443
rect -6221 26397 -6121 26443
rect -5878 26374 -5678 26420
rect -5640 26221 -5612 27147
rect -5567 26388 -5539 27327
rect -5493 26755 -5465 27453
rect -5428 27164 -5400 27640
rect -5272 27551 -5072 27597
rect -5272 27242 -5072 27288
rect -5436 27025 -5382 27164
rect -5272 26932 -5072 26978
rect -5510 26616 -5456 26755
rect -5272 26736 -5072 26782
rect -5584 26249 -5530 26388
rect -5272 26374 -5072 26420
rect -5272 26276 -5072 26322
rect -5640 26193 -5439 26221
rect -5467 26006 -5439 26193
rect -5272 26178 -5072 26224
rect -5272 26058 -5072 26104
rect -5878 25960 -5678 26006
rect -5480 25867 -5426 26006
rect -5272 25960 -5072 26006
rect -5272 25862 -5072 25908
rect -6932 25717 -6886 25853
rect -8060 25573 -7997 25590
rect -16664 25447 -16528 25451
rect -14173 25447 -13998 25467
rect -16664 25315 -5526 25447
rect -14173 25304 -13998 25315
rect -10410 25078 -9810 25124
rect -5476 25051 -4876 25097
rect -11022 24980 -10722 25026
rect -6088 24953 -5788 24999
rect -10410 24867 -9810 24913
rect -5476 24840 -4876 24886
rect -10410 24769 -9810 24815
rect -5476 24742 -4876 24788
rect -10410 24671 -9810 24717
rect -5476 24644 -4876 24690
rect -11022 24542 -10722 24588
rect -6088 24515 -5788 24561
rect -10410 24459 -9810 24505
rect -5476 24432 -4876 24478
rect -13911 24356 -13740 24367
rect -13911 24180 -7225 24356
rect -13911 24167 -13740 24180
rect -11311 23885 -11111 23931
rect -10931 23885 -10831 23931
rect -6384 23885 -6184 23931
rect -6004 23885 -5904 23931
rect -11311 23689 -11111 23735
rect -10931 23689 -10831 23735
rect -6384 23689 -6184 23735
rect -6004 23689 -5904 23735
rect -11311 23493 -11111 23539
rect -10931 23493 -10831 23539
rect -10672 23405 -10612 23446
rect -11032 23347 -10612 23405
rect -11032 23345 -10900 23347
rect -10672 23314 -10612 23347
rect -11436 23207 -11001 23264
rect -10471 23234 -10091 23242
rect -11436 19643 -11379 23207
rect -11311 23003 -11111 23049
rect -11311 22807 -11111 22853
rect -11311 22611 -11111 22657
rect -11296 22392 -11196 22438
rect -11058 22435 -11001 23207
rect -10472 23196 -10091 23234
rect -10931 23003 -10831 23049
rect -10931 22807 -10831 22853
rect -10931 22611 -10831 22657
rect -10472 22469 -10426 23196
rect -10323 23100 -10223 23146
rect -10151 23088 -10091 23196
rect -9908 23100 -9808 23146
rect -10323 23002 -10223 23048
rect -9908 23002 -9808 23048
rect -10323 22904 -10223 22950
rect -9908 22904 -9808 22950
rect -10323 22806 -10223 22852
rect -9908 22806 -9808 22852
rect -10323 22708 -10223 22754
rect -9908 22708 -9808 22754
rect -10323 22610 -10223 22656
rect -9908 22610 -9808 22656
rect -10323 22512 -10223 22558
rect -11296 22294 -11196 22340
rect -11068 22266 -10994 22435
rect -10881 22392 -10781 22438
rect -10684 22423 -10426 22469
rect -10881 22337 -10781 22340
rect -10684 22337 -10638 22423
rect -10323 22414 -10223 22460
rect -10110 22417 -10036 22586
rect -9908 22512 -9808 22558
rect -10881 22295 -10638 22337
rect -10881 22294 -10781 22295
rect -11296 22196 -11196 22242
rect -10881 22196 -10781 22242
rect -11296 22098 -11196 22144
rect -10881 22141 -10781 22144
rect -10684 22141 -10638 22295
rect -10273 22195 -10173 22241
rect -10881 22099 -10638 22141
rect -10881 22098 -10781 22099
rect -11296 22000 -11196 22046
rect -10881 22000 -10781 22046
rect -11296 21902 -11196 21948
rect -10881 21946 -10781 21948
rect -10684 21946 -10638 22099
rect -10273 21999 -10173 22045
rect -10881 21904 -10638 21946
rect -10881 21902 -10781 21904
rect -11296 21804 -11196 21850
rect -10881 21804 -10781 21850
rect -10684 21755 -10638 21904
rect -10273 21803 -10173 21849
rect -11296 21706 -11196 21752
rect -10881 21709 -10638 21755
rect -10881 21706 -10781 21709
rect -10103 21645 -10046 22417
rect -9908 22414 -9808 22460
rect -9993 22195 -9793 22241
rect -9993 21999 -9793 22045
rect -6384 23493 -6184 23539
rect -6004 23493 -5904 23539
rect -5745 23405 -5685 23446
rect -6105 23347 -5685 23405
rect -6105 23345 -5973 23347
rect -5745 23314 -5685 23347
rect -9993 21803 -9793 21849
rect -10586 21599 -10526 21642
rect -10586 21539 -10162 21599
rect -10103 21588 -9811 21645
rect -10586 21510 -10526 21539
rect -10273 21358 -10173 21404
rect -9993 21358 -9793 21404
rect -11311 21260 -11111 21306
rect -10931 21260 -10831 21306
rect -7443 21659 -7371 21693
rect -7443 21594 -7223 21659
rect -7443 21588 -7371 21594
rect -8814 21337 -8768 21536
rect -8102 21357 -7502 21403
rect -8814 21291 -8612 21337
rect -8814 21239 -8768 21291
rect -10273 21162 -10173 21208
rect -9993 21162 -9793 21208
rect -8943 21193 -8766 21239
rect -8814 21141 -8766 21193
rect -8102 21145 -7502 21191
rect -11311 21064 -11111 21110
rect -10931 21064 -10831 21110
rect -8814 21095 -8612 21141
rect -8814 21043 -8766 21095
rect -8102 21047 -7502 21093
rect -10273 20966 -10173 21012
rect -9993 20966 -9793 21012
rect -8943 20997 -8766 21043
rect -8814 20945 -8768 20997
rect -8102 20949 -7502 20995
rect -11311 20868 -11111 20914
rect -10931 20868 -10831 20914
rect -10128 20789 -10068 20872
rect -8814 20899 -8612 20945
rect -10921 20788 -10062 20789
rect -11008 20729 -10062 20788
rect -8102 20738 -7502 20784
rect -11008 20728 -10876 20729
rect -10585 20673 -10525 20701
rect -11033 20613 -10525 20673
rect -7288 20639 -7223 21594
rect -7190 21274 -6890 21320
rect -6509 23207 -6074 23264
rect -5544 23234 -5164 23242
rect -7190 20836 -6890 20882
rect -10585 20564 -10525 20613
rect -9533 20584 -9150 20630
rect -11293 20507 -11001 20564
rect -10149 20535 -10089 20536
rect -11311 20303 -11111 20349
rect -11311 20107 -11111 20153
rect -11311 19911 -11111 19957
rect -11296 19692 -11196 19738
rect -11058 19735 -11001 20507
rect -10682 20494 -10088 20535
rect -10931 20303 -10831 20349
rect -10931 20107 -10831 20153
rect -10931 19911 -10831 19957
rect -11436 19640 -11258 19643
rect -11436 19594 -11196 19640
rect -11436 19592 -11258 19594
rect -11436 19449 -11379 19592
rect -11068 19566 -10994 19735
rect -10881 19692 -10781 19738
rect -10682 19644 -10634 20494
rect -10323 20400 -10223 20446
rect -10149 20399 -10089 20494
rect -9908 20400 -9808 20446
rect -9533 20434 -9486 20584
rect -9450 20486 -8613 20532
rect -9533 20388 -9150 20434
rect -10323 20302 -10223 20348
rect -9908 20302 -9808 20348
rect -10323 20204 -10223 20250
rect -9908 20204 -9808 20250
rect -9533 20238 -9486 20388
rect -7858 20338 -7812 20537
rect -8913 20290 -8613 20336
rect -8014 20292 -7812 20338
rect -9533 20192 -9150 20238
rect -9533 20191 -9449 20192
rect -9017 20176 -8959 20255
rect -7858 20240 -7812 20292
rect -7860 20194 -7683 20240
rect -10323 20106 -10223 20152
rect -9908 20106 -9808 20152
rect -9126 20122 -8959 20176
rect -7860 20142 -7812 20194
rect -10323 20008 -10223 20054
rect -9908 20008 -9808 20054
rect -10323 19910 -10223 19956
rect -9908 19910 -9808 19956
rect -9126 19902 -9072 20122
rect -9017 20096 -8959 20122
rect -8014 20096 -7812 20142
rect -7860 20044 -7812 20096
rect -7860 19998 -7683 20044
rect -10323 19812 -10223 19858
rect -10323 19714 -10223 19760
rect -10110 19717 -10036 19886
rect -9908 19812 -9808 19858
rect -9470 19848 -9072 19902
rect -10800 19640 -10634 19644
rect -10881 19594 -10634 19640
rect -10800 19583 -10634 19594
rect -11296 19496 -11196 19542
rect -10881 19496 -10781 19542
rect -10682 19453 -10634 19583
rect -10273 19495 -10173 19541
rect -11436 19444 -11258 19449
rect -10802 19444 -10634 19453
rect -11436 19398 -11196 19444
rect -10881 19398 -10634 19444
rect -11436 19249 -11379 19398
rect -10802 19392 -10634 19398
rect -11296 19300 -11196 19346
rect -10881 19300 -10781 19346
rect -10682 19257 -10634 19392
rect -10273 19299 -10173 19345
rect -11436 19248 -11239 19249
rect -10800 19248 -10634 19257
rect -11436 19202 -11196 19248
rect -10881 19202 -10634 19248
rect -11436 19198 -11239 19202
rect -11436 19057 -11379 19198
rect -10800 19196 -10634 19202
rect -11296 19104 -11196 19150
rect -10881 19104 -10781 19150
rect -11436 19052 -11264 19057
rect -10682 19052 -10634 19196
rect -10273 19103 -10173 19149
rect -11436 19007 -11196 19052
rect -11296 19006 -11196 19007
rect -10881 19006 -10634 19052
rect -10836 19004 -10634 19006
rect -10103 18945 -10046 19717
rect -9908 19714 -9808 19760
rect -9993 19495 -9793 19541
rect -9993 19299 -9793 19345
rect -9993 19103 -9793 19149
rect -10674 18887 -10614 18923
rect -10103 18888 -9811 18945
rect -10674 18827 -10147 18887
rect -10674 18791 -10614 18827
rect -10273 18658 -10173 18704
rect -9993 18658 -9793 18704
rect -11311 18560 -11111 18606
rect -10931 18560 -10831 18606
rect -10273 18462 -10173 18508
rect -9993 18462 -9793 18508
rect -11311 18364 -11111 18410
rect -10931 18364 -10831 18410
rect -10273 18266 -10173 18312
rect -9993 18266 -9793 18312
rect -11311 18168 -11111 18214
rect -10931 18168 -10831 18214
rect -10644 18054 -10507 18114
rect -10618 17788 -10554 18054
rect -9470 17788 -9416 19848
rect -9044 19755 -8998 19954
rect -7858 19946 -7812 19998
rect -8014 19900 -7812 19946
rect -9044 19709 -8742 19755
rect -9044 19657 -8998 19709
rect -9272 19611 -8996 19657
rect -6509 19643 -6452 23207
rect -6384 23003 -6184 23049
rect -6384 22807 -6184 22853
rect -6384 22611 -6184 22657
rect -6369 22392 -6269 22438
rect -6131 22435 -6074 23207
rect -5545 23196 -5164 23234
rect -6004 23003 -5904 23049
rect -6004 22807 -5904 22853
rect -6004 22611 -5904 22657
rect -5545 22469 -5499 23196
rect -5396 23100 -5296 23146
rect -5224 23088 -5164 23196
rect -4981 23100 -4881 23146
rect -5396 23002 -5296 23048
rect -4981 23002 -4881 23048
rect -5396 22904 -5296 22950
rect -4981 22904 -4881 22950
rect -5396 22806 -5296 22852
rect -4981 22806 -4881 22852
rect -5396 22708 -5296 22754
rect -4981 22708 -4881 22754
rect -5396 22610 -5296 22656
rect -4981 22610 -4881 22656
rect -5396 22512 -5296 22558
rect -6369 22294 -6269 22340
rect -6141 22266 -6067 22435
rect -5954 22392 -5854 22438
rect -5757 22423 -5499 22469
rect -5954 22337 -5854 22340
rect -5757 22337 -5711 22423
rect -5396 22414 -5296 22460
rect -5183 22417 -5109 22586
rect -4981 22512 -4881 22558
rect -5954 22295 -5711 22337
rect -5954 22294 -5854 22295
rect -6369 22196 -6269 22242
rect -5954 22196 -5854 22242
rect -6369 22098 -6269 22144
rect -5954 22141 -5854 22144
rect -5757 22141 -5711 22295
rect -5346 22195 -5246 22241
rect -5954 22099 -5711 22141
rect -5954 22098 -5854 22099
rect -6369 22000 -6269 22046
rect -5954 22000 -5854 22046
rect -6369 21902 -6269 21948
rect -5954 21946 -5854 21948
rect -5757 21946 -5711 22099
rect -5346 21999 -5246 22045
rect -5954 21904 -5711 21946
rect -5954 21902 -5854 21904
rect -6369 21804 -6269 21850
rect -5954 21804 -5854 21850
rect -5757 21755 -5711 21904
rect -5346 21803 -5246 21849
rect -6369 21706 -6269 21752
rect -5954 21709 -5711 21755
rect -5954 21706 -5854 21709
rect -5176 21645 -5119 22417
rect -4981 22414 -4881 22460
rect -5066 22195 -4866 22241
rect -5066 21999 -4866 22045
rect -5066 21803 -4866 21849
rect -5659 21599 -5599 21642
rect -5659 21539 -5235 21599
rect -5176 21588 -4884 21645
rect -5659 21510 -5599 21539
rect -5346 21358 -5246 21404
rect -5066 21358 -4866 21404
rect -6384 21260 -6184 21306
rect -6004 21260 -5904 21306
rect -5346 21162 -5246 21208
rect -5066 21162 -4866 21208
rect -6384 21064 -6184 21110
rect -6004 21064 -5904 21110
rect -5346 20966 -5246 21012
rect -5066 20966 -4866 21012
rect -6384 20868 -6184 20914
rect -6004 20868 -5904 20914
rect -5201 20789 -5141 20872
rect -5994 20788 -5135 20789
rect -6081 20729 -5135 20788
rect -6081 20728 -5949 20729
rect -5658 20673 -5598 20701
rect -6106 20613 -5598 20673
rect -5658 20564 -5598 20613
rect -6366 20507 -6074 20564
rect -5222 20535 -5162 20536
rect -6384 20303 -6184 20349
rect -6384 20107 -6184 20153
rect -6384 19911 -6184 19957
rect -6369 19692 -6269 19738
rect -6131 19735 -6074 20507
rect -5755 20494 -5161 20535
rect -6004 20303 -5904 20349
rect -6004 20107 -5904 20153
rect -6004 19911 -5904 19957
rect -6509 19640 -6331 19643
rect -9044 19559 -8996 19611
rect -7476 19585 -7093 19631
rect -9044 19513 -8742 19559
rect -9044 19461 -8996 19513
rect -8013 19487 -7176 19533
rect -9272 19415 -8996 19461
rect -7140 19435 -7093 19585
rect -9044 19363 -8998 19415
rect -7476 19389 -7093 19435
rect -9044 19317 -8742 19363
rect -8013 19291 -7713 19337
rect -7140 19239 -7093 19389
rect -7476 19193 -7093 19239
rect -7177 19192 -7093 19193
rect -6509 19594 -6269 19640
rect -6509 19592 -6331 19594
rect -6509 19449 -6452 19592
rect -6141 19566 -6067 19735
rect -5954 19692 -5854 19738
rect -5755 19644 -5707 20494
rect -5396 20400 -5296 20446
rect -5222 20399 -5162 20494
rect -4981 20400 -4881 20446
rect -5396 20302 -5296 20348
rect -4981 20302 -4881 20348
rect -5396 20204 -5296 20250
rect -4981 20204 -4881 20250
rect -5396 20106 -5296 20152
rect -4981 20106 -4881 20152
rect -5396 20008 -5296 20054
rect -4981 20008 -4881 20054
rect -5396 19910 -5296 19956
rect -4981 19910 -4881 19956
rect -5396 19812 -5296 19858
rect -5396 19714 -5296 19760
rect -5183 19717 -5109 19886
rect -4981 19812 -4881 19858
rect -5873 19640 -5707 19644
rect -5954 19594 -5707 19640
rect -5873 19583 -5707 19594
rect -6369 19496 -6269 19542
rect -5954 19496 -5854 19542
rect -5755 19453 -5707 19583
rect -5346 19495 -5246 19541
rect -6509 19444 -6331 19449
rect -5875 19444 -5707 19453
rect -6509 19398 -6269 19444
rect -5954 19398 -5707 19444
rect -6509 19249 -6452 19398
rect -5875 19392 -5707 19398
rect -6369 19300 -6269 19346
rect -5954 19300 -5854 19346
rect -5755 19257 -5707 19392
rect -5346 19299 -5246 19345
rect -6509 19248 -6312 19249
rect -5873 19248 -5707 19257
rect -6509 19202 -6269 19248
rect -5954 19202 -5707 19248
rect -6509 19198 -6312 19202
rect -10618 17734 -9416 17788
rect -6509 19057 -6452 19198
rect -5873 19196 -5707 19202
rect -6369 19104 -6269 19150
rect -5954 19104 -5854 19150
rect -6509 19052 -6337 19057
rect -5755 19052 -5707 19196
rect -5346 19103 -5246 19149
rect -6509 19007 -6269 19052
rect -6369 19006 -6269 19007
rect -5954 19006 -5707 19052
rect -5909 19004 -5707 19006
rect -5176 18945 -5119 19717
rect -4981 19714 -4881 19760
rect -5066 19495 -4866 19541
rect -5066 19299 -4866 19345
rect -5066 19103 -4866 19149
rect -5747 18887 -5687 18923
rect -5176 18888 -4884 18945
rect -7719 18654 -7565 18840
rect -5747 18827 -5220 18887
rect -5747 18791 -5687 18827
rect -5346 18658 -5246 18704
rect -5066 18658 -4866 18704
rect -7671 17856 -7607 18654
rect -6384 18560 -6184 18606
rect -6004 18560 -5904 18606
rect -5346 18462 -5246 18508
rect -5066 18462 -4866 18508
rect -6384 18364 -6184 18410
rect -6004 18364 -5904 18410
rect -5346 18266 -5246 18312
rect -5066 18266 -4866 18312
rect -6384 18168 -6184 18214
rect -6004 18168 -5904 18214
rect -5717 18054 -5580 18114
rect -5691 17856 -5627 18054
rect -7671 17792 -5627 17856
rect -11398 17158 -9002 17366
rect -11467 16670 -11395 16704
rect -11467 16605 -11247 16670
rect -11467 16599 -11395 16605
rect -12838 16348 -12792 16547
rect -12126 16368 -11526 16414
rect -12838 16302 -12636 16348
rect -12838 16250 -12792 16302
rect -12967 16204 -12790 16250
rect -12838 16152 -12790 16204
rect -12126 16156 -11526 16202
rect -12838 16106 -12636 16152
rect -12838 16054 -12790 16106
rect -12126 16058 -11526 16104
rect -12967 16008 -12790 16054
rect -12838 15956 -12792 16008
rect -12126 15960 -11526 16006
rect -12838 15910 -12636 15956
rect -12126 15749 -11526 15795
rect -11312 15650 -11247 16605
rect -11214 16285 -10914 16331
rect -9686 16451 -9421 16487
rect -8866 16451 -8601 16482
rect -9686 16263 -8601 16451
rect -6467 16670 -6395 16704
rect -6467 16605 -6247 16670
rect -6467 16599 -6395 16605
rect -7838 16348 -7792 16547
rect -7126 16368 -6526 16414
rect -7838 16302 -7636 16348
rect -9686 16219 -9421 16263
rect -8866 16214 -8601 16263
rect -7838 16250 -7792 16302
rect -7967 16204 -7790 16250
rect -7838 16152 -7790 16204
rect -7126 16156 -6526 16202
rect -7838 16106 -7636 16152
rect -7838 16054 -7790 16106
rect -7126 16058 -6526 16104
rect -7967 16008 -7790 16054
rect -7838 15956 -7792 16008
rect -7126 15960 -6526 16006
rect -7838 15910 -7636 15956
rect -11214 15847 -10914 15893
rect -7126 15749 -6526 15795
rect -6312 15650 -6247 16605
rect -6214 16285 -5914 16331
rect -6214 15847 -5914 15893
rect -13557 15595 -13174 15641
rect -8557 15595 -8174 15641
rect -13557 15445 -13510 15595
rect -13474 15497 -12637 15543
rect -13557 15399 -13174 15445
rect -13557 15249 -13510 15399
rect -11882 15349 -11836 15548
rect -12937 15301 -12637 15347
rect -12038 15303 -11836 15349
rect -13557 15203 -13174 15249
rect -13557 15202 -13473 15203
rect -13041 15187 -12983 15266
rect -11882 15251 -11836 15303
rect -8557 15445 -8510 15595
rect -8474 15497 -7637 15543
rect -8557 15399 -8174 15445
rect -11884 15205 -11707 15251
rect -8557 15249 -8510 15399
rect -6882 15349 -6836 15548
rect -7937 15301 -7637 15347
rect -7038 15303 -6836 15349
rect -13150 15133 -12983 15187
rect -11884 15153 -11836 15205
rect -8557 15203 -8174 15249
rect -8557 15202 -8473 15203
rect -8041 15187 -7983 15266
rect -6882 15251 -6836 15303
rect -6884 15205 -6707 15251
rect -13150 14913 -13096 15133
rect -13041 15107 -12983 15133
rect -12038 15107 -11836 15153
rect -8150 15133 -7983 15187
rect -6884 15153 -6836 15205
rect -11884 15055 -11836 15107
rect -11884 15009 -11707 15055
rect -13494 14859 -13096 14913
rect -13900 13870 -13764 13930
rect -13494 13870 -13440 14859
rect -13068 14766 -13022 14965
rect -11882 14957 -11836 15009
rect -12038 14911 -11836 14957
rect -8150 14913 -8096 15133
rect -8041 15107 -7983 15133
rect -7038 15107 -6836 15153
rect -6884 15055 -6836 15107
rect -6884 15009 -6707 15055
rect -8494 14859 -8096 14913
rect -13068 14720 -12766 14766
rect -13068 14668 -13022 14720
rect -13296 14622 -13020 14668
rect -13068 14570 -13020 14622
rect -11500 14596 -11117 14642
rect -13068 14524 -12766 14570
rect -13068 14472 -13020 14524
rect -12037 14498 -11200 14544
rect -13296 14426 -13020 14472
rect -11164 14446 -11117 14596
rect -13068 14374 -13022 14426
rect -11500 14400 -11117 14446
rect -13068 14328 -12766 14374
rect -12037 14302 -11737 14348
rect -11164 14250 -11117 14400
rect -11500 14204 -11117 14250
rect -11201 14203 -11117 14204
rect -13150 14146 -13000 14172
rect -13150 14092 -11542 14146
rect -13150 14042 -13000 14092
rect -13900 13816 -13440 13870
rect -11596 13949 -11542 14092
rect -8494 14068 -8440 14859
rect -8068 14766 -8022 14965
rect -6882 14957 -6836 15009
rect -7038 14911 -6836 14957
rect -8068 14720 -7766 14766
rect -8068 14668 -8022 14720
rect -8296 14622 -8020 14668
rect -8068 14570 -8020 14622
rect -6500 14596 -6117 14642
rect -8068 14524 -7766 14570
rect -8068 14472 -8020 14524
rect -7037 14498 -6200 14544
rect -8296 14426 -8020 14472
rect -6164 14446 -6117 14596
rect -8068 14374 -8022 14426
rect -6500 14400 -6117 14446
rect -8068 14328 -7766 14374
rect -7037 14302 -6737 14348
rect -6164 14250 -6117 14400
rect -6500 14204 -6117 14250
rect -6201 14203 -6117 14204
rect -13900 13786 -13764 13816
rect -9208 13828 -8440 14068
rect -8150 14146 -8000 14172
rect -8150 14092 -6542 14146
rect -8150 14042 -8000 14092
rect -6596 13949 -6542 14092
rect -6001 14076 -5943 14141
rect -6062 13995 -5943 14076
rect -8494 13816 -8440 13828
rect -14155 13701 -14018 13747
rect -11754 13701 -11631 13723
rect -6062 13718 -6027 13995
rect -14155 13609 -11631 13701
rect -7167 13683 -6027 13718
rect -5976 13713 -5930 13912
rect -8497 13627 -8297 13673
rect -7789 13627 -7589 13673
rect -14253 13547 -14195 13608
rect -11754 13606 -11631 13609
rect -13159 13547 -13022 13565
rect -14253 13508 -13022 13547
rect -14253 13471 -14195 13508
rect -13159 13507 -13022 13508
rect -13648 13465 -13511 13480
rect -11456 13465 -11398 13482
rect -13648 13430 -11398 13465
rect -13648 13422 -13511 13430
rect -11456 13345 -11398 13430
rect -11208 13307 -10808 13353
rect -11208 13209 -10808 13255
rect -8497 13214 -8197 13260
rect -11208 13111 -10808 13157
rect -8497 13116 -8197 13162
rect -11700 12998 -11500 13044
rect -8497 13018 -8197 13064
rect -11208 12900 -10808 12946
rect -8497 12905 -8197 12951
rect -7789 12889 -7589 12935
rect -8497 12807 -8197 12853
rect -8497 12709 -8197 12755
rect -7789 12693 -7589 12739
rect -8496 12595 -8196 12641
rect -13562 12540 -13425 12555
rect -11455 12540 -11397 12551
rect -13562 12505 -11397 12540
rect -13562 12497 -13425 12505
rect -11455 12414 -11397 12505
rect -7789 12497 -7589 12543
rect -11207 12402 -10807 12448
rect -8496 12399 -8196 12445
rect -11207 12304 -10807 12350
rect -11207 12206 -10807 12252
rect -8052 12222 -7915 12271
rect -7167 12222 -7132 13683
rect -5976 13667 -5774 13713
rect -5976 13615 -5930 13667
rect -6105 13569 -5928 13615
rect -5976 13517 -5928 13569
rect -5976 13471 -5774 13517
rect -5976 13419 -5928 13471
rect -6105 13373 -5928 13419
rect -5976 13321 -5930 13373
rect -5976 13275 -5774 13321
rect -6695 12960 -6312 13006
rect -6695 12810 -6648 12960
rect -6612 12862 -5775 12908
rect -6695 12764 -6312 12810
rect -6695 12614 -6648 12764
rect -6075 12666 -5775 12712
rect -6695 12568 -6312 12614
rect -6695 12567 -6611 12568
rect -8052 12213 -7132 12222
rect -7961 12187 -7132 12213
rect -8183 12156 -8046 12174
rect -11699 12093 -11499 12139
rect -8183 12121 -6477 12156
rect -8183 12116 -8046 12121
rect -11207 11995 -10807 12041
rect -8280 11902 -8143 11960
rect -13480 11766 -12802 11856
rect -13289 11680 -12989 11726
rect -12892 11629 -12802 11766
rect -7885 11771 -7839 11970
rect -6512 11843 -6477 12121
rect -6561 11797 -6361 11843
rect -5853 11797 -5653 11843
rect -7885 11725 -7683 11771
rect -7885 11673 -7839 11725
rect -11804 11629 -11746 11664
rect -13896 11582 -13696 11628
rect -12892 11539 -11746 11629
rect -8014 11627 -7837 11673
rect -7885 11575 -7837 11627
rect -13289 11484 -12989 11530
rect -11804 11527 -11746 11539
rect -11478 11506 -10878 11552
rect -7885 11529 -7683 11575
rect -7885 11477 -7837 11529
rect -13896 11386 -13696 11432
rect -13288 11370 -12988 11416
rect -11478 11408 -10878 11454
rect -8014 11431 -7837 11477
rect -7885 11379 -7839 11431
rect -6561 11384 -6261 11430
rect -13288 11272 -12988 11318
rect -11478 11310 -10878 11356
rect -7885 11333 -7683 11379
rect -13896 11190 -13696 11236
rect -13288 11174 -12988 11220
rect -6561 11286 -6261 11332
rect -11478 11197 -10878 11243
rect -6561 11188 -6261 11234
rect -13288 11061 -12988 11107
rect -12042 11083 -11842 11129
rect -11478 11099 -10878 11145
rect -6561 11075 -6261 11121
rect -13288 10963 -12988 11009
rect -11478 11001 -10878 11047
rect -8604 11018 -8221 11064
rect -5853 11059 -5653 11105
rect -13288 10865 -12988 10911
rect -12042 10887 -11842 10933
rect -8604 10868 -8557 11018
rect -6561 10977 -6261 11023
rect -8521 10920 -7684 10966
rect -6561 10879 -6261 10925
rect -11478 10789 -10878 10835
rect -8604 10822 -8221 10868
rect -5853 10863 -5653 10909
rect -14283 10496 -14167 10561
rect -13896 10496 -13696 10498
rect -14283 10453 -13696 10496
rect -14283 10403 -14167 10453
rect -13896 10452 -13696 10453
rect -13188 10452 -12988 10498
rect -8604 10672 -8557 10822
rect -7984 10724 -7684 10770
rect -6560 10765 -6260 10811
rect -8604 10626 -8221 10672
rect -5853 10667 -5653 10713
rect -8604 10625 -8520 10626
rect -6560 10569 -6260 10615
rect -157 10922 87 12457
rect 93931 12460 95152 38495
rect -66 10473 -13 10922
rect 15082 10499 18555 10502
rect 15069 10473 18555 10499
rect -66 10420 18555 10473
rect 15069 10340 18555 10420
rect 15069 10288 18556 10340
rect 15069 10173 15122 10288
rect 16304 10178 16350 10288
rect 17686 10272 18556 10288
rect 14785 10127 14985 10173
rect 15069 10127 15388 10173
rect 16299 10132 16618 10178
rect 15069 9657 15115 10127
rect 15188 9869 15388 9915
rect 15588 9869 15788 9915
rect 16018 9874 16218 9920
rect 16299 9662 16345 10132
rect 16418 9874 16618 9920
rect 16818 9874 17018 9920
rect 14785 9611 14985 9657
rect 15069 9611 15388 9657
rect 16299 9616 16618 9662
rect 15069 9141 15115 9611
rect 15188 9353 15388 9399
rect 15588 9353 15788 9399
rect 16018 9358 16218 9404
rect 16299 9146 16345 9616
rect 17686 9560 69834 10272
rect 94130 10098 94998 12460
rect 91756 9540 94998 10098
rect 16418 9358 16618 9404
rect 16818 9358 17018 9404
rect 14785 9095 14985 9141
rect 15069 9095 15388 9141
rect 16299 9100 16618 9146
rect 13898 8915 14773 8919
rect 6966 8466 7312 8756
rect 13898 8737 14775 8915
rect -5845 2483 -5539 2764
rect -613 2710 1457 2816
rect -9391 1504 -9345 1975
rect -9155 1504 -9109 1975
rect -8919 1504 -8873 1975
rect -8683 1504 -8637 1975
rect -8447 1504 -8401 1975
rect -8211 1504 -8165 1975
rect -7975 1504 -7929 1975
rect -7739 1504 -7693 1975
rect -7373 1504 -7327 1975
rect -7137 1504 -7091 1975
rect -6901 1504 -6855 1975
rect -6665 1504 -6619 1975
rect -6299 1504 -6253 1975
rect -6063 1504 -6017 1975
rect -5742 1521 -5581 2483
rect -3492 1837 -3446 2037
rect -3296 1837 -3250 2037
rect -3100 1837 -3054 2037
rect -2642 1837 -2596 2037
rect -2446 1837 -2400 2037
rect -2250 1837 -2204 2037
rect -2094 1837 -2048 2037
rect -1996 1793 -1950 2037
rect -1898 1837 -1852 2037
rect -1800 1793 -1754 2037
rect -1702 1837 -1656 2037
rect -1604 1793 -1558 2037
rect -1506 1837 -1460 2037
rect -1408 1793 -1362 2037
rect -1310 1837 -1264 2037
rect -1996 1747 -1162 1793
rect -3590 1557 -3544 1657
rect -3492 1557 -3446 1657
rect -3394 1557 -3348 1657
rect -3296 1557 -3250 1657
rect -3198 1557 -3152 1657
rect -3100 1557 -3054 1657
rect -2937 1621 -2805 1665
rect -9506 1430 -7561 1504
rect -7500 1430 -6490 1504
rect -6429 1430 -6012 1504
rect -7732 1302 -7686 1430
rect -13317 767 -13271 1167
rect -13199 767 -13153 1167
rect -13081 767 -13035 1167
rect -12963 767 -12917 1167
rect -12845 767 -12799 1167
rect -12727 767 -12681 1167
rect -12609 767 -12563 1167
rect -12491 767 -12445 1167
rect -12373 767 -12327 1167
rect -12255 767 -12209 1167
rect -12137 767 -12091 1167
rect -12019 767 -11973 1167
rect -11901 767 -11855 1167
rect -11783 767 -11737 1167
rect -11665 767 -11619 1167
rect -11547 767 -11501 1167
rect -11429 767 -11383 1167
rect -11311 767 -11265 1167
rect -11193 767 -11147 1167
rect -11075 767 -11029 1167
rect -10957 767 -10911 1167
rect -10839 767 -10793 1167
rect -10721 767 -10675 1167
rect -10603 767 -10557 1167
rect -10485 767 -10439 1167
rect -10367 767 -10321 1167
rect -10249 767 -10203 1167
rect -10131 767 -10085 1167
rect -10013 767 -9967 1167
rect -9895 767 -9849 1167
rect -9777 767 -9731 1167
rect -9541 767 -9495 1167
rect -9305 767 -9259 1167
rect -9069 767 -9023 1167
rect -8833 767 -8787 1167
rect -8597 767 -8551 1167
rect -8361 767 -8315 1167
rect -8125 767 -8079 1167
rect -7771 1256 -7017 1302
rect -6750 1290 -6704 1430
rect -7889 767 -7843 1167
rect -7771 767 -7725 1256
rect -7653 767 -7607 1167
rect -7535 767 -7489 1256
rect -7417 767 -7371 1167
rect -7299 767 -7253 1256
rect -7181 767 -7135 1167
rect -7063 767 -7017 1256
rect -6827 1244 -6545 1290
rect -6945 767 -6899 1167
rect -6827 767 -6781 1244
rect -6709 767 -6663 1167
rect -6591 767 -6545 1244
rect -6473 767 -6427 1167
rect -6355 767 -6309 1430
rect -5774 1415 -5574 1521
rect -4212 1498 -4099 1535
rect -2849 1521 -2805 1621
rect -2740 1557 -2694 1657
rect -2642 1557 -2596 1657
rect -2544 1557 -2498 1657
rect -2446 1557 -2400 1657
rect -2348 1557 -2302 1657
rect -2250 1557 -2204 1657
rect -2094 1521 -2048 1691
rect -3572 1498 -3060 1502
rect -4212 1461 -3060 1498
rect -3572 1449 -3060 1461
rect -2849 1477 -2047 1521
rect -1996 1491 -1950 1747
rect -1898 1491 -1852 1691
rect -1800 1491 -1754 1747
rect -1702 1491 -1656 1691
rect -1604 1491 -1558 1747
rect -1506 1491 -1460 1691
rect -1408 1491 -1362 1747
rect -1310 1491 -1264 1691
rect -1208 1575 -1162 1747
rect -613 1575 -456 2710
rect 738 2401 975 2497
rect 870 2139 975 2401
rect 1021 2405 1257 2501
rect 1021 2145 1112 2405
rect 1351 2139 1457 2710
rect 1823 2405 2012 2501
rect 1921 2238 2012 2405
rect 1852 2160 2285 2238
rect 619 2001 665 2085
rect 865 1915 911 2110
rect 983 1990 1029 2110
rect 1101 1990 1147 2110
rect 1307 1990 1353 2110
rect 1395 1990 1441 2110
rect 1597 1995 1643 2115
rect 1685 2081 1731 2115
rect 1823 2081 1869 2122
rect 1685 2010 1869 2081
rect 1685 1995 1731 2010
rect 865 1869 1001 1915
rect 619 1769 665 1821
rect -2849 1415 -2805 1477
rect -5774 1371 -2805 1415
rect -1208 1423 -456 1575
rect 411 1692 665 1769
rect -5774 1352 -5574 1371
rect -6237 767 -6191 1167
rect -2740 1142 -2694 1242
rect -2642 1142 -2596 1242
rect -2544 1142 -2498 1242
rect -2446 1142 -2400 1242
rect -2348 1142 -2302 1242
rect -2250 1142 -2204 1242
rect -13350 548 -6080 721
rect -12759 -135 -12272 548
rect -11199 -135 -10712 548
rect -10006 -135 -9519 548
rect -8823 -135 -8336 548
rect -7809 -135 -7322 548
rect -1996 1052 -1950 1308
rect -1800 1052 -1754 1308
rect -1604 1052 -1558 1308
rect -1408 1052 -1362 1308
rect -1208 1052 -1162 1423
rect -1996 1006 -1162 1052
rect -2642 762 -2596 962
rect -2446 762 -2400 962
rect -2250 762 -2204 962
rect -1996 762 -1950 1006
rect -1800 762 -1754 1006
rect -1604 762 -1558 1006
rect -1408 762 -1362 1006
rect 411 308 488 1692
rect 619 1653 665 1692
rect 955 1625 1001 1869
rect 1499 1854 1590 1933
rect 1638 1899 1733 1925
rect 1823 1905 1869 2010
rect 2059 2002 2105 2122
rect 2295 2002 2341 2122
rect 2582 2001 2628 2085
rect 2891 2001 2937 2085
rect 1638 1857 1794 1899
rect 1823 1859 1994 1905
rect 1131 1699 1177 1819
rect 1307 1699 1353 1819
rect 1117 1625 1189 1655
rect 1294 1625 1366 1654
rect 1508 1639 1554 1819
rect 1596 1639 1642 1819
rect 955 1579 1366 1625
rect 1117 1574 1189 1579
rect 1120 1571 1186 1574
rect 1294 1573 1366 1579
rect 1297 1570 1363 1573
rect 1760 1453 1794 1857
rect 1948 1639 1994 1859
rect 2582 1653 2628 1821
rect 2891 1653 2937 1821
rect 1508 1407 1794 1453
rect 1120 1288 1186 1291
rect 1297 1289 1363 1292
rect 1117 1283 1189 1288
rect 1294 1283 1366 1289
rect 955 1237 1366 1283
rect 619 1041 665 1209
rect 955 993 1001 1237
rect 1117 1207 1189 1237
rect 1294 1208 1366 1237
rect 1131 1043 1177 1163
rect 1307 1043 1353 1163
rect 1508 1043 1554 1407
rect 1596 1043 1642 1223
rect 865 947 1001 993
rect 619 777 665 861
rect 865 752 911 947
rect 1638 937 1733 1005
rect 1948 1003 1994 1223
rect 2582 1041 2628 1209
rect 2891 1041 2937 1209
rect 4607 2013 4653 2213
rect 4803 2013 4849 2213
rect 4999 2013 5045 2213
rect 5457 2013 5503 2213
rect 5653 2013 5699 2213
rect 5849 2013 5895 2213
rect 6005 2013 6051 2213
rect 6103 1969 6149 2213
rect 6201 2013 6247 2213
rect 6299 1969 6345 2213
rect 6397 2013 6443 2213
rect 6495 1969 6541 2213
rect 6593 2013 6639 2213
rect 6691 1969 6737 2213
rect 6789 2013 6835 2213
rect 7080 2079 7229 8466
rect 7289 8017 7635 8307
rect 6103 1923 6937 1969
rect 4607 1733 4653 1833
rect 4803 1733 4849 1833
rect 4999 1733 5045 1833
rect 5162 1797 5294 1841
rect 5250 1697 5294 1797
rect 5457 1733 5503 1833
rect 5653 1733 5699 1833
rect 5849 1733 5895 1833
rect 6005 1697 6051 1867
rect 5250 1653 6052 1697
rect 6103 1667 6149 1923
rect 6201 1667 6247 1867
rect 6299 1667 6345 1923
rect 6397 1667 6443 1867
rect 6495 1667 6541 1923
rect 6593 1667 6639 1867
rect 6691 1667 6737 1923
rect 6789 1667 6835 1867
rect 6891 1670 6937 1923
rect 7054 1845 7303 2079
rect 7341 1680 7460 8017
rect 8996 6696 9042 7496
rect 10712 6696 10758 7496
rect 12158 6696 12204 7496
rect 9032 5643 9078 6443
rect 10748 5643 10794 6443
rect 13898 5964 14080 8737
rect 14547 8736 14775 8737
rect 15079 6970 15125 9095
rect 15726 8848 16117 8894
rect 16226 8605 16396 8743
rect 14997 6756 15211 6970
rect 16250 6623 16388 8605
rect 16227 6444 16406 6623
rect 13866 5703 14130 5964
rect 12464 4643 12510 5443
rect 7730 1786 7776 2257
rect 7966 1786 8012 2257
rect 8332 1786 8378 2257
rect 8568 1786 8614 2257
rect 8804 1786 8850 2257
rect 9040 1786 9086 2257
rect 9406 1786 9452 2257
rect 9642 1786 9688 2257
rect 9878 1786 9924 2257
rect 10114 1786 10160 2257
rect 10350 1786 10396 2257
rect 10586 1786 10632 2257
rect 10822 1786 10868 2257
rect 11058 1786 11104 2257
rect 7725 1712 8142 1786
rect 8203 1712 9213 1786
rect 9274 1712 11219 1786
rect 7337 1670 7470 1680
rect 3990 1591 4106 1638
rect 5250 1591 5294 1653
rect 3990 1547 5294 1591
rect 6891 1624 7470 1670
rect 3990 1499 4106 1547
rect 5457 1318 5503 1418
rect 5653 1318 5699 1418
rect 5849 1318 5895 1418
rect 1823 957 1994 1003
rect 983 752 1029 872
rect 1101 752 1147 872
rect 1307 752 1353 872
rect 1395 752 1441 872
rect 1597 747 1643 867
rect 1685 852 1731 867
rect 1823 852 1869 957
rect 1685 781 1869 852
rect 1685 747 1731 781
rect 1823 740 1869 781
rect 2059 740 2105 860
rect 2295 740 2341 860
rect 870 461 975 723
rect 738 365 975 461
rect 1021 457 1112 717
rect 1021 362 1257 457
rect 1020 361 1257 362
rect 1020 308 1112 361
rect 411 231 1112 308
rect -13197 -453 -7163 -135
rect -25553 -1050 -25165 -654
rect -26907 -11153 -25983 -10980
rect -27809 -11705 -25983 -11153
rect -27809 -42856 -27257 -11705
rect -26907 -11904 -25983 -11705
rect -25501 -14108 -25219 -1050
rect -12865 -10939 -11924 -453
rect -24248 -11880 -11923 -10939
rect -25931 -14876 -24870 -14108
rect -25501 -22779 -25219 -14876
rect -12865 -14969 -11924 -11880
rect -10614 -14969 -9673 -453
rect -8935 -14969 -7994 -453
rect 1351 106 1457 723
rect 1852 624 2285 702
rect 1921 457 2012 624
rect 2582 777 2628 861
rect 2891 777 2937 861
rect 3563 973 3725 1039
rect 3563 929 3812 973
rect 3563 885 3725 929
rect 1823 361 2012 457
rect -2521 0 1457 106
rect -6059 -378 -5507 -276
rect -5976 -957 -5800 -784
rect -5544 -873 -5507 -378
rect -4960 -535 -4914 -335
rect -4764 -535 -4718 -335
rect -4568 -535 -4522 -335
rect -4110 -535 -4064 -335
rect -3914 -535 -3868 -335
rect -3718 -535 -3672 -335
rect -3562 -535 -3516 -335
rect -3464 -579 -3418 -335
rect -3366 -535 -3320 -335
rect -3268 -579 -3222 -335
rect -3170 -535 -3124 -335
rect -3072 -579 -3026 -335
rect -2974 -535 -2928 -335
rect -2876 -579 -2830 -335
rect -2778 -535 -2732 -335
rect -3464 -625 -2630 -579
rect -5058 -815 -5012 -715
rect -4960 -815 -4914 -715
rect -4862 -815 -4816 -715
rect -4764 -815 -4718 -715
rect -4666 -815 -4620 -715
rect -4568 -815 -4522 -715
rect -4405 -751 -4273 -707
rect -4317 -851 -4273 -751
rect -4208 -815 -4162 -715
rect -4110 -815 -4064 -715
rect -4012 -815 -3966 -715
rect -3914 -815 -3868 -715
rect -3816 -815 -3770 -715
rect -3718 -815 -3672 -715
rect -3562 -851 -3516 -681
rect -5056 -873 -4533 -861
rect -5544 -910 -4533 -873
rect -5056 -922 -4533 -910
rect -4317 -895 -3515 -851
rect -3464 -881 -3418 -625
rect -3366 -881 -3320 -681
rect -3268 -881 -3222 -625
rect -3170 -881 -3124 -681
rect -3072 -881 -3026 -625
rect -2974 -881 -2928 -681
rect -2876 -881 -2830 -625
rect -2778 -881 -2732 -681
rect -2676 -779 -2630 -625
rect -2521 -665 -2415 0
rect -2521 -779 -2422 -665
rect -4317 -957 -4273 -895
rect -5976 -1001 -4273 -957
rect -2676 -924 -2422 -779
rect -5976 -1005 -5800 -1001
rect -4185 -1050 -4062 -989
rect -4317 -1094 -3515 -1050
rect -4317 -1194 -4273 -1094
rect -5249 -1238 -4273 -1194
rect -4208 -1230 -4162 -1130
rect -4110 -1230 -4064 -1130
rect -4012 -1230 -3966 -1130
rect -3914 -1230 -3868 -1130
rect -3816 -1230 -3770 -1130
rect -3718 -1230 -3672 -1130
rect -3562 -1264 -3516 -1094
rect -3464 -1320 -3418 -1064
rect -3366 -1264 -3320 -1064
rect -3268 -1320 -3222 -1064
rect -3170 -1264 -3124 -1064
rect -3072 -1320 -3026 -1064
rect -2974 -1264 -2928 -1064
rect -2876 -1320 -2830 -1064
rect -2778 -1264 -2732 -1064
rect -2676 -1320 -2630 -924
rect -3464 -1366 -2630 -1320
rect -4110 -1610 -4064 -1410
rect -3914 -1610 -3868 -1410
rect -3718 -1610 -3672 -1410
rect -3562 -1610 -3516 -1410
rect -3464 -1610 -3418 -1366
rect -3366 -1610 -3320 -1410
rect -3268 -1610 -3222 -1366
rect -3170 -1610 -3124 -1410
rect -3072 -1610 -3026 -1366
rect -2974 -1610 -2928 -1410
rect -2876 -1610 -2830 -1366
rect -2778 -1610 -2732 -1410
rect 3768 -1099 3812 929
rect 6103 1228 6149 1484
rect 6299 1228 6345 1484
rect 6495 1228 6541 1484
rect 6691 1228 6737 1484
rect 6891 1228 6937 1624
rect 7337 1562 7470 1624
rect 7061 1355 7270 1554
rect 6103 1182 6937 1228
rect 5457 938 5503 1138
rect 5653 938 5699 1138
rect 5849 938 5895 1138
rect 6103 938 6149 1182
rect 6299 938 6345 1182
rect 6495 938 6541 1182
rect 6691 938 6737 1182
rect 4622 -677 4668 -477
rect 4818 -677 4864 -477
rect 5014 -677 5060 -477
rect 5472 -677 5518 -477
rect 5668 -677 5714 -477
rect 5864 -677 5910 -477
rect 6020 -677 6066 -477
rect 6118 -721 6164 -477
rect 6216 -677 6262 -477
rect 6314 -721 6360 -477
rect 6412 -677 6458 -477
rect 6510 -721 6556 -477
rect 6608 -677 6654 -477
rect 6706 -721 6752 -477
rect 6804 -677 6850 -477
rect 6118 -767 6952 -721
rect 4622 -957 4668 -857
rect 4818 -957 4864 -857
rect 5014 -957 5060 -857
rect 5177 -893 5309 -849
rect 5265 -993 5309 -893
rect 5472 -957 5518 -857
rect 5668 -957 5714 -857
rect 5864 -957 5910 -857
rect 6020 -993 6066 -823
rect 5265 -1037 6067 -993
rect 6118 -1023 6164 -767
rect 6216 -1023 6262 -823
rect 6314 -1023 6360 -767
rect 6412 -1023 6458 -823
rect 6510 -1023 6556 -767
rect 6608 -1023 6654 -823
rect 6706 -1023 6752 -767
rect 6804 -1023 6850 -823
rect 6906 -1020 6952 -767
rect 7131 -1020 7230 1355
rect 8022 1049 8068 1712
rect 8417 1572 8463 1712
rect 9399 1584 9445 1712
rect 8258 1526 8540 1572
rect 8258 1049 8304 1526
rect 8494 1049 8540 1526
rect 8730 1538 9484 1584
rect 8730 1049 8776 1538
rect 8966 1049 9012 1538
rect 9202 1049 9248 1538
rect 9438 1049 9484 1538
rect 7689 -970 7735 -499
rect 7925 -970 7971 -499
rect 8291 -970 8337 -499
rect 8527 -970 8573 -499
rect 8763 -970 8809 -499
rect 8999 -970 9045 -499
rect 9365 -970 9411 -499
rect 9601 -970 9647 -499
rect 9837 -970 9883 -499
rect 10073 -970 10119 -499
rect 10309 -970 10355 -499
rect 10545 -970 10591 -499
rect 10781 -970 10827 -499
rect 11017 -970 11063 -499
rect 5265 -1099 5309 -1037
rect 3768 -1143 5309 -1099
rect 6906 -1066 7412 -1020
rect 7684 -1044 8101 -970
rect 8162 -1044 9172 -970
rect 9233 -1044 11178 -970
rect 5472 -1372 5518 -1272
rect 5668 -1372 5714 -1272
rect 5864 -1372 5910 -1272
rect 6118 -1462 6164 -1206
rect 6314 -1462 6360 -1206
rect 6510 -1462 6556 -1206
rect 6706 -1462 6752 -1206
rect 6906 -1462 6952 -1066
rect 7334 -1093 7412 -1066
rect 7334 -1207 7443 -1093
rect 6118 -1508 6952 -1462
rect 5472 -1752 5518 -1552
rect 5668 -1752 5714 -1552
rect 5864 -1752 5910 -1552
rect 6118 -1752 6164 -1508
rect 6314 -1752 6360 -1508
rect 6510 -1752 6556 -1508
rect 6706 -1752 6752 -1508
rect 7981 -1707 8027 -1044
rect 8376 -1184 8422 -1044
rect 9358 -1172 9404 -1044
rect 8217 -1230 8499 -1184
rect 8217 -1707 8263 -1230
rect 8453 -1707 8499 -1230
rect 8689 -1218 9443 -1172
rect 8689 -1707 8735 -1218
rect 8925 -1707 8971 -1218
rect 9161 -1707 9207 -1218
rect 9397 -1707 9443 -1218
rect 19201 6620 19643 7085
rect 22939 6666 23303 7116
rect 18791 5216 19168 5573
rect 18861 -594 19153 5216
rect 19341 2756 19470 6620
rect 19886 3178 19932 3378
rect 20082 3178 20128 3378
rect 20278 3178 20324 3378
rect 20736 3178 20782 3378
rect 20932 3178 20978 3378
rect 21128 3178 21174 3378
rect 21284 3178 21330 3378
rect 21382 3134 21428 3378
rect 21480 3178 21526 3378
rect 21578 3134 21624 3378
rect 21676 3178 21722 3378
rect 21774 3134 21820 3378
rect 21872 3178 21918 3378
rect 21970 3134 22016 3378
rect 22068 3178 22114 3378
rect 21382 3088 22216 3134
rect 19886 2898 19932 2998
rect 20082 2898 20128 2998
rect 20278 2898 20324 2998
rect 20441 2962 20573 3006
rect 20529 2862 20573 2962
rect 20736 2898 20782 2998
rect 20932 2898 20978 2998
rect 21128 2898 21174 2998
rect 21284 2862 21330 3032
rect 20529 2818 21331 2862
rect 21382 2832 21428 3088
rect 21480 2832 21526 3032
rect 21578 2832 21624 3088
rect 21676 2832 21722 3032
rect 21774 2832 21820 3088
rect 21872 2832 21918 3032
rect 21970 2832 22016 3088
rect 22068 2832 22114 3032
rect 22170 2875 22216 3088
rect 22316 2875 22554 2900
rect 20529 2756 20573 2818
rect 19341 2712 20573 2756
rect 22170 2745 22554 2875
rect 19341 2700 19470 2712
rect 20736 2483 20782 2583
rect 20932 2483 20978 2583
rect 21128 2483 21174 2583
rect 21382 2393 21428 2649
rect 21578 2393 21624 2649
rect 21774 2393 21820 2649
rect 21970 2393 22016 2649
rect 22170 2393 22216 2745
rect 22316 2711 22554 2745
rect 21382 2347 22216 2393
rect 20736 2103 20782 2303
rect 20932 2103 20978 2303
rect 21128 2103 21174 2303
rect 21382 2103 21428 2347
rect 21578 2103 21624 2347
rect 21774 2103 21820 2347
rect 21970 2103 22016 2347
rect 20058 -172 20104 28
rect 20254 -172 20300 28
rect 20450 -172 20496 28
rect 20908 -172 20954 28
rect 21104 -172 21150 28
rect 21300 -172 21346 28
rect 21456 -172 21502 28
rect 21554 -216 21600 28
rect 21652 -172 21698 28
rect 21750 -216 21796 28
rect 21848 -172 21894 28
rect 21946 -216 21992 28
rect 22044 -172 22090 28
rect 22142 -216 22188 28
rect 22240 -172 22286 28
rect 21554 -262 22388 -216
rect 20058 -452 20104 -352
rect 20254 -452 20300 -352
rect 20450 -452 20496 -352
rect 20613 -388 20745 -344
rect 20701 -488 20745 -388
rect 20908 -452 20954 -352
rect 21104 -452 21150 -352
rect 21300 -452 21346 -352
rect 21456 -488 21502 -318
rect 20701 -532 21503 -488
rect 21554 -518 21600 -262
rect 21652 -518 21698 -318
rect 21750 -518 21796 -262
rect 21848 -518 21894 -318
rect 21946 -518 21992 -262
rect 22044 -518 22090 -318
rect 22142 -518 22188 -262
rect 22240 -518 22286 -318
rect 22342 -345 22388 -262
rect 22342 -353 22513 -345
rect 23046 -353 23217 6666
rect 26324 3017 38590 3153
rect 25061 2295 25333 2372
rect 25947 2295 26150 2357
rect 25061 2124 26150 2295
rect 25061 2085 25333 2124
rect 25947 2092 26150 2124
rect 26324 1094 26460 3017
rect 26278 836 26470 1094
rect 27601 2571 32111 2652
rect 27601 2278 27682 2571
rect 27272 2226 27682 2278
rect 27791 2226 27952 2240
rect 27272 2171 27952 2226
rect 29191 2179 29269 2195
rect 27272 2145 27652 2171
rect 27791 2161 27952 2171
rect 29075 2153 29269 2179
rect 28016 2124 29269 2153
rect 28016 1405 28054 2124
rect 28103 1857 28149 2057
rect 28103 1405 28149 1668
rect 28419 1857 28465 2124
rect 28419 1468 28465 1668
rect 28735 1857 28781 2057
rect 28865 1862 28911 2124
rect 30482 2096 30528 2496
rect 30798 2096 30844 2496
rect 32030 2233 32111 2571
rect 32030 2153 32809 2233
rect 34046 2172 34124 2188
rect 32030 2152 32680 2153
rect 33930 2146 34124 2172
rect 32871 2117 34124 2146
rect 35217 2118 35263 2518
rect 35533 2118 35579 2518
rect 28735 1405 28781 1668
rect 28865 1468 28911 1668
rect 29181 1862 29227 2062
rect 29181 1407 29227 1668
rect 29260 1407 29415 1422
rect 29181 1405 29415 1407
rect 28016 1368 29415 1405
rect 28016 1296 29216 1368
rect 29260 1356 29415 1368
rect 30482 1440 30528 1840
rect 30798 1440 30844 1840
rect 31114 1440 31160 1840
rect 31430 1440 31476 1840
rect 32871 1398 32909 2117
rect 32958 1850 33004 2050
rect 32958 1398 33004 1661
rect 33274 1850 33320 2117
rect 33274 1461 33320 1661
rect 33590 1850 33636 2050
rect 33720 1855 33766 2117
rect 36938 2075 36984 2475
rect 37254 2075 37300 2475
rect 33590 1398 33636 1661
rect 33720 1461 33766 1661
rect 34036 1855 34082 2055
rect 38454 2013 38590 3017
rect 39945 3003 44202 3060
rect 39278 2735 39324 2935
rect 39474 2735 39520 2935
rect 39670 2735 39716 2935
rect 39945 2682 40002 3003
rect 40160 2735 40206 2935
rect 40356 2735 40402 2935
rect 40552 2735 40598 2935
rect 40771 2820 40817 2920
rect 40869 2820 40915 2920
rect 40967 2820 41013 2920
rect 41065 2820 41111 2920
rect 41163 2820 41209 2920
rect 41261 2820 41307 2920
rect 41359 2820 41405 2920
rect 41457 2820 41503 2920
rect 41903 2735 41949 2935
rect 42099 2735 42145 2935
rect 42295 2735 42341 2935
rect 40774 2682 40943 2692
rect 39278 2455 39324 2555
rect 39474 2455 39520 2555
rect 39670 2455 39716 2555
rect 39804 2524 39864 2656
rect 39945 2625 40943 2682
rect 42645 2682 42702 2917
rect 42860 2735 42906 2935
rect 43056 2735 43102 2935
rect 43252 2735 43298 2935
rect 43471 2820 43517 2920
rect 43566 2882 43617 3003
rect 43569 2820 43615 2882
rect 43667 2820 43713 2920
rect 43760 2882 43811 3003
rect 43765 2820 43811 2882
rect 43863 2820 43909 2920
rect 43960 2863 44011 3003
rect 44152 2920 44202 3003
rect 43961 2820 44007 2863
rect 44059 2820 44105 2920
rect 44152 2888 44203 2920
rect 44157 2820 44203 2888
rect 44603 2735 44649 2935
rect 44799 2735 44845 2935
rect 44995 2735 45041 2935
rect 43474 2682 43643 2692
rect 40774 2618 40943 2625
rect 39804 2296 39862 2524
rect 40160 2455 40206 2555
rect 40356 2455 40402 2555
rect 40552 2455 40598 2555
rect 40771 2405 40817 2505
rect 40869 2405 40915 2505
rect 40967 2405 41013 2505
rect 41065 2405 41111 2505
rect 41163 2405 41209 2505
rect 41261 2405 41307 2505
rect 41359 2405 41405 2505
rect 41454 2405 41503 2505
rect 41903 2455 41949 2555
rect 42099 2455 42145 2555
rect 42295 2455 42341 2555
rect 42421 2545 42481 2632
rect 42420 2500 42481 2545
rect 40872 2308 40914 2405
rect 41068 2308 41110 2405
rect 41263 2308 41305 2405
rect 41454 2308 41500 2405
rect 39763 2236 39895 2296
rect 40740 2262 41500 2308
rect 40740 2096 40786 2262
rect 41567 2150 41699 2210
rect 39975 2095 40786 2096
rect 39967 2050 40786 2095
rect 34036 1400 34082 1661
rect 34115 1400 34270 1415
rect 34036 1398 34270 1400
rect 32871 1361 34270 1398
rect 27132 986 27450 1006
rect 27655 986 27727 1035
rect 27132 921 27727 986
rect 27132 906 27450 921
rect 27655 866 27727 921
rect 26241 288 26433 546
rect 22342 -524 23217 -353
rect 20701 -594 20745 -532
rect 18861 -638 20745 -594
rect 22342 -561 22513 -524
rect 20908 -867 20954 -767
rect 21104 -867 21150 -767
rect 21300 -867 21346 -767
rect 21554 -957 21600 -701
rect 21750 -957 21796 -701
rect 21946 -957 21992 -701
rect 22142 -957 22188 -701
rect 22342 -957 22388 -561
rect 26279 -620 26415 288
rect 28090 939 28136 1139
rect 28090 489 28136 689
rect 28248 370 28294 1139
rect 28406 939 28452 1296
rect 28406 489 28452 689
rect 28564 370 28610 1139
rect 28722 939 28768 1139
rect 28840 939 28886 1296
rect 29124 1226 29446 1296
rect 32871 1289 34071 1361
rect 34115 1349 34270 1361
rect 28722 489 28768 689
rect 28840 489 28886 689
rect 28998 370 29044 1139
rect 29371 721 29446 1226
rect 31987 979 32305 999
rect 32510 979 32582 1028
rect 31987 914 32582 979
rect 31987 899 32305 914
rect 32510 859 32582 914
rect 28062 324 29056 370
rect 30482 440 30528 840
rect 30798 440 30844 840
rect 31114 440 31160 840
rect 31430 440 31476 840
rect 32945 932 32991 1132
rect 32945 482 32991 682
rect 28247 244 28293 324
rect 28564 244 28610 324
rect 28995 244 29041 324
rect 27800 215 29435 244
rect 27803 -21 27849 215
rect 28119 -21 28165 215
rect 28247 211 28293 215
rect 28435 -21 28481 215
rect 28751 -21 28797 215
rect 29067 -21 29113 215
rect 29383 -21 29429 215
rect 33103 363 33149 1132
rect 33261 932 33307 1289
rect 33261 482 33307 682
rect 33419 363 33465 1132
rect 33577 932 33623 1132
rect 33695 932 33741 1289
rect 33979 1219 34301 1289
rect 33577 482 33623 682
rect 33695 482 33741 682
rect 33853 363 33899 1132
rect 34226 714 34301 1219
rect 35217 1462 35263 1862
rect 35533 1462 35579 1862
rect 35849 1462 35895 1862
rect 36165 1462 36211 1862
rect 36938 1419 36984 1819
rect 37254 1419 37300 1819
rect 37570 1419 37616 1819
rect 37886 1419 37932 1819
rect 38429 1755 38621 2013
rect 39967 1775 40013 2050
rect 40063 1847 40109 1947
rect 40161 1847 40207 1947
rect 40259 1847 40305 1947
rect 40357 1847 40403 1947
rect 40455 1847 40501 1947
rect 40553 1847 40599 1947
rect 40651 1847 40697 1947
rect 40749 1847 40795 1947
rect 40968 1797 41014 1897
rect 41164 1797 41210 1897
rect 41360 1797 41406 1897
rect 41610 1786 41670 2150
rect 41805 1797 41851 1897
rect 42001 1797 42047 1897
rect 42197 1797 42243 1897
rect 39967 1715 40121 1775
rect 42420 1752 42480 2500
rect 42536 2209 42596 2657
rect 42645 2625 43643 2682
rect 43474 2618 43643 2625
rect 51008 2563 51054 3034
rect 51244 2563 51290 3034
rect 51610 2563 51656 3034
rect 51846 2563 51892 3034
rect 52082 2563 52128 3034
rect 52318 2563 52364 3034
rect 52684 2563 52730 3034
rect 52920 2563 52966 3034
rect 53156 2563 53202 3034
rect 53392 2563 53438 3034
rect 53628 2563 53674 3034
rect 53864 2563 53910 3034
rect 54100 2563 54146 3034
rect 54336 2563 54382 3034
rect 42860 2455 42906 2555
rect 43056 2455 43102 2555
rect 43252 2455 43298 2555
rect 43471 2405 43517 2505
rect 43569 2424 43615 2505
rect 43565 2306 43626 2424
rect 43667 2405 43713 2505
rect 43765 2426 43811 2505
rect 43756 2306 43817 2426
rect 43863 2405 43909 2505
rect 43961 2424 44007 2505
rect 43952 2306 44013 2424
rect 44059 2405 44105 2505
rect 44157 2460 44203 2505
rect 44157 2306 44205 2460
rect 44603 2455 44649 2555
rect 44799 2455 44845 2555
rect 44995 2455 45041 2555
rect 51003 2489 51420 2563
rect 51481 2489 52491 2563
rect 52552 2489 54497 2563
rect 42674 2258 44205 2306
rect 42508 2149 42645 2209
rect 42674 1773 42715 2258
rect 44286 2238 44418 2298
rect 42763 1847 42809 1947
rect 42861 1847 42907 1947
rect 42959 1847 43005 1947
rect 43057 1847 43103 1947
rect 43155 1847 43201 1947
rect 43253 1847 43299 1947
rect 43351 1847 43397 1947
rect 43449 1847 43495 1947
rect 43668 1797 43714 1897
rect 43864 1797 43910 1897
rect 44060 1797 44106 1897
rect 40623 1727 40792 1734
rect 40623 1670 41621 1727
rect 42337 1692 42480 1752
rect 42673 1713 42810 1773
rect 44322 1771 44382 2238
rect 45095 2242 45155 2268
rect 45095 2178 45449 2242
rect 50510 2215 50749 2467
rect 45095 2131 45155 2178
rect 45385 2121 45449 2178
rect 45351 1935 45497 2121
rect 44505 1797 44551 1897
rect 44701 1797 44747 1897
rect 44897 1797 44943 1897
rect 45385 1849 45449 1935
rect 45671 1887 45717 1987
rect 45867 1887 45913 1987
rect 46063 1887 46109 1987
rect 46637 1917 46961 1997
rect 47896 1917 48216 1992
rect 50542 1917 50721 2215
rect 46637 1884 48216 1917
rect 45385 1775 45505 1849
rect 43323 1727 43492 1734
rect 42674 1712 42715 1713
rect 42420 1686 42480 1692
rect 40623 1660 40792 1670
rect 40063 1432 40109 1532
rect 40161 1432 40207 1532
rect 40259 1432 40305 1532
rect 40357 1432 40403 1532
rect 40455 1432 40501 1532
rect 40553 1432 40599 1532
rect 40651 1432 40697 1532
rect 40749 1432 40795 1532
rect 40968 1417 41014 1617
rect 41164 1417 41210 1617
rect 41360 1417 41406 1617
rect 41564 1435 41621 1670
rect 43323 1670 44321 1727
rect 43323 1660 43492 1670
rect 41805 1417 41851 1617
rect 42001 1417 42047 1617
rect 42197 1417 42243 1617
rect 42763 1432 42809 1532
rect 42861 1432 42907 1532
rect 42959 1432 43005 1532
rect 43057 1432 43103 1532
rect 43155 1432 43201 1532
rect 43253 1432 43299 1532
rect 43351 1432 43397 1532
rect 43449 1432 43495 1532
rect 43668 1417 43714 1617
rect 43864 1417 43910 1617
rect 44060 1417 44106 1617
rect 44264 1435 44321 1670
rect 44505 1417 44551 1617
rect 44701 1417 44747 1617
rect 44897 1417 44943 1617
rect 45385 1314 45459 1775
rect 46637 1738 49256 1884
rect 51300 1826 51346 2489
rect 51695 2349 51741 2489
rect 52677 2361 52723 2489
rect 51536 2303 51818 2349
rect 51536 1826 51582 2303
rect 51772 1826 51818 2303
rect 52008 2315 52762 2361
rect 52008 1826 52054 2315
rect 52244 1826 52290 2315
rect 52480 1826 52526 2315
rect 52716 1826 52762 2315
rect 45671 1507 45717 1707
rect 45867 1507 45913 1707
rect 46063 1507 46109 1707
rect 46637 1686 46961 1738
rect 47896 1705 49256 1738
rect 47896 1636 48216 1705
rect 46361 1314 46507 1357
rect 45385 1240 46507 1314
rect 30482 -216 30528 184
rect 30798 -216 30844 184
rect 32917 317 33911 363
rect 35217 463 35263 863
rect 35533 463 35579 863
rect 35849 463 35895 863
rect 36165 463 36211 863
rect 36938 506 36984 906
rect 37254 506 37300 906
rect 37570 506 37616 906
rect 37886 506 37932 906
rect 33102 237 33148 317
rect 33419 237 33465 317
rect 33850 237 33896 317
rect 32655 208 34290 237
rect 32658 -28 32704 208
rect 32974 -28 33020 208
rect 33102 204 33148 208
rect 33290 -28 33336 208
rect 33606 -28 33652 208
rect 33922 -28 33968 208
rect 34238 -28 34284 208
rect 38451 307 38643 565
rect 35217 -193 35263 207
rect 35533 -193 35579 207
rect 36938 -150 36984 250
rect 37254 -150 37300 250
rect 38481 -620 38617 307
rect 26279 -756 38617 -620
rect 46227 -632 46301 1240
rect 46361 1171 46507 1240
rect 47758 -632 47953 -572
rect 46227 -706 47953 -632
rect 47758 -752 47953 -706
rect 21554 -1003 22388 -957
rect 20908 -1247 20954 -1047
rect 21104 -1247 21150 -1047
rect 21300 -1247 21346 -1047
rect 21554 -1247 21600 -1003
rect 21750 -1247 21796 -1003
rect 21946 -1247 21992 -1003
rect 22142 -1247 22188 -1003
rect 49077 -3371 49256 1705
rect 50805 -348 50851 123
rect 51041 -348 51087 123
rect 51407 -348 51453 123
rect 51643 -348 51689 123
rect 51879 -348 51925 123
rect 52115 -348 52161 123
rect 52481 -348 52527 123
rect 52717 -348 52763 123
rect 52953 -348 52999 123
rect 53189 -348 53235 123
rect 53425 -348 53471 123
rect 53661 -348 53707 123
rect 53897 -348 53943 123
rect 54133 -348 54179 123
rect 50800 -422 51217 -348
rect 51278 -422 52288 -348
rect 52349 -422 54294 -348
rect 51097 -1085 51143 -422
rect 51492 -562 51538 -422
rect 52474 -550 52520 -422
rect 51333 -608 51615 -562
rect 51333 -1085 51379 -608
rect 51569 -1085 51615 -608
rect 51805 -596 52559 -550
rect 51805 -1085 51851 -596
rect 52041 -1085 52087 -596
rect 52277 -1085 52323 -596
rect 52513 -1085 52559 -596
rect 48966 -3697 49277 -3371
rect 50805 -3395 50851 -2924
rect 51041 -3395 51087 -2924
rect 51407 -3395 51453 -2924
rect 51643 -3395 51689 -2924
rect 51879 -3395 51925 -2924
rect 52115 -3395 52161 -2924
rect 52481 -3395 52527 -2924
rect 52717 -3395 52763 -2924
rect 52953 -3395 52999 -2924
rect 53189 -3395 53235 -2924
rect 53425 -3395 53471 -2924
rect 53661 -3395 53707 -2924
rect 53897 -3395 53943 -2924
rect 54133 -3395 54179 -2924
rect 54381 -3395 54427 -2924
rect 54617 -3395 54663 -2924
rect 54853 -3395 54899 -2924
rect 55089 -3395 55135 -2924
rect 55325 -3395 55371 -2924
rect 55561 -3395 55607 -2924
rect 55797 -3395 55843 -2924
rect 56033 -3395 56079 -2924
rect 56269 -3395 56315 -2924
rect 56505 -3395 56551 -2924
rect 56741 -3395 56787 -2924
rect 56977 -3395 57023 -2924
rect 57213 -3395 57259 -2924
rect 57449 -3395 57495 -2924
rect 57685 -3395 57731 -2924
rect 57921 -3395 57967 -2924
rect 58157 -3395 58203 -2924
rect 50800 -3469 51217 -3395
rect 51278 -3469 52288 -3395
rect 52349 -3469 54294 -3395
rect 54355 -3469 58232 -3395
rect 51097 -4132 51143 -3469
rect 51492 -3609 51538 -3469
rect 52474 -3597 52520 -3469
rect 54401 -3585 54447 -3469
rect 51333 -3655 51615 -3609
rect 51333 -4132 51379 -3655
rect 51569 -4132 51615 -3655
rect 51805 -3643 52559 -3597
rect 51805 -4132 51851 -3643
rect 52041 -4132 52087 -3643
rect 52277 -4132 52323 -3643
rect 52513 -4132 52559 -3643
rect 52749 -3631 54447 -3585
rect 52749 -4132 52795 -3631
rect 52985 -4132 53031 -3631
rect 53221 -4132 53267 -3631
rect 53457 -4132 53503 -3631
rect 53693 -4132 53739 -3631
rect 53929 -4132 53975 -3631
rect 54165 -4132 54211 -3631
rect 54401 -4132 54447 -3631
rect 62485 -3038 62531 -2838
rect 62681 -3038 62727 -2838
rect 62877 -3038 62923 -2838
rect 63335 -3038 63381 -2838
rect 63531 -3038 63577 -2838
rect 63727 -3038 63773 -2838
rect 63883 -3038 63929 -2838
rect 63981 -3082 64027 -2838
rect 64079 -3038 64125 -2838
rect 64177 -3082 64223 -2838
rect 64275 -3038 64321 -2838
rect 64373 -3082 64419 -2838
rect 64471 -3038 64517 -2838
rect 64569 -3082 64615 -2838
rect 64667 -3038 64713 -2838
rect 63981 -3128 64815 -3082
rect 62485 -3318 62531 -3218
rect 62681 -3318 62727 -3218
rect 62877 -3318 62923 -3218
rect 63040 -3254 63172 -3210
rect 63128 -3354 63172 -3254
rect 63335 -3318 63381 -3218
rect 63531 -3318 63577 -3218
rect 63727 -3318 63773 -3218
rect 63883 -3354 63929 -3184
rect 61873 -3460 62067 -3407
rect 63128 -3398 63930 -3354
rect 63981 -3384 64027 -3128
rect 64079 -3384 64125 -3184
rect 64177 -3384 64223 -3128
rect 64275 -3384 64321 -3184
rect 64373 -3384 64419 -3128
rect 64471 -3384 64517 -3184
rect 64569 -3384 64615 -3128
rect 64667 -3384 64713 -3184
rect 64769 -3381 64815 -3128
rect 65187 -3381 65330 -3337
rect 63128 -3460 63172 -3398
rect 61873 -3504 63172 -3460
rect 64769 -3427 65330 -3381
rect 61873 -3516 62067 -3504
rect 63335 -3733 63381 -3633
rect 63531 -3733 63577 -3633
rect 63727 -3733 63773 -3633
rect 63981 -3823 64027 -3567
rect 64177 -3823 64223 -3567
rect 64373 -3823 64419 -3567
rect 64569 -3823 64615 -3567
rect 64769 -3823 64815 -3427
rect 65187 -3468 65330 -3427
rect 87785 -3581 88210 -3189
rect 63981 -3869 64815 -3823
rect 63335 -4113 63381 -3913
rect 63531 -4113 63577 -3913
rect 63727 -4113 63773 -3913
rect 63981 -4113 64027 -3869
rect 64177 -4113 64223 -3869
rect 64373 -4113 64419 -3869
rect 64569 -4113 64615 -3869
rect -12874 -15238 -7870 -14969
rect -12865 -15240 -11924 -15238
rect -14957 -15728 -14911 -15328
rect -14839 -15728 -14793 -15328
rect -14721 -15728 -14675 -15328
rect -14603 -15728 -14557 -15328
rect -14485 -15728 -14439 -15328
rect -14367 -15728 -14321 -15328
rect -14249 -15728 -14203 -15328
rect -14131 -15728 -14085 -15328
rect -14013 -15728 -13967 -15328
rect -13895 -15728 -13849 -15328
rect -13777 -15728 -13731 -15328
rect -13659 -15728 -13613 -15328
rect -13541 -15728 -13495 -15328
rect -13423 -15728 -13377 -15328
rect -13305 -15728 -13259 -15328
rect -13187 -15728 -13141 -15328
rect -13069 -15728 -13023 -15328
rect -12951 -15728 -12905 -15328
rect -12833 -15728 -12787 -15328
rect -12715 -15728 -12669 -15328
rect -12597 -15728 -12551 -15328
rect -12479 -15728 -12433 -15328
rect -12361 -15728 -12315 -15328
rect -12243 -15728 -12197 -15328
rect -12125 -15728 -12079 -15328
rect -12007 -15728 -11961 -15328
rect -11889 -15728 -11843 -15328
rect -11771 -15728 -11725 -15328
rect -11653 -15728 -11607 -15328
rect -11535 -15728 -11489 -15328
rect -11417 -15728 -11371 -15328
rect -11181 -15728 -11135 -15328
rect -10945 -15728 -10899 -15328
rect -10709 -15728 -10663 -15328
rect -10473 -15728 -10427 -15328
rect -10237 -15728 -10191 -15328
rect -10001 -15728 -9955 -15328
rect -9765 -15728 -9719 -15328
rect -9529 -15728 -9483 -15328
rect -9411 -15817 -9365 -15328
rect -9293 -15728 -9247 -15328
rect -9175 -15817 -9129 -15328
rect -9057 -15728 -9011 -15328
rect -8939 -15817 -8893 -15328
rect -8821 -15728 -8775 -15328
rect -8703 -15817 -8657 -15328
rect -8585 -15728 -8539 -15328
rect -9411 -15863 -8657 -15817
rect -8467 -15805 -8421 -15328
rect -8349 -15728 -8303 -15328
rect -8231 -15805 -8185 -15328
rect -8113 -15728 -8067 -15328
rect -8467 -15851 -8185 -15805
rect -9372 -15991 -9326 -15863
rect -8390 -15991 -8344 -15851
rect -7995 -15991 -7949 -15328
rect -7877 -15728 -7831 -15328
rect 12075 -15445 87696 -15161
rect -11146 -16065 -9201 -15991
rect -9140 -16065 -8130 -15991
rect -8069 -16065 -7652 -15991
rect -11031 -16536 -10985 -16065
rect -10795 -16536 -10749 -16065
rect -10559 -16536 -10513 -16065
rect -10323 -16536 -10277 -16065
rect -10087 -16536 -10041 -16065
rect -9851 -16536 -9805 -16065
rect -9615 -16536 -9569 -16065
rect -9379 -16536 -9333 -16065
rect -9013 -16536 -8967 -16065
rect -8777 -16536 -8731 -16065
rect -8541 -16536 -8495 -16065
rect -8305 -16536 -8259 -16065
rect -7939 -16536 -7893 -16065
rect -7703 -16536 -7657 -16065
rect -16604 -18135 7804 -17945
rect -24032 -20611 -23931 -20556
rect -24184 -20799 -23931 -20611
rect -24184 -20842 -23944 -20799
rect -25664 -23404 -25039 -22779
rect -24184 -29767 -24048 -20842
rect -22646 -19384 -22600 -19184
rect -22450 -19384 -22404 -19184
rect -22254 -19384 -22208 -19184
rect -21516 -19384 -21470 -19184
rect -16604 -19224 -16414 -18135
rect -15047 -18597 -15001 -18397
rect -14851 -18597 -14805 -18397
rect -14655 -18597 -14609 -18397
rect -14425 -18650 -14368 -18415
rect -14210 -18597 -14164 -18397
rect -14014 -18597 -13968 -18397
rect -13818 -18597 -13772 -18397
rect -13599 -18512 -13553 -18412
rect -13501 -18512 -13455 -18412
rect -13403 -18512 -13357 -18412
rect -13305 -18512 -13259 -18412
rect -13207 -18512 -13161 -18412
rect -13109 -18512 -13063 -18412
rect -13011 -18512 -12965 -18412
rect -12913 -18512 -12867 -18412
rect -12347 -18597 -12301 -18397
rect -12151 -18597 -12105 -18397
rect -11955 -18597 -11909 -18397
rect -13596 -18650 -13427 -18640
rect -14425 -18707 -13427 -18650
rect -11725 -18650 -11668 -18415
rect -11510 -18597 -11464 -18397
rect -11314 -18597 -11268 -18397
rect -11118 -18597 -11072 -18397
rect -10899 -18512 -10853 -18412
rect -10801 -18512 -10755 -18412
rect -10703 -18512 -10657 -18412
rect -10605 -18512 -10559 -18412
rect -10507 -18512 -10461 -18412
rect -10409 -18512 -10363 -18412
rect -10311 -18512 -10265 -18412
rect -10213 -18512 -10167 -18412
rect -10896 -18650 -10727 -18640
rect -12584 -18672 -12524 -18666
rect -12819 -18693 -12778 -18692
rect -13596 -18714 -13427 -18707
rect -15145 -18877 -15099 -18777
rect -15047 -18877 -15001 -18777
rect -14949 -18877 -14903 -18777
rect -14851 -18877 -14805 -18777
rect -14753 -18877 -14707 -18777
rect -14655 -18877 -14609 -18777
rect -14911 -19100 -14774 -19040
rect -15259 -19158 -15199 -19111
rect -15521 -19222 -15199 -19158
rect -20647 -19606 -20601 -19306
rect -22744 -20091 -22698 -19791
rect -22646 -20091 -22600 -19791
rect -22548 -20091 -22502 -19791
rect -22434 -20092 -22388 -19792
rect -22336 -20092 -22290 -19792
rect -22238 -20092 -22192 -19792
rect -22125 -20092 -22079 -19792
rect -22027 -20092 -21981 -19792
rect -21929 -20092 -21883 -19792
rect -21614 -20092 -21568 -19892
rect -21516 -20008 -21470 -19892
rect -21516 -20043 -21157 -20008
rect -21516 -20092 -21470 -20043
rect -22589 -21515 -22543 -21215
rect -22687 -22051 -22641 -21752
rect -22688 -22088 -22641 -22051
rect -22589 -22052 -22543 -21752
rect -22491 -22088 -22445 -21752
rect -22393 -22052 -22347 -21215
rect -21980 -21370 -21934 -21214
rect -21784 -21368 -21738 -21214
rect -21882 -21370 -21640 -21368
rect -21588 -21370 -21542 -21214
rect -21980 -21416 -21343 -21370
rect -21980 -21545 -21934 -21445
rect -21882 -21545 -21836 -21416
rect -21784 -21545 -21738 -21445
rect -21686 -21545 -21640 -21416
rect -21192 -21577 -21157 -20043
rect -20745 -20142 -20699 -19843
rect -20746 -20179 -20699 -20142
rect -20647 -20143 -20601 -19843
rect -20549 -20179 -20503 -19843
rect -20451 -20143 -20405 -19306
rect -20038 -19461 -19992 -19305
rect -19842 -19459 -19796 -19305
rect -19940 -19461 -19698 -19459
rect -19646 -19461 -19600 -19305
rect -16985 -19337 -16308 -19224
rect -20038 -19507 -19401 -19461
rect -20038 -19636 -19992 -19536
rect -19940 -19636 -19894 -19507
rect -19842 -19636 -19796 -19536
rect -19744 -19636 -19698 -19507
rect -19318 -19532 -19172 -19474
rect -19318 -19558 -19237 -19532
rect -19630 -19593 -19237 -19558
rect -20353 -20179 -20307 -19843
rect -20746 -20226 -20307 -20179
rect -19630 -20663 -19595 -19593
rect -19110 -19695 -18671 -19648
rect -19110 -19732 -19063 -19695
rect -19109 -20031 -19063 -19732
rect -19011 -20031 -18965 -19731
rect -18913 -20031 -18867 -19695
rect -19364 -20127 -19167 -20073
rect -21126 -20698 -19595 -20663
rect -21126 -21446 -21091 -20698
rect -20816 -21320 -20770 -21120
rect -20620 -21320 -20574 -21120
rect -20424 -21320 -20378 -21120
rect -19686 -21320 -19640 -21120
rect -21126 -21492 -21042 -21446
rect -22295 -22088 -22249 -21752
rect -21411 -21811 -21353 -21674
rect -21197 -21714 -21139 -21577
rect -21100 -21583 -21042 -21492
rect -19221 -21531 -19167 -20127
rect -19011 -20568 -18965 -20268
rect -18815 -20568 -18769 -19731
rect -18717 -20031 -18671 -19695
rect -17564 -19745 -17518 -19445
rect -17466 -19745 -17420 -19445
rect -17368 -19745 -17322 -19445
rect -17126 -19745 -17080 -19445
rect -17028 -19745 -16982 -19445
rect -17663 -19843 -16643 -19778
rect -16708 -19926 -16643 -19843
rect -16714 -19998 -16609 -19926
rect -18402 -20338 -18356 -20238
rect -18304 -20367 -18258 -20238
rect -18206 -20338 -18160 -20238
rect -18108 -20367 -18062 -20238
rect -18402 -20413 -17765 -20367
rect -18402 -20569 -18356 -20413
rect -18304 -20415 -18062 -20413
rect -18206 -20569 -18160 -20415
rect -18010 -20569 -17964 -20413
rect -17564 -20657 -17518 -20057
rect -17353 -20657 -17307 -20057
rect -17255 -20657 -17209 -20057
rect -17157 -20657 -17111 -20057
rect -16945 -20657 -16899 -20057
rect -19271 -21681 -19141 -21531
rect -18985 -21553 -18939 -21297
rect -18789 -21551 -18743 -21297
rect -18887 -21553 -18645 -21551
rect -18593 -21553 -18547 -21297
rect -18012 -21468 -17966 -21168
rect -18985 -21599 -18348 -21553
rect -18206 -21572 -18047 -21514
rect -20914 -22027 -20868 -21727
rect -20816 -22027 -20770 -21727
rect -20718 -22027 -20672 -21727
rect -20604 -22028 -20558 -21728
rect -20506 -22028 -20460 -21728
rect -20408 -22028 -20362 -21728
rect -20295 -22028 -20249 -21728
rect -20197 -22028 -20151 -21728
rect -20099 -22028 -20053 -21728
rect -18985 -21827 -18939 -21627
rect -18887 -21827 -18841 -21599
rect -18789 -21827 -18743 -21627
rect -18691 -21827 -18645 -21599
rect -18180 -21627 -18126 -21572
rect -18454 -21681 -18126 -21627
rect -19784 -22028 -19738 -21828
rect -19686 -22028 -19640 -21828
rect -18454 -21971 -18400 -21681
rect -19497 -22025 -18400 -21971
rect -18110 -22004 -18064 -21705
rect -22688 -22135 -22249 -22088
rect -19485 -22739 -19245 -22025
rect -18111 -22041 -18064 -22004
rect -18012 -22005 -17966 -21705
rect -17914 -22041 -17868 -21705
rect -17816 -22005 -17770 -21168
rect -17403 -21323 -17357 -21167
rect -17207 -21321 -17161 -21167
rect -17305 -21323 -17063 -21321
rect -17011 -21323 -16965 -21167
rect -17403 -21369 -16766 -21323
rect -17403 -21498 -17357 -21398
rect -17305 -21498 -17259 -21369
rect -17207 -21498 -17161 -21398
rect -17109 -21498 -17063 -21369
rect -16421 -21533 -16308 -19337
rect -15521 -21138 -15457 -19222
rect -15259 -19248 -15199 -19222
rect -14896 -19318 -14801 -19100
rect -14486 -19218 -14426 -18751
rect -12914 -18753 -12777 -18693
rect -12584 -18732 -12441 -18672
rect -11725 -18707 -10727 -18650
rect -10896 -18714 -10727 -18707
rect -14308 -18877 -14262 -18777
rect -14210 -18877 -14164 -18777
rect -14112 -18877 -14066 -18777
rect -14014 -18877 -13968 -18777
rect -13916 -18877 -13870 -18777
rect -13818 -18877 -13772 -18777
rect -13599 -18927 -13553 -18827
rect -13501 -18927 -13455 -18827
rect -13403 -18927 -13357 -18827
rect -13305 -18927 -13259 -18827
rect -13207 -18927 -13161 -18827
rect -13109 -18927 -13063 -18827
rect -13011 -18927 -12965 -18827
rect -12913 -18927 -12867 -18827
rect -14522 -19278 -14390 -19218
rect -12819 -19238 -12778 -18753
rect -12749 -19189 -12612 -19129
rect -14309 -19286 -12778 -19238
rect -14920 -19378 -14788 -19318
rect -15145 -19535 -15099 -19435
rect -15047 -19535 -15001 -19435
rect -14949 -19535 -14903 -19435
rect -14851 -19535 -14805 -19435
rect -14753 -19535 -14707 -19435
rect -14655 -19535 -14609 -19435
rect -14309 -19440 -14261 -19286
rect -14307 -19485 -14261 -19440
rect -14209 -19485 -14163 -19385
rect -14117 -19404 -14056 -19286
rect -14111 -19485 -14065 -19404
rect -14013 -19485 -13967 -19385
rect -13921 -19406 -13860 -19286
rect -13915 -19485 -13869 -19406
rect -13817 -19485 -13771 -19385
rect -13730 -19404 -13669 -19286
rect -13719 -19485 -13673 -19404
rect -13621 -19485 -13575 -19385
rect -13402 -19535 -13356 -19435
rect -13304 -19535 -13258 -19435
rect -13206 -19535 -13160 -19435
rect -13108 -19535 -13062 -19435
rect -13010 -19535 -12964 -19435
rect -12912 -19535 -12866 -19435
rect -13747 -19605 -13578 -19598
rect -13747 -19662 -12749 -19605
rect -12700 -19637 -12640 -19189
rect -12584 -19480 -12524 -18732
rect -10225 -18755 -10071 -18695
rect -12445 -18877 -12399 -18777
rect -12347 -18877 -12301 -18777
rect -12249 -18877 -12203 -18777
rect -12151 -18877 -12105 -18777
rect -12053 -18877 -12007 -18777
rect -11955 -18877 -11909 -18777
rect -12314 -19106 -12177 -19046
rect -12303 -19314 -12208 -19106
rect -11774 -19130 -11714 -18766
rect -11608 -18877 -11562 -18777
rect -11510 -18877 -11464 -18777
rect -11412 -18877 -11366 -18777
rect -11314 -18877 -11268 -18777
rect -11216 -18877 -11170 -18777
rect -11118 -18877 -11072 -18777
rect -10899 -18927 -10853 -18827
rect -10801 -18927 -10755 -18827
rect -10703 -18927 -10657 -18827
rect -10605 -18927 -10559 -18827
rect -10507 -18927 -10461 -18827
rect -10409 -18927 -10363 -18827
rect -10311 -18927 -10265 -18827
rect -10213 -18927 -10167 -18827
rect -10117 -19030 -10071 -18755
rect -10890 -19075 -10071 -19030
rect -10890 -19076 -10079 -19075
rect -11803 -19190 -11671 -19130
rect -10890 -19242 -10844 -19076
rect -9676 -19106 -9544 -19046
rect -9659 -19171 -9564 -19106
rect -9124 -19171 -9029 -18135
rect -8881 -19007 -8835 -18407
rect -8669 -19007 -8623 -18407
rect -8571 -19007 -8525 -18407
rect -8473 -19007 -8427 -18407
rect -8262 -19007 -8216 -18407
rect -7451 -18803 -7405 -18603
rect -7353 -18803 -7307 -18603
rect -7255 -18803 -7209 -18603
rect -7135 -18803 -7089 -18603
rect -7037 -18803 -6991 -18603
rect -6939 -18803 -6893 -18603
rect -6577 -18803 -6531 -18603
rect -6381 -18803 -6335 -18603
rect -6071 -18803 -6025 -18603
rect -5762 -18803 -5716 -18603
rect -4951 -18803 -4905 -18603
rect -4853 -18803 -4807 -18603
rect -4755 -18803 -4709 -18603
rect -4635 -18803 -4589 -18603
rect -4537 -18803 -4491 -18603
rect -4439 -18803 -4393 -18603
rect -4077 -18803 -4031 -18603
rect -3881 -18803 -3835 -18603
rect -3571 -18803 -3525 -18603
rect -3262 -18803 -3216 -18603
rect -2451 -18803 -2405 -18603
rect -2353 -18803 -2307 -18603
rect -2255 -18803 -2209 -18603
rect -2135 -18803 -2089 -18603
rect -2037 -18803 -1991 -18603
rect -1939 -18803 -1893 -18603
rect -1577 -18803 -1531 -18603
rect -1381 -18803 -1335 -18603
rect -1071 -18803 -1025 -18603
rect -762 -18803 -716 -18603
rect 49 -18803 95 -18603
rect 147 -18803 193 -18603
rect 245 -18803 291 -18603
rect 365 -18803 411 -18603
rect 463 -18803 509 -18603
rect 561 -18803 607 -18603
rect 923 -18803 969 -18603
rect 1119 -18803 1165 -18603
rect 1429 -18803 1475 -18603
rect 1738 -18803 1784 -18603
rect 2549 -18803 2595 -18603
rect 2647 -18803 2693 -18603
rect 2745 -18803 2791 -18603
rect 2865 -18803 2911 -18603
rect 2963 -18803 3009 -18603
rect 3061 -18803 3107 -18603
rect 3423 -18803 3469 -18603
rect 3619 -18803 3665 -18603
rect 3929 -18803 3975 -18603
rect 4238 -18803 4284 -18603
rect 5549 -18803 5595 -18603
rect 5647 -18803 5693 -18603
rect 5745 -18803 5791 -18603
rect 5865 -18803 5911 -18603
rect 5963 -18803 6009 -18603
rect 6061 -18803 6107 -18603
rect 6423 -18803 6469 -18603
rect 6619 -18803 6665 -18603
rect 6929 -18803 6975 -18603
rect 7238 -18803 7284 -18603
rect -6288 -18931 -6149 -18913
rect -5673 -18931 -5534 -18919
rect -3788 -18931 -3649 -18913
rect -3173 -18931 -3034 -18919
rect -1288 -18931 -1149 -18913
rect -673 -18931 -534 -18919
rect 1212 -18931 1351 -18913
rect 1827 -18931 1966 -18919
rect 3712 -18931 3851 -18913
rect 4327 -18931 4466 -18919
rect 6712 -18931 6851 -18913
rect 7327 -18931 7466 -18919
rect 8028 -18931 8228 -18579
rect -7446 -18970 -7307 -18957
rect -6288 -18959 -5383 -18931
rect -6288 -18967 -6149 -18959
rect -7446 -18998 -7092 -18970
rect -5673 -18973 -5534 -18959
rect -7446 -19011 -7307 -18998
rect -11604 -19288 -10844 -19242
rect -9999 -19276 -9867 -19216
rect -9659 -19266 -9029 -19171
rect -12321 -19374 -12184 -19314
rect -11604 -19385 -11558 -19288
rect -11409 -19385 -11367 -19288
rect -11214 -19385 -11172 -19288
rect -11018 -19385 -10976 -19288
rect -12585 -19525 -12524 -19480
rect -12585 -19612 -12525 -19525
rect -12445 -19535 -12399 -19435
rect -12347 -19535 -12301 -19435
rect -12249 -19535 -12203 -19435
rect -12151 -19535 -12105 -19435
rect -12053 -19535 -12007 -19435
rect -11955 -19535 -11909 -19435
rect -11607 -19485 -11558 -19385
rect -11509 -19485 -11463 -19385
rect -11411 -19485 -11365 -19385
rect -11313 -19485 -11267 -19385
rect -11215 -19485 -11169 -19385
rect -11117 -19485 -11071 -19385
rect -11019 -19485 -10973 -19385
rect -10921 -19485 -10875 -19385
rect -10702 -19535 -10656 -19435
rect -10604 -19535 -10558 -19435
rect -10506 -19535 -10460 -19435
rect -10408 -19535 -10362 -19435
rect -10310 -19535 -10264 -19435
rect -10212 -19535 -10166 -19435
rect -9966 -19504 -9908 -19276
rect -9659 -19315 -9564 -19266
rect -9694 -19375 -9557 -19315
rect -11047 -19605 -10878 -19598
rect -13747 -19672 -13578 -19662
rect -15145 -19915 -15099 -19715
rect -14949 -19915 -14903 -19715
rect -14753 -19915 -14707 -19715
rect -14307 -19868 -14261 -19800
rect -14307 -19900 -14256 -19868
rect -14209 -19900 -14163 -19800
rect -14111 -19843 -14065 -19800
rect -14306 -19983 -14256 -19900
rect -14115 -19983 -14064 -19843
rect -14013 -19900 -13967 -19800
rect -13915 -19862 -13869 -19800
rect -13915 -19983 -13864 -19862
rect -13817 -19900 -13771 -19800
rect -13719 -19862 -13673 -19800
rect -13721 -19983 -13670 -19862
rect -13621 -19900 -13575 -19800
rect -13402 -19915 -13356 -19715
rect -13206 -19915 -13160 -19715
rect -13010 -19915 -12964 -19715
rect -12806 -19897 -12749 -19662
rect -11047 -19662 -10049 -19605
rect -9968 -19636 -9908 -19504
rect -9820 -19535 -9774 -19435
rect -9722 -19535 -9676 -19435
rect -9624 -19535 -9578 -19435
rect -9526 -19535 -9480 -19435
rect -9428 -19535 -9382 -19435
rect -9330 -19535 -9284 -19435
rect -11047 -19672 -10878 -19662
rect -12445 -19915 -12399 -19715
rect -12249 -19915 -12203 -19715
rect -12053 -19915 -12007 -19715
rect -11607 -19900 -11561 -19800
rect -11509 -19900 -11463 -19800
rect -11411 -19900 -11365 -19800
rect -11313 -19900 -11267 -19800
rect -11215 -19900 -11169 -19800
rect -11117 -19900 -11071 -19800
rect -11019 -19900 -10973 -19800
rect -10921 -19900 -10875 -19800
rect -10702 -19915 -10656 -19715
rect -10506 -19915 -10460 -19715
rect -10310 -19915 -10264 -19715
rect -10106 -19983 -10049 -19662
rect -9820 -19915 -9774 -19715
rect -9624 -19915 -9578 -19715
rect -9428 -19915 -9382 -19715
rect -14306 -20040 -10049 -19983
rect -9124 -20200 -9029 -19266
rect -8798 -19619 -8752 -19319
rect -8700 -19619 -8654 -19319
rect -8458 -19619 -8412 -19319
rect -8360 -19619 -8314 -19319
rect -8262 -19619 -8216 -19319
rect -11996 -20313 -9028 -20200
rect -14121 -20671 -13682 -20624
rect -14121 -20708 -14074 -20671
rect -14120 -21007 -14074 -20708
rect -14022 -21007 -13976 -20707
rect -13924 -21007 -13878 -20671
rect -14659 -21138 -14473 -21096
rect -15521 -21202 -14473 -21138
rect -14659 -21250 -14473 -21202
rect -17016 -21646 -16308 -21533
rect -17718 -22041 -17672 -21705
rect -18111 -22088 -17672 -22041
rect -17099 -22397 -16831 -22132
rect -17050 -22952 -16862 -22397
rect -17094 -23217 -16826 -22952
rect -22524 -25009 -22478 -24409
rect -22312 -25009 -22266 -24409
rect -22214 -25009 -22168 -24409
rect -22116 -25009 -22070 -24409
rect -22003 -25009 -21957 -24409
rect -21905 -25009 -21859 -24409
rect -21807 -25009 -21761 -24409
rect -21318 -24738 -21272 -24338
rect -21107 -24738 -21061 -24338
rect -21009 -24738 -20963 -24338
rect -20911 -24738 -20865 -24338
rect -20413 -24739 -20367 -24339
rect -20202 -24739 -20156 -24339
rect -20104 -24739 -20058 -24339
rect -20006 -24739 -19960 -24339
rect -21786 -25335 -21649 -25277
rect -22524 -25573 -22478 -25373
rect -22426 -25573 -22380 -25373
rect -22328 -25573 -22282 -25373
rect -22230 -25573 -22184 -25373
rect -22658 -25819 -21854 -25669
rect -22646 -26231 -22559 -25819
rect -22466 -26231 -22379 -25819
rect -22293 -26231 -22206 -25819
rect -22109 -26231 -22022 -25819
rect -21984 -26231 -21897 -25819
rect -22871 -26346 -21888 -26231
rect -21774 -26333 -21684 -25335
rect -20899 -24986 -20762 -24928
rect -21318 -25230 -21272 -25030
rect -21220 -25230 -21174 -25030
rect -21122 -25230 -21076 -25030
rect -21774 -26423 -21457 -26333
rect -22861 -26719 -22815 -26519
rect -22763 -26719 -22717 -26519
rect -22448 -26819 -22402 -26519
rect -22350 -26819 -22304 -26519
rect -22252 -26819 -22206 -26519
rect -22139 -26819 -22093 -26519
rect -22041 -26819 -21995 -26519
rect -21943 -26819 -21897 -26519
rect -21829 -26820 -21783 -26520
rect -21731 -26820 -21685 -26520
rect -21633 -26820 -21587 -26520
rect -21547 -27011 -21457 -26423
rect -20808 -26956 -20773 -24986
rect -19968 -24987 -19831 -24929
rect -20413 -25231 -20367 -25031
rect -20315 -25231 -20269 -25031
rect -20217 -25231 -20171 -25031
rect -20816 -27093 -20758 -26956
rect -22861 -27427 -22815 -27227
rect -22123 -27427 -22077 -27227
rect -21927 -27427 -21881 -27227
rect -21731 -27427 -21685 -27227
rect -22860 -27698 -22817 -27427
rect -19883 -27042 -19848 -24987
rect -19707 -25285 -19590 -25162
rect -19806 -26690 -19748 -26553
rect -19891 -27179 -19833 -27042
rect -22910 -27814 -22752 -27698
rect -19805 -27726 -19766 -26690
rect -19704 -27549 -19612 -25285
rect -16421 -24224 -16308 -21646
rect -14022 -21544 -13976 -21244
rect -13826 -21544 -13780 -20707
rect -13728 -21007 -13682 -20671
rect -12575 -20721 -12529 -20421
rect -12477 -20721 -12431 -20421
rect -12379 -20721 -12333 -20421
rect -12137 -20721 -12091 -20421
rect -12039 -20721 -11993 -20421
rect -12674 -20819 -11654 -20754
rect -11719 -20902 -11654 -20819
rect -11725 -20974 -11620 -20902
rect -13413 -21314 -13367 -21214
rect -13315 -21343 -13269 -21214
rect -13217 -21314 -13171 -21214
rect -13119 -21343 -13073 -21214
rect -13413 -21389 -12776 -21343
rect -13413 -21545 -13367 -21389
rect -13315 -21391 -13073 -21389
rect -13217 -21545 -13171 -21391
rect -13021 -21545 -12975 -21389
rect -12575 -21633 -12529 -21033
rect -12364 -21633 -12318 -21033
rect -12266 -21633 -12220 -21033
rect -12168 -21633 -12122 -21033
rect -11956 -21633 -11910 -21033
rect -16985 -24337 -16308 -24224
rect -19110 -24695 -18671 -24648
rect -19110 -24732 -19063 -24695
rect -19109 -25031 -19063 -24732
rect -19011 -25031 -18965 -24731
rect -18913 -25031 -18867 -24695
rect -19364 -25127 -19167 -25073
rect -19221 -26531 -19167 -25127
rect -19011 -25568 -18965 -25268
rect -18815 -25568 -18769 -24731
rect -18717 -25031 -18671 -24695
rect -17564 -24745 -17518 -24445
rect -17466 -24745 -17420 -24445
rect -17368 -24745 -17322 -24445
rect -17126 -24745 -17080 -24445
rect -17028 -24745 -16982 -24445
rect -17663 -24843 -16643 -24778
rect -16708 -24926 -16643 -24843
rect -16714 -24998 -16609 -24926
rect -18402 -25338 -18356 -25238
rect -18304 -25367 -18258 -25238
rect -18206 -25338 -18160 -25238
rect -18108 -25367 -18062 -25238
rect -18402 -25413 -17765 -25367
rect -18402 -25569 -18356 -25413
rect -18304 -25415 -18062 -25413
rect -18206 -25569 -18160 -25415
rect -18010 -25569 -17964 -25413
rect -17564 -25657 -17518 -25057
rect -17353 -25657 -17307 -25057
rect -17255 -25657 -17209 -25057
rect -17157 -25657 -17111 -25057
rect -16945 -25657 -16899 -25057
rect -19271 -26681 -19141 -26531
rect -18985 -26553 -18939 -26297
rect -18789 -26551 -18743 -26297
rect -18887 -26553 -18645 -26551
rect -18593 -26553 -18547 -26297
rect -18012 -26468 -17966 -26168
rect -18985 -26599 -18348 -26553
rect -18206 -26572 -18047 -26514
rect -18985 -26827 -18939 -26627
rect -18887 -26827 -18841 -26599
rect -18789 -26827 -18743 -26627
rect -18691 -26827 -18645 -26599
rect -18180 -26627 -18126 -26572
rect -18454 -26681 -18126 -26627
rect -18454 -26971 -18400 -26681
rect -19497 -27025 -18400 -26971
rect -18110 -27004 -18064 -26705
rect -19497 -27295 -19443 -27025
rect -18111 -27041 -18064 -27004
rect -18012 -27005 -17966 -26705
rect -17914 -27041 -17868 -26705
rect -17816 -27005 -17770 -26168
rect -17403 -26323 -17357 -26167
rect -17207 -26321 -17161 -26167
rect -17305 -26323 -17063 -26321
rect -17011 -26323 -16965 -26167
rect -17403 -26369 -16766 -26323
rect -17403 -26498 -17357 -26398
rect -17305 -26498 -17259 -26369
rect -17207 -26498 -17161 -26398
rect -17109 -26498 -17063 -26369
rect -16421 -26533 -16308 -24337
rect -16155 -24929 -15947 -22533
rect -17016 -26646 -16308 -26533
rect -17718 -27041 -17672 -26705
rect -18111 -27088 -17672 -27041
rect -19527 -27431 -19383 -27295
rect -19704 -27686 -19566 -27549
rect -19842 -27784 -19705 -27726
rect -13996 -22529 -13950 -22273
rect -13800 -22527 -13754 -22273
rect -13898 -22529 -13656 -22527
rect -13604 -22529 -13558 -22273
rect -13023 -22444 -12977 -22144
rect -13996 -22575 -13359 -22529
rect -13217 -22548 -13058 -22490
rect -13996 -22803 -13950 -22603
rect -13898 -22803 -13852 -22575
rect -13800 -22803 -13754 -22603
rect -13702 -22803 -13656 -22575
rect -13191 -22603 -13137 -22548
rect -13465 -22657 -13137 -22603
rect -13465 -22947 -13411 -22657
rect -15579 -23001 -13411 -22947
rect -13121 -22980 -13075 -22681
rect -15579 -24085 -15525 -23001
rect -13122 -23017 -13075 -22980
rect -13023 -22981 -12977 -22681
rect -12925 -23017 -12879 -22681
rect -12827 -22981 -12781 -22144
rect -12414 -22299 -12368 -22143
rect -12218 -22297 -12172 -22143
rect -12316 -22299 -12074 -22297
rect -12022 -22299 -11976 -22143
rect -12414 -22345 -11777 -22299
rect -12414 -22474 -12368 -22374
rect -12316 -22474 -12270 -22345
rect -12218 -22474 -12172 -22374
rect -12120 -22474 -12074 -22345
rect -11432 -22509 -11319 -20313
rect -12027 -22622 -11319 -22509
rect -12729 -23017 -12683 -22681
rect -13122 -23064 -12683 -23017
rect -15047 -23524 -15001 -23324
rect -14851 -23524 -14805 -23324
rect -14655 -23524 -14609 -23324
rect -14425 -23577 -14368 -23342
rect -14210 -23524 -14164 -23324
rect -14014 -23524 -13968 -23324
rect -13818 -23524 -13772 -23324
rect -13599 -23439 -13553 -23339
rect -13501 -23439 -13455 -23339
rect -13403 -23439 -13357 -23339
rect -13305 -23439 -13259 -23339
rect -13207 -23439 -13161 -23339
rect -13109 -23439 -13063 -23339
rect -13011 -23439 -12965 -23339
rect -12913 -23439 -12867 -23339
rect -12347 -23524 -12301 -23324
rect -12151 -23524 -12105 -23324
rect -11955 -23524 -11909 -23324
rect -13596 -23577 -13427 -23567
rect -14425 -23634 -13427 -23577
rect -11725 -23577 -11668 -23342
rect -11510 -23524 -11464 -23324
rect -11314 -23524 -11268 -23324
rect -11118 -23524 -11072 -23324
rect -10899 -23439 -10853 -23339
rect -10801 -23439 -10755 -23339
rect -10703 -23439 -10657 -23339
rect -10605 -23439 -10559 -23339
rect -10507 -23439 -10461 -23339
rect -10409 -23439 -10363 -23339
rect -10311 -23439 -10265 -23339
rect -10213 -23439 -10167 -23339
rect -10896 -23577 -10727 -23567
rect -12584 -23599 -12524 -23593
rect -12819 -23620 -12778 -23619
rect -13596 -23641 -13427 -23634
rect -15145 -23804 -15099 -23704
rect -15047 -23804 -15001 -23704
rect -14949 -23804 -14903 -23704
rect -14851 -23804 -14805 -23704
rect -14753 -23804 -14707 -23704
rect -14655 -23804 -14609 -23704
rect -14911 -24027 -14774 -23967
rect -15259 -24085 -15199 -24038
rect -15579 -24149 -15199 -24085
rect -15259 -24175 -15199 -24149
rect -14896 -24245 -14801 -24027
rect -14486 -24145 -14426 -23678
rect -12914 -23680 -12777 -23620
rect -12584 -23659 -12441 -23599
rect -11725 -23634 -10727 -23577
rect -10896 -23641 -10727 -23634
rect -14308 -23804 -14262 -23704
rect -14210 -23804 -14164 -23704
rect -14112 -23804 -14066 -23704
rect -14014 -23804 -13968 -23704
rect -13916 -23804 -13870 -23704
rect -13818 -23804 -13772 -23704
rect -13599 -23854 -13553 -23754
rect -13501 -23854 -13455 -23754
rect -13403 -23854 -13357 -23754
rect -13305 -23854 -13259 -23754
rect -13207 -23854 -13161 -23754
rect -13109 -23854 -13063 -23754
rect -13011 -23854 -12965 -23754
rect -12913 -23854 -12867 -23754
rect -14522 -24205 -14390 -24145
rect -12819 -24165 -12778 -23680
rect -12749 -24116 -12612 -24056
rect -14309 -24213 -12778 -24165
rect -14920 -24305 -14788 -24245
rect -15145 -24462 -15099 -24362
rect -15047 -24462 -15001 -24362
rect -14949 -24462 -14903 -24362
rect -14851 -24462 -14805 -24362
rect -14753 -24462 -14707 -24362
rect -14655 -24462 -14609 -24362
rect -14309 -24367 -14261 -24213
rect -14307 -24412 -14261 -24367
rect -14209 -24412 -14163 -24312
rect -14117 -24331 -14056 -24213
rect -14111 -24412 -14065 -24331
rect -14013 -24412 -13967 -24312
rect -13921 -24333 -13860 -24213
rect -13915 -24412 -13869 -24333
rect -13817 -24412 -13771 -24312
rect -13730 -24331 -13669 -24213
rect -13719 -24412 -13673 -24331
rect -13621 -24412 -13575 -24312
rect -13402 -24462 -13356 -24362
rect -13304 -24462 -13258 -24362
rect -13206 -24462 -13160 -24362
rect -13108 -24462 -13062 -24362
rect -13010 -24462 -12964 -24362
rect -12912 -24462 -12866 -24362
rect -13747 -24532 -13578 -24525
rect -13747 -24589 -12749 -24532
rect -12700 -24564 -12640 -24116
rect -12584 -24407 -12524 -23659
rect -10225 -23682 -10071 -23622
rect -12445 -23804 -12399 -23704
rect -12347 -23804 -12301 -23704
rect -12249 -23804 -12203 -23704
rect -12151 -23804 -12105 -23704
rect -12053 -23804 -12007 -23704
rect -11955 -23804 -11909 -23704
rect -12314 -24033 -12177 -23973
rect -12303 -24241 -12208 -24033
rect -11774 -24057 -11714 -23693
rect -11608 -23804 -11562 -23704
rect -11510 -23804 -11464 -23704
rect -11412 -23804 -11366 -23704
rect -11314 -23804 -11268 -23704
rect -11216 -23804 -11170 -23704
rect -11118 -23804 -11072 -23704
rect -10899 -23854 -10853 -23754
rect -10801 -23854 -10755 -23754
rect -10703 -23854 -10657 -23754
rect -10605 -23854 -10559 -23754
rect -10507 -23854 -10461 -23754
rect -10409 -23854 -10363 -23754
rect -10311 -23854 -10265 -23754
rect -10213 -23854 -10167 -23754
rect -10117 -23957 -10071 -23682
rect -10890 -24002 -10071 -23957
rect -9659 -23973 -9564 -20313
rect -10890 -24003 -10079 -24002
rect -11803 -24117 -11671 -24057
rect -10890 -24169 -10844 -24003
rect -9676 -24033 -9544 -23973
rect -11604 -24215 -10844 -24169
rect -9999 -24203 -9867 -24143
rect -12321 -24301 -12184 -24241
rect -11604 -24312 -11558 -24215
rect -11409 -24312 -11367 -24215
rect -11214 -24312 -11172 -24215
rect -11018 -24312 -10976 -24215
rect -12585 -24452 -12524 -24407
rect -12585 -24539 -12525 -24452
rect -12445 -24462 -12399 -24362
rect -12347 -24462 -12301 -24362
rect -12249 -24462 -12203 -24362
rect -12151 -24462 -12105 -24362
rect -12053 -24462 -12007 -24362
rect -11955 -24462 -11909 -24362
rect -11607 -24412 -11558 -24312
rect -11509 -24412 -11463 -24312
rect -11411 -24412 -11365 -24312
rect -11313 -24412 -11267 -24312
rect -11215 -24412 -11169 -24312
rect -11117 -24412 -11071 -24312
rect -11019 -24412 -10973 -24312
rect -10921 -24412 -10875 -24312
rect -10702 -24462 -10656 -24362
rect -10604 -24462 -10558 -24362
rect -10506 -24462 -10460 -24362
rect -10408 -24462 -10362 -24362
rect -10310 -24462 -10264 -24362
rect -10212 -24462 -10166 -24362
rect -9966 -24431 -9908 -24203
rect -9659 -24242 -9564 -24033
rect -9694 -24302 -9557 -24242
rect -11047 -24532 -10878 -24525
rect -13747 -24599 -13578 -24589
rect -15145 -24842 -15099 -24642
rect -14949 -24842 -14903 -24642
rect -14753 -24842 -14707 -24642
rect -14307 -24795 -14261 -24727
rect -14307 -24827 -14256 -24795
rect -14209 -24827 -14163 -24727
rect -14111 -24770 -14065 -24727
rect -14306 -24910 -14256 -24827
rect -14115 -24910 -14064 -24770
rect -14013 -24827 -13967 -24727
rect -13915 -24789 -13869 -24727
rect -13915 -24910 -13864 -24789
rect -13817 -24827 -13771 -24727
rect -13719 -24789 -13673 -24727
rect -13721 -24910 -13670 -24789
rect -13621 -24827 -13575 -24727
rect -13402 -24842 -13356 -24642
rect -13206 -24842 -13160 -24642
rect -13010 -24842 -12964 -24642
rect -12806 -24824 -12749 -24589
rect -11047 -24589 -10049 -24532
rect -9968 -24563 -9908 -24431
rect -9820 -24462 -9774 -24362
rect -9722 -24462 -9676 -24362
rect -9624 -24462 -9578 -24362
rect -9526 -24462 -9480 -24362
rect -9428 -24462 -9382 -24362
rect -9330 -24462 -9284 -24362
rect -11047 -24599 -10878 -24589
rect -12445 -24842 -12399 -24642
rect -12249 -24842 -12203 -24642
rect -12053 -24842 -12007 -24642
rect -11607 -24827 -11561 -24727
rect -11509 -24827 -11463 -24727
rect -11411 -24827 -11365 -24727
rect -11313 -24827 -11267 -24727
rect -11215 -24827 -11169 -24727
rect -11117 -24827 -11071 -24727
rect -11019 -24827 -10973 -24727
rect -10921 -24827 -10875 -24727
rect -10702 -24842 -10656 -24642
rect -10506 -24842 -10460 -24642
rect -10310 -24842 -10264 -24642
rect -10106 -24910 -10049 -24589
rect -9820 -24842 -9774 -24642
rect -9624 -24842 -9578 -24642
rect -9428 -24842 -9382 -24642
rect -14306 -24967 -10049 -24910
rect -9133 -27271 -8957 -20756
rect -8854 -23941 -8808 -23341
rect -8642 -23941 -8596 -23341
rect -8544 -23941 -8498 -23341
rect -8446 -23941 -8400 -23341
rect -8235 -23941 -8189 -23341
rect -8771 -24553 -8725 -24253
rect -8673 -24553 -8627 -24253
rect -8431 -24553 -8385 -24253
rect -8333 -24553 -8287 -24253
rect -8235 -24553 -8189 -24253
rect -9146 -27442 -8946 -27271
rect -7998 -27529 -7866 -19057
rect -7120 -19143 -7092 -18998
rect -6697 -18996 -6558 -18987
rect -5860 -18996 -5724 -18987
rect -6697 -19024 -5724 -18996
rect -6697 -19041 -6558 -19024
rect -5860 -19033 -5724 -19024
rect -7064 -19070 -6925 -19061
rect -5986 -19068 -5847 -19067
rect -5986 -19070 -5455 -19068
rect -7064 -19096 -5455 -19070
rect -7064 -19098 -5847 -19096
rect -7064 -19115 -6925 -19098
rect -5986 -19121 -5847 -19098
rect -6166 -19143 -6035 -19131
rect -7120 -19171 -6035 -19143
rect -6166 -19177 -6035 -19171
rect -7451 -19409 -7405 -19209
rect -7353 -19409 -7307 -19209
rect -7037 -19409 -6991 -19209
rect -6939 -19409 -6893 -19209
rect -6675 -19409 -6629 -19209
rect -6577 -19409 -6531 -19209
rect -6381 -19409 -6335 -19209
rect -6283 -19409 -6237 -19209
rect -6071 -19409 -6025 -19209
rect -5973 -19409 -5927 -19209
rect -5762 -19409 -5716 -19209
rect -5664 -19409 -5618 -19209
rect -7014 -19752 -6968 -19652
rect -6916 -19752 -6870 -19652
rect -6818 -19752 -6772 -19652
rect -6720 -19752 -6674 -19652
rect -6622 -19752 -6576 -19652
rect -6524 -19752 -6478 -19652
rect -5483 -19735 -5455 -19096
rect -5501 -19871 -5455 -19735
rect -6916 -20132 -6870 -19932
rect -6720 -20132 -6674 -19932
rect -6524 -20132 -6478 -19932
rect -5411 -20167 -5383 -18959
rect -4946 -18970 -4807 -18957
rect -3788 -18959 -2812 -18931
rect -3788 -18967 -3649 -18959
rect -4946 -18998 -4592 -18970
rect -3173 -18973 -3034 -18959
rect -4946 -19011 -4807 -18998
rect -4620 -19143 -4592 -18998
rect -4197 -18996 -4058 -18987
rect -3360 -18996 -3224 -18987
rect -4197 -19024 -3224 -18996
rect -4197 -19041 -4058 -19024
rect -3360 -19033 -3224 -19024
rect -3666 -19143 -3535 -19131
rect -4620 -19171 -3535 -19143
rect -3666 -19177 -3535 -19171
rect -5119 -19376 -5073 -19240
rect -5118 -19946 -5074 -19376
rect -4951 -19409 -4905 -19209
rect -4853 -19409 -4807 -19209
rect -4537 -19409 -4491 -19209
rect -4439 -19409 -4393 -19209
rect -4175 -19409 -4129 -19209
rect -4077 -19409 -4031 -19209
rect -3881 -19409 -3835 -19209
rect -3783 -19409 -3737 -19209
rect -3571 -19409 -3525 -19209
rect -3473 -19409 -3427 -19209
rect -3262 -19409 -3216 -19209
rect -3164 -19409 -3118 -19209
rect -5119 -20082 -5073 -19946
rect -2840 -20017 -2812 -18959
rect -2446 -18970 -2307 -18957
rect -1288 -18959 -340 -18931
rect -1288 -18967 -1149 -18959
rect -2446 -18998 -2092 -18970
rect -673 -18973 -534 -18959
rect -2446 -19011 -2307 -18998
rect -2120 -19143 -2092 -18998
rect -1697 -18996 -1558 -18987
rect -860 -18996 -724 -18987
rect -1697 -19024 -724 -18996
rect -1697 -19041 -1558 -19024
rect -860 -19033 -724 -19024
rect -1166 -19143 -1035 -19131
rect -2120 -19171 -1035 -19143
rect -1166 -19177 -1035 -19171
rect -2571 -19380 -2525 -19244
rect -2570 -19617 -2526 -19380
rect -2451 -19409 -2405 -19209
rect -2353 -19409 -2307 -19209
rect -2037 -19409 -1991 -19209
rect -1939 -19409 -1893 -19209
rect -1675 -19409 -1629 -19209
rect -1577 -19409 -1531 -19209
rect -1381 -19409 -1335 -19209
rect -1283 -19409 -1237 -19209
rect -1071 -19409 -1025 -19209
rect -973 -19409 -927 -19209
rect -762 -19409 -716 -19209
rect -664 -19409 -618 -19209
rect -2406 -19617 -2270 -19616
rect -2571 -19661 -2270 -19617
rect -2406 -19662 -2270 -19661
rect -368 -19904 -340 -18959
rect 54 -18970 193 -18957
rect 1212 -18959 2135 -18931
rect 1212 -18967 1351 -18959
rect 54 -18998 408 -18970
rect 1827 -18973 1966 -18959
rect 54 -19011 193 -18998
rect 380 -19143 408 -18998
rect 803 -18996 942 -18987
rect 1640 -18996 1776 -18987
rect 803 -19024 1776 -18996
rect 803 -19041 942 -19024
rect 1640 -19033 1776 -19024
rect 1334 -19143 1465 -19131
rect 380 -19171 1465 -19143
rect 1334 -19177 1465 -19171
rect -91 -19380 -45 -19244
rect -90 -19630 -46 -19380
rect 49 -19409 95 -19209
rect 147 -19409 193 -19209
rect 463 -19409 509 -19209
rect 561 -19409 607 -19209
rect 825 -19409 871 -19209
rect 923 -19409 969 -19209
rect 1119 -19409 1165 -19209
rect 1217 -19409 1263 -19209
rect 1429 -19409 1475 -19209
rect 1527 -19409 1573 -19209
rect 1738 -19409 1784 -19209
rect 1836 -19409 1882 -19209
rect 91 -19630 227 -19629
rect -90 -19674 227 -19630
rect 91 -19675 227 -19674
rect 2107 -19767 2135 -18959
rect 2554 -18970 2693 -18957
rect 3712 -18959 5440 -18931
rect 3712 -18967 3851 -18959
rect 2554 -18998 2908 -18970
rect 4327 -18973 4466 -18959
rect 2554 -19011 2693 -18998
rect 2880 -19143 2908 -18998
rect 3303 -18996 3442 -18987
rect 4140 -18996 4276 -18987
rect 3303 -19024 4276 -18996
rect 3303 -19041 3442 -19024
rect 4140 -19033 4276 -19024
rect 3834 -19143 3965 -19131
rect 2880 -19171 3965 -19143
rect 3834 -19177 3965 -19171
rect 2326 -19380 2372 -19244
rect 2327 -19692 2371 -19380
rect 2549 -19409 2595 -19209
rect 2647 -19409 2693 -19209
rect 2963 -19409 3009 -19209
rect 3061 -19409 3107 -19209
rect 3325 -19409 3371 -19209
rect 3423 -19409 3469 -19209
rect 3619 -19409 3665 -19209
rect 3717 -19409 3763 -19209
rect 3929 -19409 3975 -19209
rect 4027 -19409 4073 -19209
rect 4238 -19409 4284 -19209
rect 4336 -19409 4382 -19209
rect 5231 -19380 5277 -19244
rect 5232 -19676 5276 -19380
rect 2274 -19738 2410 -19692
rect 5179 -19722 5315 -19676
rect 5412 -19634 5440 -18959
rect 5554 -18970 5693 -18957
rect 6712 -18959 9597 -18931
rect 6712 -18967 6851 -18959
rect 5554 -18998 5908 -18970
rect 7327 -18973 7466 -18959
rect 5554 -19011 5693 -18998
rect 5880 -19143 5908 -18998
rect 6303 -18996 6442 -18987
rect 7140 -18996 7276 -18987
rect 6303 -19024 7276 -18996
rect 6303 -19041 6442 -19024
rect 7140 -19033 7276 -19024
rect 6834 -19143 6965 -19131
rect 5880 -19171 6965 -19143
rect 6834 -19177 6965 -19171
rect 5549 -19409 5595 -19209
rect 5647 -19409 5693 -19209
rect 5963 -19409 6009 -19209
rect 6061 -19409 6107 -19209
rect 6325 -19409 6371 -19209
rect 6423 -19409 6469 -19209
rect 6619 -19409 6665 -19209
rect 6717 -19409 6763 -19209
rect 6929 -19409 6975 -19209
rect 7027 -19409 7073 -19209
rect 7238 -19409 7284 -19209
rect 7336 -19409 7382 -19209
rect 8240 -19634 9432 -19517
rect 5412 -19662 9441 -19634
rect 2107 -19805 9288 -19767
rect -368 -19932 9136 -19904
rect -2840 -20068 8977 -20017
rect -5411 -20218 8821 -20167
rect -5116 -20337 -4980 -20335
rect 1933 -20337 2069 -20333
rect -5116 -20379 2069 -20337
rect -5116 -20381 -4980 -20379
rect -7596 -20419 -7460 -20417
rect 1829 -20419 1984 -20417
rect -7596 -20461 1984 -20419
rect -7596 -20463 -7460 -20461
rect 1829 -20463 1984 -20461
rect -1363 -20554 8600 -20503
rect -7271 -21035 -7225 -20835
rect -7075 -21035 -7029 -20835
rect -6879 -21035 -6833 -20835
rect -6433 -20950 -6387 -20850
rect -6335 -20950 -6289 -20850
rect -6237 -20950 -6191 -20850
rect -6139 -20950 -6093 -20850
rect -6041 -20950 -5995 -20850
rect -5943 -20950 -5897 -20850
rect -5845 -20950 -5799 -20850
rect -5747 -20950 -5701 -20850
rect -5528 -21035 -5482 -20835
rect -5332 -21035 -5286 -20835
rect -5136 -21035 -5090 -20835
rect -5873 -21088 -5704 -21078
rect -4932 -21088 -4875 -20853
rect -4571 -21035 -4525 -20835
rect -4375 -21035 -4329 -20835
rect -4179 -21035 -4133 -20835
rect -3733 -20950 -3687 -20850
rect -3635 -20950 -3589 -20850
rect -3537 -20950 -3491 -20850
rect -3439 -20950 -3393 -20850
rect -3341 -20950 -3295 -20850
rect -3243 -20950 -3197 -20850
rect -3145 -20950 -3099 -20850
rect -3047 -20950 -3001 -20850
rect -2828 -21035 -2782 -20835
rect -2632 -21035 -2586 -20835
rect -2436 -21035 -2390 -20835
rect -5873 -21145 -4875 -21088
rect -3173 -21088 -3004 -21078
rect -2232 -21088 -2175 -20853
rect -1946 -21035 -1900 -20835
rect -1750 -21035 -1704 -20835
rect -1554 -21035 -1508 -20835
rect -1016 -21052 -970 -20852
rect -278 -21052 -232 -20852
rect -82 -21052 -36 -20852
rect 114 -21052 160 -20852
rect 340 -21013 386 -21011
rect -5873 -21152 -5704 -21145
rect -7271 -21315 -7225 -21215
rect -7173 -21315 -7127 -21215
rect -7075 -21315 -7029 -21215
rect -6977 -21315 -6931 -21215
rect -6879 -21315 -6833 -21215
rect -6781 -21315 -6735 -21215
rect -6433 -21310 -6387 -21265
rect -7046 -21432 -6914 -21372
rect -7385 -21528 -7325 -21502
rect -7740 -21591 -7325 -21528
rect -7723 -21592 -7325 -21591
rect -7385 -21639 -7325 -21592
rect -7022 -21650 -6927 -21432
rect -6435 -21464 -6387 -21310
rect -6335 -21365 -6289 -21265
rect -6237 -21346 -6191 -21265
rect -6243 -21464 -6182 -21346
rect -6139 -21365 -6093 -21265
rect -6041 -21344 -5995 -21265
rect -6047 -21464 -5986 -21344
rect -5943 -21365 -5897 -21265
rect -5845 -21346 -5799 -21265
rect -5856 -21464 -5795 -21346
rect -5747 -21365 -5701 -21265
rect -5528 -21315 -5482 -21215
rect -5430 -21315 -5384 -21215
rect -5332 -21315 -5286 -21215
rect -5234 -21315 -5188 -21215
rect -5136 -21315 -5090 -21215
rect -5038 -21315 -4992 -21215
rect -6648 -21532 -6516 -21472
rect -6435 -21512 -4904 -21464
rect -7037 -21710 -6900 -21650
rect -7271 -21973 -7225 -21873
rect -7173 -21973 -7127 -21873
rect -7075 -21973 -7029 -21873
rect -6977 -21973 -6931 -21873
rect -6879 -21973 -6833 -21873
rect -6781 -21973 -6735 -21873
rect -6612 -21999 -6552 -21532
rect -6434 -21973 -6388 -21873
rect -6336 -21973 -6290 -21873
rect -6238 -21973 -6192 -21873
rect -6140 -21973 -6094 -21873
rect -6042 -21973 -5996 -21873
rect -5944 -21973 -5898 -21873
rect -5725 -21923 -5679 -21823
rect -5627 -21923 -5581 -21823
rect -5529 -21923 -5483 -21823
rect -5431 -21923 -5385 -21823
rect -5333 -21923 -5287 -21823
rect -5235 -21923 -5189 -21823
rect -5137 -21923 -5091 -21823
rect -5039 -21923 -4993 -21823
rect -4945 -21997 -4904 -21512
rect -4826 -21561 -4766 -21113
rect -4711 -21225 -4651 -21138
rect -3173 -21145 -2175 -21088
rect -3173 -21152 -3004 -21145
rect -4711 -21270 -4650 -21225
rect -4875 -21621 -4738 -21561
rect -5722 -22043 -5553 -22036
rect -6551 -22100 -5553 -22043
rect -5040 -22057 -4903 -21997
rect -4710 -22018 -4650 -21270
rect -4571 -21315 -4525 -21215
rect -4473 -21315 -4427 -21215
rect -4375 -21315 -4329 -21215
rect -4277 -21315 -4231 -21215
rect -4179 -21315 -4133 -21215
rect -4081 -21315 -4035 -21215
rect -3733 -21365 -3684 -21265
rect -3635 -21365 -3589 -21265
rect -3537 -21365 -3491 -21265
rect -3439 -21365 -3393 -21265
rect -3341 -21365 -3295 -21265
rect -3243 -21365 -3197 -21265
rect -3145 -21365 -3099 -21265
rect -3047 -21365 -3001 -21265
rect -2828 -21315 -2782 -21215
rect -2730 -21315 -2684 -21215
rect -2632 -21315 -2586 -21215
rect -2534 -21315 -2488 -21215
rect -2436 -21315 -2390 -21215
rect -2338 -21315 -2292 -21215
rect -4447 -21436 -4310 -21376
rect -4429 -21644 -4334 -21436
rect -3730 -21462 -3684 -21365
rect -3535 -21462 -3493 -21365
rect -3340 -21462 -3298 -21365
rect -3144 -21462 -3102 -21365
rect -3730 -21508 -2970 -21462
rect -3929 -21620 -3797 -21560
rect -4440 -21704 -4303 -21644
rect -4571 -21973 -4525 -21873
rect -4473 -21973 -4427 -21873
rect -4375 -21973 -4329 -21873
rect -4277 -21973 -4231 -21873
rect -4179 -21973 -4133 -21873
rect -4081 -21973 -4035 -21873
rect -3900 -21984 -3840 -21620
rect -3016 -21674 -2970 -21508
rect -2232 -21582 -2175 -21145
rect -2094 -21246 -2034 -21114
rect 332 -21147 386 -21013
rect 717 -21021 763 -20865
rect 913 -21019 959 -20865
rect 815 -21021 1057 -21019
rect 1109 -21021 1155 -20865
rect 692 -21067 1155 -21021
rect -2092 -21474 -2034 -21246
rect -1946 -21315 -1900 -21215
rect -1848 -21315 -1802 -21215
rect -1750 -21315 -1704 -21215
rect -1652 -21315 -1606 -21215
rect -1554 -21315 -1508 -21215
rect -1456 -21315 -1410 -21215
rect -1161 -21311 -1020 -21258
rect -1690 -21435 -1553 -21375
rect -2092 -21532 -1853 -21474
rect -1911 -21561 -1853 -21532
rect -2232 -21639 -1966 -21582
rect -1915 -21621 -1783 -21561
rect -3016 -21675 -2205 -21674
rect -3016 -21720 -2197 -21675
rect -3734 -21973 -3688 -21873
rect -3636 -21973 -3590 -21873
rect -3538 -21973 -3492 -21873
rect -3440 -21973 -3394 -21873
rect -3342 -21973 -3296 -21873
rect -3244 -21973 -3198 -21873
rect -3025 -21923 -2979 -21823
rect -2927 -21923 -2881 -21823
rect -2829 -21923 -2783 -21823
rect -2731 -21923 -2685 -21823
rect -2633 -21923 -2587 -21823
rect -2535 -21923 -2489 -21823
rect -2437 -21923 -2391 -21823
rect -2339 -21923 -2293 -21823
rect -2243 -21995 -2197 -21720
rect -2023 -21760 -1966 -21639
rect -1655 -21644 -1560 -21435
rect -1672 -21704 -1540 -21644
rect -1161 -21760 -1104 -21311
rect -1016 -21760 -970 -21560
rect -918 -21760 -872 -21560
rect -603 -21760 -557 -21460
rect -505 -21760 -459 -21460
rect -407 -21760 -361 -21460
rect -294 -21760 -248 -21460
rect -196 -21760 -150 -21460
rect -98 -21760 -52 -21460
rect 16 -21759 62 -21459
rect 114 -21759 160 -21459
rect 212 -21759 258 -21459
rect -2023 -21817 -1104 -21760
rect -4945 -22058 -4904 -22057
rect -4710 -22078 -4567 -22018
rect -3022 -22043 -2853 -22036
rect -4710 -22084 -4650 -22078
rect -7173 -22353 -7127 -22153
rect -6977 -22353 -6931 -22153
rect -6781 -22353 -6735 -22153
rect -6551 -22335 -6494 -22100
rect -5722 -22110 -5553 -22100
rect -3851 -22100 -2853 -22043
rect -2351 -22055 -2197 -21995
rect 332 -21952 378 -21147
rect 421 -21231 557 -21185
rect 815 -21196 861 -21067
rect 913 -21196 959 -21096
rect 1011 -21196 1057 -21067
rect 1109 -21196 1155 -21096
rect 485 -21840 531 -21231
rect 1424 -21739 1470 -21403
rect 1522 -21703 1568 -20866
rect 1718 -21166 1764 -20866
rect 2322 -21023 2368 -20867
rect 2518 -21021 2564 -20867
rect 2420 -21023 2662 -21021
rect 2714 -21023 2760 -20867
rect 2297 -21069 2760 -21023
rect 2420 -21198 2466 -21069
rect 2518 -21198 2564 -21098
rect 2616 -21198 2662 -21069
rect 2714 -21198 2760 -21098
rect 1620 -21739 1666 -21403
rect 1718 -21703 1764 -21403
rect 1816 -21702 1862 -21403
rect 1816 -21739 1863 -21702
rect 1424 -21786 1863 -21739
rect 3029 -21741 3075 -21405
rect 3127 -21705 3173 -20868
rect 3323 -21168 3369 -20868
rect 3946 -21043 3992 -20843
rect 4684 -21043 4730 -20843
rect 4880 -21043 4926 -20843
rect 5076 -21043 5122 -20843
rect 5559 -21054 5605 -20854
rect 5657 -21085 5703 -20854
rect 5755 -21054 5801 -20854
rect 5875 -21054 5921 -20854
rect 5973 -21054 6019 -20854
rect 6071 -21054 6117 -20854
rect 6433 -21054 6479 -20854
rect 6629 -21054 6675 -20854
rect 6939 -21054 6985 -20854
rect 7248 -21054 7294 -20854
rect 5151 -21131 5703 -21085
rect 5155 -21140 5291 -21131
rect 6722 -21182 6861 -21164
rect 7337 -21175 7476 -21170
rect 8268 -21175 8486 -21116
rect 7337 -21182 8486 -21175
rect 6722 -21203 8486 -21182
rect 5564 -21221 5703 -21208
rect 6722 -21210 7577 -21203
rect 8268 -21205 8486 -21203
rect 6722 -21218 6861 -21210
rect 5564 -21249 5918 -21221
rect 7337 -21224 7476 -21210
rect 5564 -21262 5703 -21249
rect 5890 -21394 5918 -21249
rect 6313 -21247 6452 -21238
rect 7150 -21247 7286 -21238
rect 6313 -21275 7286 -21247
rect 6313 -21292 6452 -21275
rect 7150 -21284 7286 -21275
rect 6844 -21394 6975 -21382
rect 3225 -21741 3271 -21405
rect 3323 -21705 3369 -21405
rect 3421 -21704 3467 -21405
rect 5890 -21422 6975 -21394
rect 6844 -21428 6975 -21422
rect 3421 -21741 3468 -21704
rect 3029 -21788 3468 -21741
rect 3946 -21751 3992 -21551
rect 4044 -21751 4090 -21551
rect 4359 -21751 4405 -21451
rect 4457 -21751 4503 -21451
rect 4555 -21751 4601 -21451
rect 4668 -21751 4714 -21451
rect 4766 -21751 4812 -21451
rect 4864 -21751 4910 -21451
rect 4978 -21750 5024 -21450
rect 5076 -21750 5122 -21450
rect 5174 -21750 5220 -21450
rect 5559 -21660 5605 -21460
rect 5657 -21660 5703 -21460
rect 5973 -21660 6019 -21460
rect 6071 -21660 6117 -21460
rect 6335 -21660 6381 -21460
rect 6433 -21660 6479 -21460
rect 6629 -21660 6675 -21460
rect 6727 -21660 6773 -21460
rect 6939 -21660 6985 -21460
rect 7037 -21660 7083 -21460
rect 7248 -21660 7294 -21460
rect 7346 -21660 7392 -21460
rect 485 -21886 2234 -21840
rect 332 -21998 3802 -21952
rect -6336 -22353 -6290 -22153
rect -6140 -22353 -6094 -22153
rect -5944 -22353 -5898 -22153
rect -5725 -22338 -5679 -22238
rect -5627 -22338 -5581 -22238
rect -5529 -22338 -5483 -22238
rect -5431 -22338 -5385 -22238
rect -5333 -22338 -5287 -22238
rect -5235 -22338 -5189 -22238
rect -5137 -22338 -5091 -22238
rect -5039 -22338 -4993 -22238
rect -4473 -22353 -4427 -22153
rect -4277 -22353 -4231 -22153
rect -4081 -22353 -4035 -22153
rect -3851 -22335 -3794 -22100
rect -3022 -22110 -2853 -22100
rect -3636 -22353 -3590 -22153
rect -3440 -22353 -3394 -22153
rect -3244 -22353 -3198 -22153
rect -3025 -22338 -2979 -22238
rect -2927 -22338 -2881 -22238
rect -2829 -22338 -2783 -22238
rect -2731 -22338 -2685 -22238
rect -2633 -22338 -2587 -22238
rect -2535 -22338 -2489 -22238
rect -2437 -22338 -2391 -22238
rect -2339 -22338 -2293 -22238
rect -7173 -23791 -7127 -23591
rect -6977 -23791 -6931 -23591
rect -6781 -23791 -6735 -23591
rect -6551 -23844 -6494 -23609
rect -6336 -23791 -6290 -23591
rect -6140 -23791 -6094 -23591
rect -5944 -23791 -5898 -23591
rect -5725 -23706 -5679 -23606
rect -5627 -23706 -5581 -23606
rect -5529 -23706 -5483 -23606
rect -5431 -23706 -5385 -23606
rect -5333 -23706 -5287 -23606
rect -5235 -23706 -5189 -23606
rect -5137 -23706 -5091 -23606
rect -5039 -23706 -4993 -23606
rect -4473 -23791 -4427 -23591
rect -4277 -23791 -4231 -23591
rect -4081 -23791 -4035 -23591
rect -5722 -23844 -5553 -23834
rect -6551 -23901 -5553 -23844
rect -3851 -23844 -3794 -23609
rect -3636 -23791 -3590 -23591
rect -3440 -23791 -3394 -23591
rect -3244 -23791 -3198 -23591
rect -3025 -23706 -2979 -23606
rect -2927 -23706 -2881 -23606
rect -2829 -23706 -2783 -23606
rect -2731 -23706 -2685 -23606
rect -2633 -23706 -2587 -23606
rect -2535 -23706 -2489 -23606
rect -2437 -23706 -2391 -23606
rect -2339 -23706 -2293 -23606
rect -3022 -23844 -2853 -23834
rect -4710 -23866 -4650 -23860
rect -4945 -23887 -4904 -23886
rect -5722 -23908 -5553 -23901
rect -7271 -24071 -7225 -23971
rect -7173 -24071 -7127 -23971
rect -7075 -24071 -7029 -23971
rect -6977 -24071 -6931 -23971
rect -6879 -24071 -6833 -23971
rect -6781 -24071 -6735 -23971
rect -7731 -24352 -7556 -24133
rect -7037 -24294 -6900 -24234
rect -7385 -24352 -7325 -24305
rect -7731 -24416 -7325 -24352
rect -7731 -24447 -7556 -24416
rect -7385 -24442 -7325 -24416
rect -7022 -24482 -6927 -24294
rect -6612 -24412 -6552 -23945
rect -5040 -23947 -4903 -23887
rect -4710 -23926 -4567 -23866
rect -3851 -23901 -2853 -23844
rect -3022 -23908 -2853 -23901
rect -6434 -24071 -6388 -23971
rect -6336 -24071 -6290 -23971
rect -6238 -24071 -6192 -23971
rect -6140 -24071 -6094 -23971
rect -6042 -24071 -5996 -23971
rect -5944 -24071 -5898 -23971
rect -5725 -24121 -5679 -24021
rect -5627 -24121 -5581 -24021
rect -5529 -24121 -5483 -24021
rect -5431 -24121 -5385 -24021
rect -5333 -24121 -5287 -24021
rect -5235 -24121 -5189 -24021
rect -5137 -24121 -5091 -24021
rect -5039 -24121 -4993 -24021
rect -6648 -24472 -6516 -24412
rect -4945 -24432 -4904 -23947
rect -4875 -24383 -4738 -24323
rect -7509 -24512 -6927 -24482
rect -6435 -24480 -4904 -24432
rect -7509 -24572 -6914 -24512
rect -7509 -24577 -6927 -24572
rect -7509 -24656 -7414 -24577
rect -7724 -24751 -7414 -24656
rect -7271 -24729 -7225 -24629
rect -7173 -24729 -7127 -24629
rect -7075 -24729 -7029 -24629
rect -6977 -24729 -6931 -24629
rect -6879 -24729 -6833 -24629
rect -6781 -24729 -6735 -24629
rect -6435 -24634 -6387 -24480
rect -6433 -24679 -6387 -24634
rect -6335 -24679 -6289 -24579
rect -6243 -24598 -6182 -24480
rect -6237 -24679 -6191 -24598
rect -6139 -24679 -6093 -24579
rect -6047 -24600 -5986 -24480
rect -6041 -24679 -5995 -24600
rect -5943 -24679 -5897 -24579
rect -5856 -24598 -5795 -24480
rect -5845 -24679 -5799 -24598
rect -5747 -24679 -5701 -24579
rect -5528 -24729 -5482 -24629
rect -5430 -24729 -5384 -24629
rect -5332 -24729 -5286 -24629
rect -5234 -24729 -5188 -24629
rect -5136 -24729 -5090 -24629
rect -5038 -24729 -4992 -24629
rect -5873 -24799 -5704 -24792
rect -5873 -24856 -4875 -24799
rect -4826 -24831 -4766 -24383
rect -4710 -24674 -4650 -23926
rect -2351 -23949 -2197 -23889
rect -4571 -24071 -4525 -23971
rect -4473 -24071 -4427 -23971
rect -4375 -24071 -4329 -23971
rect -4277 -24071 -4231 -23971
rect -4179 -24071 -4133 -23971
rect -4081 -24071 -4035 -23971
rect -4440 -24300 -4303 -24240
rect -4429 -24508 -4334 -24300
rect -3900 -24324 -3840 -23960
rect -3734 -24071 -3688 -23971
rect -3636 -24071 -3590 -23971
rect -3538 -24071 -3492 -23971
rect -3440 -24071 -3394 -23971
rect -3342 -24071 -3296 -23971
rect -3244 -24071 -3198 -23971
rect -3025 -24121 -2979 -24021
rect -2927 -24121 -2881 -24021
rect -2829 -24121 -2783 -24021
rect -2731 -24121 -2685 -24021
rect -2633 -24121 -2587 -24021
rect -2535 -24121 -2489 -24021
rect -2437 -24121 -2391 -24021
rect -2339 -24121 -2293 -24021
rect -2243 -24224 -2197 -23949
rect 332 -23992 3802 -23946
rect -3016 -24269 -2197 -24224
rect -2023 -24184 -1104 -24127
rect -3016 -24270 -2205 -24269
rect -3929 -24384 -3797 -24324
rect -3016 -24436 -2970 -24270
rect -2023 -24305 -1966 -24184
rect -1802 -24300 -1670 -24240
rect -3730 -24482 -2970 -24436
rect -2232 -24362 -1966 -24305
rect -4447 -24568 -4310 -24508
rect -3730 -24579 -3684 -24482
rect -3535 -24579 -3493 -24482
rect -3340 -24579 -3298 -24482
rect -3144 -24579 -3102 -24482
rect -4711 -24719 -4650 -24674
rect -4711 -24806 -4651 -24719
rect -4571 -24729 -4525 -24629
rect -4473 -24729 -4427 -24629
rect -4375 -24729 -4329 -24629
rect -4277 -24729 -4231 -24629
rect -4179 -24729 -4133 -24629
rect -4081 -24729 -4035 -24629
rect -3733 -24679 -3684 -24579
rect -3635 -24679 -3589 -24579
rect -3537 -24679 -3491 -24579
rect -3439 -24679 -3393 -24579
rect -3341 -24679 -3295 -24579
rect -3243 -24679 -3197 -24579
rect -3145 -24679 -3099 -24579
rect -3047 -24679 -3001 -24579
rect -2828 -24729 -2782 -24629
rect -2730 -24729 -2684 -24629
rect -2632 -24729 -2586 -24629
rect -2534 -24729 -2488 -24629
rect -2436 -24729 -2390 -24629
rect -2338 -24729 -2292 -24629
rect -3173 -24799 -3004 -24792
rect -2232 -24799 -2175 -24362
rect -2125 -24470 -1993 -24410
rect -2092 -24698 -2034 -24470
rect -1785 -24509 -1690 -24300
rect -1820 -24569 -1683 -24509
rect -5873 -24866 -5704 -24856
rect -7271 -25109 -7225 -24909
rect -7075 -25109 -7029 -24909
rect -6879 -25109 -6833 -24909
rect -6433 -25094 -6387 -24994
rect -6335 -25094 -6289 -24994
rect -6237 -25094 -6191 -24994
rect -6139 -25094 -6093 -24994
rect -6041 -25094 -5995 -24994
rect -5943 -25094 -5897 -24994
rect -5845 -25094 -5799 -24994
rect -5747 -25094 -5701 -24994
rect -5528 -25109 -5482 -24909
rect -5332 -25109 -5286 -24909
rect -5136 -25109 -5090 -24909
rect -4932 -25091 -4875 -24856
rect -3173 -24856 -2175 -24799
rect -2094 -24830 -2034 -24698
rect -1946 -24729 -1900 -24629
rect -1848 -24729 -1802 -24629
rect -1750 -24729 -1704 -24629
rect -1652 -24729 -1606 -24629
rect -1554 -24729 -1508 -24629
rect -1456 -24729 -1410 -24629
rect -1161 -24633 -1104 -24184
rect -1016 -24384 -970 -24184
rect -918 -24384 -872 -24184
rect -603 -24484 -557 -24184
rect -505 -24484 -459 -24184
rect -407 -24484 -361 -24184
rect -294 -24484 -248 -24184
rect -196 -24484 -150 -24184
rect -98 -24484 -52 -24184
rect 16 -24485 62 -24185
rect 114 -24485 160 -24185
rect 212 -24485 258 -24185
rect -1161 -24686 -1020 -24633
rect 332 -24797 378 -23992
rect 485 -24104 2234 -24058
rect 485 -24713 531 -24104
rect 1424 -24205 1863 -24158
rect 1424 -24541 1470 -24205
rect 421 -24759 557 -24713
rect -3173 -24866 -3004 -24856
rect -4571 -25109 -4525 -24909
rect -4375 -25109 -4329 -24909
rect -4179 -25109 -4133 -24909
rect -3733 -25094 -3687 -24994
rect -3635 -25094 -3589 -24994
rect -3537 -25094 -3491 -24994
rect -3439 -25094 -3393 -24994
rect -3341 -25094 -3295 -24994
rect -3243 -25094 -3197 -24994
rect -3145 -25094 -3099 -24994
rect -3047 -25094 -3001 -24994
rect -2828 -25109 -2782 -24909
rect -2632 -25109 -2586 -24909
rect -2436 -25109 -2390 -24909
rect -2232 -25091 -2175 -24856
rect -1946 -25109 -1900 -24909
rect -1750 -25109 -1704 -24909
rect -1554 -25109 -1508 -24909
rect -1016 -25092 -970 -24892
rect -278 -25092 -232 -24892
rect -82 -25092 -36 -24892
rect 114 -25092 160 -24892
rect 332 -24931 386 -24797
rect 815 -24877 861 -24748
rect 913 -24848 959 -24748
rect 1011 -24877 1057 -24748
rect 1109 -24848 1155 -24748
rect 692 -24923 1155 -24877
rect 340 -24933 386 -24931
rect 717 -25079 763 -24923
rect 815 -24925 1057 -24923
rect 913 -25079 959 -24925
rect 1109 -25079 1155 -24923
rect 1522 -25078 1568 -24241
rect 1620 -24541 1666 -24205
rect 1718 -24541 1764 -24241
rect 1816 -24242 1863 -24205
rect 3029 -24203 3468 -24156
rect 1816 -24541 1862 -24242
rect 3029 -24539 3075 -24203
rect 1718 -25078 1764 -24778
rect 2420 -24875 2466 -24746
rect 2518 -24846 2564 -24746
rect 2616 -24875 2662 -24746
rect 2714 -24846 2760 -24746
rect 2297 -24921 2760 -24875
rect 2322 -25077 2368 -24921
rect 2420 -24923 2662 -24921
rect 2518 -25077 2564 -24923
rect 2714 -25077 2760 -24921
rect 3127 -25076 3173 -24239
rect 3225 -24539 3271 -24203
rect 3323 -24539 3369 -24239
rect 3421 -24240 3468 -24203
rect 3421 -24539 3467 -24240
rect 3946 -24393 3992 -24193
rect 4044 -24393 4090 -24193
rect 4359 -24493 4405 -24193
rect 4457 -24493 4503 -24193
rect 4555 -24493 4601 -24193
rect 4668 -24493 4714 -24193
rect 4766 -24493 4812 -24193
rect 4864 -24493 4910 -24193
rect 4978 -24494 5024 -24194
rect 5076 -24494 5122 -24194
rect 5174 -24494 5220 -24194
rect 5559 -24484 5605 -24284
rect 5657 -24484 5703 -24284
rect 5973 -24484 6019 -24284
rect 6071 -24484 6117 -24284
rect 6335 -24484 6381 -24284
rect 6433 -24484 6479 -24284
rect 6629 -24484 6675 -24284
rect 6727 -24484 6773 -24284
rect 6939 -24484 6985 -24284
rect 7037 -24484 7083 -24284
rect 7248 -24484 7294 -24284
rect 7346 -24484 7392 -24284
rect 6844 -24522 6975 -24516
rect 5890 -24550 6975 -24522
rect 5564 -24695 5703 -24682
rect 5890 -24695 5918 -24550
rect 6844 -24562 6975 -24550
rect 5564 -24723 5918 -24695
rect 6313 -24669 6452 -24652
rect 7150 -24669 7286 -24660
rect 6313 -24697 7286 -24669
rect 6313 -24706 6452 -24697
rect 7150 -24706 7286 -24697
rect 5564 -24736 5703 -24723
rect 6722 -24734 6861 -24726
rect 7337 -24734 7476 -24720
rect 6722 -24741 7577 -24734
rect 8435 -24741 8463 -21205
rect 6722 -24762 8463 -24741
rect 3323 -25076 3369 -24776
rect 6722 -24780 6861 -24762
rect 7337 -24769 8463 -24762
rect 7337 -24774 7476 -24769
rect 5155 -24813 5291 -24804
rect 5151 -24859 5703 -24813
rect 3946 -25101 3992 -24901
rect 4684 -25101 4730 -24901
rect 4880 -25101 4926 -24901
rect 5076 -25101 5122 -24901
rect 5559 -25090 5605 -24890
rect 5657 -25090 5703 -24859
rect 5755 -25090 5801 -24890
rect 5875 -25090 5921 -24890
rect 5973 -25090 6019 -24890
rect 6071 -25090 6117 -24890
rect 6433 -25090 6479 -24890
rect 6629 -25090 6675 -24890
rect 6939 -25090 6985 -24890
rect 7248 -25090 7294 -24890
rect 8549 -25390 8600 -20554
rect -1363 -25441 8600 -25390
rect 1829 -25483 1984 -25481
rect -7472 -25490 1984 -25483
rect -7596 -25525 1984 -25490
rect 8549 -25512 8600 -25441
rect -7596 -25536 -7460 -25525
rect 1829 -25527 1984 -25525
rect -5116 -25565 -4980 -25563
rect -5116 -25607 2069 -25565
rect -5116 -25609 -4980 -25607
rect 1933 -25611 2069 -25607
rect 8429 -25619 8620 -25512
rect 8770 -23896 8821 -20218
rect 8767 -23991 8826 -23896
rect -7451 -26735 -7405 -26535
rect -7353 -26735 -7307 -26535
rect -7037 -26735 -6991 -26535
rect -6939 -26735 -6893 -26535
rect -6675 -26735 -6629 -26535
rect -6577 -26735 -6531 -26535
rect -6381 -26735 -6335 -26535
rect -6283 -26735 -6237 -26535
rect -6071 -26735 -6025 -26535
rect -5973 -26735 -5927 -26535
rect -5762 -26735 -5716 -26535
rect -5664 -26735 -5618 -26535
rect -6166 -26773 -6035 -26767
rect -7120 -26801 -6035 -26773
rect -7446 -26946 -7307 -26933
rect -7120 -26946 -7092 -26801
rect -6166 -26813 -6035 -26801
rect 8770 -25726 8821 -23991
rect -5411 -25772 8821 -25726
rect -5411 -25777 8397 -25772
rect -7446 -26974 -7092 -26946
rect -6697 -26920 -6558 -26903
rect -5860 -26920 -5724 -26911
rect -6697 -26948 -5724 -26920
rect -6697 -26957 -6558 -26948
rect -5860 -26957 -5724 -26948
rect -7446 -26987 -7307 -26974
rect -6288 -26985 -6149 -26977
rect -5673 -26985 -5534 -26971
rect -5411 -26985 -5383 -25777
rect 8926 -24688 8977 -20068
rect 8920 -24827 8989 -24688
rect -5119 -25998 -5073 -25862
rect -5118 -26568 -5074 -25998
rect -5119 -26704 -5073 -26568
rect -4951 -26735 -4905 -26535
rect -4853 -26735 -4807 -26535
rect -4537 -26735 -4491 -26535
rect -4439 -26735 -4393 -26535
rect -4175 -26735 -4129 -26535
rect -4077 -26735 -4031 -26535
rect -3881 -26735 -3835 -26535
rect -3783 -26735 -3737 -26535
rect -3571 -26735 -3525 -26535
rect -3473 -26735 -3427 -26535
rect -3262 -26735 -3216 -26535
rect -3164 -26735 -3118 -26535
rect -3666 -26773 -3535 -26767
rect -4620 -26801 -3535 -26773
rect -6288 -27013 -5383 -26985
rect -4946 -26946 -4807 -26933
rect -4620 -26946 -4592 -26801
rect -3666 -26813 -3535 -26801
rect 8926 -25876 8977 -24827
rect -2840 -25907 8977 -25876
rect -2840 -25927 8397 -25907
rect 8590 -25914 8977 -25907
rect -4946 -26974 -4592 -26946
rect -4197 -26920 -4058 -26903
rect -3360 -26920 -3224 -26911
rect -4197 -26948 -3224 -26920
rect -4197 -26957 -4058 -26948
rect -3360 -26957 -3224 -26948
rect -4946 -26987 -4807 -26974
rect -3788 -26985 -3649 -26977
rect -3173 -26985 -3034 -26971
rect -2840 -26985 -2812 -25927
rect 9108 -23576 9136 -19932
rect 9088 -23694 9152 -23576
rect -2406 -26283 -2270 -26282
rect -2571 -26327 -2270 -26283
rect -2570 -26564 -2526 -26327
rect -2406 -26328 -2270 -26327
rect -2571 -26700 -2525 -26564
rect -2451 -26735 -2405 -26535
rect -2353 -26735 -2307 -26535
rect -2037 -26735 -1991 -26535
rect -1939 -26735 -1893 -26535
rect -1675 -26735 -1629 -26535
rect -1577 -26735 -1531 -26535
rect -1381 -26735 -1335 -26535
rect -1283 -26735 -1237 -26535
rect -1071 -26735 -1025 -26535
rect -973 -26735 -927 -26535
rect -762 -26735 -716 -26535
rect -664 -26735 -618 -26535
rect -1166 -26773 -1035 -26767
rect -2120 -26801 -1035 -26773
rect -3788 -27013 -2812 -26985
rect -2446 -26946 -2307 -26933
rect -2120 -26946 -2092 -26801
rect -1166 -26813 -1035 -26801
rect 9108 -26012 9136 -23694
rect -368 -26040 9136 -26012
rect -2446 -26974 -2092 -26946
rect -1697 -26920 -1558 -26903
rect -860 -26920 -724 -26911
rect -1697 -26948 -724 -26920
rect -1697 -26957 -1558 -26948
rect -860 -26957 -724 -26948
rect -2446 -26987 -2307 -26974
rect -1288 -26985 -1149 -26977
rect -673 -26985 -534 -26971
rect -368 -26985 -340 -26040
rect 9250 -21339 9288 -19805
rect 9250 -21472 9300 -21339
rect 91 -26270 227 -26269
rect -90 -26314 227 -26270
rect -90 -26564 -46 -26314
rect 91 -26315 227 -26314
rect -91 -26700 -45 -26564
rect 49 -26735 95 -26535
rect 147 -26735 193 -26535
rect 463 -26735 509 -26535
rect 561 -26735 607 -26535
rect 825 -26735 871 -26535
rect 923 -26735 969 -26535
rect 1119 -26735 1165 -26535
rect 1217 -26735 1263 -26535
rect 1429 -26735 1475 -26535
rect 1527 -26735 1573 -26535
rect 1738 -26735 1784 -26535
rect 1836 -26735 1882 -26535
rect 1334 -26773 1465 -26767
rect 380 -26801 1465 -26773
rect -1288 -27013 -340 -26985
rect 54 -26946 193 -26933
rect 380 -26946 408 -26801
rect 1334 -26813 1465 -26801
rect 9250 -26139 9288 -21472
rect 2107 -26149 7805 -26139
rect 8485 -26149 9288 -26139
rect 2107 -26177 9288 -26149
rect 54 -26974 408 -26946
rect 803 -26920 942 -26903
rect 1640 -26920 1776 -26911
rect 803 -26948 1776 -26920
rect 803 -26957 942 -26948
rect 1640 -26957 1776 -26948
rect 54 -26987 193 -26974
rect 1212 -26985 1351 -26977
rect 1827 -26985 1966 -26971
rect 2107 -26985 2135 -26177
rect 2274 -26252 2410 -26206
rect 2327 -26564 2371 -26252
rect 5179 -26268 5315 -26222
rect 2326 -26700 2372 -26564
rect 2549 -26735 2595 -26535
rect 2647 -26735 2693 -26535
rect 2963 -26735 3009 -26535
rect 3061 -26735 3107 -26535
rect 3325 -26735 3371 -26535
rect 3423 -26735 3469 -26535
rect 3619 -26735 3665 -26535
rect 3717 -26735 3763 -26535
rect 3929 -26735 3975 -26535
rect 4027 -26735 4073 -26535
rect 4238 -26735 4284 -26535
rect 4336 -26735 4382 -26535
rect 5232 -26564 5276 -26268
rect 5231 -26700 5277 -26564
rect 3834 -26773 3965 -26767
rect 2880 -26801 3965 -26773
rect 1212 -27013 2135 -26985
rect 2554 -26946 2693 -26933
rect 2880 -26946 2908 -26801
rect 3834 -26813 3965 -26801
rect 9413 -26282 9441 -19662
rect 5412 -26310 9441 -26282
rect 2554 -26974 2908 -26946
rect 3303 -26920 3442 -26903
rect 4140 -26920 4276 -26911
rect 3303 -26948 4276 -26920
rect 3303 -26957 3442 -26948
rect 4140 -26957 4276 -26948
rect 2554 -26987 2693 -26974
rect 3712 -26985 3851 -26977
rect 4327 -26985 4466 -26971
rect 5412 -26985 5440 -26310
rect 5549 -26735 5595 -26535
rect 5647 -26735 5693 -26535
rect 5963 -26735 6009 -26535
rect 6061 -26735 6107 -26535
rect 6325 -26735 6371 -26535
rect 6423 -26735 6469 -26535
rect 6619 -26735 6665 -26535
rect 6717 -26735 6763 -26535
rect 6929 -26735 6975 -26535
rect 7027 -26735 7073 -26535
rect 7238 -26735 7284 -26535
rect 7336 -26735 7382 -26535
rect 6834 -26773 6965 -26767
rect 5880 -26801 6965 -26773
rect 3712 -27013 5440 -26985
rect 5554 -26946 5693 -26933
rect 5880 -26946 5908 -26801
rect 6834 -26813 6965 -26801
rect 5554 -26974 5908 -26946
rect 6303 -26920 6442 -26903
rect 7140 -26920 7276 -26911
rect 6303 -26948 7276 -26920
rect 6303 -26957 6442 -26948
rect 7140 -26957 7276 -26948
rect 5554 -26987 5693 -26974
rect 6712 -26985 6851 -26977
rect 7327 -26985 7466 -26971
rect 9569 -26985 9597 -18959
rect 6712 -27013 9597 -26985
rect -6288 -27031 -6149 -27013
rect -5673 -27025 -5534 -27013
rect -3788 -27031 -3649 -27013
rect -3173 -27025 -3034 -27013
rect -1288 -27031 -1149 -27013
rect -673 -27025 -534 -27013
rect 1212 -27031 1351 -27013
rect 1827 -27025 1966 -27013
rect 3712 -27031 3851 -27013
rect 4327 -27025 4466 -27013
rect 6712 -27031 6851 -27013
rect 7327 -27025 7466 -27013
rect -7451 -27341 -7405 -27141
rect -7353 -27341 -7307 -27141
rect -7255 -27341 -7209 -27141
rect -7135 -27341 -7089 -27141
rect -7037 -27341 -6991 -27141
rect -6939 -27341 -6893 -27141
rect -6577 -27341 -6531 -27141
rect -6381 -27341 -6335 -27141
rect -6071 -27341 -6025 -27141
rect -5762 -27341 -5716 -27141
rect -4951 -27341 -4905 -27141
rect -4853 -27341 -4807 -27141
rect -4755 -27341 -4709 -27141
rect -4635 -27341 -4589 -27141
rect -4537 -27341 -4491 -27141
rect -4439 -27341 -4393 -27141
rect -4077 -27341 -4031 -27141
rect -3881 -27341 -3835 -27141
rect -3571 -27341 -3525 -27141
rect -3262 -27341 -3216 -27141
rect -2451 -27341 -2405 -27141
rect -2353 -27341 -2307 -27141
rect -2255 -27341 -2209 -27141
rect -2135 -27341 -2089 -27141
rect -2037 -27341 -1991 -27141
rect -1939 -27341 -1893 -27141
rect -1577 -27341 -1531 -27141
rect -1381 -27341 -1335 -27141
rect -1071 -27341 -1025 -27141
rect -762 -27341 -716 -27141
rect 49 -27341 95 -27141
rect 147 -27341 193 -27141
rect 245 -27341 291 -27141
rect 365 -27341 411 -27141
rect 463 -27341 509 -27141
rect 561 -27341 607 -27141
rect 923 -27341 969 -27141
rect 1119 -27341 1165 -27141
rect 1429 -27341 1475 -27141
rect 1738 -27341 1784 -27141
rect 2549 -27341 2595 -27141
rect 2647 -27341 2693 -27141
rect 2745 -27341 2791 -27141
rect 2865 -27341 2911 -27141
rect 2963 -27341 3009 -27141
rect 3061 -27341 3107 -27141
rect 3423 -27341 3469 -27141
rect 3619 -27341 3665 -27141
rect 3929 -27341 3975 -27141
rect 4238 -27341 4284 -27141
rect 5549 -27341 5595 -27141
rect 5647 -27341 5693 -27141
rect 5745 -27341 5791 -27141
rect 5865 -27341 5911 -27141
rect 5963 -27341 6009 -27141
rect 6061 -27341 6107 -27141
rect 6423 -27341 6469 -27141
rect 6619 -27341 6665 -27141
rect 6929 -27341 6975 -27141
rect 7238 -27341 7284 -27141
rect 9859 -27404 10154 -20114
rect -8009 -27704 -7846 -27529
rect -24201 -29945 -23988 -29767
rect -7998 -30059 -7866 -27704
rect 8807 -27673 10154 -27404
rect 9859 -29935 10154 -27673
rect 10211 -26585 10411 -20529
rect 12075 -24071 12344 -15445
rect 13067 -16378 78192 -16067
rect 12014 -24412 12400 -24071
rect 13067 -24361 13318 -16378
rect 13654 -16828 68924 -16651
rect 13654 -23111 13985 -16828
rect 14766 -17387 60215 -17166
rect 14766 -21331 14856 -17387
rect 16147 -17944 51026 -17718
rect 15755 -18424 42201 -18159
rect 15473 -18830 33720 -18581
rect 15499 -19510 16064 -19509
rect 15214 -19650 16064 -19510
rect 25899 -19942 32364 -19773
rect 15196 -20071 25429 -20031
rect 15196 -20365 25609 -20071
rect 15196 -20383 25574 -20365
rect 15181 -20572 15448 -20494
rect 15181 -20727 25095 -20572
rect 15181 -20792 15448 -20727
rect 15444 -21236 16271 -21085
rect 17040 -21227 17219 -21151
rect 19577 -21219 19623 -21119
rect 19675 -21219 19721 -21119
rect 19773 -21219 19819 -21119
rect 19871 -21219 19917 -21119
rect 19969 -21219 20015 -21119
rect 20067 -21219 20113 -21119
rect 20165 -21219 20211 -21119
rect 20263 -21219 20309 -21119
rect 17040 -21302 18710 -21227
rect 14762 -21495 14860 -21331
rect 17040 -21340 17219 -21302
rect 13550 -23536 14064 -23111
rect 14766 -23660 14856 -21495
rect 17471 -21538 17517 -21338
rect 17569 -21538 17615 -21338
rect 17667 -21538 17713 -21338
rect 17765 -21538 17811 -21338
rect 18635 -21377 18710 -21302
rect 20482 -21304 20528 -21104
rect 20678 -21304 20724 -21104
rect 20874 -21304 20920 -21104
rect 20137 -21357 20306 -21347
rect 21078 -21357 21135 -21122
rect 21319 -21304 21365 -21104
rect 21515 -21304 21561 -21104
rect 21711 -21304 21757 -21104
rect 22277 -21219 22323 -21119
rect 22375 -21219 22421 -21119
rect 22473 -21219 22519 -21119
rect 22571 -21219 22617 -21119
rect 22669 -21219 22715 -21119
rect 22767 -21219 22813 -21119
rect 22865 -21219 22911 -21119
rect 22963 -21219 23009 -21119
rect 23182 -21304 23228 -21104
rect 23378 -21304 23424 -21104
rect 23574 -21304 23620 -21104
rect 18608 -21512 18740 -21377
rect 19481 -21462 19635 -21402
rect 20137 -21414 21135 -21357
rect 22837 -21357 23006 -21347
rect 23778 -21357 23835 -21122
rect 24019 -21304 24065 -21104
rect 24215 -21304 24261 -21104
rect 24411 -21304 24457 -21104
rect 21934 -21379 21994 -21373
rect 20137 -21421 20306 -21414
rect 21851 -21439 21994 -21379
rect 22188 -21400 22229 -21399
rect 18307 -21576 18349 -21572
rect 18225 -21636 18357 -21576
rect 17471 -22502 17517 -21902
rect 17683 -22502 17729 -21902
rect 17781 -22502 17827 -21902
rect 17879 -22502 17925 -21902
rect 17992 -22502 18038 -21902
rect 18090 -22502 18136 -21902
rect 18188 -22502 18234 -21902
rect 15306 -23439 17416 -23243
rect 17220 -23445 17416 -23439
rect 17220 -23599 17418 -23445
rect 17213 -23641 18250 -23599
rect 14766 -23673 16749 -23660
rect 14766 -23715 18160 -23673
rect 14766 -23750 16749 -23715
rect 17466 -24156 17512 -23956
rect 17564 -24156 17610 -23956
rect 17662 -24156 17708 -23956
rect 17876 -24261 18008 -24201
rect 13051 -24591 13339 -24361
rect 17963 -24374 18005 -24261
rect 18118 -24286 18160 -23715
rect 18208 -24202 18250 -23641
rect 18307 -23670 18349 -21636
rect 18397 -21697 19307 -21640
rect 18397 -23048 18454 -21697
rect 18954 -21813 19086 -21753
rect 18974 -22022 19069 -21813
rect 19250 -21818 19307 -21697
rect 19481 -21737 19527 -21462
rect 19577 -21634 19623 -21534
rect 19675 -21634 19721 -21534
rect 19773 -21634 19819 -21534
rect 19871 -21634 19917 -21534
rect 19969 -21634 20015 -21534
rect 20067 -21634 20113 -21534
rect 20165 -21634 20211 -21534
rect 20263 -21634 20309 -21534
rect 20482 -21584 20528 -21484
rect 20580 -21584 20626 -21484
rect 20678 -21584 20724 -21484
rect 20776 -21584 20822 -21484
rect 20874 -21584 20920 -21484
rect 20972 -21584 21018 -21484
rect 19481 -21782 20300 -21737
rect 19489 -21783 20300 -21782
rect 19250 -21875 19516 -21818
rect 19277 -21983 19409 -21923
rect 18967 -22082 19104 -22022
rect 18694 -22242 18740 -22142
rect 18792 -22242 18838 -22142
rect 18890 -22242 18936 -22142
rect 18988 -22242 19034 -22142
rect 19086 -22242 19132 -22142
rect 19184 -22242 19230 -22142
rect 19318 -22211 19376 -21983
rect 19318 -22343 19378 -22211
rect 19459 -22312 19516 -21875
rect 20254 -21949 20300 -21783
rect 21124 -21837 21184 -21473
rect 21319 -21584 21365 -21484
rect 21417 -21584 21463 -21484
rect 21515 -21584 21561 -21484
rect 21613 -21584 21659 -21484
rect 21711 -21584 21757 -21484
rect 21809 -21584 21855 -21484
rect 21587 -21813 21724 -21753
rect 21081 -21897 21213 -21837
rect 20254 -21995 21014 -21949
rect 20386 -22092 20428 -21995
rect 20582 -22092 20624 -21995
rect 20777 -22092 20819 -21995
rect 20968 -22092 21014 -21995
rect 21618 -22021 21713 -21813
rect 21594 -22081 21731 -22021
rect 19576 -22242 19622 -22142
rect 19674 -22242 19720 -22142
rect 19772 -22242 19818 -22142
rect 19870 -22242 19916 -22142
rect 19968 -22242 20014 -22142
rect 20066 -22242 20112 -22142
rect 20285 -22192 20331 -22092
rect 20383 -22192 20429 -22092
rect 20481 -22192 20527 -22092
rect 20579 -22192 20625 -22092
rect 20677 -22192 20723 -22092
rect 20775 -22192 20821 -22092
rect 20873 -22192 20919 -22092
rect 20968 -22192 21017 -22092
rect 21319 -22242 21365 -22142
rect 21417 -22242 21463 -22142
rect 21515 -22242 21561 -22142
rect 21613 -22242 21659 -22142
rect 21711 -22242 21757 -22142
rect 21809 -22242 21855 -22142
rect 21934 -22187 21994 -21439
rect 22187 -21460 22324 -21400
rect 22837 -21414 23835 -21357
rect 22837 -21421 23006 -21414
rect 22022 -21896 22159 -21836
rect 21934 -22232 21995 -22187
rect 20288 -22312 20457 -22305
rect 19459 -22369 20457 -22312
rect 21935 -22319 21995 -22232
rect 22050 -22344 22110 -21896
rect 22188 -21945 22229 -21460
rect 22277 -21634 22323 -21534
rect 22375 -21634 22421 -21534
rect 22473 -21634 22519 -21534
rect 22571 -21634 22617 -21534
rect 22669 -21634 22715 -21534
rect 22767 -21634 22813 -21534
rect 22865 -21634 22911 -21534
rect 22963 -21634 23009 -21534
rect 23182 -21584 23228 -21484
rect 23280 -21584 23326 -21484
rect 23378 -21584 23424 -21484
rect 23476 -21584 23522 -21484
rect 23574 -21584 23620 -21484
rect 23672 -21584 23718 -21484
rect 23836 -21925 23896 -21458
rect 24019 -21584 24065 -21484
rect 24117 -21584 24163 -21484
rect 24215 -21584 24261 -21484
rect 24313 -21584 24359 -21484
rect 24411 -21584 24457 -21484
rect 24509 -21584 24555 -21484
rect 24184 -21807 24321 -21747
rect 22188 -21993 23719 -21945
rect 23800 -21985 23932 -21925
rect 22276 -22242 22322 -22142
rect 22374 -22242 22420 -22142
rect 22472 -22242 22518 -22142
rect 22570 -22242 22616 -22142
rect 22668 -22242 22714 -22142
rect 22766 -22242 22812 -22142
rect 22985 -22192 23031 -22092
rect 23079 -22111 23140 -21993
rect 23083 -22192 23129 -22111
rect 23181 -22192 23227 -22092
rect 23270 -22113 23331 -21993
rect 23279 -22192 23325 -22113
rect 23377 -22192 23423 -22092
rect 23466 -22111 23527 -21993
rect 23475 -22192 23521 -22111
rect 23573 -22192 23619 -22092
rect 23671 -22147 23719 -21993
rect 24211 -22025 24306 -21807
rect 24609 -21865 24669 -21818
rect 24609 -21929 24878 -21865
rect 24609 -21955 24755 -21929
rect 24198 -22085 24330 -22025
rect 23671 -22192 23717 -22147
rect 24019 -22242 24065 -22142
rect 24117 -22242 24163 -22142
rect 24215 -22242 24261 -22142
rect 24313 -22242 24359 -22142
rect 24411 -22242 24457 -22142
rect 24509 -22242 24555 -22142
rect 22988 -22312 23157 -22305
rect 18792 -22622 18838 -22422
rect 18988 -22622 19034 -22422
rect 19184 -22622 19230 -22422
rect 19459 -22604 19516 -22369
rect 20288 -22379 20457 -22369
rect 22159 -22369 23157 -22312
rect 19674 -22622 19720 -22422
rect 19870 -22622 19916 -22422
rect 20066 -22622 20112 -22422
rect 20285 -22607 20331 -22507
rect 20383 -22607 20429 -22507
rect 20481 -22607 20527 -22507
rect 20579 -22607 20625 -22507
rect 20677 -22607 20723 -22507
rect 20775 -22607 20821 -22507
rect 20873 -22607 20919 -22507
rect 20971 -22607 21017 -22507
rect 21417 -22622 21463 -22422
rect 21613 -22622 21659 -22422
rect 21809 -22622 21855 -22422
rect 22159 -22604 22216 -22369
rect 22988 -22379 23157 -22369
rect 22374 -22622 22420 -22422
rect 22570 -22622 22616 -22422
rect 22766 -22622 22812 -22422
rect 22985 -22607 23031 -22507
rect 23083 -22607 23129 -22507
rect 23181 -22607 23227 -22507
rect 23279 -22607 23325 -22507
rect 23377 -22607 23423 -22507
rect 23475 -22607 23521 -22507
rect 23573 -22607 23619 -22507
rect 23671 -22607 23717 -22507
rect 24117 -22622 24163 -22422
rect 24313 -22622 24359 -22422
rect 24509 -22622 24555 -22422
rect 24665 -22799 24755 -21955
rect 20723 -22889 24755 -22799
rect 20723 -22980 20883 -22889
rect 18397 -23105 21669 -23048
rect 20720 -23295 20880 -23163
rect 18307 -23712 19077 -23670
rect 20617 -23678 20749 -23618
rect 18412 -24156 18458 -23956
rect 18510 -24156 18556 -23956
rect 18608 -24156 18654 -23956
rect 18324 -24202 18456 -24195
rect 18208 -24244 18456 -24202
rect 18324 -24255 18456 -24244
rect 18547 -24286 18679 -24275
rect 18118 -24328 18679 -24286
rect 18547 -24335 18679 -24328
rect 18912 -24374 18972 -24344
rect 17963 -24416 18972 -24374
rect 17466 -24848 17512 -24448
rect 17677 -24848 17723 -24448
rect 17775 -24848 17821 -24448
rect 17873 -24848 17919 -24448
rect 18412 -24848 18458 -24448
rect 18623 -24848 18669 -24448
rect 18721 -24848 18767 -24448
rect 18819 -24848 18865 -24448
rect 18912 -24476 18972 -24416
rect 19035 -24594 19077 -23712
rect 19230 -24275 19276 -23975
rect 19328 -24275 19374 -23975
rect 19426 -24275 19472 -23975
rect 19540 -24274 19586 -23974
rect 19638 -24274 19684 -23974
rect 19736 -24274 19782 -23974
rect 19849 -24274 19895 -23974
rect 19947 -24274 19993 -23974
rect 20045 -24274 20091 -23974
rect 20360 -24174 20406 -23974
rect 20458 -24174 20504 -23974
rect 20649 -24363 20709 -23678
rect 20788 -23719 20848 -23295
rect 21237 -23574 21283 -23174
rect 21433 -23574 21479 -23174
rect 21612 -23627 21669 -23105
rect 24940 -23116 25095 -20727
rect 21808 -23186 25095 -23116
rect 21808 -23365 21878 -23186
rect 20788 -23720 21129 -23719
rect 20788 -23778 21130 -23720
rect 21583 -23761 21669 -23627
rect 20788 -23779 21129 -23778
rect 20610 -24423 20741 -24363
rect 20788 -24533 20848 -23779
rect 21139 -24028 21185 -23828
rect 21237 -24028 21283 -23828
rect 21349 -24028 21395 -23828
rect 21447 -24028 21493 -23828
rect 21969 -23919 22015 -23219
rect 22067 -23919 22113 -23219
rect 22369 -23919 22415 -23219
rect 22467 -23919 22513 -23219
rect 22852 -23916 22922 -23186
rect 22969 -23919 23015 -23219
rect 23067 -23919 23113 -23219
rect 23369 -23919 23415 -23219
rect 23467 -23919 23513 -23219
rect 23843 -23917 23913 -23186
rect 23969 -23919 24015 -23219
rect 24067 -23919 24113 -23219
rect 24369 -23919 24415 -23219
rect 24467 -23919 24513 -23219
rect 22581 -23969 22699 -23957
rect 22581 -24003 22788 -23969
rect 24554 -23976 24672 -23972
rect 25105 -23976 25226 -23953
rect 22581 -24015 22699 -24003
rect 21089 -24495 21135 -24395
rect 21187 -24495 21233 -24395
rect 21285 -24495 21331 -24395
rect 21383 -24495 21429 -24395
rect 21481 -24495 21527 -24395
rect 21579 -24495 21625 -24395
rect 20788 -24593 21115 -24533
rect 19027 -24726 19087 -24594
rect 19328 -24882 19374 -24682
rect 19524 -24882 19570 -24682
rect 19720 -24882 19766 -24682
rect 20458 -24882 20504 -24682
rect 21187 -24875 21233 -24675
rect 21383 -24875 21429 -24675
rect 21579 -24875 21625 -24675
rect 22067 -24804 22113 -24104
rect 22467 -24804 22513 -24104
rect 22754 -24904 22788 -24003
rect 23658 -24042 23776 -23984
rect 24554 -24021 25226 -23976
rect 24554 -24030 24672 -24021
rect 23067 -24804 23113 -24104
rect 23467 -24804 23513 -24104
rect 23664 -24839 23698 -24042
rect 24067 -24804 24113 -24104
rect 24467 -24804 24513 -24104
rect 23664 -24873 24972 -24839
rect 22754 -24938 24884 -24904
rect 10664 -25860 10710 -25660
rect 10860 -25860 10906 -25660
rect 11056 -25860 11102 -25660
rect 11331 -25913 11388 -25678
rect 11546 -25860 11592 -25660
rect 11742 -25860 11788 -25660
rect 11938 -25860 11984 -25660
rect 12157 -25775 12203 -25675
rect 12255 -25775 12301 -25675
rect 12353 -25775 12399 -25675
rect 12451 -25775 12497 -25675
rect 12549 -25775 12595 -25675
rect 12647 -25775 12693 -25675
rect 12745 -25775 12791 -25675
rect 12843 -25775 12889 -25675
rect 13289 -25860 13335 -25660
rect 13485 -25860 13531 -25660
rect 13681 -25860 13727 -25660
rect 12160 -25913 12329 -25903
rect 10566 -26140 10612 -26040
rect 10664 -26140 10710 -26040
rect 10762 -26140 10808 -26040
rect 10860 -26140 10906 -26040
rect 10958 -26140 11004 -26040
rect 11056 -26140 11102 -26040
rect 11190 -26071 11250 -25939
rect 11331 -25970 12329 -25913
rect 14031 -25913 14088 -25678
rect 14246 -25860 14292 -25660
rect 14442 -25860 14488 -25660
rect 14638 -25860 14684 -25660
rect 14857 -25775 14903 -25675
rect 14955 -25775 15001 -25675
rect 15053 -25775 15099 -25675
rect 15151 -25775 15197 -25675
rect 15249 -25775 15295 -25675
rect 15347 -25775 15393 -25675
rect 15445 -25775 15491 -25675
rect 15543 -25775 15589 -25675
rect 15989 -25860 16035 -25660
rect 16185 -25860 16231 -25660
rect 16381 -25860 16427 -25660
rect 14860 -25913 15029 -25903
rect 10839 -26260 10976 -26200
rect 10846 -26469 10941 -26260
rect 11190 -26299 11248 -26071
rect 11149 -26359 11281 -26299
rect 11331 -26407 11388 -25970
rect 12160 -25977 12329 -25970
rect 11448 -26140 11494 -26040
rect 11546 -26140 11592 -26040
rect 11644 -26140 11690 -26040
rect 11742 -26140 11788 -26040
rect 11840 -26140 11886 -26040
rect 11938 -26140 11984 -26040
rect 12157 -26190 12203 -26090
rect 12255 -26190 12301 -26090
rect 12353 -26190 12399 -26090
rect 12451 -26190 12497 -26090
rect 12549 -26190 12595 -26090
rect 12647 -26190 12693 -26090
rect 12745 -26190 12791 -26090
rect 12840 -26190 12889 -26090
rect 13191 -26140 13237 -26040
rect 13289 -26140 13335 -26040
rect 13387 -26140 13433 -26040
rect 13485 -26140 13531 -26040
rect 13583 -26140 13629 -26040
rect 13681 -26140 13727 -26040
rect 13807 -26050 13867 -25963
rect 13806 -26095 13867 -26050
rect 12258 -26287 12300 -26190
rect 12454 -26287 12496 -26190
rect 12649 -26287 12691 -26190
rect 12840 -26287 12886 -26190
rect 13466 -26261 13603 -26201
rect 11122 -26464 11388 -26407
rect 12126 -26333 12886 -26287
rect 10826 -26529 10958 -26469
rect 11122 -26585 11179 -26464
rect 12126 -26499 12172 -26333
rect 12953 -26445 13085 -26385
rect 11361 -26500 12172 -26499
rect 10211 -26642 11179 -26585
rect 11353 -26545 12172 -26500
rect -7998 -30195 -7862 -30059
rect 10211 -30432 10411 -26642
rect 11353 -26820 11399 -26545
rect 11449 -26748 11495 -26648
rect 11547 -26748 11593 -26648
rect 11645 -26748 11691 -26648
rect 11743 -26748 11789 -26648
rect 11841 -26748 11887 -26648
rect 11939 -26748 11985 -26648
rect 12037 -26748 12083 -26648
rect 12135 -26748 12181 -26648
rect 12354 -26798 12400 -26698
rect 12452 -26798 12498 -26698
rect 12550 -26798 12596 -26698
rect 12648 -26798 12694 -26698
rect 12746 -26798 12792 -26698
rect 12844 -26798 12890 -26698
rect 12996 -26809 13056 -26445
rect 13490 -26469 13585 -26261
rect 13459 -26529 13596 -26469
rect 13191 -26798 13237 -26698
rect 13289 -26798 13335 -26698
rect 13387 -26798 13433 -26698
rect 13485 -26798 13531 -26698
rect 13583 -26798 13629 -26698
rect 13681 -26798 13727 -26698
rect 11353 -26880 11507 -26820
rect 13806 -26843 13866 -26095
rect 13922 -26386 13982 -25938
rect 14031 -25970 15029 -25913
rect 14860 -25977 15029 -25970
rect 14148 -26140 14194 -26040
rect 14246 -26140 14292 -26040
rect 14344 -26140 14390 -26040
rect 14442 -26140 14488 -26040
rect 14540 -26140 14586 -26040
rect 14638 -26140 14684 -26040
rect 14857 -26190 14903 -26090
rect 14955 -26171 15001 -26090
rect 14951 -26289 15012 -26171
rect 15053 -26190 15099 -26090
rect 15151 -26169 15197 -26090
rect 15142 -26289 15203 -26169
rect 15249 -26190 15295 -26090
rect 15347 -26171 15393 -26090
rect 15338 -26289 15399 -26171
rect 15445 -26190 15491 -26090
rect 15543 -26135 15589 -26090
rect 15543 -26289 15591 -26135
rect 15891 -26140 15937 -26040
rect 15989 -26140 16035 -26040
rect 16087 -26140 16133 -26040
rect 16185 -26140 16231 -26040
rect 16283 -26140 16329 -26040
rect 16381 -26140 16427 -26040
rect 16070 -26257 16202 -26197
rect 14060 -26337 15591 -26289
rect 13894 -26446 14031 -26386
rect 14060 -26822 14101 -26337
rect 15672 -26357 15804 -26297
rect 14149 -26748 14195 -26648
rect 14247 -26748 14293 -26648
rect 14345 -26748 14391 -26648
rect 14443 -26748 14489 -26648
rect 14541 -26748 14587 -26648
rect 14639 -26748 14685 -26648
rect 14737 -26748 14783 -26648
rect 14835 -26748 14881 -26648
rect 15054 -26798 15100 -26698
rect 15152 -26798 15198 -26698
rect 15250 -26798 15296 -26698
rect 15348 -26798 15394 -26698
rect 15446 -26798 15492 -26698
rect 15544 -26798 15590 -26698
rect 12009 -26868 12178 -26861
rect 12009 -26925 13007 -26868
rect 13723 -26903 13866 -26843
rect 14059 -26882 14196 -26822
rect 15708 -26824 15768 -26357
rect 16083 -26475 16178 -26257
rect 16481 -26353 16541 -26327
rect 16481 -26417 16937 -26353
rect 16481 -26464 16541 -26417
rect 16056 -26535 16193 -26475
rect 15891 -26798 15937 -26698
rect 15989 -26798 16035 -26698
rect 16087 -26798 16133 -26698
rect 16185 -26798 16231 -26698
rect 16283 -26798 16329 -26698
rect 16381 -26798 16427 -26698
rect 14709 -26868 14878 -26861
rect 14060 -26883 14101 -26882
rect 13806 -26909 13866 -26903
rect 12009 -26935 12178 -26925
rect 11449 -27163 11495 -27063
rect 11547 -27163 11593 -27063
rect 11645 -27163 11691 -27063
rect 11743 -27163 11789 -27063
rect 11841 -27163 11887 -27063
rect 11939 -27163 11985 -27063
rect 12037 -27163 12083 -27063
rect 12135 -27163 12181 -27063
rect 12354 -27178 12400 -26978
rect 12550 -27178 12596 -26978
rect 12746 -27178 12792 -26978
rect 12950 -27160 13007 -26925
rect 14709 -26925 15707 -26868
rect 14709 -26935 14878 -26925
rect 13191 -27178 13237 -26978
rect 13387 -27178 13433 -26978
rect 13583 -27178 13629 -26978
rect 14149 -27163 14195 -27063
rect 14247 -27163 14293 -27063
rect 14345 -27163 14391 -27063
rect 14443 -27163 14489 -27063
rect 14541 -27163 14587 -27063
rect 14639 -27163 14685 -27063
rect 14737 -27163 14783 -27063
rect 14835 -27163 14881 -27063
rect 15054 -27178 15100 -26978
rect 15250 -27178 15296 -26978
rect 15446 -27178 15492 -26978
rect 15650 -27160 15707 -26925
rect 15891 -27178 15937 -26978
rect 16087 -27178 16133 -26978
rect 16283 -27178 16329 -26978
rect 16809 -30059 16937 -26417
rect 24311 -27109 24381 -24938
rect 24938 -25001 24972 -24873
rect 24192 -27329 24563 -27109
rect 24877 -27658 24998 -25001
rect 16804 -30195 16937 -30059
rect 23597 -27779 24998 -27658
rect 23597 -30622 23718 -27779
rect 25105 -30020 25226 -24021
rect 25329 -27482 25574 -20383
rect 25899 -23590 26068 -19942
rect 26197 -20223 26410 -20184
rect 27924 -20207 28363 -20160
rect 26197 -20277 27635 -20223
rect 27924 -20244 27971 -20207
rect 26197 -20317 26410 -20277
rect 26764 -20717 26894 -20567
rect 27050 -20621 27096 -20421
rect 27148 -20649 27194 -20421
rect 27246 -20621 27292 -20421
rect 27344 -20649 27390 -20421
rect 27581 -20567 27635 -20277
rect 27925 -20543 27971 -20244
rect 28023 -20543 28069 -20243
rect 28121 -20543 28167 -20207
rect 27581 -20621 27909 -20567
rect 27050 -20695 27687 -20649
rect 27855 -20676 27909 -20621
rect 26198 -22144 26457 -21881
rect 26814 -22121 26868 -20717
rect 27050 -20951 27096 -20695
rect 27148 -20697 27390 -20695
rect 27246 -20951 27292 -20697
rect 27442 -20951 27488 -20695
rect 27829 -20734 27988 -20676
rect 28023 -21080 28069 -20780
rect 28219 -21080 28265 -20243
rect 28317 -20543 28363 -20207
rect 29019 -20715 29727 -20602
rect 28632 -20850 28678 -20750
rect 28730 -20879 28776 -20750
rect 28828 -20850 28874 -20750
rect 28926 -20879 28972 -20750
rect 28632 -20925 29269 -20879
rect 28632 -21081 28678 -20925
rect 28730 -20927 28972 -20925
rect 28828 -21081 28874 -20927
rect 29024 -21081 29070 -20925
rect 27024 -21980 27070 -21680
rect 26671 -22175 26868 -22121
rect 26926 -22516 26972 -22217
rect 26925 -22553 26972 -22516
rect 27024 -22517 27070 -22217
rect 27122 -22553 27168 -22217
rect 27220 -22517 27266 -21680
rect 27633 -21835 27679 -21679
rect 27829 -21833 27875 -21679
rect 27731 -21835 27973 -21833
rect 28025 -21835 28071 -21679
rect 27633 -21881 28270 -21835
rect 27633 -22010 27679 -21910
rect 27731 -22010 27777 -21881
rect 27829 -22010 27875 -21910
rect 27927 -22010 27973 -21881
rect 28471 -22191 28517 -21591
rect 28682 -22191 28728 -21591
rect 28780 -22191 28826 -21591
rect 28878 -22191 28924 -21591
rect 29090 -22191 29136 -21591
rect 27318 -22553 27364 -22217
rect 29321 -22322 29426 -22250
rect 29327 -22405 29392 -22322
rect 28372 -22470 29392 -22405
rect 26925 -22600 27364 -22553
rect 28471 -22803 28517 -22503
rect 28569 -22803 28615 -22503
rect 28667 -22803 28713 -22503
rect 28909 -22803 28955 -22503
rect 29007 -22803 29053 -22503
rect 29240 -22911 29353 -22910
rect 29614 -22911 29727 -20715
rect 30463 -21949 30509 -21449
rect 30732 -21949 30778 -21449
rect 30830 -21949 30876 -21449
rect 30928 -21949 30974 -21449
rect 31058 -21949 31104 -21449
rect 31384 -21949 31430 -21449
rect 31612 -21749 31658 -21449
rect 30232 -22109 30370 -22105
rect 31038 -22109 31176 -22105
rect 31423 -22109 31477 -22036
rect 30232 -22153 31477 -22109
rect 30232 -22159 30370 -22153
rect 31038 -22159 31176 -22153
rect 31423 -22174 31477 -22153
rect 31595 -22189 31661 -22177
rect 32195 -22189 32364 -19942
rect 33471 -20064 33720 -18830
rect 33882 -19890 40964 -19699
rect 33380 -20200 33737 -20064
rect 33380 -20254 33743 -20200
rect 33380 -20331 33737 -20254
rect 30071 -22496 30174 -22405
rect 29050 -23024 29727 -22911
rect 25899 -23676 26249 -23590
rect 27916 -23660 28355 -23613
rect 25899 -23730 27627 -23676
rect 27916 -23697 27963 -23660
rect 25899 -23759 26249 -23730
rect 26756 -24170 26886 -24020
rect 27042 -24074 27088 -23874
rect 27140 -24102 27186 -23874
rect 27238 -24074 27284 -23874
rect 27336 -24102 27382 -23874
rect 27573 -24020 27627 -23730
rect 27917 -23996 27963 -23697
rect 28015 -23996 28061 -23696
rect 28113 -23996 28159 -23660
rect 27573 -24074 27901 -24020
rect 27042 -24148 27679 -24102
rect 27847 -24129 27901 -24074
rect 26806 -25574 26860 -24170
rect 27042 -24404 27088 -24148
rect 27140 -24150 27382 -24148
rect 27238 -24404 27284 -24150
rect 27434 -24404 27480 -24148
rect 27821 -24187 27980 -24129
rect 28015 -24533 28061 -24233
rect 28211 -24533 28257 -23696
rect 28309 -23996 28355 -23660
rect 29240 -24055 29353 -23024
rect 30083 -23129 30162 -22496
rect 30365 -22745 30411 -22445
rect 30463 -22745 30509 -22445
rect 30835 -22745 30881 -22245
rect 30933 -22745 30979 -22245
rect 31058 -22745 31104 -22245
rect 31156 -22745 31202 -22245
rect 31286 -22745 31332 -22245
rect 31384 -22745 31430 -22245
rect 31482 -22745 31528 -22245
rect 31595 -22251 33217 -22189
rect 31595 -22260 31661 -22251
rect 31612 -22745 31658 -22445
rect 31710 -22745 31756 -22445
rect 29583 -23208 30162 -23129
rect 29583 -23563 29662 -23208
rect 29557 -23660 29673 -23563
rect 31584 -23691 32023 -23644
rect 30186 -23707 30283 -23701
rect 30186 -23761 31295 -23707
rect 31584 -23728 31631 -23691
rect 30186 -23767 30283 -23761
rect 29011 -24168 29719 -24055
rect 28624 -24303 28670 -24203
rect 28722 -24332 28768 -24203
rect 28820 -24303 28866 -24203
rect 28918 -24332 28964 -24203
rect 28624 -24378 29261 -24332
rect 28624 -24534 28670 -24378
rect 28722 -24380 28964 -24378
rect 28820 -24534 28866 -24380
rect 29016 -24534 29062 -24378
rect 27016 -25433 27062 -25133
rect 26663 -25628 26860 -25574
rect 26918 -25969 26964 -25670
rect 26917 -26006 26964 -25969
rect 27016 -25970 27062 -25670
rect 27114 -26006 27160 -25670
rect 27212 -25970 27258 -25133
rect 27625 -25288 27671 -25132
rect 27821 -25286 27867 -25132
rect 27723 -25288 27965 -25286
rect 28017 -25288 28063 -25132
rect 27625 -25334 28262 -25288
rect 27625 -25463 27671 -25363
rect 27723 -25463 27769 -25334
rect 27821 -25463 27867 -25363
rect 27919 -25463 27965 -25334
rect 28463 -25644 28509 -25044
rect 28674 -25644 28720 -25044
rect 28772 -25644 28818 -25044
rect 28870 -25644 28916 -25044
rect 29082 -25644 29128 -25044
rect 27310 -26006 27356 -25670
rect 29313 -25775 29418 -25703
rect 29319 -25858 29384 -25775
rect 28364 -25923 29384 -25858
rect 26917 -26053 27356 -26006
rect 28463 -26256 28509 -25956
rect 28561 -26256 28607 -25956
rect 28659 -26256 28705 -25956
rect 28901 -26256 28947 -25956
rect 28999 -26256 29045 -25956
rect 29606 -26364 29719 -24168
rect 30424 -24201 30554 -24051
rect 30710 -24105 30756 -23905
rect 30808 -24133 30854 -23905
rect 30906 -24105 30952 -23905
rect 31004 -24133 31050 -23905
rect 31241 -24051 31295 -23761
rect 31585 -24027 31631 -23728
rect 31683 -24027 31729 -23727
rect 31781 -24027 31827 -23691
rect 31241 -24105 31569 -24051
rect 30710 -24179 31347 -24133
rect 31515 -24160 31569 -24105
rect 30474 -25605 30528 -24201
rect 30710 -24435 30756 -24179
rect 30808 -24181 31050 -24179
rect 30906 -24435 30952 -24181
rect 31102 -24435 31148 -24179
rect 31489 -24218 31648 -24160
rect 31683 -24564 31729 -24264
rect 31879 -24564 31925 -23727
rect 31977 -24027 32023 -23691
rect 32679 -24199 33387 -24086
rect 32292 -24334 32338 -24234
rect 32390 -24363 32436 -24234
rect 32488 -24334 32534 -24234
rect 32586 -24363 32632 -24234
rect 32292 -24409 32929 -24363
rect 32292 -24565 32338 -24409
rect 32390 -24411 32632 -24409
rect 32488 -24565 32534 -24411
rect 32684 -24565 32730 -24409
rect 30684 -25464 30730 -25164
rect 30331 -25659 30528 -25605
rect 30586 -26000 30632 -25701
rect 30585 -26037 30632 -26000
rect 30684 -26001 30730 -25701
rect 30782 -26037 30828 -25701
rect 30880 -26001 30926 -25164
rect 31293 -25319 31339 -25163
rect 31489 -25317 31535 -25163
rect 31391 -25319 31633 -25317
rect 31685 -25319 31731 -25163
rect 31293 -25365 31930 -25319
rect 31293 -25494 31339 -25394
rect 31391 -25494 31437 -25365
rect 31489 -25494 31535 -25394
rect 31587 -25494 31633 -25365
rect 32131 -25675 32177 -25075
rect 32342 -25675 32388 -25075
rect 32440 -25675 32486 -25075
rect 32538 -25675 32584 -25075
rect 32750 -25675 32796 -25075
rect 30978 -26037 31024 -25701
rect 32981 -25806 33086 -25734
rect 32987 -25889 33052 -25806
rect 32032 -25954 33052 -25889
rect 30585 -26084 31024 -26037
rect 32131 -26287 32177 -25987
rect 32229 -26287 32275 -25987
rect 32327 -26287 32373 -25987
rect 32569 -26287 32615 -25987
rect 32667 -26287 32713 -25987
rect 29042 -26395 29719 -26364
rect 33274 -26395 33387 -24199
rect 33471 -25820 33720 -20331
rect 33882 -23604 34073 -19890
rect 34558 -20234 34915 -20098
rect 36364 -20218 36803 -20171
rect 34558 -20288 36075 -20234
rect 36364 -20255 36411 -20218
rect 34558 -20365 34915 -20288
rect 35204 -20728 35334 -20578
rect 35490 -20632 35536 -20432
rect 35588 -20660 35634 -20432
rect 35686 -20632 35732 -20432
rect 35784 -20660 35830 -20432
rect 36021 -20578 36075 -20288
rect 36365 -20554 36411 -20255
rect 36463 -20554 36509 -20254
rect 36561 -20554 36607 -20218
rect 36021 -20632 36349 -20578
rect 35490 -20706 36127 -20660
rect 36295 -20687 36349 -20632
rect 35254 -22132 35308 -20728
rect 35490 -20962 35536 -20706
rect 35588 -20708 35830 -20706
rect 35686 -20962 35732 -20708
rect 35882 -20962 35928 -20706
rect 36269 -20745 36428 -20687
rect 36463 -21091 36509 -20791
rect 36659 -21091 36705 -20254
rect 36757 -20554 36803 -20218
rect 37459 -20726 38167 -20613
rect 37072 -20861 37118 -20761
rect 37170 -20890 37216 -20761
rect 37268 -20861 37314 -20761
rect 37366 -20890 37412 -20761
rect 37072 -20936 37709 -20890
rect 37072 -21092 37118 -20936
rect 37170 -20938 37412 -20936
rect 37268 -21092 37314 -20938
rect 37464 -21092 37510 -20936
rect 35464 -21991 35510 -21691
rect 35111 -22186 35308 -22132
rect 35366 -22527 35412 -22228
rect 35365 -22564 35412 -22527
rect 35464 -22528 35510 -22228
rect 35562 -22564 35608 -22228
rect 35660 -22528 35706 -21691
rect 36073 -21846 36119 -21690
rect 36269 -21844 36315 -21690
rect 36171 -21846 36413 -21844
rect 36465 -21846 36511 -21690
rect 36073 -21892 36710 -21846
rect 36073 -22021 36119 -21921
rect 36171 -22021 36217 -21892
rect 36269 -22021 36315 -21921
rect 36367 -22021 36413 -21892
rect 36911 -22202 36957 -21602
rect 37122 -22202 37168 -21602
rect 37220 -22202 37266 -21602
rect 37318 -22202 37364 -21602
rect 37530 -22202 37576 -21602
rect 35758 -22564 35804 -22228
rect 37761 -22333 37866 -22261
rect 37767 -22416 37832 -22333
rect 36812 -22481 37832 -22416
rect 35365 -22611 35804 -22564
rect 36911 -22814 36957 -22514
rect 37009 -22814 37055 -22514
rect 37107 -22814 37153 -22514
rect 37349 -22814 37395 -22514
rect 37447 -22814 37493 -22514
rect 37680 -22922 37793 -22921
rect 38054 -22922 38167 -20726
rect 38903 -21960 38949 -21460
rect 39172 -21960 39218 -21460
rect 39270 -21960 39316 -21460
rect 39368 -21960 39414 -21460
rect 39498 -21960 39544 -21460
rect 39824 -21960 39870 -21460
rect 40052 -21760 40098 -21460
rect 38672 -22120 38810 -22116
rect 39478 -22120 39616 -22116
rect 39863 -22120 39917 -22047
rect 38672 -22164 39917 -22120
rect 38672 -22170 38810 -22164
rect 39478 -22170 39616 -22164
rect 39863 -22185 39917 -22164
rect 40035 -22200 40101 -22188
rect 40748 -22200 40964 -19890
rect 38511 -22507 38614 -22416
rect 37490 -23035 38167 -22922
rect 33882 -23687 34732 -23604
rect 36356 -23671 36795 -23624
rect 33882 -23741 36067 -23687
rect 36356 -23708 36403 -23671
rect 33882 -23795 34732 -23741
rect 35196 -24181 35326 -24031
rect 35482 -24085 35528 -23885
rect 35580 -24113 35626 -23885
rect 35678 -24085 35724 -23885
rect 35776 -24113 35822 -23885
rect 36013 -24031 36067 -23741
rect 36357 -24007 36403 -23708
rect 36455 -24007 36501 -23707
rect 36553 -24007 36599 -23671
rect 36013 -24085 36341 -24031
rect 35482 -24159 36119 -24113
rect 36287 -24140 36341 -24085
rect 35246 -25585 35300 -24181
rect 35482 -24415 35528 -24159
rect 35580 -24161 35822 -24159
rect 35678 -24415 35724 -24161
rect 35874 -24415 35920 -24159
rect 36261 -24198 36420 -24140
rect 36455 -24544 36501 -24244
rect 36651 -24544 36697 -23707
rect 36749 -24007 36795 -23671
rect 37680 -24066 37793 -23035
rect 38523 -23140 38602 -22507
rect 38805 -22756 38851 -22456
rect 38903 -22756 38949 -22456
rect 39275 -22756 39321 -22256
rect 39373 -22756 39419 -22256
rect 39498 -22756 39544 -22256
rect 39596 -22756 39642 -22256
rect 39726 -22756 39772 -22256
rect 39824 -22756 39870 -22256
rect 39922 -22756 39968 -22256
rect 40035 -22262 41657 -22200
rect 40035 -22271 40101 -22262
rect 40052 -22756 40098 -22456
rect 40150 -22756 40196 -22456
rect 38023 -23219 38602 -23140
rect 38023 -23574 38102 -23219
rect 37997 -23671 38113 -23574
rect 40024 -23702 40463 -23655
rect 38626 -23718 38723 -23712
rect 38626 -23772 39735 -23718
rect 40024 -23739 40071 -23702
rect 38626 -23778 38723 -23772
rect 37451 -24179 38159 -24066
rect 37064 -24314 37110 -24214
rect 37162 -24343 37208 -24214
rect 37260 -24314 37306 -24214
rect 37358 -24343 37404 -24214
rect 37064 -24389 37701 -24343
rect 37064 -24545 37110 -24389
rect 37162 -24391 37404 -24389
rect 37260 -24545 37306 -24391
rect 37456 -24545 37502 -24389
rect 35456 -25444 35502 -25144
rect 35103 -25639 35300 -25585
rect 33487 -25989 33710 -25820
rect 35358 -25980 35404 -25681
rect 35357 -26017 35404 -25980
rect 35456 -25981 35502 -25681
rect 35554 -26017 35600 -25681
rect 35652 -25981 35698 -25144
rect 36065 -25299 36111 -25143
rect 36261 -25297 36307 -25143
rect 36163 -25299 36405 -25297
rect 36457 -25299 36503 -25143
rect 36065 -25345 36702 -25299
rect 36065 -25474 36111 -25374
rect 36163 -25474 36209 -25345
rect 36261 -25474 36307 -25374
rect 36359 -25474 36405 -25345
rect 36903 -25655 36949 -25055
rect 37114 -25655 37160 -25055
rect 37212 -25655 37258 -25055
rect 37310 -25655 37356 -25055
rect 37522 -25655 37568 -25055
rect 35750 -26017 35796 -25681
rect 37753 -25786 37858 -25714
rect 37759 -25869 37824 -25786
rect 36804 -25934 37824 -25869
rect 35357 -26064 35796 -26017
rect 36903 -26267 36949 -25967
rect 37001 -26267 37047 -25967
rect 37099 -26267 37145 -25967
rect 37341 -26267 37387 -25967
rect 37439 -26267 37485 -25967
rect 38046 -26375 38159 -24179
rect 38864 -24212 38994 -24062
rect 39150 -24116 39196 -23916
rect 39248 -24144 39294 -23916
rect 39346 -24116 39392 -23916
rect 39444 -24144 39490 -23916
rect 39681 -24062 39735 -23772
rect 40025 -24038 40071 -23739
rect 40123 -24038 40169 -23738
rect 40221 -24038 40267 -23702
rect 39681 -24116 40009 -24062
rect 39150 -24190 39787 -24144
rect 39955 -24171 40009 -24116
rect 38914 -25616 38968 -24212
rect 39150 -24446 39196 -24190
rect 39248 -24192 39490 -24190
rect 39346 -24446 39392 -24192
rect 39542 -24446 39588 -24190
rect 39929 -24229 40088 -24171
rect 40123 -24575 40169 -24275
rect 40319 -24575 40365 -23738
rect 40417 -24038 40463 -23702
rect 41119 -24210 41827 -24097
rect 40732 -24345 40778 -24245
rect 40830 -24374 40876 -24245
rect 40928 -24345 40974 -24245
rect 41026 -24374 41072 -24245
rect 40732 -24420 41369 -24374
rect 40732 -24576 40778 -24420
rect 40830 -24422 41072 -24420
rect 40928 -24576 40974 -24422
rect 41124 -24576 41170 -24420
rect 39124 -25475 39170 -25175
rect 38771 -25670 38968 -25616
rect 39026 -26011 39072 -25712
rect 39025 -26048 39072 -26011
rect 39124 -26012 39170 -25712
rect 39222 -26048 39268 -25712
rect 39320 -26012 39366 -25175
rect 39733 -25330 39779 -25174
rect 39929 -25328 39975 -25174
rect 39831 -25330 40073 -25328
rect 40125 -25330 40171 -25174
rect 39733 -25376 40370 -25330
rect 39733 -25505 39779 -25405
rect 39831 -25505 39877 -25376
rect 39929 -25505 39975 -25405
rect 40027 -25505 40073 -25376
rect 40571 -25686 40617 -25086
rect 40782 -25686 40828 -25086
rect 40880 -25686 40926 -25086
rect 40978 -25686 41024 -25086
rect 41190 -25686 41236 -25086
rect 39418 -26048 39464 -25712
rect 41421 -25817 41526 -25745
rect 41427 -25900 41492 -25817
rect 40472 -25965 41492 -25900
rect 39025 -26095 39464 -26048
rect 40571 -26298 40617 -25998
rect 40669 -26298 40715 -25998
rect 40767 -26298 40813 -25998
rect 41009 -26298 41055 -25998
rect 41107 -26298 41153 -25998
rect 29042 -26477 33387 -26395
rect 29046 -26508 33387 -26477
rect 37482 -26406 38159 -26375
rect 41714 -26406 41827 -24210
rect 41936 -25757 42201 -18424
rect 42378 -19883 50339 -19681
rect 42378 -23673 42580 -19883
rect 43462 -20273 43759 -20187
rect 45227 -20257 45666 -20210
rect 43462 -20327 44938 -20273
rect 45227 -20294 45274 -20257
rect 43462 -20409 43759 -20327
rect 44067 -20767 44197 -20617
rect 44353 -20671 44399 -20471
rect 44451 -20699 44497 -20471
rect 44549 -20671 44595 -20471
rect 44647 -20699 44693 -20471
rect 44884 -20617 44938 -20327
rect 45228 -20593 45274 -20294
rect 45326 -20593 45372 -20293
rect 45424 -20593 45470 -20257
rect 44884 -20671 45212 -20617
rect 44353 -20745 44990 -20699
rect 45158 -20726 45212 -20671
rect 44117 -22171 44171 -20767
rect 44353 -21001 44399 -20745
rect 44451 -20747 44693 -20745
rect 44549 -21001 44595 -20747
rect 44745 -21001 44791 -20745
rect 45132 -20784 45291 -20726
rect 45326 -21130 45372 -20830
rect 45522 -21130 45568 -20293
rect 45620 -20593 45666 -20257
rect 46322 -20765 47030 -20652
rect 45935 -20900 45981 -20800
rect 46033 -20929 46079 -20800
rect 46131 -20900 46177 -20800
rect 46229 -20929 46275 -20800
rect 45935 -20975 46572 -20929
rect 45935 -21131 45981 -20975
rect 46033 -20977 46275 -20975
rect 46131 -21131 46177 -20977
rect 46327 -21131 46373 -20975
rect 44327 -22030 44373 -21730
rect 43974 -22225 44171 -22171
rect 44229 -22566 44275 -22267
rect 44228 -22603 44275 -22566
rect 44327 -22567 44373 -22267
rect 44425 -22603 44471 -22267
rect 44523 -22567 44569 -21730
rect 44936 -21885 44982 -21729
rect 45132 -21883 45178 -21729
rect 45034 -21885 45276 -21883
rect 45328 -21885 45374 -21729
rect 44936 -21931 45573 -21885
rect 44936 -22060 44982 -21960
rect 45034 -22060 45080 -21931
rect 45132 -22060 45178 -21960
rect 45230 -22060 45276 -21931
rect 45774 -22241 45820 -21641
rect 45985 -22241 46031 -21641
rect 46083 -22241 46129 -21641
rect 46181 -22241 46227 -21641
rect 46393 -22241 46439 -21641
rect 44621 -22603 44667 -22267
rect 46624 -22372 46729 -22300
rect 46630 -22455 46695 -22372
rect 45675 -22520 46695 -22455
rect 44228 -22650 44667 -22603
rect 45774 -22853 45820 -22553
rect 45872 -22853 45918 -22553
rect 45970 -22853 46016 -22553
rect 46212 -22853 46258 -22553
rect 46310 -22853 46356 -22553
rect 46543 -22961 46656 -22960
rect 46917 -22961 47030 -20765
rect 47766 -21999 47812 -21499
rect 48035 -21999 48081 -21499
rect 48133 -21999 48179 -21499
rect 48231 -21999 48277 -21499
rect 48361 -21999 48407 -21499
rect 48687 -21999 48733 -21499
rect 48915 -21799 48961 -21499
rect 47535 -22159 47673 -22155
rect 48341 -22159 48479 -22155
rect 48726 -22159 48780 -22086
rect 47535 -22203 48780 -22159
rect 47535 -22209 47673 -22203
rect 48341 -22209 48479 -22203
rect 48726 -22224 48780 -22203
rect 48898 -22239 48964 -22227
rect 50137 -22239 50339 -19883
rect 47374 -22546 47477 -22455
rect 46353 -23074 47030 -22961
rect 42378 -23726 43708 -23673
rect 45219 -23710 45658 -23663
rect 42378 -23780 44930 -23726
rect 45219 -23747 45266 -23710
rect 42378 -23875 43708 -23780
rect 44059 -24220 44189 -24070
rect 44345 -24124 44391 -23924
rect 44443 -24152 44489 -23924
rect 44541 -24124 44587 -23924
rect 44639 -24152 44685 -23924
rect 44876 -24070 44930 -23780
rect 45220 -24046 45266 -23747
rect 45318 -24046 45364 -23746
rect 45416 -24046 45462 -23710
rect 44876 -24124 45204 -24070
rect 44345 -24198 44982 -24152
rect 45150 -24179 45204 -24124
rect 44109 -25624 44163 -24220
rect 44345 -24454 44391 -24198
rect 44443 -24200 44685 -24198
rect 44541 -24454 44587 -24200
rect 44737 -24454 44783 -24198
rect 45124 -24237 45283 -24179
rect 45318 -24583 45364 -24283
rect 45514 -24583 45560 -23746
rect 45612 -24046 45658 -23710
rect 46543 -24105 46656 -23074
rect 47386 -23179 47465 -22546
rect 47668 -22795 47714 -22495
rect 47766 -22795 47812 -22495
rect 48138 -22795 48184 -22295
rect 48236 -22795 48282 -22295
rect 48361 -22795 48407 -22295
rect 48459 -22795 48505 -22295
rect 48589 -22795 48635 -22295
rect 48687 -22795 48733 -22295
rect 48785 -22795 48831 -22295
rect 48898 -22301 50520 -22239
rect 48898 -22310 48964 -22301
rect 48915 -22795 48961 -22495
rect 49013 -22795 49059 -22495
rect 46886 -23258 47465 -23179
rect 46886 -23613 46965 -23258
rect 46860 -23710 46976 -23613
rect 48887 -23741 49326 -23694
rect 47489 -23757 47586 -23751
rect 47489 -23811 48598 -23757
rect 48887 -23778 48934 -23741
rect 47489 -23817 47586 -23811
rect 46314 -24218 47022 -24105
rect 45927 -24353 45973 -24253
rect 46025 -24382 46071 -24253
rect 46123 -24353 46169 -24253
rect 46221 -24382 46267 -24253
rect 45927 -24428 46564 -24382
rect 45927 -24584 45973 -24428
rect 46025 -24430 46267 -24428
rect 46123 -24584 46169 -24430
rect 46319 -24584 46365 -24428
rect 44319 -25483 44365 -25183
rect 43966 -25678 44163 -25624
rect 41936 -26088 42273 -25757
rect 44221 -26019 44267 -25720
rect 44220 -26056 44267 -26019
rect 44319 -26020 44365 -25720
rect 44417 -26056 44463 -25720
rect 44515 -26020 44561 -25183
rect 44928 -25338 44974 -25182
rect 45124 -25336 45170 -25182
rect 45026 -25338 45268 -25336
rect 45320 -25338 45366 -25182
rect 44928 -25384 45565 -25338
rect 44928 -25513 44974 -25413
rect 45026 -25513 45072 -25384
rect 45124 -25513 45170 -25413
rect 45222 -25513 45268 -25384
rect 45766 -25694 45812 -25094
rect 45977 -25694 46023 -25094
rect 46075 -25694 46121 -25094
rect 46173 -25694 46219 -25094
rect 46385 -25694 46431 -25094
rect 44613 -26056 44659 -25720
rect 46616 -25825 46721 -25753
rect 46622 -25908 46687 -25825
rect 45667 -25973 46687 -25908
rect 44220 -26103 44659 -26056
rect 45766 -26306 45812 -26006
rect 45864 -26306 45910 -26006
rect 45962 -26306 46008 -26006
rect 46204 -26306 46250 -26006
rect 46302 -26306 46348 -26006
rect 37482 -26488 41827 -26406
rect 46909 -26414 47022 -24218
rect 47727 -24251 47857 -24101
rect 48013 -24155 48059 -23955
rect 48111 -24183 48157 -23955
rect 48209 -24155 48255 -23955
rect 48307 -24183 48353 -23955
rect 48544 -24101 48598 -23811
rect 48888 -24077 48934 -23778
rect 48986 -24077 49032 -23777
rect 49084 -24077 49130 -23741
rect 48544 -24155 48872 -24101
rect 48013 -24229 48650 -24183
rect 48818 -24210 48872 -24155
rect 47777 -25655 47831 -24251
rect 48013 -24485 48059 -24229
rect 48111 -24231 48353 -24229
rect 48209 -24485 48255 -24231
rect 48405 -24485 48451 -24229
rect 48792 -24268 48951 -24210
rect 48986 -24614 49032 -24314
rect 49182 -24614 49228 -23777
rect 49280 -24077 49326 -23741
rect 49982 -24249 50690 -24136
rect 49595 -24384 49641 -24284
rect 49693 -24413 49739 -24284
rect 49791 -24384 49837 -24284
rect 49889 -24413 49935 -24284
rect 49595 -24459 50232 -24413
rect 49595 -24615 49641 -24459
rect 49693 -24461 49935 -24459
rect 49791 -24615 49837 -24461
rect 49987 -24615 50033 -24459
rect 47987 -25514 48033 -25214
rect 47634 -25709 47831 -25655
rect 47889 -26050 47935 -25751
rect 47888 -26087 47935 -26050
rect 47987 -26051 48033 -25751
rect 48085 -26087 48131 -25751
rect 48183 -26051 48229 -25214
rect 48596 -25369 48642 -25213
rect 48792 -25367 48838 -25213
rect 48694 -25369 48936 -25367
rect 48988 -25369 49034 -25213
rect 48596 -25415 49233 -25369
rect 48596 -25544 48642 -25444
rect 48694 -25544 48740 -25415
rect 48792 -25544 48838 -25444
rect 48890 -25544 48936 -25415
rect 49434 -25725 49480 -25125
rect 49645 -25725 49691 -25125
rect 49743 -25725 49789 -25125
rect 49841 -25725 49887 -25125
rect 50053 -25725 50099 -25125
rect 48281 -26087 48327 -25751
rect 50284 -25856 50389 -25784
rect 50290 -25939 50355 -25856
rect 49335 -26004 50355 -25939
rect 47888 -26134 48327 -26087
rect 49434 -26337 49480 -26037
rect 49532 -26337 49578 -26037
rect 49630 -26337 49676 -26037
rect 49872 -26337 49918 -26037
rect 49970 -26337 50016 -26037
rect 37486 -26519 41827 -26488
rect 46345 -26445 47022 -26414
rect 50577 -26445 50690 -24249
rect 50800 -25618 51026 -17944
rect 51657 -19948 59643 -19689
rect 51657 -23552 51916 -19948
rect 52453 -20239 52699 -20143
rect 54425 -20223 54864 -20176
rect 52453 -20293 54136 -20239
rect 54425 -20260 54472 -20223
rect 52453 -20363 52699 -20293
rect 53265 -20733 53395 -20583
rect 53551 -20637 53597 -20437
rect 53649 -20665 53695 -20437
rect 53747 -20637 53793 -20437
rect 53845 -20665 53891 -20437
rect 54082 -20583 54136 -20293
rect 54426 -20559 54472 -20260
rect 54524 -20559 54570 -20259
rect 54622 -20559 54668 -20223
rect 54082 -20637 54410 -20583
rect 53551 -20711 54188 -20665
rect 54356 -20692 54410 -20637
rect 53315 -22137 53369 -20733
rect 53551 -20967 53597 -20711
rect 53649 -20713 53891 -20711
rect 53747 -20967 53793 -20713
rect 53943 -20967 53989 -20711
rect 54330 -20750 54489 -20692
rect 54524 -21096 54570 -20796
rect 54720 -21096 54766 -20259
rect 54818 -20559 54864 -20223
rect 55520 -20731 56228 -20618
rect 55133 -20866 55179 -20766
rect 55231 -20895 55277 -20766
rect 55329 -20866 55375 -20766
rect 55427 -20895 55473 -20766
rect 55133 -20941 55770 -20895
rect 55133 -21097 55179 -20941
rect 55231 -20943 55473 -20941
rect 55329 -21097 55375 -20943
rect 55525 -21097 55571 -20941
rect 53525 -21996 53571 -21696
rect 53172 -22191 53369 -22137
rect 53427 -22532 53473 -22233
rect 53426 -22569 53473 -22532
rect 53525 -22533 53571 -22233
rect 53623 -22569 53669 -22233
rect 53721 -22533 53767 -21696
rect 54134 -21851 54180 -21695
rect 54330 -21849 54376 -21695
rect 54232 -21851 54474 -21849
rect 54526 -21851 54572 -21695
rect 54134 -21897 54771 -21851
rect 54134 -22026 54180 -21926
rect 54232 -22026 54278 -21897
rect 54330 -22026 54376 -21926
rect 54428 -22026 54474 -21897
rect 54972 -22207 55018 -21607
rect 55183 -22207 55229 -21607
rect 55281 -22207 55327 -21607
rect 55379 -22207 55425 -21607
rect 55591 -22207 55637 -21607
rect 53819 -22569 53865 -22233
rect 55822 -22338 55927 -22266
rect 55828 -22421 55893 -22338
rect 54873 -22486 55893 -22421
rect 53426 -22616 53865 -22569
rect 54972 -22819 55018 -22519
rect 55070 -22819 55116 -22519
rect 55168 -22819 55214 -22519
rect 55410 -22819 55456 -22519
rect 55508 -22819 55554 -22519
rect 55741 -22927 55854 -22926
rect 56115 -22927 56228 -20731
rect 56964 -21965 57010 -21465
rect 57233 -21965 57279 -21465
rect 57331 -21965 57377 -21465
rect 57429 -21965 57475 -21465
rect 57559 -21965 57605 -21465
rect 57885 -21965 57931 -21465
rect 58113 -21765 58159 -21465
rect 56733 -22125 56871 -22121
rect 57539 -22125 57677 -22121
rect 57924 -22125 57978 -22052
rect 56733 -22169 57978 -22125
rect 56733 -22175 56871 -22169
rect 57539 -22175 57677 -22169
rect 57924 -22190 57978 -22169
rect 58096 -22205 58162 -22193
rect 59384 -22205 59643 -19948
rect 59994 -20005 60215 -17387
rect 60446 -19968 68430 -19730
rect 59891 -20319 60267 -20005
rect 56572 -22512 56675 -22421
rect 55551 -23040 56228 -22927
rect 51657 -23692 52865 -23552
rect 54417 -23676 54856 -23629
rect 51657 -23746 54128 -23692
rect 54417 -23713 54464 -23676
rect 51657 -23811 52865 -23746
rect 53257 -24186 53387 -24036
rect 53543 -24090 53589 -23890
rect 53641 -24118 53687 -23890
rect 53739 -24090 53785 -23890
rect 53837 -24118 53883 -23890
rect 54074 -24036 54128 -23746
rect 54418 -24012 54464 -23713
rect 54516 -24012 54562 -23712
rect 54614 -24012 54660 -23676
rect 54074 -24090 54402 -24036
rect 53543 -24164 54180 -24118
rect 54348 -24145 54402 -24090
rect 53307 -25590 53361 -24186
rect 53543 -24420 53589 -24164
rect 53641 -24166 53883 -24164
rect 53739 -24420 53785 -24166
rect 53935 -24420 53981 -24164
rect 54322 -24203 54481 -24145
rect 54516 -24549 54562 -24249
rect 54712 -24549 54758 -23712
rect 54810 -24012 54856 -23676
rect 55741 -24071 55854 -23040
rect 56584 -23145 56663 -22512
rect 56866 -22761 56912 -22461
rect 56964 -22761 57010 -22461
rect 57336 -22761 57382 -22261
rect 57434 -22761 57480 -22261
rect 57559 -22761 57605 -22261
rect 57657 -22761 57703 -22261
rect 57787 -22761 57833 -22261
rect 57885 -22761 57931 -22261
rect 57983 -22761 58029 -22261
rect 58096 -22267 59718 -22205
rect 58096 -22276 58162 -22267
rect 58113 -22761 58159 -22461
rect 58211 -22761 58257 -22461
rect 56084 -23224 56663 -23145
rect 56084 -23579 56163 -23224
rect 56058 -23676 56174 -23579
rect 58085 -23707 58524 -23660
rect 56687 -23723 56784 -23717
rect 56687 -23777 57796 -23723
rect 58085 -23744 58132 -23707
rect 56687 -23783 56784 -23777
rect 55512 -24184 56220 -24071
rect 55125 -24319 55171 -24219
rect 55223 -24348 55269 -24219
rect 55321 -24319 55367 -24219
rect 55419 -24348 55465 -24219
rect 55125 -24394 55762 -24348
rect 55125 -24550 55171 -24394
rect 55223 -24396 55465 -24394
rect 55321 -24550 55367 -24396
rect 55517 -24550 55563 -24394
rect 53517 -25449 53563 -25149
rect 50778 -26118 51076 -25618
rect 53164 -25644 53361 -25590
rect 53419 -25985 53465 -25686
rect 53418 -26022 53465 -25985
rect 53517 -25986 53563 -25686
rect 53615 -26022 53661 -25686
rect 53713 -25986 53759 -25149
rect 54126 -25304 54172 -25148
rect 54322 -25302 54368 -25148
rect 54224 -25304 54466 -25302
rect 54518 -25304 54564 -25148
rect 54126 -25350 54763 -25304
rect 54126 -25479 54172 -25379
rect 54224 -25479 54270 -25350
rect 54322 -25479 54368 -25379
rect 54420 -25479 54466 -25350
rect 54964 -25660 55010 -25060
rect 55175 -25660 55221 -25060
rect 55273 -25660 55319 -25060
rect 55371 -25660 55417 -25060
rect 55583 -25660 55629 -25060
rect 53811 -26022 53857 -25686
rect 55814 -25791 55919 -25719
rect 55820 -25874 55885 -25791
rect 54865 -25939 55885 -25874
rect 53418 -26069 53857 -26022
rect 54964 -26272 55010 -25972
rect 55062 -26272 55108 -25972
rect 55160 -26272 55206 -25972
rect 55402 -26272 55448 -25972
rect 55500 -26272 55546 -25972
rect 56107 -26380 56220 -24184
rect 56925 -24217 57055 -24067
rect 57211 -24121 57257 -23921
rect 57309 -24149 57355 -23921
rect 57407 -24121 57453 -23921
rect 57505 -24149 57551 -23921
rect 57742 -24067 57796 -23777
rect 58086 -24043 58132 -23744
rect 58184 -24043 58230 -23743
rect 58282 -24043 58328 -23707
rect 57742 -24121 58070 -24067
rect 57211 -24195 57848 -24149
rect 58016 -24176 58070 -24121
rect 56975 -25621 57029 -24217
rect 57211 -24451 57257 -24195
rect 57309 -24197 57551 -24195
rect 57407 -24451 57453 -24197
rect 57603 -24451 57649 -24195
rect 57990 -24234 58149 -24176
rect 58184 -24580 58230 -24280
rect 58380 -24580 58426 -23743
rect 58478 -24043 58524 -23707
rect 59180 -24215 59888 -24102
rect 58793 -24350 58839 -24250
rect 58891 -24379 58937 -24250
rect 58989 -24350 59035 -24250
rect 59087 -24379 59133 -24250
rect 58793 -24425 59430 -24379
rect 58793 -24581 58839 -24425
rect 58891 -24427 59133 -24425
rect 58989 -24581 59035 -24427
rect 59185 -24581 59231 -24425
rect 57185 -25480 57231 -25180
rect 56832 -25675 57029 -25621
rect 57087 -26016 57133 -25717
rect 57086 -26053 57133 -26016
rect 57185 -26017 57231 -25717
rect 57283 -26053 57329 -25717
rect 57381 -26017 57427 -25180
rect 57794 -25335 57840 -25179
rect 57990 -25333 58036 -25179
rect 57892 -25335 58134 -25333
rect 58186 -25335 58232 -25179
rect 57794 -25381 58431 -25335
rect 57794 -25510 57840 -25410
rect 57892 -25510 57938 -25381
rect 57990 -25510 58036 -25410
rect 58088 -25510 58134 -25381
rect 58632 -25691 58678 -25091
rect 58843 -25691 58889 -25091
rect 58941 -25691 58987 -25091
rect 59039 -25691 59085 -25091
rect 59251 -25691 59297 -25091
rect 57479 -26053 57525 -25717
rect 59482 -25822 59587 -25750
rect 59488 -25905 59553 -25822
rect 58533 -25970 59553 -25905
rect 57086 -26100 57525 -26053
rect 58632 -26303 58678 -26003
rect 58730 -26303 58776 -26003
rect 58828 -26303 58874 -26003
rect 59070 -26303 59116 -26003
rect 59168 -26303 59214 -26003
rect 46345 -26527 50690 -26445
rect 55543 -26411 56220 -26380
rect 59775 -26411 59888 -24215
rect 59994 -25756 60215 -20319
rect 60446 -23492 60684 -19968
rect 61492 -20173 61742 -20073
rect 63179 -20157 63618 -20110
rect 61492 -20227 62890 -20173
rect 63179 -20194 63226 -20157
rect 61492 -20302 61742 -20227
rect 62019 -20667 62149 -20517
rect 62305 -20571 62351 -20371
rect 62403 -20599 62449 -20371
rect 62501 -20571 62547 -20371
rect 62599 -20599 62645 -20371
rect 62836 -20517 62890 -20227
rect 63180 -20493 63226 -20194
rect 63278 -20493 63324 -20193
rect 63376 -20493 63422 -20157
rect 62836 -20571 63164 -20517
rect 62305 -20645 62942 -20599
rect 63110 -20626 63164 -20571
rect 62069 -22071 62123 -20667
rect 62305 -20901 62351 -20645
rect 62403 -20647 62645 -20645
rect 62501 -20901 62547 -20647
rect 62697 -20901 62743 -20645
rect 63084 -20684 63243 -20626
rect 63278 -21030 63324 -20730
rect 63474 -21030 63520 -20193
rect 63572 -20493 63618 -20157
rect 64274 -20665 64982 -20552
rect 63887 -20800 63933 -20700
rect 63985 -20829 64031 -20700
rect 64083 -20800 64129 -20700
rect 64181 -20829 64227 -20700
rect 63887 -20875 64524 -20829
rect 63887 -21031 63933 -20875
rect 63985 -20877 64227 -20875
rect 64083 -21031 64129 -20877
rect 64279 -21031 64325 -20875
rect 62279 -21930 62325 -21630
rect 61926 -22125 62123 -22071
rect 62181 -22466 62227 -22167
rect 62180 -22503 62227 -22466
rect 62279 -22467 62325 -22167
rect 62377 -22503 62423 -22167
rect 62475 -22467 62521 -21630
rect 62888 -21785 62934 -21629
rect 63084 -21783 63130 -21629
rect 62986 -21785 63228 -21783
rect 63280 -21785 63326 -21629
rect 62888 -21831 63525 -21785
rect 62888 -21960 62934 -21860
rect 62986 -21960 63032 -21831
rect 63084 -21960 63130 -21860
rect 63182 -21960 63228 -21831
rect 63726 -22141 63772 -21541
rect 63937 -22141 63983 -21541
rect 64035 -22141 64081 -21541
rect 64133 -22141 64179 -21541
rect 64345 -22141 64391 -21541
rect 62573 -22503 62619 -22167
rect 64576 -22272 64681 -22200
rect 64582 -22355 64647 -22272
rect 63627 -22420 64647 -22355
rect 62180 -22550 62619 -22503
rect 63726 -22753 63772 -22453
rect 63824 -22753 63870 -22453
rect 63922 -22753 63968 -22453
rect 64164 -22753 64210 -22453
rect 64262 -22753 64308 -22453
rect 64495 -22861 64608 -22860
rect 64869 -22861 64982 -20665
rect 65718 -21899 65764 -21399
rect 65987 -21899 66033 -21399
rect 66085 -21899 66131 -21399
rect 66183 -21899 66229 -21399
rect 66313 -21899 66359 -21399
rect 66639 -21899 66685 -21399
rect 66867 -21699 66913 -21399
rect 65487 -22059 65625 -22055
rect 66293 -22059 66431 -22055
rect 66678 -22059 66732 -21986
rect 65487 -22103 66732 -22059
rect 65487 -22109 65625 -22103
rect 66293 -22109 66431 -22103
rect 66678 -22124 66732 -22103
rect 66850 -22139 66916 -22127
rect 68192 -22139 68430 -19968
rect 68747 -20010 68924 -16828
rect 69232 -19976 77620 -19676
rect 68667 -20301 69005 -20010
rect 65326 -22446 65429 -22355
rect 64305 -22974 64982 -22861
rect 60446 -23626 61582 -23492
rect 63171 -23610 63610 -23563
rect 60446 -23680 62882 -23626
rect 63171 -23647 63218 -23610
rect 60446 -23730 61582 -23680
rect 62011 -24120 62141 -23970
rect 62297 -24024 62343 -23824
rect 62395 -24052 62441 -23824
rect 62493 -24024 62539 -23824
rect 62591 -24052 62637 -23824
rect 62828 -23970 62882 -23680
rect 63172 -23946 63218 -23647
rect 63270 -23946 63316 -23646
rect 63368 -23946 63414 -23610
rect 62828 -24024 63156 -23970
rect 62297 -24098 62934 -24052
rect 63102 -24079 63156 -24024
rect 62061 -25524 62115 -24120
rect 62297 -24354 62343 -24098
rect 62395 -24100 62637 -24098
rect 62493 -24354 62539 -24100
rect 62689 -24354 62735 -24098
rect 63076 -24137 63235 -24079
rect 63270 -24483 63316 -24183
rect 63466 -24483 63512 -23646
rect 63564 -23946 63610 -23610
rect 64495 -24005 64608 -22974
rect 65338 -23079 65417 -22446
rect 65620 -22695 65666 -22395
rect 65718 -22695 65764 -22395
rect 66090 -22695 66136 -22195
rect 66188 -22695 66234 -22195
rect 66313 -22695 66359 -22195
rect 66411 -22695 66457 -22195
rect 66541 -22695 66587 -22195
rect 66639 -22695 66685 -22195
rect 66737 -22695 66783 -22195
rect 66850 -22201 68472 -22139
rect 66850 -22210 66916 -22201
rect 66867 -22695 66913 -22395
rect 66965 -22695 67011 -22395
rect 64838 -23158 65417 -23079
rect 64838 -23513 64917 -23158
rect 64812 -23610 64928 -23513
rect 66839 -23641 67278 -23594
rect 65441 -23657 65538 -23651
rect 65441 -23711 66550 -23657
rect 66839 -23678 66886 -23641
rect 65441 -23717 65538 -23711
rect 64266 -24118 64974 -24005
rect 63879 -24253 63925 -24153
rect 63977 -24282 64023 -24153
rect 64075 -24253 64121 -24153
rect 64173 -24282 64219 -24153
rect 63879 -24328 64516 -24282
rect 63879 -24484 63925 -24328
rect 63977 -24330 64219 -24328
rect 64075 -24484 64121 -24330
rect 64271 -24484 64317 -24328
rect 62271 -25383 62317 -25083
rect 61918 -25578 62115 -25524
rect 59940 -26055 60232 -25756
rect 62173 -25919 62219 -25620
rect 62172 -25956 62219 -25919
rect 62271 -25920 62317 -25620
rect 62369 -25956 62415 -25620
rect 62467 -25920 62513 -25083
rect 62880 -25238 62926 -25082
rect 63076 -25236 63122 -25082
rect 62978 -25238 63220 -25236
rect 63272 -25238 63318 -25082
rect 62880 -25284 63517 -25238
rect 62880 -25413 62926 -25313
rect 62978 -25413 63024 -25284
rect 63076 -25413 63122 -25313
rect 63174 -25413 63220 -25284
rect 63718 -25594 63764 -24994
rect 63929 -25594 63975 -24994
rect 64027 -25594 64073 -24994
rect 64125 -25594 64171 -24994
rect 64337 -25594 64383 -24994
rect 62565 -25956 62611 -25620
rect 64568 -25725 64673 -25653
rect 64574 -25808 64639 -25725
rect 63619 -25873 64639 -25808
rect 62172 -26003 62611 -25956
rect 63718 -26206 63764 -25906
rect 63816 -26206 63862 -25906
rect 63914 -26206 63960 -25906
rect 64156 -26206 64202 -25906
rect 64254 -26206 64300 -25906
rect 64861 -26314 64974 -24118
rect 65679 -24151 65809 -24001
rect 65965 -24055 66011 -23855
rect 66063 -24083 66109 -23855
rect 66161 -24055 66207 -23855
rect 66259 -24083 66305 -23855
rect 66496 -24001 66550 -23711
rect 66840 -23977 66886 -23678
rect 66938 -23977 66984 -23677
rect 67036 -23977 67082 -23641
rect 66496 -24055 66824 -24001
rect 65965 -24129 66602 -24083
rect 66770 -24110 66824 -24055
rect 65729 -25555 65783 -24151
rect 65965 -24385 66011 -24129
rect 66063 -24131 66305 -24129
rect 66161 -24385 66207 -24131
rect 66357 -24385 66403 -24129
rect 66744 -24168 66903 -24110
rect 66938 -24514 66984 -24214
rect 67134 -24514 67180 -23677
rect 67232 -23977 67278 -23641
rect 67934 -24149 68642 -24036
rect 67547 -24284 67593 -24184
rect 67645 -24313 67691 -24184
rect 67743 -24284 67789 -24184
rect 67841 -24313 67887 -24184
rect 67547 -24359 68184 -24313
rect 67547 -24515 67593 -24359
rect 67645 -24361 67887 -24359
rect 67743 -24515 67789 -24361
rect 67939 -24515 67985 -24359
rect 65939 -25414 65985 -25114
rect 65586 -25609 65783 -25555
rect 65841 -25950 65887 -25651
rect 65840 -25987 65887 -25950
rect 65939 -25951 65985 -25651
rect 66037 -25987 66083 -25651
rect 66135 -25951 66181 -25114
rect 66548 -25269 66594 -25113
rect 66744 -25267 66790 -25113
rect 66646 -25269 66888 -25267
rect 66940 -25269 66986 -25113
rect 66548 -25315 67185 -25269
rect 66548 -25444 66594 -25344
rect 66646 -25444 66692 -25315
rect 66744 -25444 66790 -25344
rect 66842 -25444 66888 -25315
rect 67386 -25625 67432 -25025
rect 67597 -25625 67643 -25025
rect 67695 -25625 67741 -25025
rect 67793 -25625 67839 -25025
rect 68005 -25625 68051 -25025
rect 66233 -25987 66279 -25651
rect 68236 -25756 68341 -25684
rect 68242 -25839 68307 -25756
rect 67287 -25904 68307 -25839
rect 65840 -26034 66279 -25987
rect 67386 -26237 67432 -25937
rect 67484 -26237 67530 -25937
rect 67582 -26237 67628 -25937
rect 67824 -26237 67870 -25937
rect 67922 -26237 67968 -25937
rect 55543 -26493 59888 -26411
rect 64297 -26345 64974 -26314
rect 68529 -26345 68642 -24149
rect 68747 -25698 68924 -20301
rect 69232 -23426 69532 -19976
rect 70655 -20156 70923 -20065
rect 72332 -20140 72771 -20093
rect 70655 -20210 72043 -20156
rect 72332 -20177 72379 -20140
rect 70655 -20305 70923 -20210
rect 71172 -20650 71302 -20500
rect 71458 -20554 71504 -20354
rect 71556 -20582 71602 -20354
rect 71654 -20554 71700 -20354
rect 71752 -20582 71798 -20354
rect 71989 -20500 72043 -20210
rect 72333 -20476 72379 -20177
rect 72431 -20476 72477 -20176
rect 72529 -20476 72575 -20140
rect 71989 -20554 72317 -20500
rect 71458 -20628 72095 -20582
rect 72263 -20609 72317 -20554
rect 71222 -22054 71276 -20650
rect 71458 -20884 71504 -20628
rect 71556 -20630 71798 -20628
rect 71654 -20884 71700 -20630
rect 71850 -20884 71896 -20628
rect 72237 -20667 72396 -20609
rect 72431 -21013 72477 -20713
rect 72627 -21013 72673 -20176
rect 72725 -20476 72771 -20140
rect 73427 -20648 74135 -20535
rect 73040 -20783 73086 -20683
rect 73138 -20812 73184 -20683
rect 73236 -20783 73282 -20683
rect 73334 -20812 73380 -20683
rect 73040 -20858 73677 -20812
rect 73040 -21014 73086 -20858
rect 73138 -20860 73380 -20858
rect 73236 -21014 73282 -20860
rect 73432 -21014 73478 -20858
rect 71432 -21913 71478 -21613
rect 71079 -22108 71276 -22054
rect 71334 -22449 71380 -22150
rect 71333 -22486 71380 -22449
rect 71432 -22450 71478 -22150
rect 71530 -22486 71576 -22150
rect 71628 -22450 71674 -21613
rect 72041 -21768 72087 -21612
rect 72237 -21766 72283 -21612
rect 72139 -21768 72381 -21766
rect 72433 -21768 72479 -21612
rect 72041 -21814 72678 -21768
rect 72041 -21943 72087 -21843
rect 72139 -21943 72185 -21814
rect 72237 -21943 72283 -21843
rect 72335 -21943 72381 -21814
rect 72879 -22124 72925 -21524
rect 73090 -22124 73136 -21524
rect 73188 -22124 73234 -21524
rect 73286 -22124 73332 -21524
rect 73498 -22124 73544 -21524
rect 71726 -22486 71772 -22150
rect 73729 -22255 73834 -22183
rect 73735 -22338 73800 -22255
rect 72780 -22403 73800 -22338
rect 71333 -22533 71772 -22486
rect 72879 -22736 72925 -22436
rect 72977 -22736 73023 -22436
rect 73075 -22736 73121 -22436
rect 73317 -22736 73363 -22436
rect 73415 -22736 73461 -22436
rect 73648 -22844 73761 -22843
rect 74022 -22844 74135 -20648
rect 74871 -21882 74917 -21382
rect 75140 -21882 75186 -21382
rect 75238 -21882 75284 -21382
rect 75336 -21882 75382 -21382
rect 75466 -21882 75512 -21382
rect 75792 -21882 75838 -21382
rect 76020 -21682 76066 -21382
rect 74640 -22042 74778 -22038
rect 75446 -22042 75584 -22038
rect 75831 -22042 75885 -21969
rect 74640 -22086 75885 -22042
rect 74640 -22092 74778 -22086
rect 75446 -22092 75584 -22086
rect 75831 -22107 75885 -22086
rect 76003 -22122 76069 -22110
rect 77313 -22122 77620 -19976
rect 74479 -22429 74582 -22338
rect 73458 -22957 74135 -22844
rect 69232 -23609 70722 -23426
rect 72324 -23593 72763 -23546
rect 69232 -23663 72035 -23609
rect 72324 -23630 72371 -23593
rect 69232 -23726 70722 -23663
rect 71164 -24103 71294 -23953
rect 71450 -24007 71496 -23807
rect 71548 -24035 71594 -23807
rect 71646 -24007 71692 -23807
rect 71744 -24035 71790 -23807
rect 71981 -23953 72035 -23663
rect 72325 -23929 72371 -23630
rect 72423 -23929 72469 -23629
rect 72521 -23929 72567 -23593
rect 71981 -24007 72309 -23953
rect 71450 -24081 72087 -24035
rect 72255 -24062 72309 -24007
rect 71214 -25507 71268 -24103
rect 71450 -24337 71496 -24081
rect 71548 -24083 71790 -24081
rect 71646 -24337 71692 -24083
rect 71842 -24337 71888 -24081
rect 72229 -24120 72388 -24062
rect 72423 -24466 72469 -24166
rect 72619 -24466 72665 -23629
rect 72717 -23929 72763 -23593
rect 73648 -23988 73761 -22957
rect 74491 -23062 74570 -22429
rect 74773 -22678 74819 -22378
rect 74871 -22678 74917 -22378
rect 75243 -22678 75289 -22178
rect 75341 -22678 75387 -22178
rect 75466 -22678 75512 -22178
rect 75564 -22678 75610 -22178
rect 75694 -22678 75740 -22178
rect 75792 -22678 75838 -22178
rect 75890 -22678 75936 -22178
rect 76003 -22184 77625 -22122
rect 76003 -22193 76069 -22184
rect 76020 -22678 76066 -22378
rect 76118 -22678 76164 -22378
rect 73991 -23141 74570 -23062
rect 73991 -23496 74070 -23141
rect 73965 -23593 74081 -23496
rect 75992 -23624 76431 -23577
rect 74594 -23640 74691 -23634
rect 74594 -23694 75703 -23640
rect 75992 -23661 76039 -23624
rect 74594 -23700 74691 -23694
rect 73419 -24101 74127 -23988
rect 73032 -24236 73078 -24136
rect 73130 -24265 73176 -24136
rect 73228 -24236 73274 -24136
rect 73326 -24265 73372 -24136
rect 73032 -24311 73669 -24265
rect 73032 -24467 73078 -24311
rect 73130 -24313 73372 -24311
rect 73228 -24467 73274 -24313
rect 73424 -24467 73470 -24311
rect 71424 -25366 71470 -25066
rect 71071 -25561 71268 -25507
rect 68705 -26002 68966 -25698
rect 71326 -25902 71372 -25603
rect 71325 -25939 71372 -25902
rect 71424 -25903 71470 -25603
rect 71522 -25939 71568 -25603
rect 71620 -25903 71666 -25066
rect 72033 -25221 72079 -25065
rect 72229 -25219 72275 -25065
rect 72131 -25221 72373 -25219
rect 72425 -25221 72471 -25065
rect 72033 -25267 72670 -25221
rect 72033 -25396 72079 -25296
rect 72131 -25396 72177 -25267
rect 72229 -25396 72275 -25296
rect 72327 -25396 72373 -25267
rect 72871 -25577 72917 -24977
rect 73082 -25577 73128 -24977
rect 73180 -25577 73226 -24977
rect 73278 -25577 73324 -24977
rect 73490 -25577 73536 -24977
rect 71718 -25939 71764 -25603
rect 73721 -25708 73826 -25636
rect 73727 -25791 73792 -25708
rect 72772 -25856 73792 -25791
rect 71325 -25986 71764 -25939
rect 72871 -26189 72917 -25889
rect 72969 -26189 73015 -25889
rect 73067 -26189 73113 -25889
rect 73309 -26189 73355 -25889
rect 73407 -26189 73453 -25889
rect 74014 -26297 74127 -24101
rect 74832 -24134 74962 -23984
rect 75118 -24038 75164 -23838
rect 75216 -24066 75262 -23838
rect 75314 -24038 75360 -23838
rect 75412 -24066 75458 -23838
rect 75649 -23984 75703 -23694
rect 75993 -23960 76039 -23661
rect 76091 -23960 76137 -23660
rect 76189 -23960 76235 -23624
rect 75649 -24038 75977 -23984
rect 75118 -24112 75755 -24066
rect 75923 -24093 75977 -24038
rect 74882 -25538 74936 -24134
rect 75118 -24368 75164 -24112
rect 75216 -24114 75458 -24112
rect 75314 -24368 75360 -24114
rect 75510 -24368 75556 -24112
rect 75897 -24151 76056 -24093
rect 76091 -24497 76137 -24197
rect 76287 -24497 76333 -23660
rect 76385 -23960 76431 -23624
rect 77087 -24132 77795 -24019
rect 76700 -24267 76746 -24167
rect 76798 -24296 76844 -24167
rect 76896 -24267 76942 -24167
rect 76994 -24296 77040 -24167
rect 76700 -24342 77337 -24296
rect 76700 -24498 76746 -24342
rect 76798 -24344 77040 -24342
rect 76896 -24498 76942 -24344
rect 77092 -24498 77138 -24342
rect 75092 -25397 75138 -25097
rect 74739 -25592 74936 -25538
rect 74994 -25933 75040 -25634
rect 74993 -25970 75040 -25933
rect 75092 -25934 75138 -25634
rect 75190 -25970 75236 -25634
rect 75288 -25934 75334 -25097
rect 75701 -25252 75747 -25096
rect 75897 -25250 75943 -25096
rect 75799 -25252 76041 -25250
rect 76093 -25252 76139 -25096
rect 75701 -25298 76338 -25252
rect 75701 -25427 75747 -25327
rect 75799 -25427 75845 -25298
rect 75897 -25427 75943 -25327
rect 75995 -25427 76041 -25298
rect 76539 -25608 76585 -25008
rect 76750 -25608 76796 -25008
rect 76848 -25608 76894 -25008
rect 76946 -25608 76992 -25008
rect 77158 -25608 77204 -25008
rect 75386 -25970 75432 -25634
rect 77389 -25739 77494 -25667
rect 77395 -25822 77460 -25739
rect 76440 -25887 77460 -25822
rect 74993 -26017 75432 -25970
rect 76539 -26220 76585 -25920
rect 76637 -26220 76683 -25920
rect 76735 -26220 76781 -25920
rect 76977 -26220 77023 -25920
rect 77075 -26220 77121 -25920
rect 64297 -26427 68642 -26345
rect 73450 -26328 74127 -26297
rect 77682 -26328 77795 -24132
rect 77881 -26022 78192 -16378
rect 78457 -19894 86976 -19675
rect 78457 -23532 78676 -19894
rect 79910 -20118 80205 -20003
rect 81696 -20102 82135 -20055
rect 79910 -20172 81407 -20118
rect 81696 -20139 81743 -20102
rect 79910 -20276 80205 -20172
rect 80536 -20612 80666 -20462
rect 80822 -20516 80868 -20316
rect 80920 -20544 80966 -20316
rect 81018 -20516 81064 -20316
rect 81116 -20544 81162 -20316
rect 81353 -20462 81407 -20172
rect 81697 -20438 81743 -20139
rect 81795 -20438 81841 -20138
rect 81893 -20438 81939 -20102
rect 81353 -20516 81681 -20462
rect 80822 -20590 81459 -20544
rect 81627 -20571 81681 -20516
rect 80586 -22016 80640 -20612
rect 80822 -20846 80868 -20590
rect 80920 -20592 81162 -20590
rect 81018 -20846 81064 -20592
rect 81214 -20846 81260 -20590
rect 81601 -20629 81760 -20571
rect 81795 -20975 81841 -20675
rect 81991 -20975 82037 -20138
rect 82089 -20438 82135 -20102
rect 82791 -20610 83499 -20497
rect 82404 -20745 82450 -20645
rect 82502 -20774 82548 -20645
rect 82600 -20745 82646 -20645
rect 82698 -20774 82744 -20645
rect 82404 -20820 83041 -20774
rect 82404 -20976 82450 -20820
rect 82502 -20822 82744 -20820
rect 82600 -20976 82646 -20822
rect 82796 -20976 82842 -20820
rect 80796 -21875 80842 -21575
rect 80443 -22070 80640 -22016
rect 80698 -22411 80744 -22112
rect 80697 -22448 80744 -22411
rect 80796 -22412 80842 -22112
rect 80894 -22448 80940 -22112
rect 80992 -22412 81038 -21575
rect 81405 -21730 81451 -21574
rect 81601 -21728 81647 -21574
rect 81503 -21730 81745 -21728
rect 81797 -21730 81843 -21574
rect 81405 -21776 82042 -21730
rect 81405 -21905 81451 -21805
rect 81503 -21905 81549 -21776
rect 81601 -21905 81647 -21805
rect 81699 -21905 81745 -21776
rect 82243 -22086 82289 -21486
rect 82454 -22086 82500 -21486
rect 82552 -22086 82598 -21486
rect 82650 -22086 82696 -21486
rect 82862 -22086 82908 -21486
rect 81090 -22448 81136 -22112
rect 83093 -22217 83198 -22145
rect 83099 -22300 83164 -22217
rect 82144 -22365 83164 -22300
rect 80697 -22495 81136 -22448
rect 82243 -22698 82289 -22398
rect 82341 -22698 82387 -22398
rect 82439 -22698 82485 -22398
rect 82681 -22698 82727 -22398
rect 82779 -22698 82825 -22398
rect 83012 -22806 83125 -22805
rect 83386 -22806 83499 -20610
rect 84235 -21844 84281 -21344
rect 84504 -21844 84550 -21344
rect 84602 -21844 84648 -21344
rect 84700 -21844 84746 -21344
rect 84830 -21844 84876 -21344
rect 85156 -21844 85202 -21344
rect 85384 -21644 85430 -21344
rect 84004 -22004 84142 -22000
rect 84810 -22004 84948 -22000
rect 85195 -22004 85249 -21931
rect 84004 -22048 85249 -22004
rect 84004 -22054 84142 -22048
rect 84810 -22054 84948 -22048
rect 85195 -22069 85249 -22048
rect 85367 -22084 85433 -22072
rect 86757 -22084 86976 -19894
rect 83843 -22391 83946 -22300
rect 82822 -22919 83499 -22806
rect 78457 -23571 80236 -23532
rect 81688 -23555 82127 -23508
rect 78457 -23625 81399 -23571
rect 81688 -23592 81735 -23555
rect 78457 -23751 80236 -23625
rect 80528 -24065 80658 -23915
rect 80814 -23969 80860 -23769
rect 80912 -23997 80958 -23769
rect 81010 -23969 81056 -23769
rect 81108 -23997 81154 -23769
rect 81345 -23915 81399 -23625
rect 81689 -23891 81735 -23592
rect 81787 -23891 81833 -23591
rect 81885 -23891 81931 -23555
rect 81345 -23969 81673 -23915
rect 80814 -24043 81451 -23997
rect 81619 -24024 81673 -23969
rect 80578 -25469 80632 -24065
rect 80814 -24299 80860 -24043
rect 80912 -24045 81154 -24043
rect 81010 -24299 81056 -24045
rect 81206 -24299 81252 -24043
rect 81593 -24082 81752 -24024
rect 81787 -24428 81833 -24128
rect 81983 -24428 82029 -23591
rect 82081 -23891 82127 -23555
rect 83012 -23950 83125 -22919
rect 83855 -23024 83934 -22391
rect 84137 -22640 84183 -22340
rect 84235 -22640 84281 -22340
rect 84607 -22640 84653 -22140
rect 84705 -22640 84751 -22140
rect 84830 -22640 84876 -22140
rect 84928 -22640 84974 -22140
rect 85058 -22640 85104 -22140
rect 85156 -22640 85202 -22140
rect 85254 -22640 85300 -22140
rect 85367 -22146 86989 -22084
rect 85367 -22155 85433 -22146
rect 85384 -22640 85430 -22340
rect 85482 -22640 85528 -22340
rect 83355 -23103 83934 -23024
rect 83355 -23458 83434 -23103
rect 83329 -23555 83445 -23458
rect 85356 -23586 85795 -23539
rect 83958 -23602 84055 -23596
rect 83958 -23656 85067 -23602
rect 85356 -23623 85403 -23586
rect 83958 -23662 84055 -23656
rect 82783 -24063 83491 -23950
rect 82396 -24198 82442 -24098
rect 82494 -24227 82540 -24098
rect 82592 -24198 82638 -24098
rect 82690 -24227 82736 -24098
rect 82396 -24273 83033 -24227
rect 82396 -24429 82442 -24273
rect 82494 -24275 82736 -24273
rect 82592 -24429 82638 -24275
rect 82788 -24429 82834 -24273
rect 80788 -25328 80834 -25028
rect 80435 -25523 80632 -25469
rect 80690 -25864 80736 -25565
rect 80689 -25901 80736 -25864
rect 80788 -25865 80834 -25565
rect 80886 -25901 80932 -25565
rect 80984 -25865 81030 -25028
rect 81397 -25183 81443 -25027
rect 81593 -25181 81639 -25027
rect 81495 -25183 81737 -25181
rect 81789 -25183 81835 -25027
rect 81397 -25229 82034 -25183
rect 81397 -25358 81443 -25258
rect 81495 -25358 81541 -25229
rect 81593 -25358 81639 -25258
rect 81691 -25358 81737 -25229
rect 82235 -25539 82281 -24939
rect 82446 -25539 82492 -24939
rect 82544 -25539 82590 -24939
rect 82642 -25539 82688 -24939
rect 82854 -25539 82900 -24939
rect 81082 -25901 81128 -25565
rect 83085 -25670 83190 -25598
rect 83091 -25753 83156 -25670
rect 82136 -25818 83156 -25753
rect 80689 -25948 81128 -25901
rect 82235 -26151 82281 -25851
rect 82333 -26151 82379 -25851
rect 82431 -26151 82477 -25851
rect 82673 -26151 82719 -25851
rect 82771 -26151 82817 -25851
rect 83378 -26259 83491 -24063
rect 84196 -24096 84326 -23946
rect 84482 -24000 84528 -23800
rect 84580 -24028 84626 -23800
rect 84678 -24000 84724 -23800
rect 84776 -24028 84822 -23800
rect 85013 -23946 85067 -23656
rect 85357 -23922 85403 -23623
rect 85455 -23922 85501 -23622
rect 85553 -23922 85599 -23586
rect 85013 -24000 85341 -23946
rect 84482 -24074 85119 -24028
rect 85287 -24055 85341 -24000
rect 84246 -25500 84300 -24096
rect 84482 -24330 84528 -24074
rect 84580 -24076 84822 -24074
rect 84678 -24330 84724 -24076
rect 84874 -24330 84920 -24074
rect 85261 -24113 85420 -24055
rect 85455 -24459 85501 -24159
rect 85651 -24459 85697 -23622
rect 85749 -23922 85795 -23586
rect 86451 -24094 87159 -23981
rect 86064 -24229 86110 -24129
rect 86162 -24258 86208 -24129
rect 86260 -24229 86306 -24129
rect 86358 -24258 86404 -24129
rect 86064 -24304 86701 -24258
rect 86064 -24460 86110 -24304
rect 86162 -24306 86404 -24304
rect 86260 -24460 86306 -24306
rect 86456 -24460 86502 -24304
rect 84456 -25359 84502 -25059
rect 84103 -25554 84300 -25500
rect 84358 -25895 84404 -25596
rect 84357 -25932 84404 -25895
rect 84456 -25896 84502 -25596
rect 84554 -25932 84600 -25596
rect 84652 -25896 84698 -25059
rect 85065 -25214 85111 -25058
rect 85261 -25212 85307 -25058
rect 85163 -25214 85405 -25212
rect 85457 -25214 85503 -25058
rect 85065 -25260 85702 -25214
rect 85065 -25389 85111 -25289
rect 85163 -25389 85209 -25260
rect 85261 -25389 85307 -25289
rect 85359 -25389 85405 -25260
rect 85903 -25570 85949 -24970
rect 86114 -25570 86160 -24970
rect 86212 -25570 86258 -24970
rect 86310 -25570 86356 -24970
rect 86522 -25570 86568 -24970
rect 84750 -25932 84796 -25596
rect 86753 -25701 86858 -25629
rect 86759 -25784 86824 -25701
rect 85804 -25849 86824 -25784
rect 84357 -25979 84796 -25932
rect 85903 -26182 85949 -25882
rect 86001 -26182 86047 -25882
rect 86099 -26182 86145 -25882
rect 86341 -26182 86387 -25882
rect 86439 -26182 86485 -25882
rect 73450 -26410 77795 -26328
rect 82814 -26290 83491 -26259
rect 87046 -26290 87159 -24094
rect 87412 -25654 87696 -15445
rect 87382 -25997 87741 -25654
rect 82814 -26372 87159 -26290
rect 82818 -26403 87159 -26372
rect 64301 -26458 68642 -26427
rect 73454 -26441 77795 -26410
rect 55547 -26524 59888 -26493
rect 46349 -26558 50690 -26527
rect 87916 -26943 88161 -3581
rect 41577 -27132 41894 -27049
rect 25877 -27313 34677 -27132
rect 41577 -27313 81327 -27132
rect 84040 -27188 88161 -26943
rect 41577 -27340 41894 -27313
rect 84612 -27482 84857 -27188
rect 25329 -27727 84857 -27482
rect 41534 -28232 41903 -27855
rect 42854 -28153 81327 -27868
rect 41543 -30020 41843 -28232
rect 24065 -30320 41843 -30020
rect 42854 -30563 43139 -28153
rect 23860 -30622 43139 -30563
rect 23597 -30743 43139 -30622
rect 23860 -30848 43139 -30743
rect 12773 -32036 88394 -31752
rect -26820 -34157 -26420 -34111
rect -26820 -34275 -26420 -34229
rect -26820 -34393 -26420 -34347
rect -26820 -34511 -26420 -34465
rect -26820 -34629 -26420 -34583
rect -26820 -34747 -26420 -34701
rect -15906 -34726 8502 -34536
rect -26820 -34865 -26420 -34819
rect -26820 -34983 -26420 -34937
rect -26820 -35101 -26420 -35055
rect -26820 -35219 -26420 -35173
rect -26820 -35337 -26420 -35291
rect -26820 -35455 -26420 -35409
rect -26820 -35573 -26420 -35527
rect -26820 -35691 -26420 -35645
rect -26820 -35809 -26420 -35763
rect -26820 -35927 -26420 -35881
rect -26820 -36045 -26420 -35999
rect -26820 -36163 -26420 -36117
rect -26820 -36281 -26420 -36235
rect -26820 -36399 -26420 -36353
rect -26820 -36517 -26420 -36471
rect -26820 -36635 -26420 -36589
rect -26820 -36753 -26420 -36707
rect -26820 -36871 -26420 -36825
rect -26820 -36989 -26420 -36943
rect -26820 -37107 -26420 -37061
rect -26820 -37225 -26420 -37179
rect -26820 -37343 -26420 -37297
rect -26820 -37461 -26420 -37415
rect -26820 -37579 -26420 -37533
rect -26820 -37697 -26420 -37651
rect -26820 -37933 -26420 -37887
rect -26820 -38169 -26420 -38123
rect -26820 -38405 -26420 -38359
rect -26820 -38641 -26420 -38595
rect -26820 -38877 -26420 -38831
rect -26820 -39113 -26420 -39067
rect -26820 -39349 -26420 -39303
rect -26157 -38037 -26083 -37922
rect -26157 -38083 -25612 -38037
rect -26157 -38273 -26083 -38083
rect -26157 -38319 -25612 -38273
rect -26157 -38509 -26083 -38319
rect -26157 -38555 -25612 -38509
rect -26157 -38745 -26083 -38555
rect -26157 -38791 -25612 -38745
rect -26157 -38981 -26083 -38791
rect -26157 -39027 -25612 -38981
rect -26157 -39217 -26083 -39027
rect -26157 -39263 -25612 -39217
rect -26157 -39453 -26083 -39263
rect -26157 -39499 -25612 -39453
rect -26820 -39585 -26420 -39539
rect -26820 -39696 -26285 -39657
rect -26157 -39689 -26083 -39499
rect -26157 -39696 -25612 -39689
rect -26820 -39703 -25612 -39696
rect -26331 -39735 -25612 -39703
rect -26331 -39742 -26083 -39735
rect -26820 -39821 -26420 -39775
rect -26331 -39893 -26285 -39742
rect -26157 -39867 -26083 -39742
rect -26820 -39939 -26285 -39893
rect -26820 -40057 -26420 -40011
rect -26331 -40129 -26285 -39939
rect -26820 -40175 -26285 -40129
rect -26820 -40293 -26420 -40247
rect -26331 -40365 -26285 -40175
rect -26820 -40411 -26285 -40365
rect -26157 -40055 -26083 -39928
rect -26157 -40101 -25612 -40055
rect -26157 -40291 -26083 -40101
rect -26157 -40337 -25612 -40291
rect -26820 -40529 -26420 -40483
rect -26157 -40527 -26083 -40337
rect -26157 -40573 -25612 -40527
rect -26820 -40647 -26297 -40601
rect -26343 -40678 -26297 -40647
rect -26157 -40678 -26083 -40573
rect -26820 -40765 -26420 -40719
rect -26343 -40724 -26083 -40678
rect -26343 -40837 -26297 -40724
rect -26820 -40883 -26297 -40837
rect -26157 -40763 -26083 -40724
rect -26157 -40809 -25612 -40763
rect -26157 -40938 -26083 -40809
rect -26820 -41001 -26420 -40955
rect -26157 -41073 -26083 -40999
rect -26820 -41119 -26083 -41073
rect -26157 -41129 -26083 -41119
rect -26157 -41175 -25612 -41129
rect -26820 -41237 -26420 -41191
rect -26157 -41365 -26083 -41175
rect -26157 -41411 -25612 -41365
rect -26157 -41416 -26083 -41411
rect -25977 -42856 -25639 -42789
rect -27809 -43047 -25639 -42856
rect -27809 -43351 -27257 -43047
rect -25977 -43127 -25639 -43047
rect -21948 -35975 -21902 -35775
rect -21752 -35975 -21706 -35775
rect -21556 -35975 -21510 -35775
rect -20818 -35975 -20772 -35775
rect -15906 -35815 -15716 -34726
rect -14349 -35188 -14303 -34988
rect -14153 -35188 -14107 -34988
rect -13957 -35188 -13911 -34988
rect -13727 -35241 -13670 -35006
rect -13512 -35188 -13466 -34988
rect -13316 -35188 -13270 -34988
rect -13120 -35188 -13074 -34988
rect -12901 -35103 -12855 -35003
rect -12803 -35103 -12757 -35003
rect -12705 -35103 -12659 -35003
rect -12607 -35103 -12561 -35003
rect -12509 -35103 -12463 -35003
rect -12411 -35103 -12365 -35003
rect -12313 -35103 -12267 -35003
rect -12215 -35103 -12169 -35003
rect -11649 -35188 -11603 -34988
rect -11453 -35188 -11407 -34988
rect -11257 -35188 -11211 -34988
rect -12898 -35241 -12729 -35231
rect -13727 -35298 -12729 -35241
rect -11027 -35241 -10970 -35006
rect -10812 -35188 -10766 -34988
rect -10616 -35188 -10570 -34988
rect -10420 -35188 -10374 -34988
rect -10201 -35103 -10155 -35003
rect -10103 -35103 -10057 -35003
rect -10005 -35103 -9959 -35003
rect -9907 -35103 -9861 -35003
rect -9809 -35103 -9763 -35003
rect -9711 -35103 -9665 -35003
rect -9613 -35103 -9567 -35003
rect -9515 -35103 -9469 -35003
rect -10198 -35241 -10029 -35231
rect -11886 -35263 -11826 -35257
rect -12121 -35284 -12080 -35283
rect -12898 -35305 -12729 -35298
rect -14447 -35468 -14401 -35368
rect -14349 -35468 -14303 -35368
rect -14251 -35468 -14205 -35368
rect -14153 -35468 -14107 -35368
rect -14055 -35468 -14009 -35368
rect -13957 -35468 -13911 -35368
rect -14213 -35691 -14076 -35631
rect -14561 -35749 -14501 -35702
rect -14823 -35813 -14501 -35749
rect -19949 -36197 -19903 -35897
rect -20356 -36252 -20219 -36235
rect -20384 -36293 -20219 -36252
rect -22046 -36682 -22000 -36382
rect -21948 -36682 -21902 -36382
rect -21850 -36682 -21804 -36382
rect -21736 -36683 -21690 -36383
rect -21638 -36683 -21592 -36383
rect -21540 -36683 -21494 -36383
rect -21427 -36683 -21381 -36383
rect -21329 -36683 -21283 -36383
rect -21231 -36683 -21185 -36383
rect -20916 -36683 -20870 -36483
rect -20818 -36599 -20772 -36483
rect -20818 -36634 -20459 -36599
rect -20818 -36683 -20772 -36634
rect -22674 -45488 -22613 -36921
rect -22743 -45489 -22613 -45488
rect -22743 -45522 -22612 -45489
rect -22742 -45607 -22612 -45522
rect -22560 -45616 -22496 -38393
rect -22562 -45788 -22496 -45616
rect -22583 -45789 -22496 -45788
rect -22415 -42864 -22355 -37962
rect -21891 -38106 -21845 -37806
rect -21989 -38642 -21943 -38343
rect -21990 -38679 -21943 -38642
rect -21891 -38643 -21845 -38343
rect -21793 -38679 -21747 -38343
rect -21695 -38643 -21649 -37806
rect -21282 -37961 -21236 -37805
rect -21086 -37959 -21040 -37805
rect -21184 -37961 -20942 -37959
rect -20890 -37961 -20844 -37805
rect -21282 -38007 -20645 -37961
rect -21282 -38136 -21236 -38036
rect -21184 -38136 -21138 -38007
rect -21086 -38136 -21040 -38036
rect -20988 -38136 -20942 -38007
rect -20494 -38168 -20459 -36634
rect -20384 -37003 -20348 -36293
rect -20386 -37135 -20333 -37003
rect -20047 -36733 -20001 -36434
rect -20048 -36770 -20001 -36733
rect -19949 -36734 -19903 -36434
rect -19851 -36770 -19805 -36434
rect -19753 -36734 -19707 -35897
rect -19340 -36052 -19294 -35896
rect -19144 -36050 -19098 -35896
rect -19242 -36052 -19000 -36050
rect -18948 -36052 -18902 -35896
rect -16287 -35928 -15610 -35815
rect -19340 -36098 -18703 -36052
rect -19340 -36227 -19294 -36127
rect -19242 -36227 -19196 -36098
rect -19144 -36227 -19098 -36127
rect -19046 -36227 -19000 -36098
rect -18620 -36123 -18474 -36065
rect -18620 -36149 -18539 -36123
rect -18932 -36184 -18539 -36149
rect -19655 -36770 -19609 -36434
rect -20048 -36817 -19609 -36770
rect -18932 -37254 -18897 -36184
rect -18412 -36286 -17973 -36239
rect -18412 -36323 -18365 -36286
rect -18411 -36622 -18365 -36323
rect -18313 -36622 -18267 -36322
rect -18215 -36622 -18169 -36286
rect -18666 -36718 -18469 -36664
rect -20428 -37289 -18897 -37254
rect -20428 -38037 -20393 -37289
rect -20118 -37911 -20072 -37711
rect -19922 -37911 -19876 -37711
rect -19726 -37911 -19680 -37711
rect -18988 -37911 -18942 -37711
rect -20428 -38083 -20344 -38037
rect -21597 -38679 -21551 -38343
rect -20713 -38402 -20655 -38265
rect -20499 -38305 -20441 -38168
rect -20402 -38174 -20344 -38083
rect -18523 -38122 -18469 -36718
rect -18313 -37159 -18267 -36859
rect -18117 -37159 -18071 -36322
rect -18019 -36622 -17973 -36286
rect -16866 -36336 -16820 -36036
rect -16768 -36336 -16722 -36036
rect -16670 -36336 -16624 -36036
rect -16428 -36336 -16382 -36036
rect -16330 -36336 -16284 -36036
rect -16965 -36434 -15945 -36369
rect -16010 -36517 -15945 -36434
rect -16016 -36589 -15911 -36517
rect -17704 -36929 -17658 -36829
rect -17606 -36958 -17560 -36829
rect -17508 -36929 -17462 -36829
rect -17410 -36958 -17364 -36829
rect -17704 -37004 -17067 -36958
rect -17704 -37160 -17658 -37004
rect -17606 -37006 -17364 -37004
rect -17508 -37160 -17462 -37006
rect -17312 -37160 -17266 -37004
rect -16866 -37248 -16820 -36648
rect -16655 -37248 -16609 -36648
rect -16557 -37248 -16511 -36648
rect -16459 -37248 -16413 -36648
rect -16247 -37248 -16201 -36648
rect -18573 -38272 -18443 -38122
rect -18287 -38144 -18241 -37888
rect -18091 -38142 -18045 -37888
rect -18189 -38144 -17947 -38142
rect -17895 -38144 -17849 -37888
rect -17314 -38059 -17268 -37759
rect -18287 -38190 -17650 -38144
rect -17508 -38163 -17349 -38105
rect -20216 -38618 -20170 -38318
rect -20118 -38618 -20072 -38318
rect -20020 -38618 -19974 -38318
rect -19906 -38619 -19860 -38319
rect -19808 -38619 -19762 -38319
rect -19710 -38619 -19664 -38319
rect -19597 -38619 -19551 -38319
rect -19499 -38619 -19453 -38319
rect -19401 -38619 -19355 -38319
rect -18287 -38418 -18241 -38218
rect -18189 -38418 -18143 -38190
rect -18091 -38418 -18045 -38218
rect -17993 -38418 -17947 -38190
rect -17482 -38218 -17428 -38163
rect -17756 -38272 -17428 -38218
rect -19086 -38619 -19040 -38419
rect -18988 -38619 -18942 -38419
rect -17756 -38562 -17702 -38272
rect -18799 -38616 -17702 -38562
rect -17412 -38595 -17366 -38296
rect -21990 -38726 -21551 -38679
rect -18787 -39330 -18547 -38616
rect -17413 -38632 -17366 -38595
rect -17314 -38596 -17268 -38296
rect -17216 -38632 -17170 -38296
rect -17118 -38596 -17072 -37759
rect -16705 -37914 -16659 -37758
rect -16509 -37912 -16463 -37758
rect -16607 -37914 -16365 -37912
rect -16313 -37914 -16267 -37758
rect -16705 -37960 -16068 -37914
rect -16705 -38089 -16659 -37989
rect -16607 -38089 -16561 -37960
rect -16509 -38089 -16463 -37989
rect -16411 -38089 -16365 -37960
rect -15723 -38124 -15610 -35928
rect -14823 -37729 -14759 -35813
rect -14561 -35839 -14501 -35813
rect -14198 -35909 -14103 -35691
rect -13788 -35809 -13728 -35342
rect -12216 -35344 -12079 -35284
rect -11886 -35323 -11743 -35263
rect -11027 -35298 -10029 -35241
rect -10198 -35305 -10029 -35298
rect -13610 -35468 -13564 -35368
rect -13512 -35468 -13466 -35368
rect -13414 -35468 -13368 -35368
rect -13316 -35468 -13270 -35368
rect -13218 -35468 -13172 -35368
rect -13120 -35468 -13074 -35368
rect -12901 -35518 -12855 -35418
rect -12803 -35518 -12757 -35418
rect -12705 -35518 -12659 -35418
rect -12607 -35518 -12561 -35418
rect -12509 -35518 -12463 -35418
rect -12411 -35518 -12365 -35418
rect -12313 -35518 -12267 -35418
rect -12215 -35518 -12169 -35418
rect -13824 -35869 -13692 -35809
rect -12121 -35829 -12080 -35344
rect -12051 -35780 -11914 -35720
rect -13611 -35877 -12080 -35829
rect -14222 -35969 -14090 -35909
rect -14447 -36126 -14401 -36026
rect -14349 -36126 -14303 -36026
rect -14251 -36126 -14205 -36026
rect -14153 -36126 -14107 -36026
rect -14055 -36126 -14009 -36026
rect -13957 -36126 -13911 -36026
rect -13611 -36031 -13563 -35877
rect -13609 -36076 -13563 -36031
rect -13511 -36076 -13465 -35976
rect -13419 -35995 -13358 -35877
rect -13413 -36076 -13367 -35995
rect -13315 -36076 -13269 -35976
rect -13223 -35997 -13162 -35877
rect -13217 -36076 -13171 -35997
rect -13119 -36076 -13073 -35976
rect -13032 -35995 -12971 -35877
rect -13021 -36076 -12975 -35995
rect -12923 -36076 -12877 -35976
rect -12704 -36126 -12658 -36026
rect -12606 -36126 -12560 -36026
rect -12508 -36126 -12462 -36026
rect -12410 -36126 -12364 -36026
rect -12312 -36126 -12266 -36026
rect -12214 -36126 -12168 -36026
rect -13049 -36196 -12880 -36189
rect -13049 -36253 -12051 -36196
rect -12002 -36228 -11942 -35780
rect -11886 -36071 -11826 -35323
rect -9527 -35346 -9373 -35286
rect -11747 -35468 -11701 -35368
rect -11649 -35468 -11603 -35368
rect -11551 -35468 -11505 -35368
rect -11453 -35468 -11407 -35368
rect -11355 -35468 -11309 -35368
rect -11257 -35468 -11211 -35368
rect -11616 -35697 -11479 -35637
rect -11605 -35905 -11510 -35697
rect -11076 -35721 -11016 -35357
rect -10910 -35468 -10864 -35368
rect -10812 -35468 -10766 -35368
rect -10714 -35468 -10668 -35368
rect -10616 -35468 -10570 -35368
rect -10518 -35468 -10472 -35368
rect -10420 -35468 -10374 -35368
rect -10201 -35518 -10155 -35418
rect -10103 -35518 -10057 -35418
rect -10005 -35518 -9959 -35418
rect -9907 -35518 -9861 -35418
rect -9809 -35518 -9763 -35418
rect -9711 -35518 -9665 -35418
rect -9613 -35518 -9567 -35418
rect -9515 -35518 -9469 -35418
rect -9419 -35621 -9373 -35346
rect -10192 -35666 -9373 -35621
rect -10192 -35667 -9381 -35666
rect -11105 -35781 -10973 -35721
rect -10192 -35833 -10146 -35667
rect -8978 -35697 -8846 -35637
rect -8961 -35762 -8866 -35697
rect -8426 -35762 -8331 -34726
rect -8183 -35598 -8137 -34998
rect -7971 -35598 -7925 -34998
rect -7873 -35598 -7827 -34998
rect -7775 -35598 -7729 -34998
rect -7564 -35598 -7518 -34998
rect -6753 -35394 -6707 -35194
rect -6655 -35394 -6609 -35194
rect -6557 -35394 -6511 -35194
rect -6437 -35394 -6391 -35194
rect -6339 -35394 -6293 -35194
rect -6241 -35394 -6195 -35194
rect -5879 -35394 -5833 -35194
rect -5683 -35394 -5637 -35194
rect -5373 -35394 -5327 -35194
rect -5064 -35394 -5018 -35194
rect -4253 -35394 -4207 -35194
rect -4155 -35394 -4109 -35194
rect -4057 -35394 -4011 -35194
rect -3937 -35394 -3891 -35194
rect -3839 -35394 -3793 -35194
rect -3741 -35394 -3695 -35194
rect -3379 -35394 -3333 -35194
rect -3183 -35394 -3137 -35194
rect -2873 -35394 -2827 -35194
rect -2564 -35394 -2518 -35194
rect -1753 -35394 -1707 -35194
rect -1655 -35394 -1609 -35194
rect -1557 -35394 -1511 -35194
rect -1437 -35394 -1391 -35194
rect -1339 -35394 -1293 -35194
rect -1241 -35394 -1195 -35194
rect -879 -35394 -833 -35194
rect -683 -35394 -637 -35194
rect -373 -35394 -327 -35194
rect -64 -35394 -18 -35194
rect 747 -35394 793 -35194
rect 845 -35394 891 -35194
rect 943 -35394 989 -35194
rect 1063 -35394 1109 -35194
rect 1161 -35394 1207 -35194
rect 1259 -35394 1305 -35194
rect 1621 -35394 1667 -35194
rect 1817 -35394 1863 -35194
rect 2127 -35394 2173 -35194
rect 2436 -35394 2482 -35194
rect 3247 -35394 3293 -35194
rect 3345 -35394 3391 -35194
rect 3443 -35394 3489 -35194
rect 3563 -35394 3609 -35194
rect 3661 -35394 3707 -35194
rect 3759 -35394 3805 -35194
rect 4121 -35394 4167 -35194
rect 4317 -35394 4363 -35194
rect 4627 -35394 4673 -35194
rect 4936 -35394 4982 -35194
rect 6247 -35394 6293 -35194
rect 6345 -35394 6391 -35194
rect 6443 -35394 6489 -35194
rect 6563 -35394 6609 -35194
rect 6661 -35394 6707 -35194
rect 6759 -35394 6805 -35194
rect 7121 -35394 7167 -35194
rect 7317 -35394 7363 -35194
rect 7627 -35394 7673 -35194
rect 7936 -35394 7982 -35194
rect -5590 -35522 -5451 -35504
rect -4975 -35522 -4836 -35510
rect -3090 -35522 -2951 -35504
rect -2475 -35522 -2336 -35510
rect -590 -35522 -451 -35504
rect 25 -35522 164 -35510
rect 1910 -35522 2049 -35504
rect 2525 -35522 2664 -35510
rect 4410 -35522 4549 -35504
rect 5025 -35522 5164 -35510
rect 7410 -35522 7549 -35504
rect 8025 -35522 8164 -35510
rect 8726 -35522 8926 -35170
rect -6748 -35561 -6609 -35548
rect -5590 -35550 -4685 -35522
rect -5590 -35558 -5451 -35550
rect -6748 -35589 -6394 -35561
rect -4975 -35564 -4836 -35550
rect -6748 -35602 -6609 -35589
rect -10906 -35879 -10146 -35833
rect -9301 -35867 -9169 -35807
rect -8961 -35857 -8331 -35762
rect -11623 -35965 -11486 -35905
rect -10906 -35976 -10860 -35879
rect -10711 -35976 -10669 -35879
rect -10516 -35976 -10474 -35879
rect -10320 -35976 -10278 -35879
rect -11887 -36116 -11826 -36071
rect -11887 -36203 -11827 -36116
rect -11747 -36126 -11701 -36026
rect -11649 -36126 -11603 -36026
rect -11551 -36126 -11505 -36026
rect -11453 -36126 -11407 -36026
rect -11355 -36126 -11309 -36026
rect -11257 -36126 -11211 -36026
rect -10909 -36076 -10860 -35976
rect -10811 -36076 -10765 -35976
rect -10713 -36076 -10667 -35976
rect -10615 -36076 -10569 -35976
rect -10517 -36076 -10471 -35976
rect -10419 -36076 -10373 -35976
rect -10321 -36076 -10275 -35976
rect -10223 -36076 -10177 -35976
rect -10004 -36126 -9958 -36026
rect -9906 -36126 -9860 -36026
rect -9808 -36126 -9762 -36026
rect -9710 -36126 -9664 -36026
rect -9612 -36126 -9566 -36026
rect -9514 -36126 -9468 -36026
rect -9268 -36095 -9210 -35867
rect -8961 -35906 -8866 -35857
rect -8996 -35966 -8859 -35906
rect -10349 -36196 -10180 -36189
rect -13049 -36263 -12880 -36253
rect -14447 -36506 -14401 -36306
rect -14251 -36506 -14205 -36306
rect -14055 -36506 -14009 -36306
rect -13609 -36459 -13563 -36391
rect -13609 -36491 -13558 -36459
rect -13511 -36491 -13465 -36391
rect -13413 -36434 -13367 -36391
rect -13608 -36574 -13558 -36491
rect -13417 -36574 -13366 -36434
rect -13315 -36491 -13269 -36391
rect -13217 -36453 -13171 -36391
rect -13217 -36574 -13166 -36453
rect -13119 -36491 -13073 -36391
rect -13021 -36453 -12975 -36391
rect -13023 -36574 -12972 -36453
rect -12923 -36491 -12877 -36391
rect -12704 -36506 -12658 -36306
rect -12508 -36506 -12462 -36306
rect -12312 -36506 -12266 -36306
rect -12108 -36488 -12051 -36253
rect -10349 -36253 -9351 -36196
rect -9270 -36227 -9210 -36095
rect -9122 -36126 -9076 -36026
rect -9024 -36126 -8978 -36026
rect -8926 -36126 -8880 -36026
rect -8828 -36126 -8782 -36026
rect -8730 -36126 -8684 -36026
rect -8632 -36126 -8586 -36026
rect -10349 -36263 -10180 -36253
rect -11747 -36506 -11701 -36306
rect -11551 -36506 -11505 -36306
rect -11355 -36506 -11309 -36306
rect -10909 -36491 -10863 -36391
rect -10811 -36491 -10765 -36391
rect -10713 -36491 -10667 -36391
rect -10615 -36491 -10569 -36391
rect -10517 -36491 -10471 -36391
rect -10419 -36491 -10373 -36391
rect -10321 -36491 -10275 -36391
rect -10223 -36491 -10177 -36391
rect -10004 -36506 -9958 -36306
rect -9808 -36506 -9762 -36306
rect -9612 -36506 -9566 -36306
rect -9408 -36574 -9351 -36253
rect -9122 -36506 -9076 -36306
rect -8926 -36506 -8880 -36306
rect -8730 -36506 -8684 -36306
rect -13608 -36631 -9351 -36574
rect -8426 -36791 -8331 -35857
rect -8100 -36210 -8054 -35910
rect -8002 -36210 -7956 -35910
rect -7760 -36210 -7714 -35910
rect -7662 -36210 -7616 -35910
rect -7564 -36210 -7518 -35910
rect -11298 -36904 -8330 -36791
rect -13423 -37262 -12984 -37215
rect -13423 -37299 -13376 -37262
rect -13422 -37598 -13376 -37299
rect -13324 -37598 -13278 -37298
rect -13226 -37598 -13180 -37262
rect -13961 -37729 -13775 -37687
rect -14823 -37793 -13775 -37729
rect -13961 -37841 -13775 -37793
rect -16318 -38237 -15610 -38124
rect -17020 -38632 -16974 -38296
rect -17413 -38679 -16974 -38632
rect -16401 -38988 -16133 -38723
rect -16352 -39543 -16164 -38988
rect -16396 -39808 -16128 -39543
rect -21826 -41600 -21780 -41000
rect -21614 -41600 -21568 -41000
rect -21516 -41600 -21470 -41000
rect -21418 -41600 -21372 -41000
rect -21305 -41600 -21259 -41000
rect -21207 -41600 -21161 -41000
rect -21109 -41600 -21063 -41000
rect -20620 -41329 -20574 -40929
rect -20409 -41329 -20363 -40929
rect -20311 -41329 -20265 -40929
rect -20213 -41329 -20167 -40929
rect -19715 -41330 -19669 -40930
rect -19504 -41330 -19458 -40930
rect -19406 -41330 -19360 -40930
rect -19308 -41330 -19262 -40930
rect -21088 -41926 -20951 -41868
rect -21826 -42164 -21780 -41964
rect -21728 -42164 -21682 -41964
rect -21630 -42164 -21584 -41964
rect -21532 -42164 -21486 -41964
rect -21960 -42410 -21156 -42260
rect -21948 -42822 -21861 -42410
rect -21768 -42822 -21681 -42410
rect -21595 -42822 -21508 -42410
rect -21411 -42822 -21324 -42410
rect -21286 -42822 -21199 -42410
rect -22173 -42864 -21190 -42822
rect -22415 -42924 -21190 -42864
rect -22583 -45912 -22460 -45789
rect -22415 -46156 -22355 -42924
rect -22173 -42937 -21190 -42924
rect -21076 -42924 -20986 -41926
rect -19976 -41492 -19918 -41355
rect -20817 -41529 -20759 -41525
rect -20818 -41662 -20759 -41529
rect -20201 -41577 -20064 -41519
rect -20818 -42479 -20775 -41662
rect -20620 -41821 -20574 -41621
rect -20522 -41821 -20476 -41621
rect -20424 -41821 -20378 -41621
rect -20819 -42616 -20761 -42479
rect -21076 -43014 -20759 -42924
rect -22163 -43310 -22117 -43110
rect -22065 -43310 -22019 -43110
rect -21750 -43410 -21704 -43110
rect -21652 -43410 -21606 -43110
rect -21554 -43410 -21508 -43110
rect -21441 -43410 -21395 -43110
rect -21343 -43410 -21297 -43110
rect -21245 -43410 -21199 -43110
rect -21131 -43411 -21085 -43111
rect -21033 -43411 -20987 -43111
rect -20935 -43411 -20889 -43111
rect -20849 -43602 -20759 -43014
rect -20110 -43547 -20075 -41577
rect -19976 -42558 -19941 -41492
rect -19899 -41664 -19841 -41527
rect -19270 -41578 -19133 -41520
rect -19998 -42695 -19940 -42558
rect -19899 -42635 -19864 -41664
rect -19715 -41822 -19669 -41622
rect -19617 -41822 -19571 -41622
rect -19519 -41822 -19473 -41622
rect -19905 -42772 -19847 -42635
rect -20118 -43684 -20060 -43547
rect -22163 -44018 -22117 -43818
rect -21425 -44018 -21379 -43818
rect -21229 -44018 -21183 -43818
rect -21033 -44018 -20987 -43818
rect -22162 -44289 -22119 -44018
rect -19185 -43633 -19150 -41578
rect -19009 -41876 -18892 -41753
rect -19108 -43281 -19050 -43144
rect -19193 -43770 -19135 -43633
rect -22212 -44405 -22054 -44289
rect -19107 -44317 -19068 -43281
rect -19006 -44140 -18914 -41876
rect -15723 -40815 -15610 -38237
rect -13324 -38135 -13278 -37835
rect -13128 -38135 -13082 -37298
rect -13030 -37598 -12984 -37262
rect -11877 -37312 -11831 -37012
rect -11779 -37312 -11733 -37012
rect -11681 -37312 -11635 -37012
rect -11439 -37312 -11393 -37012
rect -11341 -37312 -11295 -37012
rect -11976 -37410 -10956 -37345
rect -11021 -37493 -10956 -37410
rect -11027 -37565 -10922 -37493
rect -12715 -37905 -12669 -37805
rect -12617 -37934 -12571 -37805
rect -12519 -37905 -12473 -37805
rect -12421 -37934 -12375 -37805
rect -12715 -37980 -12078 -37934
rect -12715 -38136 -12669 -37980
rect -12617 -37982 -12375 -37980
rect -12519 -38136 -12473 -37982
rect -12323 -38136 -12277 -37980
rect -11877 -38224 -11831 -37624
rect -11666 -38224 -11620 -37624
rect -11568 -38224 -11522 -37624
rect -11470 -38224 -11424 -37624
rect -11258 -38224 -11212 -37624
rect -16287 -40928 -15610 -40815
rect -18412 -41286 -17973 -41239
rect -18412 -41323 -18365 -41286
rect -18411 -41622 -18365 -41323
rect -18313 -41622 -18267 -41322
rect -18215 -41622 -18169 -41286
rect -18666 -41718 -18469 -41664
rect -18523 -43122 -18469 -41718
rect -18313 -42159 -18267 -41859
rect -18117 -42159 -18071 -41322
rect -18019 -41622 -17973 -41286
rect -16866 -41336 -16820 -41036
rect -16768 -41336 -16722 -41036
rect -16670 -41336 -16624 -41036
rect -16428 -41336 -16382 -41036
rect -16330 -41336 -16284 -41036
rect -16965 -41434 -15945 -41369
rect -16010 -41517 -15945 -41434
rect -16016 -41589 -15911 -41517
rect -17704 -41929 -17658 -41829
rect -17606 -41958 -17560 -41829
rect -17508 -41929 -17462 -41829
rect -17410 -41958 -17364 -41829
rect -17704 -42004 -17067 -41958
rect -17704 -42160 -17658 -42004
rect -17606 -42006 -17364 -42004
rect -17508 -42160 -17462 -42006
rect -17312 -42160 -17266 -42004
rect -16866 -42248 -16820 -41648
rect -16655 -42248 -16609 -41648
rect -16557 -42248 -16511 -41648
rect -16459 -42248 -16413 -41648
rect -16247 -42248 -16201 -41648
rect -18573 -43272 -18443 -43122
rect -18287 -43144 -18241 -42888
rect -18091 -43142 -18045 -42888
rect -18189 -43144 -17947 -43142
rect -17895 -43144 -17849 -42888
rect -17314 -43059 -17268 -42759
rect -18287 -43190 -17650 -43144
rect -17508 -43163 -17349 -43105
rect -18287 -43418 -18241 -43218
rect -18189 -43418 -18143 -43190
rect -18091 -43418 -18045 -43218
rect -17993 -43418 -17947 -43190
rect -17482 -43218 -17428 -43163
rect -17756 -43272 -17428 -43218
rect -17756 -43562 -17702 -43272
rect -18799 -43616 -17702 -43562
rect -17412 -43595 -17366 -43296
rect -18799 -43886 -18745 -43616
rect -17413 -43632 -17366 -43595
rect -17314 -43596 -17268 -43296
rect -17216 -43632 -17170 -43296
rect -17118 -43596 -17072 -42759
rect -16705 -42914 -16659 -42758
rect -16509 -42912 -16463 -42758
rect -16607 -42914 -16365 -42912
rect -16313 -42914 -16267 -42758
rect -16705 -42960 -16068 -42914
rect -16705 -43089 -16659 -42989
rect -16607 -43089 -16561 -42960
rect -16509 -43089 -16463 -42989
rect -16411 -43089 -16365 -42960
rect -15723 -43124 -15610 -40928
rect -15457 -41520 -15249 -39124
rect -16318 -43237 -15610 -43124
rect -17020 -43632 -16974 -43296
rect -17413 -43679 -16974 -43632
rect -18829 -44022 -18685 -43886
rect -19006 -44277 -18868 -44140
rect -19144 -44375 -19007 -44317
rect -13298 -39120 -13252 -38864
rect -13102 -39118 -13056 -38864
rect -13200 -39120 -12958 -39118
rect -12906 -39120 -12860 -38864
rect -12325 -39035 -12279 -38735
rect -13298 -39166 -12661 -39120
rect -12519 -39139 -12360 -39081
rect -13298 -39394 -13252 -39194
rect -13200 -39394 -13154 -39166
rect -13102 -39394 -13056 -39194
rect -13004 -39394 -12958 -39166
rect -12493 -39194 -12439 -39139
rect -12767 -39248 -12439 -39194
rect -12767 -39538 -12713 -39248
rect -14881 -39592 -12713 -39538
rect -12423 -39571 -12377 -39272
rect -14881 -40676 -14827 -39592
rect -12424 -39608 -12377 -39571
rect -12325 -39572 -12279 -39272
rect -12227 -39608 -12181 -39272
rect -12129 -39572 -12083 -38735
rect -11716 -38890 -11670 -38734
rect -11520 -38888 -11474 -38734
rect -11618 -38890 -11376 -38888
rect -11324 -38890 -11278 -38734
rect -11716 -38936 -11079 -38890
rect -11716 -39065 -11670 -38965
rect -11618 -39065 -11572 -38936
rect -11520 -39065 -11474 -38965
rect -11422 -39065 -11376 -38936
rect -10734 -39100 -10621 -36904
rect -11329 -39213 -10621 -39100
rect -12031 -39608 -11985 -39272
rect -12424 -39655 -11985 -39608
rect -14349 -40115 -14303 -39915
rect -14153 -40115 -14107 -39915
rect -13957 -40115 -13911 -39915
rect -13727 -40168 -13670 -39933
rect -13512 -40115 -13466 -39915
rect -13316 -40115 -13270 -39915
rect -13120 -40115 -13074 -39915
rect -12901 -40030 -12855 -39930
rect -12803 -40030 -12757 -39930
rect -12705 -40030 -12659 -39930
rect -12607 -40030 -12561 -39930
rect -12509 -40030 -12463 -39930
rect -12411 -40030 -12365 -39930
rect -12313 -40030 -12267 -39930
rect -12215 -40030 -12169 -39930
rect -11649 -40115 -11603 -39915
rect -11453 -40115 -11407 -39915
rect -11257 -40115 -11211 -39915
rect -12898 -40168 -12729 -40158
rect -13727 -40225 -12729 -40168
rect -11027 -40168 -10970 -39933
rect -10812 -40115 -10766 -39915
rect -10616 -40115 -10570 -39915
rect -10420 -40115 -10374 -39915
rect -10201 -40030 -10155 -39930
rect -10103 -40030 -10057 -39930
rect -10005 -40030 -9959 -39930
rect -9907 -40030 -9861 -39930
rect -9809 -40030 -9763 -39930
rect -9711 -40030 -9665 -39930
rect -9613 -40030 -9567 -39930
rect -9515 -40030 -9469 -39930
rect -10198 -40168 -10029 -40158
rect -11886 -40190 -11826 -40184
rect -12121 -40211 -12080 -40210
rect -12898 -40232 -12729 -40225
rect -14447 -40395 -14401 -40295
rect -14349 -40395 -14303 -40295
rect -14251 -40395 -14205 -40295
rect -14153 -40395 -14107 -40295
rect -14055 -40395 -14009 -40295
rect -13957 -40395 -13911 -40295
rect -14213 -40618 -14076 -40558
rect -14561 -40676 -14501 -40629
rect -14881 -40740 -14501 -40676
rect -14561 -40766 -14501 -40740
rect -14198 -40836 -14103 -40618
rect -13788 -40736 -13728 -40269
rect -12216 -40271 -12079 -40211
rect -11886 -40250 -11743 -40190
rect -11027 -40225 -10029 -40168
rect -10198 -40232 -10029 -40225
rect -13610 -40395 -13564 -40295
rect -13512 -40395 -13466 -40295
rect -13414 -40395 -13368 -40295
rect -13316 -40395 -13270 -40295
rect -13218 -40395 -13172 -40295
rect -13120 -40395 -13074 -40295
rect -12901 -40445 -12855 -40345
rect -12803 -40445 -12757 -40345
rect -12705 -40445 -12659 -40345
rect -12607 -40445 -12561 -40345
rect -12509 -40445 -12463 -40345
rect -12411 -40445 -12365 -40345
rect -12313 -40445 -12267 -40345
rect -12215 -40445 -12169 -40345
rect -13824 -40796 -13692 -40736
rect -12121 -40756 -12080 -40271
rect -12051 -40707 -11914 -40647
rect -13611 -40804 -12080 -40756
rect -14222 -40896 -14090 -40836
rect -14447 -41053 -14401 -40953
rect -14349 -41053 -14303 -40953
rect -14251 -41053 -14205 -40953
rect -14153 -41053 -14107 -40953
rect -14055 -41053 -14009 -40953
rect -13957 -41053 -13911 -40953
rect -13611 -40958 -13563 -40804
rect -13609 -41003 -13563 -40958
rect -13511 -41003 -13465 -40903
rect -13419 -40922 -13358 -40804
rect -13413 -41003 -13367 -40922
rect -13315 -41003 -13269 -40903
rect -13223 -40924 -13162 -40804
rect -13217 -41003 -13171 -40924
rect -13119 -41003 -13073 -40903
rect -13032 -40922 -12971 -40804
rect -13021 -41003 -12975 -40922
rect -12923 -41003 -12877 -40903
rect -12704 -41053 -12658 -40953
rect -12606 -41053 -12560 -40953
rect -12508 -41053 -12462 -40953
rect -12410 -41053 -12364 -40953
rect -12312 -41053 -12266 -40953
rect -12214 -41053 -12168 -40953
rect -13049 -41123 -12880 -41116
rect -13049 -41180 -12051 -41123
rect -12002 -41155 -11942 -40707
rect -11886 -40998 -11826 -40250
rect -9527 -40273 -9373 -40213
rect -11747 -40395 -11701 -40295
rect -11649 -40395 -11603 -40295
rect -11551 -40395 -11505 -40295
rect -11453 -40395 -11407 -40295
rect -11355 -40395 -11309 -40295
rect -11257 -40395 -11211 -40295
rect -11616 -40624 -11479 -40564
rect -11605 -40832 -11510 -40624
rect -11076 -40648 -11016 -40284
rect -10910 -40395 -10864 -40295
rect -10812 -40395 -10766 -40295
rect -10714 -40395 -10668 -40295
rect -10616 -40395 -10570 -40295
rect -10518 -40395 -10472 -40295
rect -10420 -40395 -10374 -40295
rect -10201 -40445 -10155 -40345
rect -10103 -40445 -10057 -40345
rect -10005 -40445 -9959 -40345
rect -9907 -40445 -9861 -40345
rect -9809 -40445 -9763 -40345
rect -9711 -40445 -9665 -40345
rect -9613 -40445 -9567 -40345
rect -9515 -40445 -9469 -40345
rect -9419 -40548 -9373 -40273
rect -10192 -40593 -9373 -40548
rect -8961 -40564 -8866 -36904
rect -10192 -40594 -9381 -40593
rect -11105 -40708 -10973 -40648
rect -10192 -40760 -10146 -40594
rect -8978 -40624 -8846 -40564
rect -10906 -40806 -10146 -40760
rect -9301 -40794 -9169 -40734
rect -11623 -40892 -11486 -40832
rect -10906 -40903 -10860 -40806
rect -10711 -40903 -10669 -40806
rect -10516 -40903 -10474 -40806
rect -10320 -40903 -10278 -40806
rect -11887 -41043 -11826 -40998
rect -11887 -41130 -11827 -41043
rect -11747 -41053 -11701 -40953
rect -11649 -41053 -11603 -40953
rect -11551 -41053 -11505 -40953
rect -11453 -41053 -11407 -40953
rect -11355 -41053 -11309 -40953
rect -11257 -41053 -11211 -40953
rect -10909 -41003 -10860 -40903
rect -10811 -41003 -10765 -40903
rect -10713 -41003 -10667 -40903
rect -10615 -41003 -10569 -40903
rect -10517 -41003 -10471 -40903
rect -10419 -41003 -10373 -40903
rect -10321 -41003 -10275 -40903
rect -10223 -41003 -10177 -40903
rect -10004 -41053 -9958 -40953
rect -9906 -41053 -9860 -40953
rect -9808 -41053 -9762 -40953
rect -9710 -41053 -9664 -40953
rect -9612 -41053 -9566 -40953
rect -9514 -41053 -9468 -40953
rect -9268 -41022 -9210 -40794
rect -8961 -40833 -8866 -40624
rect -8996 -40893 -8859 -40833
rect -10349 -41123 -10180 -41116
rect -13049 -41190 -12880 -41180
rect -14447 -41433 -14401 -41233
rect -14251 -41433 -14205 -41233
rect -14055 -41433 -14009 -41233
rect -13609 -41386 -13563 -41318
rect -13609 -41418 -13558 -41386
rect -13511 -41418 -13465 -41318
rect -13413 -41361 -13367 -41318
rect -13608 -41501 -13558 -41418
rect -13417 -41501 -13366 -41361
rect -13315 -41418 -13269 -41318
rect -13217 -41380 -13171 -41318
rect -13217 -41501 -13166 -41380
rect -13119 -41418 -13073 -41318
rect -13021 -41380 -12975 -41318
rect -13023 -41501 -12972 -41380
rect -12923 -41418 -12877 -41318
rect -12704 -41433 -12658 -41233
rect -12508 -41433 -12462 -41233
rect -12312 -41433 -12266 -41233
rect -12108 -41415 -12051 -41180
rect -10349 -41180 -9351 -41123
rect -9270 -41154 -9210 -41022
rect -9122 -41053 -9076 -40953
rect -9024 -41053 -8978 -40953
rect -8926 -41053 -8880 -40953
rect -8828 -41053 -8782 -40953
rect -8730 -41053 -8684 -40953
rect -8632 -41053 -8586 -40953
rect -10349 -41190 -10180 -41180
rect -11747 -41433 -11701 -41233
rect -11551 -41433 -11505 -41233
rect -11355 -41433 -11309 -41233
rect -10909 -41418 -10863 -41318
rect -10811 -41418 -10765 -41318
rect -10713 -41418 -10667 -41318
rect -10615 -41418 -10569 -41318
rect -10517 -41418 -10471 -41318
rect -10419 -41418 -10373 -41318
rect -10321 -41418 -10275 -41318
rect -10223 -41418 -10177 -41318
rect -10004 -41433 -9958 -41233
rect -9808 -41433 -9762 -41233
rect -9612 -41433 -9566 -41233
rect -9408 -41501 -9351 -41180
rect -9122 -41433 -9076 -41233
rect -8926 -41433 -8880 -41233
rect -8730 -41433 -8684 -41233
rect -13608 -41558 -9351 -41501
rect -8435 -43862 -8259 -37347
rect -8156 -40532 -8110 -39932
rect -7944 -40532 -7898 -39932
rect -7846 -40532 -7800 -39932
rect -7748 -40532 -7702 -39932
rect -7537 -40532 -7491 -39932
rect -8073 -41144 -8027 -40844
rect -7975 -41144 -7929 -40844
rect -7733 -41144 -7687 -40844
rect -7635 -41144 -7589 -40844
rect -7537 -41144 -7491 -40844
rect -8448 -44033 -8248 -43862
rect -7300 -44120 -7168 -35648
rect -6422 -35734 -6394 -35589
rect -5999 -35587 -5860 -35578
rect -5162 -35587 -5026 -35578
rect -5999 -35615 -5026 -35587
rect -5999 -35632 -5860 -35615
rect -5162 -35624 -5026 -35615
rect -6366 -35661 -6227 -35652
rect -5288 -35659 -5149 -35658
rect -5288 -35661 -4757 -35659
rect -6366 -35687 -4757 -35661
rect -6366 -35689 -5149 -35687
rect -6366 -35706 -6227 -35689
rect -5288 -35712 -5149 -35689
rect -5468 -35734 -5337 -35722
rect -6422 -35762 -5337 -35734
rect -5468 -35768 -5337 -35762
rect -6753 -36000 -6707 -35800
rect -6655 -36000 -6609 -35800
rect -6339 -36000 -6293 -35800
rect -6241 -36000 -6195 -35800
rect -5977 -36000 -5931 -35800
rect -5879 -36000 -5833 -35800
rect -5683 -36000 -5637 -35800
rect -5585 -36000 -5539 -35800
rect -5373 -36000 -5327 -35800
rect -5275 -36000 -5229 -35800
rect -5064 -36000 -5018 -35800
rect -4966 -36000 -4920 -35800
rect -6316 -36343 -6270 -36243
rect -6218 -36343 -6172 -36243
rect -6120 -36343 -6074 -36243
rect -6022 -36343 -5976 -36243
rect -5924 -36343 -5878 -36243
rect -5826 -36343 -5780 -36243
rect -4785 -36326 -4757 -35687
rect -4803 -36462 -4757 -36326
rect -6218 -36723 -6172 -36523
rect -6022 -36723 -5976 -36523
rect -5826 -36723 -5780 -36523
rect -4713 -36758 -4685 -35550
rect -4248 -35561 -4109 -35548
rect -3090 -35550 -2114 -35522
rect -3090 -35558 -2951 -35550
rect -4248 -35589 -3894 -35561
rect -2475 -35564 -2336 -35550
rect -4248 -35602 -4109 -35589
rect -3922 -35734 -3894 -35589
rect -3499 -35587 -3360 -35578
rect -2662 -35587 -2526 -35578
rect -3499 -35615 -2526 -35587
rect -3499 -35632 -3360 -35615
rect -2662 -35624 -2526 -35615
rect -3866 -35661 -3727 -35652
rect -2788 -35659 -2649 -35658
rect -2788 -35661 -2200 -35659
rect -3866 -35687 -2200 -35661
rect -3866 -35689 -2649 -35687
rect -3866 -35706 -3727 -35689
rect -2788 -35712 -2649 -35689
rect -2968 -35734 -2837 -35722
rect -3922 -35762 -2837 -35734
rect -2968 -35768 -2837 -35762
rect -4421 -35967 -4375 -35831
rect -4420 -36537 -4376 -35967
rect -4253 -36000 -4207 -35800
rect -4155 -36000 -4109 -35800
rect -3839 -36000 -3793 -35800
rect -3741 -36000 -3695 -35800
rect -3477 -36000 -3431 -35800
rect -3379 -36000 -3333 -35800
rect -3183 -36000 -3137 -35800
rect -3085 -36000 -3039 -35800
rect -2873 -36000 -2827 -35800
rect -2775 -36000 -2729 -35800
rect -2564 -36000 -2518 -35800
rect -2466 -36000 -2420 -35800
rect -4421 -36673 -4375 -36537
rect -2228 -36691 -2200 -35687
rect -2142 -36608 -2114 -35550
rect -1748 -35561 -1609 -35548
rect -590 -35550 358 -35522
rect -590 -35558 -451 -35550
rect -1748 -35589 -1394 -35561
rect 25 -35564 164 -35550
rect -1748 -35602 -1609 -35589
rect -1422 -35734 -1394 -35589
rect -999 -35587 -860 -35578
rect -162 -35587 -26 -35578
rect -999 -35615 -26 -35587
rect -999 -35632 -860 -35615
rect -162 -35624 -26 -35615
rect -1366 -35661 -1227 -35652
rect -288 -35659 -149 -35658
rect -288 -35661 284 -35659
rect -1366 -35687 284 -35661
rect -1366 -35689 -149 -35687
rect -1366 -35706 -1227 -35689
rect -288 -35712 -149 -35689
rect -468 -35734 -337 -35722
rect -1422 -35762 -337 -35734
rect -468 -35768 -337 -35762
rect -1873 -35971 -1827 -35835
rect -1872 -36208 -1828 -35971
rect -1753 -36000 -1707 -35800
rect -1655 -36000 -1609 -35800
rect -1339 -36000 -1293 -35800
rect -1241 -36000 -1195 -35800
rect -977 -36000 -931 -35800
rect -879 -36000 -833 -35800
rect -683 -36000 -637 -35800
rect -585 -36000 -539 -35800
rect -373 -36000 -327 -35800
rect -275 -36000 -229 -35800
rect -64 -36000 -18 -35800
rect 34 -36000 80 -35800
rect -1708 -36208 -1572 -36207
rect -1873 -36252 -1572 -36208
rect -1708 -36253 -1572 -36252
rect 256 -36552 284 -35687
rect 330 -36495 358 -35550
rect 752 -35561 891 -35548
rect 1910 -35550 2833 -35522
rect 1910 -35558 2049 -35550
rect 752 -35589 1106 -35561
rect 2525 -35564 2664 -35550
rect 752 -35602 891 -35589
rect 1078 -35734 1106 -35589
rect 1501 -35587 1640 -35578
rect 2338 -35587 2474 -35578
rect 1501 -35615 2474 -35587
rect 1501 -35632 1640 -35615
rect 2338 -35624 2474 -35615
rect 1134 -35661 1273 -35652
rect 2212 -35659 2351 -35658
rect 2212 -35661 2750 -35659
rect 1134 -35687 2750 -35661
rect 1134 -35689 2351 -35687
rect 1134 -35706 1273 -35689
rect 2212 -35712 2351 -35689
rect 2032 -35734 2163 -35722
rect 1078 -35762 2163 -35734
rect 2032 -35768 2163 -35762
rect 607 -35971 653 -35835
rect 608 -36221 652 -35971
rect 747 -36000 793 -35800
rect 845 -36000 891 -35800
rect 1161 -36000 1207 -35800
rect 1259 -36000 1305 -35800
rect 1523 -36000 1569 -35800
rect 1621 -36000 1667 -35800
rect 1817 -36000 1863 -35800
rect 1915 -36000 1961 -35800
rect 2127 -36000 2173 -35800
rect 2225 -36000 2271 -35800
rect 2436 -36000 2482 -35800
rect 2534 -36000 2580 -35800
rect 789 -36221 925 -36220
rect 608 -36265 925 -36221
rect 789 -36266 925 -36265
rect 2722 -36432 2750 -35687
rect 2805 -36358 2833 -35550
rect 3252 -35561 3391 -35548
rect 4410 -35550 6138 -35522
rect 4410 -35558 4549 -35550
rect 3252 -35589 3606 -35561
rect 5025 -35564 5164 -35550
rect 3252 -35602 3391 -35589
rect 3578 -35734 3606 -35589
rect 4001 -35587 4140 -35578
rect 4838 -35587 4974 -35578
rect 4001 -35615 4974 -35587
rect 4001 -35632 4140 -35615
rect 4838 -35624 4974 -35615
rect 4532 -35734 4663 -35722
rect 3578 -35762 4663 -35734
rect 4532 -35768 4663 -35762
rect 3024 -35971 3070 -35835
rect 3025 -36283 3069 -35971
rect 3247 -36000 3293 -35800
rect 3345 -36000 3391 -35800
rect 3661 -36000 3707 -35800
rect 3759 -36000 3805 -35800
rect 4023 -36000 4069 -35800
rect 4121 -36000 4167 -35800
rect 4317 -36000 4363 -35800
rect 4415 -36000 4461 -35800
rect 4627 -36000 4673 -35800
rect 4725 -36000 4771 -35800
rect 4936 -36000 4982 -35800
rect 5034 -36000 5080 -35800
rect 5929 -35971 5975 -35835
rect 5930 -36267 5974 -35971
rect 2972 -36329 3108 -36283
rect 5877 -36313 6013 -36267
rect 6110 -36225 6138 -35550
rect 6252 -35561 6391 -35548
rect 7410 -35550 10295 -35522
rect 7410 -35558 7549 -35550
rect 6252 -35589 6606 -35561
rect 8025 -35564 8164 -35550
rect 6252 -35602 6391 -35589
rect 6578 -35734 6606 -35589
rect 7001 -35587 7140 -35578
rect 7838 -35587 7974 -35578
rect 7001 -35615 7974 -35587
rect 7001 -35632 7140 -35615
rect 7838 -35624 7974 -35615
rect 7532 -35734 7663 -35722
rect 6578 -35762 7663 -35734
rect 7532 -35768 7663 -35762
rect 6247 -36000 6293 -35800
rect 6345 -36000 6391 -35800
rect 6661 -36000 6707 -35800
rect 6759 -36000 6805 -35800
rect 7023 -36000 7069 -35800
rect 7121 -36000 7167 -35800
rect 7317 -36000 7363 -35800
rect 7415 -36000 7461 -35800
rect 7627 -36000 7673 -35800
rect 7725 -36000 7771 -35800
rect 7936 -36000 7982 -35800
rect 8034 -36000 8080 -35800
rect 8938 -36225 10130 -36108
rect 6110 -36253 10139 -36225
rect 2805 -36396 9986 -36358
rect 2722 -36460 9911 -36432
rect 330 -36523 9834 -36495
rect 256 -36580 9749 -36552
rect -2142 -36659 9675 -36608
rect -2228 -36727 9590 -36691
rect -4713 -36809 9519 -36758
rect -4418 -36928 -4282 -36926
rect 2631 -36928 2767 -36924
rect -4418 -36970 2767 -36928
rect -4418 -36972 -4282 -36970
rect -6898 -37010 -6762 -37008
rect 2527 -37010 2682 -37008
rect -6898 -37052 2682 -37010
rect -6898 -37054 -6762 -37052
rect 2527 -37054 2682 -37052
rect -6573 -37626 -6527 -37426
rect -6377 -37626 -6331 -37426
rect -6181 -37626 -6135 -37426
rect -5735 -37541 -5689 -37441
rect -5637 -37541 -5591 -37441
rect -5539 -37541 -5493 -37441
rect -5441 -37541 -5395 -37441
rect -5343 -37541 -5297 -37441
rect -5245 -37541 -5199 -37441
rect -5147 -37541 -5101 -37441
rect -5049 -37541 -5003 -37441
rect -4830 -37626 -4784 -37426
rect -4634 -37626 -4588 -37426
rect -4438 -37626 -4392 -37426
rect -5175 -37679 -5006 -37669
rect -4234 -37679 -4177 -37444
rect -3873 -37626 -3827 -37426
rect -3677 -37626 -3631 -37426
rect -3481 -37626 -3435 -37426
rect -3035 -37541 -2989 -37441
rect -2937 -37541 -2891 -37441
rect -2839 -37541 -2793 -37441
rect -2741 -37541 -2695 -37441
rect -2643 -37541 -2597 -37441
rect -2545 -37541 -2499 -37441
rect -2447 -37541 -2401 -37441
rect -2349 -37541 -2303 -37441
rect -2130 -37626 -2084 -37426
rect -1934 -37626 -1888 -37426
rect -1738 -37626 -1692 -37426
rect -5175 -37736 -4177 -37679
rect -2475 -37679 -2306 -37669
rect -1534 -37679 -1477 -37444
rect -1248 -37626 -1202 -37426
rect -1052 -37626 -1006 -37426
rect -856 -37626 -810 -37426
rect -318 -37643 -272 -37443
rect 420 -37643 466 -37443
rect 616 -37643 662 -37443
rect 812 -37643 858 -37443
rect 1038 -37604 1084 -37602
rect -5175 -37743 -5006 -37736
rect -6573 -37906 -6527 -37806
rect -6475 -37906 -6429 -37806
rect -6377 -37906 -6331 -37806
rect -6279 -37906 -6233 -37806
rect -6181 -37906 -6135 -37806
rect -6083 -37906 -6037 -37806
rect -5735 -37901 -5689 -37856
rect -6348 -38023 -6216 -37963
rect -6687 -38119 -6627 -38093
rect -7042 -38182 -6627 -38119
rect -7025 -38183 -6627 -38182
rect -6687 -38230 -6627 -38183
rect -6324 -38241 -6229 -38023
rect -5737 -38055 -5689 -37901
rect -5637 -37956 -5591 -37856
rect -5539 -37937 -5493 -37856
rect -5545 -38055 -5484 -37937
rect -5441 -37956 -5395 -37856
rect -5343 -37935 -5297 -37856
rect -5349 -38055 -5288 -37935
rect -5245 -37956 -5199 -37856
rect -5147 -37937 -5101 -37856
rect -5158 -38055 -5097 -37937
rect -5049 -37956 -5003 -37856
rect -4830 -37906 -4784 -37806
rect -4732 -37906 -4686 -37806
rect -4634 -37906 -4588 -37806
rect -4536 -37906 -4490 -37806
rect -4438 -37906 -4392 -37806
rect -4340 -37906 -4294 -37806
rect -5737 -38103 -4206 -38055
rect -6339 -38301 -6202 -38241
rect -6573 -38564 -6527 -38464
rect -6475 -38564 -6429 -38464
rect -6377 -38564 -6331 -38464
rect -6279 -38564 -6233 -38464
rect -6181 -38564 -6135 -38464
rect -6083 -38564 -6037 -38464
rect -5736 -38564 -5690 -38464
rect -5638 -38564 -5592 -38464
rect -5540 -38564 -5494 -38464
rect -5442 -38564 -5396 -38464
rect -5344 -38564 -5298 -38464
rect -5246 -38564 -5200 -38464
rect -5027 -38514 -4981 -38414
rect -4929 -38514 -4883 -38414
rect -4831 -38514 -4785 -38414
rect -4733 -38514 -4687 -38414
rect -4635 -38514 -4589 -38414
rect -4537 -38514 -4491 -38414
rect -4439 -38514 -4393 -38414
rect -4341 -38514 -4295 -38414
rect -4247 -38588 -4206 -38103
rect -4128 -38152 -4068 -37704
rect -4013 -37816 -3953 -37729
rect -2475 -37736 -1477 -37679
rect -2475 -37743 -2306 -37736
rect -4013 -37861 -3952 -37816
rect -4177 -38212 -4040 -38152
rect -5024 -38634 -4855 -38627
rect -5853 -38691 -4855 -38634
rect -4342 -38648 -4205 -38588
rect -4012 -38609 -3952 -37861
rect -3873 -37906 -3827 -37806
rect -3775 -37906 -3729 -37806
rect -3677 -37906 -3631 -37806
rect -3579 -37906 -3533 -37806
rect -3481 -37906 -3435 -37806
rect -3383 -37906 -3337 -37806
rect -3035 -37956 -2986 -37856
rect -2937 -37956 -2891 -37856
rect -2839 -37956 -2793 -37856
rect -2741 -37956 -2695 -37856
rect -2643 -37956 -2597 -37856
rect -2545 -37956 -2499 -37856
rect -2447 -37956 -2401 -37856
rect -2349 -37956 -2303 -37856
rect -2130 -37906 -2084 -37806
rect -2032 -37906 -1986 -37806
rect -1934 -37906 -1888 -37806
rect -1836 -37906 -1790 -37806
rect -1738 -37906 -1692 -37806
rect -1640 -37906 -1594 -37806
rect -3749 -38027 -3612 -37967
rect -3731 -38235 -3636 -38027
rect -3032 -38053 -2986 -37956
rect -2837 -38053 -2795 -37956
rect -2642 -38053 -2600 -37956
rect -2446 -38053 -2404 -37956
rect -3032 -38099 -2272 -38053
rect -3231 -38211 -3099 -38151
rect -3742 -38295 -3605 -38235
rect -3873 -38564 -3827 -38464
rect -3775 -38564 -3729 -38464
rect -3677 -38564 -3631 -38464
rect -3579 -38564 -3533 -38464
rect -3481 -38564 -3435 -38464
rect -3383 -38564 -3337 -38464
rect -3202 -38575 -3142 -38211
rect -2318 -38265 -2272 -38099
rect -1534 -38173 -1477 -37736
rect -1396 -37837 -1336 -37705
rect 1030 -37738 1084 -37604
rect 1415 -37612 1461 -37456
rect 1611 -37610 1657 -37456
rect 1513 -37612 1755 -37610
rect 1807 -37612 1853 -37456
rect 1390 -37658 1853 -37612
rect -1394 -38065 -1336 -37837
rect -1248 -37906 -1202 -37806
rect -1150 -37906 -1104 -37806
rect -1052 -37906 -1006 -37806
rect -954 -37906 -908 -37806
rect -856 -37906 -810 -37806
rect -758 -37906 -712 -37806
rect -463 -37902 -322 -37849
rect -992 -38026 -855 -37966
rect -1394 -38123 -1155 -38065
rect -1213 -38152 -1155 -38123
rect -1534 -38230 -1268 -38173
rect -1217 -38212 -1085 -38152
rect -2318 -38266 -1507 -38265
rect -2318 -38311 -1499 -38266
rect -3036 -38564 -2990 -38464
rect -2938 -38564 -2892 -38464
rect -2840 -38564 -2794 -38464
rect -2742 -38564 -2696 -38464
rect -2644 -38564 -2598 -38464
rect -2546 -38564 -2500 -38464
rect -2327 -38514 -2281 -38414
rect -2229 -38514 -2183 -38414
rect -2131 -38514 -2085 -38414
rect -2033 -38514 -1987 -38414
rect -1935 -38514 -1889 -38414
rect -1837 -38514 -1791 -38414
rect -1739 -38514 -1693 -38414
rect -1641 -38514 -1595 -38414
rect -1545 -38586 -1499 -38311
rect -1325 -38351 -1268 -38230
rect -957 -38235 -862 -38026
rect -974 -38295 -842 -38235
rect -463 -38351 -406 -37902
rect -318 -38351 -272 -38151
rect -220 -38351 -174 -38151
rect 95 -38351 141 -38051
rect 193 -38351 239 -38051
rect 291 -38351 337 -38051
rect 404 -38351 450 -38051
rect 502 -38351 548 -38051
rect 600 -38351 646 -38051
rect 714 -38350 760 -38050
rect 812 -38350 858 -38050
rect 910 -38350 956 -38050
rect -1325 -38408 -406 -38351
rect -4247 -38649 -4206 -38648
rect -4012 -38669 -3869 -38609
rect -2324 -38634 -2155 -38627
rect -4012 -38675 -3952 -38669
rect -6475 -38944 -6429 -38744
rect -6279 -38944 -6233 -38744
rect -6083 -38944 -6037 -38744
rect -5853 -38926 -5796 -38691
rect -5024 -38701 -4855 -38691
rect -3153 -38691 -2155 -38634
rect -1653 -38646 -1499 -38586
rect 1030 -38543 1076 -37738
rect 1119 -37822 1255 -37776
rect 1513 -37787 1559 -37658
rect 1611 -37787 1657 -37687
rect 1709 -37787 1755 -37658
rect 1807 -37787 1853 -37687
rect 1183 -38431 1229 -37822
rect 2122 -38330 2168 -37994
rect 2220 -38294 2266 -37457
rect 2416 -37757 2462 -37457
rect 3020 -37614 3066 -37458
rect 3216 -37612 3262 -37458
rect 3118 -37614 3360 -37612
rect 3412 -37614 3458 -37458
rect 2995 -37660 3458 -37614
rect 3118 -37789 3164 -37660
rect 3216 -37789 3262 -37689
rect 3314 -37789 3360 -37660
rect 3412 -37789 3458 -37689
rect 2318 -38330 2364 -37994
rect 2416 -38294 2462 -37994
rect 2514 -38293 2560 -37994
rect 2514 -38330 2561 -38293
rect 2122 -38377 2561 -38330
rect 3727 -38332 3773 -37996
rect 3825 -38296 3871 -37459
rect 4021 -37759 4067 -37459
rect 4644 -37634 4690 -37434
rect 5382 -37634 5428 -37434
rect 5578 -37634 5624 -37434
rect 5774 -37634 5820 -37434
rect 6257 -37645 6303 -37445
rect 6355 -37676 6401 -37445
rect 6453 -37645 6499 -37445
rect 6573 -37645 6619 -37445
rect 6671 -37645 6717 -37445
rect 6769 -37645 6815 -37445
rect 7131 -37645 7177 -37445
rect 7327 -37645 7373 -37445
rect 7637 -37645 7683 -37445
rect 7946 -37645 7992 -37445
rect 5849 -37722 6401 -37676
rect 5853 -37731 5989 -37722
rect 7420 -37773 7559 -37755
rect 8035 -37766 8174 -37761
rect 8966 -37766 9184 -37707
rect 8035 -37773 9184 -37766
rect 7420 -37794 9184 -37773
rect 6262 -37812 6401 -37799
rect 7420 -37801 8275 -37794
rect 8966 -37796 9184 -37794
rect 7420 -37809 7559 -37801
rect 6262 -37840 6616 -37812
rect 8035 -37815 8174 -37801
rect 6262 -37853 6401 -37840
rect 6588 -37985 6616 -37840
rect 7011 -37838 7150 -37829
rect 7848 -37838 7984 -37829
rect 7011 -37866 7984 -37838
rect 7011 -37883 7150 -37866
rect 7848 -37875 7984 -37866
rect 7542 -37985 7673 -37973
rect 3923 -38332 3969 -37996
rect 4021 -38296 4067 -37996
rect 4119 -38295 4165 -37996
rect 6588 -38013 7673 -37985
rect 7542 -38019 7673 -38013
rect 4119 -38332 4166 -38295
rect 3727 -38379 4166 -38332
rect 4644 -38342 4690 -38142
rect 4742 -38342 4788 -38142
rect 5057 -38342 5103 -38042
rect 5155 -38342 5201 -38042
rect 5253 -38342 5299 -38042
rect 5366 -38342 5412 -38042
rect 5464 -38342 5510 -38042
rect 5562 -38342 5608 -38042
rect 5676 -38341 5722 -38041
rect 5774 -38341 5820 -38041
rect 5872 -38341 5918 -38041
rect 6257 -38251 6303 -38051
rect 6355 -38251 6401 -38051
rect 6671 -38251 6717 -38051
rect 6769 -38251 6815 -38051
rect 7033 -38251 7079 -38051
rect 7131 -38251 7177 -38051
rect 7327 -38251 7373 -38051
rect 7425 -38251 7471 -38051
rect 7637 -38251 7683 -38051
rect 7735 -38251 7781 -38051
rect 7946 -38251 7992 -38051
rect 8044 -38251 8090 -38051
rect 1183 -38477 2932 -38431
rect 1030 -38589 4500 -38543
rect -5638 -38944 -5592 -38744
rect -5442 -38944 -5396 -38744
rect -5246 -38944 -5200 -38744
rect -5027 -38929 -4981 -38829
rect -4929 -38929 -4883 -38829
rect -4831 -38929 -4785 -38829
rect -4733 -38929 -4687 -38829
rect -4635 -38929 -4589 -38829
rect -4537 -38929 -4491 -38829
rect -4439 -38929 -4393 -38829
rect -4341 -38929 -4295 -38829
rect -3775 -38944 -3729 -38744
rect -3579 -38944 -3533 -38744
rect -3383 -38944 -3337 -38744
rect -3153 -38926 -3096 -38691
rect -2324 -38701 -2155 -38691
rect -2938 -38944 -2892 -38744
rect -2742 -38944 -2696 -38744
rect -2546 -38944 -2500 -38744
rect -2327 -38929 -2281 -38829
rect -2229 -38929 -2183 -38829
rect -2131 -38929 -2085 -38829
rect -2033 -38929 -1987 -38829
rect -1935 -38929 -1889 -38829
rect -1837 -38929 -1791 -38829
rect -1739 -38929 -1693 -38829
rect -1641 -38929 -1595 -38829
rect -6475 -40382 -6429 -40182
rect -6279 -40382 -6233 -40182
rect -6083 -40382 -6037 -40182
rect -5853 -40435 -5796 -40200
rect -5638 -40382 -5592 -40182
rect -5442 -40382 -5396 -40182
rect -5246 -40382 -5200 -40182
rect -5027 -40297 -4981 -40197
rect -4929 -40297 -4883 -40197
rect -4831 -40297 -4785 -40197
rect -4733 -40297 -4687 -40197
rect -4635 -40297 -4589 -40197
rect -4537 -40297 -4491 -40197
rect -4439 -40297 -4393 -40197
rect -4341 -40297 -4295 -40197
rect -3775 -40382 -3729 -40182
rect -3579 -40382 -3533 -40182
rect -3383 -40382 -3337 -40182
rect -5024 -40435 -4855 -40425
rect -5853 -40492 -4855 -40435
rect -3153 -40435 -3096 -40200
rect -2938 -40382 -2892 -40182
rect -2742 -40382 -2696 -40182
rect -2546 -40382 -2500 -40182
rect -2327 -40297 -2281 -40197
rect -2229 -40297 -2183 -40197
rect -2131 -40297 -2085 -40197
rect -2033 -40297 -1987 -40197
rect -1935 -40297 -1889 -40197
rect -1837 -40297 -1791 -40197
rect -1739 -40297 -1693 -40197
rect -1641 -40297 -1595 -40197
rect -2324 -40435 -2155 -40425
rect -4012 -40457 -3952 -40451
rect -4247 -40478 -4206 -40477
rect -5024 -40499 -4855 -40492
rect -6573 -40662 -6527 -40562
rect -6475 -40662 -6429 -40562
rect -6377 -40662 -6331 -40562
rect -6279 -40662 -6233 -40562
rect -6181 -40662 -6135 -40562
rect -6083 -40662 -6037 -40562
rect -7033 -40943 -6858 -40724
rect -6339 -40885 -6202 -40825
rect -6687 -40943 -6627 -40896
rect -7033 -41007 -6627 -40943
rect -7033 -41038 -6858 -41007
rect -6687 -41033 -6627 -41007
rect -6324 -41073 -6229 -40885
rect -5914 -41003 -5854 -40536
rect -4342 -40538 -4205 -40478
rect -4012 -40517 -3869 -40457
rect -3153 -40492 -2155 -40435
rect -2324 -40499 -2155 -40492
rect -5736 -40662 -5690 -40562
rect -5638 -40662 -5592 -40562
rect -5540 -40662 -5494 -40562
rect -5442 -40662 -5396 -40562
rect -5344 -40662 -5298 -40562
rect -5246 -40662 -5200 -40562
rect -5027 -40712 -4981 -40612
rect -4929 -40712 -4883 -40612
rect -4831 -40712 -4785 -40612
rect -4733 -40712 -4687 -40612
rect -4635 -40712 -4589 -40612
rect -4537 -40712 -4491 -40612
rect -4439 -40712 -4393 -40612
rect -4341 -40712 -4295 -40612
rect -5950 -41063 -5818 -41003
rect -4247 -41023 -4206 -40538
rect -6811 -41103 -6229 -41073
rect -5737 -41071 -4206 -41023
rect -6811 -41163 -6216 -41103
rect -6811 -41168 -6229 -41163
rect -6811 -41247 -6716 -41168
rect -7026 -41342 -6716 -41247
rect -6573 -41320 -6527 -41220
rect -6475 -41320 -6429 -41220
rect -6377 -41320 -6331 -41220
rect -6279 -41320 -6233 -41220
rect -6181 -41320 -6135 -41220
rect -6083 -41320 -6037 -41220
rect -5737 -41225 -5689 -41071
rect -5735 -41270 -5689 -41225
rect -5637 -41270 -5591 -41170
rect -5545 -41189 -5484 -41071
rect -5539 -41270 -5493 -41189
rect -5441 -41270 -5395 -41170
rect -5349 -41191 -5288 -41071
rect -5343 -41270 -5297 -41191
rect -5245 -41270 -5199 -41170
rect -5158 -41189 -5097 -41071
rect -5147 -41270 -5101 -41189
rect -5049 -41270 -5003 -41170
rect -4830 -41320 -4784 -41220
rect -4732 -41320 -4686 -41220
rect -4634 -41320 -4588 -41220
rect -4536 -41320 -4490 -41220
rect -4438 -41320 -4392 -41220
rect -4340 -41320 -4294 -41220
rect -5175 -41390 -5006 -41383
rect -5175 -41447 -4177 -41390
rect -4012 -41265 -3952 -40517
rect -1653 -40540 -1499 -40480
rect -3873 -40662 -3827 -40562
rect -3775 -40662 -3729 -40562
rect -3677 -40662 -3631 -40562
rect -3579 -40662 -3533 -40562
rect -3481 -40662 -3435 -40562
rect -3383 -40662 -3337 -40562
rect -3742 -40891 -3605 -40831
rect -3731 -41099 -3636 -40891
rect -3036 -40662 -2990 -40562
rect -2938 -40662 -2892 -40562
rect -2840 -40662 -2794 -40562
rect -2742 -40662 -2696 -40562
rect -2644 -40662 -2598 -40562
rect -2546 -40662 -2500 -40562
rect -2327 -40712 -2281 -40612
rect -2229 -40712 -2183 -40612
rect -2131 -40712 -2085 -40612
rect -2033 -40712 -1987 -40612
rect -1935 -40712 -1889 -40612
rect -1837 -40712 -1791 -40612
rect -1739 -40712 -1693 -40612
rect -1641 -40712 -1595 -40612
rect -1545 -40815 -1499 -40540
rect 1030 -40583 4500 -40537
rect -2318 -40860 -1499 -40815
rect -1325 -40775 -406 -40718
rect -2318 -40861 -1507 -40860
rect -2318 -41027 -2272 -40861
rect -1325 -40896 -1268 -40775
rect -1104 -40891 -972 -40831
rect -3032 -41073 -2272 -41027
rect -1534 -40953 -1268 -40896
rect -3749 -41159 -3612 -41099
rect -3032 -41170 -2986 -41073
rect -2837 -41170 -2795 -41073
rect -2642 -41170 -2600 -41073
rect -2446 -41170 -2404 -41073
rect -4013 -41310 -3952 -41265
rect -4013 -41397 -3953 -41310
rect -3873 -41320 -3827 -41220
rect -3775 -41320 -3729 -41220
rect -3677 -41320 -3631 -41220
rect -3579 -41320 -3533 -41220
rect -3481 -41320 -3435 -41220
rect -3383 -41320 -3337 -41220
rect -3035 -41270 -2986 -41170
rect -2937 -41270 -2891 -41170
rect -2839 -41270 -2793 -41170
rect -2741 -41270 -2695 -41170
rect -2643 -41270 -2597 -41170
rect -2545 -41270 -2499 -41170
rect -2447 -41270 -2401 -41170
rect -2349 -41270 -2303 -41170
rect -2130 -41320 -2084 -41220
rect -2032 -41320 -1986 -41220
rect -1934 -41320 -1888 -41220
rect -1836 -41320 -1790 -41220
rect -1738 -41320 -1692 -41220
rect -1640 -41320 -1594 -41220
rect -2475 -41390 -2306 -41383
rect -1534 -41390 -1477 -40953
rect -1427 -41061 -1295 -41001
rect -1394 -41289 -1336 -41061
rect -1087 -41100 -992 -40891
rect -1122 -41160 -985 -41100
rect -5175 -41457 -5006 -41447
rect -6573 -41700 -6527 -41500
rect -6377 -41700 -6331 -41500
rect -6181 -41700 -6135 -41500
rect -5735 -41685 -5689 -41585
rect -5637 -41685 -5591 -41585
rect -5539 -41685 -5493 -41585
rect -5441 -41685 -5395 -41585
rect -5343 -41685 -5297 -41585
rect -5245 -41685 -5199 -41585
rect -5147 -41685 -5101 -41585
rect -5049 -41685 -5003 -41585
rect -4830 -41700 -4784 -41500
rect -4634 -41700 -4588 -41500
rect -4438 -41700 -4392 -41500
rect -4234 -41682 -4177 -41447
rect -2475 -41447 -1477 -41390
rect -1396 -41421 -1336 -41289
rect -1248 -41320 -1202 -41220
rect -1150 -41320 -1104 -41220
rect -1052 -41320 -1006 -41220
rect -954 -41320 -908 -41220
rect -856 -41320 -810 -41220
rect -758 -41320 -712 -41220
rect -463 -41224 -406 -40775
rect -318 -40975 -272 -40775
rect -220 -40975 -174 -40775
rect 95 -41075 141 -40775
rect 193 -41075 239 -40775
rect 291 -41075 337 -40775
rect 404 -41075 450 -40775
rect 502 -41075 548 -40775
rect 600 -41075 646 -40775
rect 714 -41076 760 -40776
rect 812 -41076 858 -40776
rect 910 -41076 956 -40776
rect -463 -41277 -322 -41224
rect 1030 -41388 1076 -40583
rect 1183 -40695 2932 -40649
rect 1183 -41304 1229 -40695
rect 2122 -40796 2561 -40749
rect 2122 -41132 2168 -40796
rect 1119 -41350 1255 -41304
rect -2475 -41457 -2306 -41447
rect -3873 -41700 -3827 -41500
rect -3677 -41700 -3631 -41500
rect -3481 -41700 -3435 -41500
rect -3035 -41685 -2989 -41585
rect -2937 -41685 -2891 -41585
rect -2839 -41685 -2793 -41585
rect -2741 -41685 -2695 -41585
rect -2643 -41685 -2597 -41585
rect -2545 -41685 -2499 -41585
rect -2447 -41685 -2401 -41585
rect -2349 -41685 -2303 -41585
rect -2130 -41700 -2084 -41500
rect -1934 -41700 -1888 -41500
rect -1738 -41700 -1692 -41500
rect -1534 -41682 -1477 -41447
rect -1248 -41700 -1202 -41500
rect -1052 -41700 -1006 -41500
rect -856 -41700 -810 -41500
rect -318 -41683 -272 -41483
rect 420 -41683 466 -41483
rect 616 -41683 662 -41483
rect 812 -41683 858 -41483
rect 1030 -41522 1084 -41388
rect 1513 -41468 1559 -41339
rect 1611 -41439 1657 -41339
rect 1709 -41468 1755 -41339
rect 1807 -41439 1853 -41339
rect 1390 -41514 1853 -41468
rect 1038 -41524 1084 -41522
rect 1415 -41670 1461 -41514
rect 1513 -41516 1755 -41514
rect 1611 -41670 1657 -41516
rect 1807 -41670 1853 -41514
rect 2220 -41669 2266 -40832
rect 2318 -41132 2364 -40796
rect 2416 -41132 2462 -40832
rect 2514 -40833 2561 -40796
rect 3727 -40794 4166 -40747
rect 2514 -41132 2560 -40833
rect 3727 -41130 3773 -40794
rect 2416 -41669 2462 -41369
rect 3118 -41466 3164 -41337
rect 3216 -41437 3262 -41337
rect 3314 -41466 3360 -41337
rect 3412 -41437 3458 -41337
rect 2995 -41512 3458 -41466
rect 3020 -41668 3066 -41512
rect 3118 -41514 3360 -41512
rect 3216 -41668 3262 -41514
rect 3412 -41668 3458 -41512
rect 3825 -41667 3871 -40830
rect 3923 -41130 3969 -40794
rect 4021 -41130 4067 -40830
rect 4119 -40831 4166 -40794
rect 4119 -41130 4165 -40831
rect 4644 -40984 4690 -40784
rect 4742 -40984 4788 -40784
rect 5057 -41084 5103 -40784
rect 5155 -41084 5201 -40784
rect 5253 -41084 5299 -40784
rect 5366 -41084 5412 -40784
rect 5464 -41084 5510 -40784
rect 5562 -41084 5608 -40784
rect 5676 -41085 5722 -40785
rect 5774 -41085 5820 -40785
rect 5872 -41085 5918 -40785
rect 6257 -41075 6303 -40875
rect 6355 -41075 6401 -40875
rect 6671 -41075 6717 -40875
rect 6769 -41075 6815 -40875
rect 7033 -41075 7079 -40875
rect 7131 -41075 7177 -40875
rect 7327 -41075 7373 -40875
rect 7425 -41075 7471 -40875
rect 7637 -41075 7683 -40875
rect 7735 -41075 7781 -40875
rect 7946 -41075 7992 -40875
rect 8044 -41075 8090 -40875
rect 7542 -41113 7673 -41107
rect 6588 -41141 7673 -41113
rect 6262 -41286 6401 -41273
rect 6588 -41286 6616 -41141
rect 7542 -41153 7673 -41141
rect 6262 -41314 6616 -41286
rect 7011 -41260 7150 -41243
rect 7848 -41260 7984 -41251
rect 7011 -41288 7984 -41260
rect 7011 -41297 7150 -41288
rect 7848 -41297 7984 -41288
rect 6262 -41327 6401 -41314
rect 7420 -41325 7559 -41317
rect 8035 -41325 8174 -41311
rect 7420 -41332 8275 -41325
rect 9133 -41332 9161 -37796
rect 7420 -41353 9161 -41332
rect 4021 -41667 4067 -41367
rect 7420 -41371 7559 -41353
rect 8035 -41360 9161 -41353
rect 8035 -41365 8174 -41360
rect 5853 -41404 5989 -41395
rect 5849 -41450 6401 -41404
rect 4644 -41692 4690 -41492
rect 5382 -41692 5428 -41492
rect 5578 -41692 5624 -41492
rect 5774 -41692 5820 -41492
rect 6257 -41681 6303 -41481
rect 6355 -41681 6401 -41450
rect 6453 -41681 6499 -41481
rect 6573 -41681 6619 -41481
rect 6671 -41681 6717 -41481
rect 6769 -41681 6815 -41481
rect 7131 -41681 7177 -41481
rect 7327 -41681 7373 -41481
rect 7637 -41681 7683 -41481
rect 7946 -41681 7992 -41481
rect 2527 -42074 2682 -42072
rect -6774 -42081 2682 -42074
rect -6898 -42116 2682 -42081
rect -6898 -42127 -6762 -42116
rect 2527 -42118 2682 -42116
rect -4418 -42156 -4282 -42154
rect -4418 -42198 2767 -42156
rect -4418 -42200 -4282 -42198
rect 2631 -42202 2767 -42198
rect 9468 -40487 9519 -36809
rect 9465 -40582 9524 -40487
rect -6753 -43326 -6707 -43126
rect -6655 -43326 -6609 -43126
rect -6339 -43326 -6293 -43126
rect -6241 -43326 -6195 -43126
rect -5977 -43326 -5931 -43126
rect -5879 -43326 -5833 -43126
rect -5683 -43326 -5637 -43126
rect -5585 -43326 -5539 -43126
rect -5373 -43326 -5327 -43126
rect -5275 -43326 -5229 -43126
rect -5064 -43326 -5018 -43126
rect -4966 -43326 -4920 -43126
rect -5468 -43364 -5337 -43358
rect -6422 -43392 -5337 -43364
rect -6748 -43537 -6609 -43524
rect -6422 -43537 -6394 -43392
rect -5468 -43404 -5337 -43392
rect 9468 -42317 9519 -40582
rect -4713 -42363 9519 -42317
rect -4713 -42368 9095 -42363
rect -6748 -43565 -6394 -43537
rect -5999 -43511 -5860 -43494
rect -5162 -43511 -5026 -43502
rect -5999 -43539 -5026 -43511
rect -5999 -43548 -5860 -43539
rect -5162 -43548 -5026 -43539
rect -6748 -43578 -6609 -43565
rect -5590 -43576 -5451 -43568
rect -4975 -43576 -4836 -43562
rect -4713 -43576 -4685 -42368
rect 9283 -42399 9431 -42391
rect 9554 -42399 9590 -36727
rect 9624 -41279 9675 -36659
rect 9618 -41418 9687 -41279
rect -2228 -42435 9590 -42399
rect -4421 -42589 -4375 -42453
rect -4420 -43159 -4376 -42589
rect -4421 -43295 -4375 -43159
rect -4253 -43326 -4207 -43126
rect -4155 -43326 -4109 -43126
rect -3839 -43326 -3793 -43126
rect -3741 -43326 -3695 -43126
rect -3477 -43326 -3431 -43126
rect -3379 -43326 -3333 -43126
rect -3183 -43326 -3137 -43126
rect -3085 -43326 -3039 -43126
rect -2873 -43326 -2827 -43126
rect -2775 -43326 -2729 -43126
rect -2564 -43326 -2518 -43126
rect -2466 -43326 -2420 -43126
rect -2968 -43364 -2837 -43358
rect -3922 -43392 -2837 -43364
rect -5590 -43604 -4685 -43576
rect -4248 -43537 -4109 -43524
rect -3922 -43537 -3894 -43392
rect -2968 -43404 -2837 -43392
rect -3866 -43437 -3727 -43420
rect -2788 -43437 -2649 -43414
rect -3866 -43439 -2649 -43437
rect -2228 -43439 -2200 -42435
rect 9283 -42439 9431 -42435
rect 9624 -42467 9675 -41418
rect -3866 -43465 -2200 -43439
rect -3866 -43474 -3727 -43465
rect -2788 -43467 -2200 -43465
rect -2142 -42498 9675 -42467
rect -2142 -42518 9095 -42498
rect 9288 -42505 9675 -42498
rect -2788 -43468 -2649 -43467
rect -4248 -43565 -3894 -43537
rect -3499 -43511 -3360 -43494
rect -2662 -43511 -2526 -43502
rect -3499 -43539 -2526 -43511
rect -3499 -43548 -3360 -43539
rect -2662 -43548 -2526 -43539
rect -4248 -43578 -4109 -43565
rect -3090 -43576 -2951 -43568
rect -2475 -43576 -2336 -43562
rect -2142 -43576 -2114 -42518
rect 9123 -42546 9266 -42528
rect 9721 -42546 9749 -36580
rect 9806 -40167 9834 -36523
rect 9786 -40285 9850 -40167
rect 256 -42574 9749 -42546
rect -1708 -42874 -1572 -42873
rect -1873 -42918 -1572 -42874
rect -1872 -43155 -1828 -42918
rect -1708 -42919 -1572 -42918
rect -1873 -43291 -1827 -43155
rect -1753 -43326 -1707 -43126
rect -1655 -43326 -1609 -43126
rect -1339 -43326 -1293 -43126
rect -1241 -43326 -1195 -43126
rect -977 -43326 -931 -43126
rect -879 -43326 -833 -43126
rect -683 -43326 -637 -43126
rect -585 -43326 -539 -43126
rect -373 -43326 -327 -43126
rect -275 -43326 -229 -43126
rect -64 -43326 -18 -43126
rect 34 -43326 80 -43126
rect -468 -43364 -337 -43358
rect -1422 -43392 -337 -43364
rect -3090 -43604 -2114 -43576
rect -1748 -43537 -1609 -43524
rect -1422 -43537 -1394 -43392
rect -468 -43404 -337 -43392
rect -1366 -43437 -1227 -43420
rect -288 -43437 -149 -43414
rect -1366 -43439 -149 -43437
rect 256 -43439 284 -42574
rect 9123 -42575 9266 -42574
rect 9806 -42603 9834 -40285
rect -1366 -43465 284 -43439
rect -1366 -43474 -1227 -43465
rect -288 -43467 284 -43465
rect 330 -42631 9834 -42603
rect -288 -43468 -149 -43467
rect -1748 -43565 -1394 -43537
rect -999 -43511 -860 -43494
rect -162 -43511 -26 -43502
rect -999 -43539 -26 -43511
rect -999 -43548 -860 -43539
rect -162 -43548 -26 -43539
rect -1748 -43578 -1609 -43565
rect -590 -43576 -451 -43568
rect 25 -43576 164 -43562
rect 330 -43576 358 -42631
rect 8997 -42666 9141 -42659
rect 9883 -42666 9911 -36460
rect 2722 -42694 9911 -42666
rect 9948 -37930 9986 -36396
rect 9948 -38063 9998 -37930
rect 789 -42861 925 -42860
rect 608 -42905 925 -42861
rect 608 -43155 652 -42905
rect 789 -42906 925 -42905
rect 607 -43291 653 -43155
rect 747 -43326 793 -43126
rect 845 -43326 891 -43126
rect 1161 -43326 1207 -43126
rect 1259 -43326 1305 -43126
rect 1523 -43326 1569 -43126
rect 1621 -43326 1667 -43126
rect 1817 -43326 1863 -43126
rect 1915 -43326 1961 -43126
rect 2127 -43326 2173 -43126
rect 2225 -43326 2271 -43126
rect 2436 -43326 2482 -43126
rect 2534 -43326 2580 -43126
rect 2032 -43364 2163 -43358
rect 1078 -43392 2163 -43364
rect -590 -43604 358 -43576
rect 752 -43537 891 -43524
rect 1078 -43537 1106 -43392
rect 2032 -43404 2163 -43392
rect 1134 -43437 1273 -43420
rect 2212 -43437 2351 -43414
rect 1134 -43439 2351 -43437
rect 2722 -43439 2750 -42694
rect 8997 -42706 9141 -42694
rect 9948 -42730 9986 -38063
rect 1134 -43465 2750 -43439
rect 1134 -43474 1273 -43465
rect 2212 -43467 2750 -43465
rect 2805 -42740 8503 -42730
rect 9183 -42740 9986 -42730
rect 2805 -42768 9986 -42740
rect 2212 -43468 2351 -43467
rect 752 -43565 1106 -43537
rect 1501 -43511 1640 -43494
rect 2338 -43511 2474 -43502
rect 1501 -43539 2474 -43511
rect 1501 -43548 1640 -43539
rect 2338 -43548 2474 -43539
rect 752 -43578 891 -43565
rect 1910 -43576 2049 -43568
rect 2525 -43576 2664 -43562
rect 2805 -43576 2833 -42768
rect 2972 -42843 3108 -42797
rect 3025 -43155 3069 -42843
rect 5877 -42859 6013 -42813
rect 3024 -43291 3070 -43155
rect 3247 -43326 3293 -43126
rect 3345 -43326 3391 -43126
rect 3661 -43326 3707 -43126
rect 3759 -43326 3805 -43126
rect 4023 -43326 4069 -43126
rect 4121 -43326 4167 -43126
rect 4317 -43326 4363 -43126
rect 4415 -43326 4461 -43126
rect 4627 -43326 4673 -43126
rect 4725 -43326 4771 -43126
rect 4936 -43326 4982 -43126
rect 5034 -43326 5080 -43126
rect 5930 -43155 5974 -42859
rect 5929 -43291 5975 -43155
rect 4532 -43364 4663 -43358
rect 3578 -43392 4663 -43364
rect 1910 -43604 2833 -43576
rect 3252 -43537 3391 -43524
rect 3578 -43537 3606 -43392
rect 4532 -43404 4663 -43392
rect 10111 -42873 10139 -36253
rect 6110 -42901 10139 -42873
rect 3252 -43565 3606 -43537
rect 4001 -43511 4140 -43494
rect 4838 -43511 4974 -43502
rect 4001 -43539 4974 -43511
rect 4001 -43548 4140 -43539
rect 4838 -43548 4974 -43539
rect 3252 -43578 3391 -43565
rect 4410 -43576 4549 -43568
rect 5025 -43576 5164 -43562
rect 6110 -43576 6138 -42901
rect 6247 -43326 6293 -43126
rect 6345 -43326 6391 -43126
rect 6661 -43326 6707 -43126
rect 6759 -43326 6805 -43126
rect 7023 -43326 7069 -43126
rect 7121 -43326 7167 -43126
rect 7317 -43326 7363 -43126
rect 7415 -43326 7461 -43126
rect 7627 -43326 7673 -43126
rect 7725 -43326 7771 -43126
rect 7936 -43326 7982 -43126
rect 8034 -43326 8080 -43126
rect 7532 -43364 7663 -43358
rect 6578 -43392 7663 -43364
rect 4410 -43604 6138 -43576
rect 6252 -43537 6391 -43524
rect 6578 -43537 6606 -43392
rect 7532 -43404 7663 -43392
rect 6252 -43565 6606 -43537
rect 7001 -43511 7140 -43494
rect 7838 -43511 7974 -43502
rect 7001 -43539 7974 -43511
rect 7001 -43548 7140 -43539
rect 7838 -43548 7974 -43539
rect 6252 -43578 6391 -43565
rect 7410 -43576 7549 -43568
rect 8025 -43576 8164 -43562
rect 10267 -43576 10295 -35550
rect 7410 -43604 10295 -43576
rect -5590 -43622 -5451 -43604
rect -4975 -43616 -4836 -43604
rect -3090 -43622 -2951 -43604
rect -2475 -43616 -2336 -43604
rect -590 -43622 -451 -43604
rect 25 -43616 164 -43604
rect 1910 -43622 2049 -43604
rect 2525 -43616 2664 -43604
rect 4410 -43622 4549 -43604
rect 5025 -43616 5164 -43604
rect 7410 -43622 7549 -43604
rect 8025 -43616 8164 -43604
rect -6753 -43932 -6707 -43732
rect -6655 -43932 -6609 -43732
rect -6557 -43932 -6511 -43732
rect -6437 -43932 -6391 -43732
rect -6339 -43932 -6293 -43732
rect -6241 -43932 -6195 -43732
rect -5879 -43932 -5833 -43732
rect -5683 -43932 -5637 -43732
rect -5373 -43932 -5327 -43732
rect -5064 -43932 -5018 -43732
rect -4253 -43932 -4207 -43732
rect -4155 -43932 -4109 -43732
rect -4057 -43932 -4011 -43732
rect -3937 -43932 -3891 -43732
rect -3839 -43932 -3793 -43732
rect -3741 -43932 -3695 -43732
rect -3379 -43932 -3333 -43732
rect -3183 -43932 -3137 -43732
rect -2873 -43932 -2827 -43732
rect -2564 -43932 -2518 -43732
rect -1753 -43932 -1707 -43732
rect -1655 -43932 -1609 -43732
rect -1557 -43932 -1511 -43732
rect -1437 -43932 -1391 -43732
rect -1339 -43932 -1293 -43732
rect -1241 -43932 -1195 -43732
rect -879 -43932 -833 -43732
rect -683 -43932 -637 -43732
rect -373 -43932 -327 -43732
rect -64 -43932 -18 -43732
rect 747 -43932 793 -43732
rect 845 -43932 891 -43732
rect 943 -43932 989 -43732
rect 1063 -43932 1109 -43732
rect 1161 -43932 1207 -43732
rect 1259 -43932 1305 -43732
rect 1621 -43932 1667 -43732
rect 1817 -43932 1863 -43732
rect 2127 -43932 2173 -43732
rect 2436 -43932 2482 -43732
rect 3247 -43932 3293 -43732
rect 3345 -43932 3391 -43732
rect 3443 -43932 3489 -43732
rect 3563 -43932 3609 -43732
rect 3661 -43932 3707 -43732
rect 3759 -43932 3805 -43732
rect 4121 -43932 4167 -43732
rect 4317 -43932 4363 -43732
rect 4627 -43932 4673 -43732
rect 4936 -43932 4982 -43732
rect 6247 -43932 6293 -43732
rect 6345 -43932 6391 -43732
rect 6443 -43932 6489 -43732
rect 6563 -43932 6609 -43732
rect 6661 -43932 6707 -43732
rect 6759 -43932 6805 -43732
rect 7121 -43932 7167 -43732
rect 7317 -43932 7363 -43732
rect 7627 -43932 7673 -43732
rect 7936 -43932 7982 -43732
rect -7311 -44295 -7148 -44120
rect -22432 -46279 -22309 -46156
rect -7300 -46650 -7168 -44295
rect 8965 -45483 9026 -44106
rect 8896 -45484 9026 -45483
rect 8896 -45517 9027 -45484
rect 8897 -45602 9027 -45517
rect 9079 -45611 9143 -44102
rect 9077 -45783 9143 -45611
rect 9056 -45784 9143 -45783
rect 9056 -45907 9179 -45784
rect 9224 -46151 9284 -44066
rect 9207 -46274 9330 -46151
rect 10909 -43176 11109 -37120
rect 12773 -40662 13042 -32036
rect 13765 -32969 78890 -32658
rect 12712 -41003 13098 -40662
rect 13765 -40952 14016 -32969
rect 14352 -33419 69622 -33242
rect 14352 -39702 14683 -33419
rect 15464 -33978 60913 -33757
rect 15464 -37922 15554 -33978
rect 16845 -34535 51724 -34309
rect 16453 -35015 42899 -34750
rect 16171 -35421 34418 -35172
rect 16197 -36101 16762 -36100
rect 15912 -36241 16762 -36101
rect 26597 -36533 33062 -36364
rect 15879 -37163 16146 -37085
rect 15879 -37318 25793 -37163
rect 15879 -37383 16146 -37318
rect 16142 -37827 16969 -37676
rect 20275 -37810 20321 -37710
rect 20373 -37810 20419 -37710
rect 20471 -37810 20517 -37710
rect 20569 -37810 20615 -37710
rect 20667 -37810 20713 -37710
rect 20765 -37810 20811 -37710
rect 20863 -37810 20909 -37710
rect 20961 -37810 21007 -37710
rect 15460 -38086 15558 -37922
rect 14248 -40127 14762 -39702
rect 15464 -40251 15554 -38086
rect 18169 -38129 18215 -37929
rect 18267 -38129 18313 -37929
rect 18365 -38129 18411 -37929
rect 18463 -38129 18509 -37929
rect 21180 -37895 21226 -37695
rect 21376 -37895 21422 -37695
rect 21572 -37895 21618 -37695
rect 20835 -37948 21004 -37938
rect 21776 -37948 21833 -37713
rect 22017 -37895 22063 -37695
rect 22213 -37895 22259 -37695
rect 22409 -37895 22455 -37695
rect 22975 -37810 23021 -37710
rect 23073 -37810 23119 -37710
rect 23171 -37810 23217 -37710
rect 23269 -37810 23315 -37710
rect 23367 -37810 23413 -37710
rect 23465 -37810 23511 -37710
rect 23563 -37810 23609 -37710
rect 23661 -37810 23707 -37710
rect 23880 -37895 23926 -37695
rect 24076 -37895 24122 -37695
rect 24272 -37895 24318 -37695
rect 20179 -38053 20333 -37993
rect 20835 -38005 21833 -37948
rect 23535 -37948 23704 -37938
rect 24476 -37948 24533 -37713
rect 24717 -37895 24763 -37695
rect 24913 -37895 24959 -37695
rect 25109 -37895 25155 -37695
rect 22632 -37970 22692 -37964
rect 20835 -38012 21004 -38005
rect 22549 -38030 22692 -37970
rect 22886 -37991 22927 -37990
rect 19005 -38167 19047 -38163
rect 18923 -38227 19055 -38167
rect 18169 -39093 18215 -38493
rect 18381 -39093 18427 -38493
rect 18479 -39093 18525 -38493
rect 18577 -39093 18623 -38493
rect 18690 -39093 18736 -38493
rect 18788 -39093 18834 -38493
rect 18886 -39093 18932 -38493
rect 16004 -40030 18114 -39834
rect 17918 -40036 18114 -40030
rect 17918 -40190 18116 -40036
rect 17911 -40232 18948 -40190
rect 15464 -40264 17447 -40251
rect 15464 -40306 18858 -40264
rect 15464 -40341 17447 -40306
rect 18164 -40747 18210 -40547
rect 18262 -40747 18308 -40547
rect 18360 -40747 18406 -40547
rect 18574 -40852 18706 -40792
rect 13749 -41182 14037 -40952
rect 18661 -40965 18703 -40852
rect 18816 -40877 18858 -40306
rect 18906 -40793 18948 -40232
rect 19005 -40261 19047 -38227
rect 19095 -38288 20005 -38231
rect 19095 -39639 19152 -38288
rect 19652 -38404 19784 -38344
rect 19672 -38613 19767 -38404
rect 19948 -38409 20005 -38288
rect 20179 -38328 20225 -38053
rect 20275 -38225 20321 -38125
rect 20373 -38225 20419 -38125
rect 20471 -38225 20517 -38125
rect 20569 -38225 20615 -38125
rect 20667 -38225 20713 -38125
rect 20765 -38225 20811 -38125
rect 20863 -38225 20909 -38125
rect 20961 -38225 21007 -38125
rect 21180 -38175 21226 -38075
rect 21278 -38175 21324 -38075
rect 21376 -38175 21422 -38075
rect 21474 -38175 21520 -38075
rect 21572 -38175 21618 -38075
rect 21670 -38175 21716 -38075
rect 20179 -38373 20998 -38328
rect 20187 -38374 20998 -38373
rect 19948 -38466 20214 -38409
rect 19975 -38574 20107 -38514
rect 19665 -38673 19802 -38613
rect 19392 -38833 19438 -38733
rect 19490 -38833 19536 -38733
rect 19588 -38833 19634 -38733
rect 19686 -38833 19732 -38733
rect 19784 -38833 19830 -38733
rect 19882 -38833 19928 -38733
rect 20016 -38802 20074 -38574
rect 20016 -38934 20076 -38802
rect 20157 -38903 20214 -38466
rect 20952 -38540 20998 -38374
rect 22017 -38175 22063 -38075
rect 22115 -38175 22161 -38075
rect 22213 -38175 22259 -38075
rect 22311 -38175 22357 -38075
rect 22409 -38175 22455 -38075
rect 22507 -38175 22553 -38075
rect 22285 -38404 22422 -38344
rect 20952 -38586 21712 -38540
rect 21084 -38683 21126 -38586
rect 21280 -38683 21322 -38586
rect 21475 -38683 21517 -38586
rect 21666 -38683 21712 -38586
rect 22316 -38612 22411 -38404
rect 22292 -38672 22429 -38612
rect 20274 -38833 20320 -38733
rect 20372 -38833 20418 -38733
rect 20470 -38833 20516 -38733
rect 20568 -38833 20614 -38733
rect 20666 -38833 20712 -38733
rect 20764 -38833 20810 -38733
rect 20983 -38783 21029 -38683
rect 21081 -38783 21127 -38683
rect 21179 -38783 21225 -38683
rect 21277 -38783 21323 -38683
rect 21375 -38783 21421 -38683
rect 21473 -38783 21519 -38683
rect 21571 -38783 21617 -38683
rect 21666 -38783 21715 -38683
rect 22017 -38833 22063 -38733
rect 22115 -38833 22161 -38733
rect 22213 -38833 22259 -38733
rect 22311 -38833 22357 -38733
rect 22409 -38833 22455 -38733
rect 22507 -38833 22553 -38733
rect 22632 -38778 22692 -38030
rect 22885 -38051 23022 -37991
rect 23535 -38005 24533 -37948
rect 23535 -38012 23704 -38005
rect 22632 -38823 22693 -38778
rect 20986 -38903 21155 -38896
rect 20157 -38960 21155 -38903
rect 22633 -38910 22693 -38823
rect 22886 -38536 22927 -38051
rect 22975 -38225 23021 -38125
rect 23073 -38225 23119 -38125
rect 23171 -38225 23217 -38125
rect 23269 -38225 23315 -38125
rect 23367 -38225 23413 -38125
rect 23465 -38225 23511 -38125
rect 23563 -38225 23609 -38125
rect 23661 -38225 23707 -38125
rect 23880 -38175 23926 -38075
rect 23978 -38175 24024 -38075
rect 24076 -38175 24122 -38075
rect 24174 -38175 24220 -38075
rect 24272 -38175 24318 -38075
rect 24370 -38175 24416 -38075
rect 24534 -38516 24594 -38049
rect 24717 -38175 24763 -38075
rect 24815 -38175 24861 -38075
rect 24913 -38175 24959 -38075
rect 25011 -38175 25057 -38075
rect 25109 -38175 25155 -38075
rect 25207 -38175 25253 -38075
rect 24882 -38398 25019 -38338
rect 22886 -38584 24417 -38536
rect 24498 -38576 24630 -38516
rect 22974 -38833 23020 -38733
rect 23072 -38833 23118 -38733
rect 23170 -38833 23216 -38733
rect 23268 -38833 23314 -38733
rect 23366 -38833 23412 -38733
rect 23464 -38833 23510 -38733
rect 23683 -38783 23729 -38683
rect 23777 -38702 23838 -38584
rect 23781 -38783 23827 -38702
rect 23879 -38783 23925 -38683
rect 23968 -38704 24029 -38584
rect 23977 -38783 24023 -38704
rect 24075 -38783 24121 -38683
rect 24164 -38702 24225 -38584
rect 24173 -38783 24219 -38702
rect 24271 -38783 24317 -38683
rect 24369 -38738 24417 -38584
rect 24909 -38616 25004 -38398
rect 25307 -38456 25367 -38409
rect 25307 -38520 25576 -38456
rect 25307 -38546 25453 -38520
rect 24896 -38676 25028 -38616
rect 24369 -38783 24415 -38738
rect 24717 -38833 24763 -38733
rect 24815 -38833 24861 -38733
rect 24913 -38833 24959 -38733
rect 25011 -38833 25057 -38733
rect 25109 -38833 25155 -38733
rect 25207 -38833 25253 -38733
rect 23686 -38903 23855 -38896
rect 19490 -39213 19536 -39013
rect 19686 -39213 19732 -39013
rect 19882 -39213 19928 -39013
rect 20157 -39195 20214 -38960
rect 20986 -38970 21155 -38960
rect 22857 -38960 23855 -38903
rect 20372 -39213 20418 -39013
rect 20568 -39213 20614 -39013
rect 20764 -39213 20810 -39013
rect 20983 -39198 21029 -39098
rect 21081 -39198 21127 -39098
rect 21179 -39198 21225 -39098
rect 21277 -39198 21323 -39098
rect 21375 -39198 21421 -39098
rect 21473 -39198 21519 -39098
rect 21571 -39198 21617 -39098
rect 21669 -39198 21715 -39098
rect 22115 -39213 22161 -39013
rect 22311 -39213 22357 -39013
rect 22507 -39213 22553 -39013
rect 22857 -39195 22914 -38960
rect 23686 -38970 23855 -38960
rect 23072 -39213 23118 -39013
rect 23268 -39213 23314 -39013
rect 23464 -39213 23510 -39013
rect 23683 -39198 23729 -39098
rect 23781 -39198 23827 -39098
rect 23879 -39198 23925 -39098
rect 23977 -39198 24023 -39098
rect 24075 -39198 24121 -39098
rect 24173 -39198 24219 -39098
rect 24271 -39198 24317 -39098
rect 24369 -39198 24415 -39098
rect 24815 -39213 24861 -39013
rect 25011 -39213 25057 -39013
rect 25207 -39213 25253 -39013
rect 25363 -39390 25453 -38546
rect 21421 -39480 25453 -39390
rect 21421 -39571 21581 -39480
rect 19095 -39696 22367 -39639
rect 21418 -39886 21578 -39754
rect 19005 -40303 19775 -40261
rect 21315 -40269 21447 -40209
rect 19110 -40747 19156 -40547
rect 19208 -40747 19254 -40547
rect 19306 -40747 19352 -40547
rect 19022 -40793 19154 -40786
rect 18906 -40835 19154 -40793
rect 19022 -40846 19154 -40835
rect 19245 -40877 19377 -40866
rect 18816 -40919 19377 -40877
rect 19245 -40926 19377 -40919
rect 19610 -40965 19670 -40935
rect 18661 -41007 19670 -40965
rect 18164 -41439 18210 -41039
rect 18375 -41439 18421 -41039
rect 18473 -41439 18519 -41039
rect 18571 -41439 18617 -41039
rect 19110 -41439 19156 -41039
rect 19321 -41439 19367 -41039
rect 19419 -41439 19465 -41039
rect 19517 -41439 19563 -41039
rect 19610 -41067 19670 -41007
rect 19733 -41185 19775 -40303
rect 19928 -40866 19974 -40566
rect 20026 -40866 20072 -40566
rect 20124 -40866 20170 -40566
rect 20238 -40865 20284 -40565
rect 20336 -40865 20382 -40565
rect 20434 -40865 20480 -40565
rect 20547 -40865 20593 -40565
rect 20645 -40865 20691 -40565
rect 20743 -40865 20789 -40565
rect 21058 -40765 21104 -40565
rect 21156 -40765 21202 -40565
rect 21347 -40954 21407 -40269
rect 21486 -40310 21546 -39886
rect 21935 -40165 21981 -39765
rect 22131 -40165 22177 -39765
rect 22310 -40218 22367 -39696
rect 25638 -39707 25793 -37318
rect 22506 -39777 25793 -39707
rect 22506 -39956 22576 -39777
rect 21486 -40311 21827 -40310
rect 21486 -40369 21828 -40311
rect 22281 -40352 22367 -40218
rect 21486 -40370 21827 -40369
rect 21308 -41014 21439 -40954
rect 21486 -41124 21546 -40370
rect 21837 -40619 21883 -40419
rect 21935 -40619 21981 -40419
rect 22047 -40619 22093 -40419
rect 22145 -40619 22191 -40419
rect 22667 -40510 22713 -39810
rect 22765 -40510 22811 -39810
rect 23067 -40510 23113 -39810
rect 23165 -40510 23211 -39810
rect 23550 -40507 23620 -39777
rect 23667 -40510 23713 -39810
rect 23765 -40510 23811 -39810
rect 24067 -40510 24113 -39810
rect 24165 -40510 24211 -39810
rect 24541 -40508 24611 -39777
rect 24667 -40510 24713 -39810
rect 24765 -40510 24811 -39810
rect 25067 -40510 25113 -39810
rect 25165 -40510 25211 -39810
rect 23279 -40560 23397 -40548
rect 23279 -40594 23486 -40560
rect 25252 -40567 25370 -40563
rect 25803 -40567 25924 -40544
rect 23279 -40606 23397 -40594
rect 21787 -41086 21833 -40986
rect 21885 -41086 21931 -40986
rect 21983 -41086 22029 -40986
rect 22081 -41086 22127 -40986
rect 22179 -41086 22225 -40986
rect 22277 -41086 22323 -40986
rect 21486 -41184 21813 -41124
rect 19725 -41317 19785 -41185
rect 20026 -41473 20072 -41273
rect 20222 -41473 20268 -41273
rect 20418 -41473 20464 -41273
rect 21156 -41473 21202 -41273
rect 21885 -41466 21931 -41266
rect 22081 -41466 22127 -41266
rect 22277 -41466 22323 -41266
rect 22765 -41395 22811 -40695
rect 23165 -41395 23211 -40695
rect 23452 -41495 23486 -40594
rect 24356 -40633 24474 -40575
rect 25252 -40612 25924 -40567
rect 25252 -40621 25370 -40612
rect 23765 -41395 23811 -40695
rect 24165 -41395 24211 -40695
rect 24362 -41430 24396 -40633
rect 24765 -41395 24811 -40695
rect 25165 -41395 25211 -40695
rect 24362 -41464 25670 -41430
rect 23452 -41529 25582 -41495
rect 11362 -42451 11408 -42251
rect 11558 -42451 11604 -42251
rect 11754 -42451 11800 -42251
rect 12029 -42504 12086 -42269
rect 12244 -42451 12290 -42251
rect 12440 -42451 12486 -42251
rect 12636 -42451 12682 -42251
rect 12855 -42366 12901 -42266
rect 12953 -42366 12999 -42266
rect 13051 -42366 13097 -42266
rect 13149 -42366 13195 -42266
rect 13247 -42366 13293 -42266
rect 13345 -42366 13391 -42266
rect 13443 -42366 13489 -42266
rect 13541 -42366 13587 -42266
rect 13987 -42451 14033 -42251
rect 14183 -42451 14229 -42251
rect 14379 -42451 14425 -42251
rect 12858 -42504 13027 -42494
rect 11264 -42731 11310 -42631
rect 11362 -42731 11408 -42631
rect 11460 -42731 11506 -42631
rect 11558 -42731 11604 -42631
rect 11656 -42731 11702 -42631
rect 11754 -42731 11800 -42631
rect 11888 -42662 11948 -42530
rect 12029 -42561 13027 -42504
rect 14729 -42504 14786 -42269
rect 14944 -42451 14990 -42251
rect 15140 -42451 15186 -42251
rect 15336 -42451 15382 -42251
rect 15555 -42366 15601 -42266
rect 15653 -42366 15699 -42266
rect 15751 -42366 15797 -42266
rect 15849 -42366 15895 -42266
rect 15947 -42366 15993 -42266
rect 16045 -42366 16091 -42266
rect 16143 -42366 16189 -42266
rect 16241 -42366 16287 -42266
rect 16687 -42451 16733 -42251
rect 16883 -42451 16929 -42251
rect 17079 -42451 17125 -42251
rect 15558 -42504 15727 -42494
rect 11537 -42851 11674 -42791
rect 11544 -43060 11639 -42851
rect 11888 -42890 11946 -42662
rect 11847 -42950 11979 -42890
rect 12029 -42998 12086 -42561
rect 12858 -42568 13027 -42561
rect 12146 -42731 12192 -42631
rect 12244 -42731 12290 -42631
rect 12342 -42731 12388 -42631
rect 12440 -42731 12486 -42631
rect 12538 -42731 12584 -42631
rect 12636 -42731 12682 -42631
rect 12855 -42781 12901 -42681
rect 12953 -42781 12999 -42681
rect 13051 -42781 13097 -42681
rect 13149 -42781 13195 -42681
rect 13247 -42781 13293 -42681
rect 13345 -42781 13391 -42681
rect 13443 -42781 13489 -42681
rect 13538 -42781 13587 -42681
rect 13889 -42731 13935 -42631
rect 13987 -42731 14033 -42631
rect 14085 -42731 14131 -42631
rect 14183 -42731 14229 -42631
rect 14281 -42731 14327 -42631
rect 14379 -42731 14425 -42631
rect 14505 -42641 14565 -42554
rect 14504 -42686 14565 -42641
rect 12956 -42878 12998 -42781
rect 13152 -42878 13194 -42781
rect 13347 -42878 13389 -42781
rect 13538 -42878 13584 -42781
rect 14164 -42852 14301 -42792
rect 11820 -43055 12086 -42998
rect 12824 -42924 13584 -42878
rect 11524 -43120 11656 -43060
rect 11820 -43176 11877 -43055
rect 12824 -43090 12870 -42924
rect 12059 -43091 12870 -43090
rect 10909 -43233 11877 -43176
rect 12051 -43136 12870 -43091
rect -7300 -46786 -7164 -46650
rect 10909 -47023 11109 -43233
rect 12051 -43411 12097 -43136
rect 12147 -43339 12193 -43239
rect 12245 -43339 12291 -43239
rect 12343 -43339 12389 -43239
rect 12441 -43339 12487 -43239
rect 12539 -43339 12585 -43239
rect 12637 -43339 12683 -43239
rect 12735 -43339 12781 -43239
rect 12833 -43339 12879 -43239
rect 13052 -43389 13098 -43289
rect 13150 -43389 13196 -43289
rect 13248 -43389 13294 -43289
rect 13346 -43389 13392 -43289
rect 13444 -43389 13490 -43289
rect 13542 -43389 13588 -43289
rect 14188 -43060 14283 -42852
rect 14157 -43120 14294 -43060
rect 13889 -43389 13935 -43289
rect 13987 -43389 14033 -43289
rect 14085 -43389 14131 -43289
rect 14183 -43389 14229 -43289
rect 14281 -43389 14327 -43289
rect 14379 -43389 14425 -43289
rect 12051 -43471 12205 -43411
rect 14504 -43434 14564 -42686
rect 14729 -42561 15727 -42504
rect 15558 -42568 15727 -42561
rect 14846 -42731 14892 -42631
rect 14944 -42731 14990 -42631
rect 15042 -42731 15088 -42631
rect 15140 -42731 15186 -42631
rect 15238 -42731 15284 -42631
rect 15336 -42731 15382 -42631
rect 15555 -42781 15601 -42681
rect 15653 -42762 15699 -42681
rect 15649 -42880 15710 -42762
rect 15751 -42781 15797 -42681
rect 15849 -42760 15895 -42681
rect 15840 -42880 15901 -42760
rect 15947 -42781 15993 -42681
rect 16045 -42762 16091 -42681
rect 16036 -42880 16097 -42762
rect 16143 -42781 16189 -42681
rect 16241 -42726 16287 -42681
rect 16241 -42880 16289 -42726
rect 16589 -42731 16635 -42631
rect 16687 -42731 16733 -42631
rect 16785 -42731 16831 -42631
rect 16883 -42731 16929 -42631
rect 16981 -42731 17027 -42631
rect 17079 -42731 17125 -42631
rect 16768 -42848 16900 -42788
rect 14758 -42928 16289 -42880
rect 14758 -43413 14799 -42928
rect 16370 -42948 16502 -42888
rect 14847 -43339 14893 -43239
rect 14945 -43339 14991 -43239
rect 15043 -43339 15089 -43239
rect 15141 -43339 15187 -43239
rect 15239 -43339 15285 -43239
rect 15337 -43339 15383 -43239
rect 15435 -43339 15481 -43239
rect 15533 -43339 15579 -43239
rect 15752 -43389 15798 -43289
rect 15850 -43389 15896 -43289
rect 15948 -43389 15994 -43289
rect 16046 -43389 16092 -43289
rect 16144 -43389 16190 -43289
rect 16242 -43389 16288 -43289
rect 12707 -43459 12876 -43452
rect 12707 -43516 13705 -43459
rect 14421 -43494 14564 -43434
rect 14757 -43473 14894 -43413
rect 16406 -43415 16466 -42948
rect 16781 -43066 16876 -42848
rect 17179 -42944 17239 -42918
rect 17179 -43008 17635 -42944
rect 17179 -43055 17239 -43008
rect 16754 -43126 16891 -43066
rect 16589 -43389 16635 -43289
rect 16687 -43389 16733 -43289
rect 16785 -43389 16831 -43289
rect 16883 -43389 16929 -43289
rect 16981 -43389 17027 -43289
rect 17079 -43389 17125 -43289
rect 15407 -43459 15576 -43452
rect 14758 -43474 14799 -43473
rect 14504 -43500 14564 -43494
rect 12707 -43526 12876 -43516
rect 12147 -43754 12193 -43654
rect 12245 -43754 12291 -43654
rect 12343 -43754 12389 -43654
rect 12441 -43754 12487 -43654
rect 12539 -43754 12585 -43654
rect 12637 -43754 12683 -43654
rect 12735 -43754 12781 -43654
rect 12833 -43754 12879 -43654
rect 13052 -43769 13098 -43569
rect 13248 -43769 13294 -43569
rect 13444 -43769 13490 -43569
rect 13648 -43751 13705 -43516
rect 15407 -43516 16405 -43459
rect 15407 -43526 15576 -43516
rect 13889 -43769 13935 -43569
rect 14085 -43769 14131 -43569
rect 14281 -43769 14327 -43569
rect 14847 -43754 14893 -43654
rect 14945 -43754 14991 -43654
rect 15043 -43754 15089 -43654
rect 15141 -43754 15187 -43654
rect 15239 -43754 15285 -43654
rect 15337 -43754 15383 -43654
rect 15435 -43754 15481 -43654
rect 15533 -43754 15579 -43654
rect 15752 -43769 15798 -43569
rect 15948 -43769 15994 -43569
rect 16144 -43769 16190 -43569
rect 16348 -43751 16405 -43516
rect 16589 -43769 16635 -43569
rect 16785 -43769 16831 -43569
rect 16981 -43769 17027 -43569
rect 17507 -46650 17635 -43008
rect 25009 -43700 25079 -41529
rect 25636 -41592 25670 -41464
rect 24890 -43920 25261 -43700
rect 25575 -44249 25696 -41592
rect 17502 -46786 17635 -46650
rect 24295 -44370 25696 -44249
rect 24295 -47213 24416 -44370
rect 25803 -46611 25924 -40612
rect 26597 -40181 26766 -36533
rect 28622 -36798 29061 -36751
rect 28622 -36835 28669 -36798
rect 27462 -37308 27592 -37158
rect 27748 -37212 27794 -37012
rect 27846 -37240 27892 -37012
rect 27944 -37212 27990 -37012
rect 28042 -37240 28088 -37012
rect 28623 -37134 28669 -36835
rect 28721 -37134 28767 -36834
rect 28819 -37134 28865 -36798
rect 27748 -37286 28385 -37240
rect 27512 -38712 27566 -37308
rect 27748 -37542 27794 -37286
rect 27846 -37288 28088 -37286
rect 27944 -37542 27990 -37288
rect 28140 -37542 28186 -37286
rect 28721 -37671 28767 -37371
rect 28917 -37671 28963 -36834
rect 29015 -37134 29061 -36798
rect 29717 -37306 30425 -37193
rect 29330 -37441 29376 -37341
rect 29428 -37470 29474 -37341
rect 29526 -37441 29572 -37341
rect 29624 -37470 29670 -37341
rect 29330 -37516 29967 -37470
rect 29330 -37672 29376 -37516
rect 29428 -37518 29670 -37516
rect 29526 -37672 29572 -37518
rect 29722 -37672 29768 -37516
rect 27722 -38571 27768 -38271
rect 27369 -38766 27566 -38712
rect 27624 -39107 27670 -38808
rect 27623 -39144 27670 -39107
rect 27722 -39108 27768 -38808
rect 27820 -39144 27866 -38808
rect 27918 -39108 27964 -38271
rect 28331 -38426 28377 -38270
rect 28527 -38424 28573 -38270
rect 28429 -38426 28671 -38424
rect 28723 -38426 28769 -38270
rect 28331 -38472 28968 -38426
rect 28331 -38601 28377 -38501
rect 28429 -38601 28475 -38472
rect 28527 -38601 28573 -38501
rect 28625 -38601 28671 -38472
rect 29169 -38782 29215 -38182
rect 29380 -38782 29426 -38182
rect 29478 -38782 29524 -38182
rect 29576 -38782 29622 -38182
rect 29788 -38782 29834 -38182
rect 28016 -39144 28062 -38808
rect 30019 -38913 30124 -38841
rect 30025 -38996 30090 -38913
rect 29070 -39061 30090 -38996
rect 27623 -39191 28062 -39144
rect 29169 -39394 29215 -39094
rect 29267 -39394 29313 -39094
rect 29365 -39394 29411 -39094
rect 29607 -39394 29653 -39094
rect 29705 -39394 29751 -39094
rect 29938 -39502 30051 -39501
rect 30312 -39502 30425 -37306
rect 31161 -38540 31207 -38040
rect 31430 -38540 31476 -38040
rect 31528 -38540 31574 -38040
rect 31626 -38540 31672 -38040
rect 31756 -38540 31802 -38040
rect 32082 -38540 32128 -38040
rect 32310 -38340 32356 -38040
rect 30930 -38700 31068 -38696
rect 31736 -38700 31874 -38696
rect 32121 -38700 32175 -38627
rect 30930 -38744 32175 -38700
rect 30930 -38750 31068 -38744
rect 31736 -38750 31874 -38744
rect 32121 -38765 32175 -38744
rect 32293 -38780 32359 -38768
rect 32893 -38780 33062 -36533
rect 34169 -36655 34418 -35421
rect 34580 -36481 41662 -36290
rect 34078 -36791 34435 -36655
rect 34078 -36845 34441 -36791
rect 34078 -36922 34435 -36845
rect 30769 -39087 30872 -38996
rect 29748 -39615 30425 -39502
rect 26597 -40267 26947 -40181
rect 28614 -40251 29053 -40204
rect 26597 -40321 28325 -40267
rect 28614 -40288 28661 -40251
rect 26597 -40350 26947 -40321
rect 27454 -40761 27584 -40611
rect 27740 -40665 27786 -40465
rect 27838 -40693 27884 -40465
rect 27936 -40665 27982 -40465
rect 28034 -40693 28080 -40465
rect 28271 -40611 28325 -40321
rect 28615 -40587 28661 -40288
rect 28713 -40587 28759 -40287
rect 28811 -40587 28857 -40251
rect 28271 -40665 28599 -40611
rect 27740 -40739 28377 -40693
rect 28545 -40720 28599 -40665
rect 27504 -42165 27558 -40761
rect 27740 -40995 27786 -40739
rect 27838 -40741 28080 -40739
rect 27936 -40995 27982 -40741
rect 28132 -40995 28178 -40739
rect 28519 -40778 28678 -40720
rect 28713 -41124 28759 -40824
rect 28909 -41124 28955 -40287
rect 29007 -40587 29053 -40251
rect 29938 -40646 30051 -39615
rect 30781 -39720 30860 -39087
rect 31063 -39336 31109 -39036
rect 31161 -39336 31207 -39036
rect 31533 -39336 31579 -38836
rect 31631 -39336 31677 -38836
rect 31756 -39336 31802 -38836
rect 31854 -39336 31900 -38836
rect 31984 -39336 32030 -38836
rect 32082 -39336 32128 -38836
rect 32180 -39336 32226 -38836
rect 32293 -38842 33915 -38780
rect 32293 -38851 32359 -38842
rect 32310 -39336 32356 -39036
rect 32408 -39336 32454 -39036
rect 30281 -39799 30860 -39720
rect 30281 -40154 30360 -39799
rect 30255 -40251 30371 -40154
rect 32282 -40282 32721 -40235
rect 30884 -40298 30981 -40292
rect 30884 -40352 31993 -40298
rect 32282 -40319 32329 -40282
rect 30884 -40358 30981 -40352
rect 29709 -40759 30417 -40646
rect 29322 -40894 29368 -40794
rect 29420 -40923 29466 -40794
rect 29518 -40894 29564 -40794
rect 29616 -40923 29662 -40794
rect 29322 -40969 29959 -40923
rect 29322 -41125 29368 -40969
rect 29420 -40971 29662 -40969
rect 29518 -41125 29564 -40971
rect 29714 -41125 29760 -40969
rect 27714 -42024 27760 -41724
rect 27361 -42219 27558 -42165
rect 27616 -42560 27662 -42261
rect 27615 -42597 27662 -42560
rect 27714 -42561 27760 -42261
rect 27812 -42597 27858 -42261
rect 27910 -42561 27956 -41724
rect 28323 -41879 28369 -41723
rect 28519 -41877 28565 -41723
rect 28421 -41879 28663 -41877
rect 28715 -41879 28761 -41723
rect 28323 -41925 28960 -41879
rect 28323 -42054 28369 -41954
rect 28421 -42054 28467 -41925
rect 28519 -42054 28565 -41954
rect 28617 -42054 28663 -41925
rect 29161 -42235 29207 -41635
rect 29372 -42235 29418 -41635
rect 29470 -42235 29516 -41635
rect 29568 -42235 29614 -41635
rect 29780 -42235 29826 -41635
rect 28008 -42597 28054 -42261
rect 30011 -42366 30116 -42294
rect 30017 -42449 30082 -42366
rect 29062 -42514 30082 -42449
rect 27615 -42644 28054 -42597
rect 29161 -42847 29207 -42547
rect 29259 -42847 29305 -42547
rect 29357 -42847 29403 -42547
rect 29599 -42847 29645 -42547
rect 29697 -42847 29743 -42547
rect 30304 -42955 30417 -40759
rect 31122 -40792 31252 -40642
rect 31408 -40696 31454 -40496
rect 31506 -40724 31552 -40496
rect 31604 -40696 31650 -40496
rect 31702 -40724 31748 -40496
rect 31939 -40642 31993 -40352
rect 32283 -40618 32329 -40319
rect 32381 -40618 32427 -40318
rect 32479 -40618 32525 -40282
rect 31939 -40696 32267 -40642
rect 31408 -40770 32045 -40724
rect 32213 -40751 32267 -40696
rect 31172 -42196 31226 -40792
rect 31408 -41026 31454 -40770
rect 31506 -40772 31748 -40770
rect 31604 -41026 31650 -40772
rect 31800 -41026 31846 -40770
rect 32187 -40809 32346 -40751
rect 32381 -41155 32427 -40855
rect 32577 -41155 32623 -40318
rect 32675 -40618 32721 -40282
rect 33377 -40790 34085 -40677
rect 32990 -40925 33036 -40825
rect 33088 -40954 33134 -40825
rect 33186 -40925 33232 -40825
rect 33284 -40954 33330 -40825
rect 32990 -41000 33627 -40954
rect 32990 -41156 33036 -41000
rect 33088 -41002 33330 -41000
rect 33186 -41156 33232 -41002
rect 33382 -41156 33428 -41000
rect 31382 -42055 31428 -41755
rect 31029 -42250 31226 -42196
rect 31284 -42591 31330 -42292
rect 31283 -42628 31330 -42591
rect 31382 -42592 31428 -42292
rect 31480 -42628 31526 -42292
rect 31578 -42592 31624 -41755
rect 31991 -41910 32037 -41754
rect 32187 -41908 32233 -41754
rect 32089 -41910 32331 -41908
rect 32383 -41910 32429 -41754
rect 31991 -41956 32628 -41910
rect 31991 -42085 32037 -41985
rect 32089 -42085 32135 -41956
rect 32187 -42085 32233 -41985
rect 32285 -42085 32331 -41956
rect 32829 -42266 32875 -41666
rect 33040 -42266 33086 -41666
rect 33138 -42266 33184 -41666
rect 33236 -42266 33282 -41666
rect 33448 -42266 33494 -41666
rect 31676 -42628 31722 -42292
rect 33679 -42397 33784 -42325
rect 33685 -42480 33750 -42397
rect 32730 -42545 33750 -42480
rect 31283 -42675 31722 -42628
rect 32829 -42878 32875 -42578
rect 32927 -42878 32973 -42578
rect 33025 -42878 33071 -42578
rect 33267 -42878 33313 -42578
rect 33365 -42878 33411 -42578
rect 29740 -42986 30417 -42955
rect 33972 -42986 34085 -40790
rect 34169 -42411 34418 -36922
rect 34580 -40195 34771 -36481
rect 35256 -36825 35613 -36689
rect 37062 -36809 37501 -36762
rect 35256 -36879 36773 -36825
rect 37062 -36846 37109 -36809
rect 35256 -36956 35613 -36879
rect 35902 -37319 36032 -37169
rect 36188 -37223 36234 -37023
rect 36286 -37251 36332 -37023
rect 36384 -37223 36430 -37023
rect 36482 -37251 36528 -37023
rect 36719 -37169 36773 -36879
rect 37063 -37145 37109 -36846
rect 37161 -37145 37207 -36845
rect 37259 -37145 37305 -36809
rect 36719 -37223 37047 -37169
rect 36188 -37297 36825 -37251
rect 36993 -37278 37047 -37223
rect 35952 -38723 36006 -37319
rect 36188 -37553 36234 -37297
rect 36286 -37299 36528 -37297
rect 36384 -37553 36430 -37299
rect 36580 -37553 36626 -37297
rect 36967 -37336 37126 -37278
rect 37161 -37682 37207 -37382
rect 37357 -37682 37403 -36845
rect 37455 -37145 37501 -36809
rect 38157 -37317 38865 -37204
rect 37770 -37452 37816 -37352
rect 37868 -37481 37914 -37352
rect 37966 -37452 38012 -37352
rect 38064 -37481 38110 -37352
rect 37770 -37527 38407 -37481
rect 37770 -37683 37816 -37527
rect 37868 -37529 38110 -37527
rect 37966 -37683 38012 -37529
rect 38162 -37683 38208 -37527
rect 36162 -38582 36208 -38282
rect 35809 -38777 36006 -38723
rect 36064 -39118 36110 -38819
rect 36063 -39155 36110 -39118
rect 36162 -39119 36208 -38819
rect 36260 -39155 36306 -38819
rect 36358 -39119 36404 -38282
rect 36771 -38437 36817 -38281
rect 36967 -38435 37013 -38281
rect 36869 -38437 37111 -38435
rect 37163 -38437 37209 -38281
rect 36771 -38483 37408 -38437
rect 36771 -38612 36817 -38512
rect 36869 -38612 36915 -38483
rect 36967 -38612 37013 -38512
rect 37065 -38612 37111 -38483
rect 37609 -38793 37655 -38193
rect 37820 -38793 37866 -38193
rect 37918 -38793 37964 -38193
rect 38016 -38793 38062 -38193
rect 38228 -38793 38274 -38193
rect 36456 -39155 36502 -38819
rect 38459 -38924 38564 -38852
rect 38465 -39007 38530 -38924
rect 37510 -39072 38530 -39007
rect 36063 -39202 36502 -39155
rect 37609 -39405 37655 -39105
rect 37707 -39405 37753 -39105
rect 37805 -39405 37851 -39105
rect 38047 -39405 38093 -39105
rect 38145 -39405 38191 -39105
rect 38378 -39513 38491 -39512
rect 38752 -39513 38865 -37317
rect 39601 -38551 39647 -38051
rect 39870 -38551 39916 -38051
rect 39968 -38551 40014 -38051
rect 40066 -38551 40112 -38051
rect 40196 -38551 40242 -38051
rect 40522 -38551 40568 -38051
rect 40750 -38351 40796 -38051
rect 39370 -38711 39508 -38707
rect 40176 -38711 40314 -38707
rect 40561 -38711 40615 -38638
rect 39370 -38755 40615 -38711
rect 39370 -38761 39508 -38755
rect 40176 -38761 40314 -38755
rect 40561 -38776 40615 -38755
rect 40733 -38791 40799 -38779
rect 41446 -38791 41662 -36481
rect 39209 -39098 39312 -39007
rect 38188 -39626 38865 -39513
rect 34580 -40278 35430 -40195
rect 37054 -40262 37493 -40215
rect 34580 -40332 36765 -40278
rect 37054 -40299 37101 -40262
rect 34580 -40386 35430 -40332
rect 35894 -40772 36024 -40622
rect 36180 -40676 36226 -40476
rect 36278 -40704 36324 -40476
rect 36376 -40676 36422 -40476
rect 36474 -40704 36520 -40476
rect 36711 -40622 36765 -40332
rect 37055 -40598 37101 -40299
rect 37153 -40598 37199 -40298
rect 37251 -40598 37297 -40262
rect 36711 -40676 37039 -40622
rect 36180 -40750 36817 -40704
rect 36985 -40731 37039 -40676
rect 35944 -42176 35998 -40772
rect 36180 -41006 36226 -40750
rect 36278 -40752 36520 -40750
rect 36376 -41006 36422 -40752
rect 36572 -41006 36618 -40750
rect 36959 -40789 37118 -40731
rect 37153 -41135 37199 -40835
rect 37349 -41135 37395 -40298
rect 37447 -40598 37493 -40262
rect 38378 -40657 38491 -39626
rect 39221 -39731 39300 -39098
rect 39503 -39347 39549 -39047
rect 39601 -39347 39647 -39047
rect 39973 -39347 40019 -38847
rect 40071 -39347 40117 -38847
rect 40196 -39347 40242 -38847
rect 40294 -39347 40340 -38847
rect 40424 -39347 40470 -38847
rect 40522 -39347 40568 -38847
rect 40620 -39347 40666 -38847
rect 40733 -38853 42355 -38791
rect 40733 -38862 40799 -38853
rect 40750 -39347 40796 -39047
rect 40848 -39347 40894 -39047
rect 38721 -39810 39300 -39731
rect 38721 -40165 38800 -39810
rect 38695 -40262 38811 -40165
rect 40722 -40293 41161 -40246
rect 39324 -40309 39421 -40303
rect 39324 -40363 40433 -40309
rect 40722 -40330 40769 -40293
rect 39324 -40369 39421 -40363
rect 38149 -40770 38857 -40657
rect 37762 -40905 37808 -40805
rect 37860 -40934 37906 -40805
rect 37958 -40905 38004 -40805
rect 38056 -40934 38102 -40805
rect 37762 -40980 38399 -40934
rect 37762 -41136 37808 -40980
rect 37860 -40982 38102 -40980
rect 37958 -41136 38004 -40982
rect 38154 -41136 38200 -40980
rect 36154 -42035 36200 -41735
rect 35801 -42230 35998 -42176
rect 34185 -42580 34408 -42411
rect 36056 -42571 36102 -42272
rect 36055 -42608 36102 -42571
rect 36154 -42572 36200 -42272
rect 36252 -42608 36298 -42272
rect 36350 -42572 36396 -41735
rect 36763 -41890 36809 -41734
rect 36959 -41888 37005 -41734
rect 36861 -41890 37103 -41888
rect 37155 -41890 37201 -41734
rect 36763 -41936 37400 -41890
rect 36763 -42065 36809 -41965
rect 36861 -42065 36907 -41936
rect 36959 -42065 37005 -41965
rect 37057 -42065 37103 -41936
rect 37601 -42246 37647 -41646
rect 37812 -42246 37858 -41646
rect 37910 -42246 37956 -41646
rect 38008 -42246 38054 -41646
rect 38220 -42246 38266 -41646
rect 36448 -42608 36494 -42272
rect 38451 -42377 38556 -42305
rect 38457 -42460 38522 -42377
rect 37502 -42525 38522 -42460
rect 36055 -42655 36494 -42608
rect 37601 -42858 37647 -42558
rect 37699 -42858 37745 -42558
rect 37797 -42858 37843 -42558
rect 38039 -42858 38085 -42558
rect 38137 -42858 38183 -42558
rect 38744 -42966 38857 -40770
rect 39562 -40803 39692 -40653
rect 39848 -40707 39894 -40507
rect 39946 -40735 39992 -40507
rect 40044 -40707 40090 -40507
rect 40142 -40735 40188 -40507
rect 40379 -40653 40433 -40363
rect 40723 -40629 40769 -40330
rect 40821 -40629 40867 -40329
rect 40919 -40629 40965 -40293
rect 40379 -40707 40707 -40653
rect 39848 -40781 40485 -40735
rect 40653 -40762 40707 -40707
rect 39612 -42207 39666 -40803
rect 39848 -41037 39894 -40781
rect 39946 -40783 40188 -40781
rect 40044 -41037 40090 -40783
rect 40240 -41037 40286 -40781
rect 40627 -40820 40786 -40762
rect 40821 -41166 40867 -40866
rect 41017 -41166 41063 -40329
rect 41115 -40629 41161 -40293
rect 41817 -40801 42525 -40688
rect 41430 -40936 41476 -40836
rect 41528 -40965 41574 -40836
rect 41626 -40936 41672 -40836
rect 41724 -40965 41770 -40836
rect 41430 -41011 42067 -40965
rect 41430 -41167 41476 -41011
rect 41528 -41013 41770 -41011
rect 41626 -41167 41672 -41013
rect 41822 -41167 41868 -41011
rect 39822 -42066 39868 -41766
rect 39469 -42261 39666 -42207
rect 39724 -42602 39770 -42303
rect 39723 -42639 39770 -42602
rect 39822 -42603 39868 -42303
rect 39920 -42639 39966 -42303
rect 40018 -42603 40064 -41766
rect 40431 -41921 40477 -41765
rect 40627 -41919 40673 -41765
rect 40529 -41921 40771 -41919
rect 40823 -41921 40869 -41765
rect 40431 -41967 41068 -41921
rect 40431 -42096 40477 -41996
rect 40529 -42096 40575 -41967
rect 40627 -42096 40673 -41996
rect 40725 -42096 40771 -41967
rect 41269 -42277 41315 -41677
rect 41480 -42277 41526 -41677
rect 41578 -42277 41624 -41677
rect 41676 -42277 41722 -41677
rect 41888 -42277 41934 -41677
rect 40116 -42639 40162 -42303
rect 42119 -42408 42224 -42336
rect 42125 -42491 42190 -42408
rect 41170 -42556 42190 -42491
rect 39723 -42686 40162 -42639
rect 41269 -42889 41315 -42589
rect 41367 -42889 41413 -42589
rect 41465 -42889 41511 -42589
rect 41707 -42889 41753 -42589
rect 41805 -42889 41851 -42589
rect 29740 -43068 34085 -42986
rect 29744 -43099 34085 -43068
rect 38180 -42997 38857 -42966
rect 42412 -42997 42525 -40801
rect 42634 -42348 42899 -35015
rect 43076 -36474 51037 -36272
rect 43076 -40264 43278 -36474
rect 44160 -36864 44457 -36778
rect 45925 -36848 46364 -36801
rect 44160 -36918 45636 -36864
rect 45925 -36885 45972 -36848
rect 44160 -37000 44457 -36918
rect 44765 -37358 44895 -37208
rect 45051 -37262 45097 -37062
rect 45149 -37290 45195 -37062
rect 45247 -37262 45293 -37062
rect 45345 -37290 45391 -37062
rect 45582 -37208 45636 -36918
rect 45926 -37184 45972 -36885
rect 46024 -37184 46070 -36884
rect 46122 -37184 46168 -36848
rect 45582 -37262 45910 -37208
rect 45051 -37336 45688 -37290
rect 45856 -37317 45910 -37262
rect 44815 -38762 44869 -37358
rect 45051 -37592 45097 -37336
rect 45149 -37338 45391 -37336
rect 45247 -37592 45293 -37338
rect 45443 -37592 45489 -37336
rect 45830 -37375 45989 -37317
rect 46024 -37721 46070 -37421
rect 46220 -37721 46266 -36884
rect 46318 -37184 46364 -36848
rect 47020 -37356 47728 -37243
rect 46633 -37491 46679 -37391
rect 46731 -37520 46777 -37391
rect 46829 -37491 46875 -37391
rect 46927 -37520 46973 -37391
rect 46633 -37566 47270 -37520
rect 46633 -37722 46679 -37566
rect 46731 -37568 46973 -37566
rect 46829 -37722 46875 -37568
rect 47025 -37722 47071 -37566
rect 45025 -38621 45071 -38321
rect 44672 -38816 44869 -38762
rect 44927 -39157 44973 -38858
rect 44926 -39194 44973 -39157
rect 45025 -39158 45071 -38858
rect 45123 -39194 45169 -38858
rect 45221 -39158 45267 -38321
rect 45634 -38476 45680 -38320
rect 45830 -38474 45876 -38320
rect 45732 -38476 45974 -38474
rect 46026 -38476 46072 -38320
rect 45634 -38522 46271 -38476
rect 45634 -38651 45680 -38551
rect 45732 -38651 45778 -38522
rect 45830 -38651 45876 -38551
rect 45928 -38651 45974 -38522
rect 46472 -38832 46518 -38232
rect 46683 -38832 46729 -38232
rect 46781 -38832 46827 -38232
rect 46879 -38832 46925 -38232
rect 47091 -38832 47137 -38232
rect 45319 -39194 45365 -38858
rect 47322 -38963 47427 -38891
rect 47328 -39046 47393 -38963
rect 46373 -39111 47393 -39046
rect 44926 -39241 45365 -39194
rect 46472 -39444 46518 -39144
rect 46570 -39444 46616 -39144
rect 46668 -39444 46714 -39144
rect 46910 -39444 46956 -39144
rect 47008 -39444 47054 -39144
rect 47241 -39552 47354 -39551
rect 47615 -39552 47728 -37356
rect 48464 -38590 48510 -38090
rect 48733 -38590 48779 -38090
rect 48831 -38590 48877 -38090
rect 48929 -38590 48975 -38090
rect 49059 -38590 49105 -38090
rect 49385 -38590 49431 -38090
rect 49613 -38390 49659 -38090
rect 48233 -38750 48371 -38746
rect 49039 -38750 49177 -38746
rect 49424 -38750 49478 -38677
rect 48233 -38794 49478 -38750
rect 48233 -38800 48371 -38794
rect 49039 -38800 49177 -38794
rect 49424 -38815 49478 -38794
rect 49596 -38830 49662 -38818
rect 50835 -38830 51037 -36474
rect 48072 -39137 48175 -39046
rect 47051 -39665 47728 -39552
rect 43076 -40317 44406 -40264
rect 45917 -40301 46356 -40254
rect 43076 -40371 45628 -40317
rect 45917 -40338 45964 -40301
rect 43076 -40466 44406 -40371
rect 44757 -40811 44887 -40661
rect 45043 -40715 45089 -40515
rect 45141 -40743 45187 -40515
rect 45239 -40715 45285 -40515
rect 45337 -40743 45383 -40515
rect 45574 -40661 45628 -40371
rect 45918 -40637 45964 -40338
rect 46016 -40637 46062 -40337
rect 46114 -40637 46160 -40301
rect 45574 -40715 45902 -40661
rect 45043 -40789 45680 -40743
rect 45848 -40770 45902 -40715
rect 44807 -42215 44861 -40811
rect 45043 -41045 45089 -40789
rect 45141 -40791 45383 -40789
rect 45239 -41045 45285 -40791
rect 45435 -41045 45481 -40789
rect 45822 -40828 45981 -40770
rect 46016 -41174 46062 -40874
rect 46212 -41174 46258 -40337
rect 46310 -40637 46356 -40301
rect 47241 -40696 47354 -39665
rect 48084 -39770 48163 -39137
rect 48366 -39386 48412 -39086
rect 48464 -39386 48510 -39086
rect 48836 -39386 48882 -38886
rect 48934 -39386 48980 -38886
rect 49059 -39386 49105 -38886
rect 49157 -39386 49203 -38886
rect 49287 -39386 49333 -38886
rect 49385 -39386 49431 -38886
rect 49483 -39386 49529 -38886
rect 49596 -38892 51218 -38830
rect 49596 -38901 49662 -38892
rect 49613 -39386 49659 -39086
rect 49711 -39386 49757 -39086
rect 47584 -39849 48163 -39770
rect 47584 -40204 47663 -39849
rect 47558 -40301 47674 -40204
rect 49585 -40332 50024 -40285
rect 48187 -40348 48284 -40342
rect 48187 -40402 49296 -40348
rect 49585 -40369 49632 -40332
rect 48187 -40408 48284 -40402
rect 47012 -40809 47720 -40696
rect 46625 -40944 46671 -40844
rect 46723 -40973 46769 -40844
rect 46821 -40944 46867 -40844
rect 46919 -40973 46965 -40844
rect 46625 -41019 47262 -40973
rect 46625 -41175 46671 -41019
rect 46723 -41021 46965 -41019
rect 46821 -41175 46867 -41021
rect 47017 -41175 47063 -41019
rect 45017 -42074 45063 -41774
rect 44664 -42269 44861 -42215
rect 42634 -42679 42971 -42348
rect 44919 -42610 44965 -42311
rect 44918 -42647 44965 -42610
rect 45017 -42611 45063 -42311
rect 45115 -42647 45161 -42311
rect 45213 -42611 45259 -41774
rect 45626 -41929 45672 -41773
rect 45822 -41927 45868 -41773
rect 45724 -41929 45966 -41927
rect 46018 -41929 46064 -41773
rect 45626 -41975 46263 -41929
rect 45626 -42104 45672 -42004
rect 45724 -42104 45770 -41975
rect 45822 -42104 45868 -42004
rect 45920 -42104 45966 -41975
rect 46464 -42285 46510 -41685
rect 46675 -42285 46721 -41685
rect 46773 -42285 46819 -41685
rect 46871 -42285 46917 -41685
rect 47083 -42285 47129 -41685
rect 45311 -42647 45357 -42311
rect 47314 -42416 47419 -42344
rect 47320 -42499 47385 -42416
rect 46365 -42564 47385 -42499
rect 44918 -42694 45357 -42647
rect 46464 -42897 46510 -42597
rect 46562 -42897 46608 -42597
rect 46660 -42897 46706 -42597
rect 46902 -42897 46948 -42597
rect 47000 -42897 47046 -42597
rect 38180 -43079 42525 -42997
rect 47607 -43005 47720 -40809
rect 48425 -40842 48555 -40692
rect 48711 -40746 48757 -40546
rect 48809 -40774 48855 -40546
rect 48907 -40746 48953 -40546
rect 49005 -40774 49051 -40546
rect 49242 -40692 49296 -40402
rect 49586 -40668 49632 -40369
rect 49684 -40668 49730 -40368
rect 49782 -40668 49828 -40332
rect 49242 -40746 49570 -40692
rect 48711 -40820 49348 -40774
rect 49516 -40801 49570 -40746
rect 48475 -42246 48529 -40842
rect 48711 -41076 48757 -40820
rect 48809 -40822 49051 -40820
rect 48907 -41076 48953 -40822
rect 49103 -41076 49149 -40820
rect 49490 -40859 49649 -40801
rect 49684 -41205 49730 -40905
rect 49880 -41205 49926 -40368
rect 49978 -40668 50024 -40332
rect 50680 -40840 51388 -40727
rect 50293 -40975 50339 -40875
rect 50391 -41004 50437 -40875
rect 50489 -40975 50535 -40875
rect 50587 -41004 50633 -40875
rect 50293 -41050 50930 -41004
rect 50293 -41206 50339 -41050
rect 50391 -41052 50633 -41050
rect 50489 -41206 50535 -41052
rect 50685 -41206 50731 -41050
rect 48685 -42105 48731 -41805
rect 48332 -42300 48529 -42246
rect 48587 -42641 48633 -42342
rect 48586 -42678 48633 -42641
rect 48685 -42642 48731 -42342
rect 48783 -42678 48829 -42342
rect 48881 -42642 48927 -41805
rect 49294 -41960 49340 -41804
rect 49490 -41958 49536 -41804
rect 49392 -41960 49634 -41958
rect 49686 -41960 49732 -41804
rect 49294 -42006 49931 -41960
rect 49294 -42135 49340 -42035
rect 49392 -42135 49438 -42006
rect 49490 -42135 49536 -42035
rect 49588 -42135 49634 -42006
rect 50132 -42316 50178 -41716
rect 50343 -42316 50389 -41716
rect 50441 -42316 50487 -41716
rect 50539 -42316 50585 -41716
rect 50751 -42316 50797 -41716
rect 48979 -42678 49025 -42342
rect 50982 -42447 51087 -42375
rect 50988 -42530 51053 -42447
rect 50033 -42595 51053 -42530
rect 48586 -42725 49025 -42678
rect 50132 -42928 50178 -42628
rect 50230 -42928 50276 -42628
rect 50328 -42928 50374 -42628
rect 50570 -42928 50616 -42628
rect 50668 -42928 50714 -42628
rect 38184 -43110 42525 -43079
rect 47043 -43036 47720 -43005
rect 51275 -43036 51388 -40840
rect 51498 -42209 51724 -34535
rect 52355 -36539 60341 -36280
rect 52355 -40143 52614 -36539
rect 53151 -36830 53397 -36734
rect 55123 -36814 55562 -36767
rect 53151 -36884 54834 -36830
rect 55123 -36851 55170 -36814
rect 53151 -36954 53397 -36884
rect 53963 -37324 54093 -37174
rect 54249 -37228 54295 -37028
rect 54347 -37256 54393 -37028
rect 54445 -37228 54491 -37028
rect 54543 -37256 54589 -37028
rect 54780 -37174 54834 -36884
rect 55124 -37150 55170 -36851
rect 55222 -37150 55268 -36850
rect 55320 -37150 55366 -36814
rect 54780 -37228 55108 -37174
rect 54249 -37302 54886 -37256
rect 55054 -37283 55108 -37228
rect 54013 -38728 54067 -37324
rect 54249 -37558 54295 -37302
rect 54347 -37304 54589 -37302
rect 54445 -37558 54491 -37304
rect 54641 -37558 54687 -37302
rect 55028 -37341 55187 -37283
rect 55222 -37687 55268 -37387
rect 55418 -37687 55464 -36850
rect 55516 -37150 55562 -36814
rect 56218 -37322 56926 -37209
rect 55831 -37457 55877 -37357
rect 55929 -37486 55975 -37357
rect 56027 -37457 56073 -37357
rect 56125 -37486 56171 -37357
rect 55831 -37532 56468 -37486
rect 55831 -37688 55877 -37532
rect 55929 -37534 56171 -37532
rect 56027 -37688 56073 -37534
rect 56223 -37688 56269 -37532
rect 54223 -38587 54269 -38287
rect 53870 -38782 54067 -38728
rect 54125 -39123 54171 -38824
rect 54124 -39160 54171 -39123
rect 54223 -39124 54269 -38824
rect 54321 -39160 54367 -38824
rect 54419 -39124 54465 -38287
rect 54832 -38442 54878 -38286
rect 55028 -38440 55074 -38286
rect 54930 -38442 55172 -38440
rect 55224 -38442 55270 -38286
rect 54832 -38488 55469 -38442
rect 54832 -38617 54878 -38517
rect 54930 -38617 54976 -38488
rect 55028 -38617 55074 -38517
rect 55126 -38617 55172 -38488
rect 55670 -38798 55716 -38198
rect 55881 -38798 55927 -38198
rect 55979 -38798 56025 -38198
rect 56077 -38798 56123 -38198
rect 56289 -38798 56335 -38198
rect 54517 -39160 54563 -38824
rect 56520 -38929 56625 -38857
rect 56526 -39012 56591 -38929
rect 55571 -39077 56591 -39012
rect 54124 -39207 54563 -39160
rect 55670 -39410 55716 -39110
rect 55768 -39410 55814 -39110
rect 55866 -39410 55912 -39110
rect 56108 -39410 56154 -39110
rect 56206 -39410 56252 -39110
rect 56439 -39518 56552 -39517
rect 56813 -39518 56926 -37322
rect 57662 -38556 57708 -38056
rect 57931 -38556 57977 -38056
rect 58029 -38556 58075 -38056
rect 58127 -38556 58173 -38056
rect 58257 -38556 58303 -38056
rect 58583 -38556 58629 -38056
rect 58811 -38356 58857 -38056
rect 57431 -38716 57569 -38712
rect 58237 -38716 58375 -38712
rect 58622 -38716 58676 -38643
rect 57431 -38760 58676 -38716
rect 57431 -38766 57569 -38760
rect 58237 -38766 58375 -38760
rect 58622 -38781 58676 -38760
rect 58794 -38796 58860 -38784
rect 60082 -38796 60341 -36539
rect 60692 -36596 60913 -33978
rect 61144 -36559 69128 -36321
rect 60589 -36910 60965 -36596
rect 57270 -39103 57373 -39012
rect 56249 -39631 56926 -39518
rect 52355 -40283 53563 -40143
rect 55115 -40267 55554 -40220
rect 52355 -40337 54826 -40283
rect 55115 -40304 55162 -40267
rect 52355 -40402 53563 -40337
rect 53955 -40777 54085 -40627
rect 54241 -40681 54287 -40481
rect 54339 -40709 54385 -40481
rect 54437 -40681 54483 -40481
rect 54535 -40709 54581 -40481
rect 54772 -40627 54826 -40337
rect 55116 -40603 55162 -40304
rect 55214 -40603 55260 -40303
rect 55312 -40603 55358 -40267
rect 54772 -40681 55100 -40627
rect 54241 -40755 54878 -40709
rect 55046 -40736 55100 -40681
rect 54005 -42181 54059 -40777
rect 54241 -41011 54287 -40755
rect 54339 -40757 54581 -40755
rect 54437 -41011 54483 -40757
rect 54633 -41011 54679 -40755
rect 55020 -40794 55179 -40736
rect 55214 -41140 55260 -40840
rect 55410 -41140 55456 -40303
rect 55508 -40603 55554 -40267
rect 56439 -40662 56552 -39631
rect 57282 -39736 57361 -39103
rect 57564 -39352 57610 -39052
rect 57662 -39352 57708 -39052
rect 58034 -39352 58080 -38852
rect 58132 -39352 58178 -38852
rect 58257 -39352 58303 -38852
rect 58355 -39352 58401 -38852
rect 58485 -39352 58531 -38852
rect 58583 -39352 58629 -38852
rect 58681 -39352 58727 -38852
rect 58794 -38858 60416 -38796
rect 58794 -38867 58860 -38858
rect 58811 -39352 58857 -39052
rect 58909 -39352 58955 -39052
rect 56782 -39815 57361 -39736
rect 56782 -40170 56861 -39815
rect 56756 -40267 56872 -40170
rect 58783 -40298 59222 -40251
rect 57385 -40314 57482 -40308
rect 57385 -40368 58494 -40314
rect 58783 -40335 58830 -40298
rect 57385 -40374 57482 -40368
rect 56210 -40775 56918 -40662
rect 55823 -40910 55869 -40810
rect 55921 -40939 55967 -40810
rect 56019 -40910 56065 -40810
rect 56117 -40939 56163 -40810
rect 55823 -40985 56460 -40939
rect 55823 -41141 55869 -40985
rect 55921 -40987 56163 -40985
rect 56019 -41141 56065 -40987
rect 56215 -41141 56261 -40985
rect 54215 -42040 54261 -41740
rect 51476 -42709 51774 -42209
rect 53862 -42235 54059 -42181
rect 54117 -42576 54163 -42277
rect 54116 -42613 54163 -42576
rect 54215 -42577 54261 -42277
rect 54313 -42613 54359 -42277
rect 54411 -42577 54457 -41740
rect 54824 -41895 54870 -41739
rect 55020 -41893 55066 -41739
rect 54922 -41895 55164 -41893
rect 55216 -41895 55262 -41739
rect 54824 -41941 55461 -41895
rect 54824 -42070 54870 -41970
rect 54922 -42070 54968 -41941
rect 55020 -42070 55066 -41970
rect 55118 -42070 55164 -41941
rect 55662 -42251 55708 -41651
rect 55873 -42251 55919 -41651
rect 55971 -42251 56017 -41651
rect 56069 -42251 56115 -41651
rect 56281 -42251 56327 -41651
rect 54509 -42613 54555 -42277
rect 56512 -42382 56617 -42310
rect 56518 -42465 56583 -42382
rect 55563 -42530 56583 -42465
rect 54116 -42660 54555 -42613
rect 55662 -42863 55708 -42563
rect 55760 -42863 55806 -42563
rect 55858 -42863 55904 -42563
rect 56100 -42863 56146 -42563
rect 56198 -42863 56244 -42563
rect 56805 -42971 56918 -40775
rect 57623 -40808 57753 -40658
rect 57909 -40712 57955 -40512
rect 58007 -40740 58053 -40512
rect 58105 -40712 58151 -40512
rect 58203 -40740 58249 -40512
rect 58440 -40658 58494 -40368
rect 58784 -40634 58830 -40335
rect 58882 -40634 58928 -40334
rect 58980 -40634 59026 -40298
rect 58440 -40712 58768 -40658
rect 57909 -40786 58546 -40740
rect 58714 -40767 58768 -40712
rect 57673 -42212 57727 -40808
rect 57909 -41042 57955 -40786
rect 58007 -40788 58249 -40786
rect 58105 -41042 58151 -40788
rect 58301 -41042 58347 -40786
rect 58688 -40825 58847 -40767
rect 58882 -41171 58928 -40871
rect 59078 -41171 59124 -40334
rect 59176 -40634 59222 -40298
rect 59878 -40806 60586 -40693
rect 59491 -40941 59537 -40841
rect 59589 -40970 59635 -40841
rect 59687 -40941 59733 -40841
rect 59785 -40970 59831 -40841
rect 59491 -41016 60128 -40970
rect 59491 -41172 59537 -41016
rect 59589 -41018 59831 -41016
rect 59687 -41172 59733 -41018
rect 59883 -41172 59929 -41016
rect 57883 -42071 57929 -41771
rect 57530 -42266 57727 -42212
rect 57785 -42607 57831 -42308
rect 57784 -42644 57831 -42607
rect 57883 -42608 57929 -42308
rect 57981 -42644 58027 -42308
rect 58079 -42608 58125 -41771
rect 58492 -41926 58538 -41770
rect 58688 -41924 58734 -41770
rect 58590 -41926 58832 -41924
rect 58884 -41926 58930 -41770
rect 58492 -41972 59129 -41926
rect 58492 -42101 58538 -42001
rect 58590 -42101 58636 -41972
rect 58688 -42101 58734 -42001
rect 58786 -42101 58832 -41972
rect 59330 -42282 59376 -41682
rect 59541 -42282 59587 -41682
rect 59639 -42282 59685 -41682
rect 59737 -42282 59783 -41682
rect 59949 -42282 59995 -41682
rect 58177 -42644 58223 -42308
rect 60180 -42413 60285 -42341
rect 60186 -42496 60251 -42413
rect 59231 -42561 60251 -42496
rect 57784 -42691 58223 -42644
rect 59330 -42894 59376 -42594
rect 59428 -42894 59474 -42594
rect 59526 -42894 59572 -42594
rect 59768 -42894 59814 -42594
rect 59866 -42894 59912 -42594
rect 47043 -43118 51388 -43036
rect 56241 -43002 56918 -42971
rect 60473 -43002 60586 -40806
rect 60692 -42347 60913 -36910
rect 61144 -40083 61382 -36559
rect 62190 -36764 62440 -36664
rect 63877 -36748 64316 -36701
rect 62190 -36818 63588 -36764
rect 63877 -36785 63924 -36748
rect 62190 -36893 62440 -36818
rect 62717 -37258 62847 -37108
rect 63003 -37162 63049 -36962
rect 63101 -37190 63147 -36962
rect 63199 -37162 63245 -36962
rect 63297 -37190 63343 -36962
rect 63534 -37108 63588 -36818
rect 63878 -37084 63924 -36785
rect 63976 -37084 64022 -36784
rect 64074 -37084 64120 -36748
rect 63534 -37162 63862 -37108
rect 63003 -37236 63640 -37190
rect 63808 -37217 63862 -37162
rect 62767 -38662 62821 -37258
rect 63003 -37492 63049 -37236
rect 63101 -37238 63343 -37236
rect 63199 -37492 63245 -37238
rect 63395 -37492 63441 -37236
rect 63782 -37275 63941 -37217
rect 63976 -37621 64022 -37321
rect 64172 -37621 64218 -36784
rect 64270 -37084 64316 -36748
rect 64972 -37256 65680 -37143
rect 64585 -37391 64631 -37291
rect 64683 -37420 64729 -37291
rect 64781 -37391 64827 -37291
rect 64879 -37420 64925 -37291
rect 64585 -37466 65222 -37420
rect 64585 -37622 64631 -37466
rect 64683 -37468 64925 -37466
rect 64781 -37622 64827 -37468
rect 64977 -37622 65023 -37466
rect 62977 -38521 63023 -38221
rect 62624 -38716 62821 -38662
rect 62879 -39057 62925 -38758
rect 62878 -39094 62925 -39057
rect 62977 -39058 63023 -38758
rect 63075 -39094 63121 -38758
rect 63173 -39058 63219 -38221
rect 63586 -38376 63632 -38220
rect 63782 -38374 63828 -38220
rect 63684 -38376 63926 -38374
rect 63978 -38376 64024 -38220
rect 63586 -38422 64223 -38376
rect 63586 -38551 63632 -38451
rect 63684 -38551 63730 -38422
rect 63782 -38551 63828 -38451
rect 63880 -38551 63926 -38422
rect 64424 -38732 64470 -38132
rect 64635 -38732 64681 -38132
rect 64733 -38732 64779 -38132
rect 64831 -38732 64877 -38132
rect 65043 -38732 65089 -38132
rect 63271 -39094 63317 -38758
rect 65274 -38863 65379 -38791
rect 65280 -38946 65345 -38863
rect 64325 -39011 65345 -38946
rect 62878 -39141 63317 -39094
rect 64424 -39344 64470 -39044
rect 64522 -39344 64568 -39044
rect 64620 -39344 64666 -39044
rect 64862 -39344 64908 -39044
rect 64960 -39344 65006 -39044
rect 65193 -39452 65306 -39451
rect 65567 -39452 65680 -37256
rect 66416 -38490 66462 -37990
rect 66685 -38490 66731 -37990
rect 66783 -38490 66829 -37990
rect 66881 -38490 66927 -37990
rect 67011 -38490 67057 -37990
rect 67337 -38490 67383 -37990
rect 67565 -38290 67611 -37990
rect 66185 -38650 66323 -38646
rect 66991 -38650 67129 -38646
rect 67376 -38650 67430 -38577
rect 66185 -38694 67430 -38650
rect 66185 -38700 66323 -38694
rect 66991 -38700 67129 -38694
rect 67376 -38715 67430 -38694
rect 67548 -38730 67614 -38718
rect 68890 -38730 69128 -36559
rect 69445 -36601 69622 -33419
rect 69930 -36567 78318 -36267
rect 69365 -36892 69703 -36601
rect 66024 -39037 66127 -38946
rect 65003 -39565 65680 -39452
rect 61144 -40217 62280 -40083
rect 63869 -40201 64308 -40154
rect 61144 -40271 63580 -40217
rect 63869 -40238 63916 -40201
rect 61144 -40321 62280 -40271
rect 62709 -40711 62839 -40561
rect 62995 -40615 63041 -40415
rect 63093 -40643 63139 -40415
rect 63191 -40615 63237 -40415
rect 63289 -40643 63335 -40415
rect 63526 -40561 63580 -40271
rect 63870 -40537 63916 -40238
rect 63968 -40537 64014 -40237
rect 64066 -40537 64112 -40201
rect 63526 -40615 63854 -40561
rect 62995 -40689 63632 -40643
rect 63800 -40670 63854 -40615
rect 62759 -42115 62813 -40711
rect 62995 -40945 63041 -40689
rect 63093 -40691 63335 -40689
rect 63191 -40945 63237 -40691
rect 63387 -40945 63433 -40689
rect 63774 -40728 63933 -40670
rect 63968 -41074 64014 -40774
rect 64164 -41074 64210 -40237
rect 64262 -40537 64308 -40201
rect 65193 -40596 65306 -39565
rect 66036 -39670 66115 -39037
rect 66318 -39286 66364 -38986
rect 66416 -39286 66462 -38986
rect 66788 -39286 66834 -38786
rect 66886 -39286 66932 -38786
rect 67011 -39286 67057 -38786
rect 67109 -39286 67155 -38786
rect 67239 -39286 67285 -38786
rect 67337 -39286 67383 -38786
rect 67435 -39286 67481 -38786
rect 67548 -38792 69170 -38730
rect 67548 -38801 67614 -38792
rect 67565 -39286 67611 -38986
rect 67663 -39286 67709 -38986
rect 65536 -39749 66115 -39670
rect 65536 -40104 65615 -39749
rect 65510 -40201 65626 -40104
rect 67537 -40232 67976 -40185
rect 66139 -40248 66236 -40242
rect 66139 -40302 67248 -40248
rect 67537 -40269 67584 -40232
rect 66139 -40308 66236 -40302
rect 64964 -40709 65672 -40596
rect 64577 -40844 64623 -40744
rect 64675 -40873 64721 -40744
rect 64773 -40844 64819 -40744
rect 64871 -40873 64917 -40744
rect 64577 -40919 65214 -40873
rect 64577 -41075 64623 -40919
rect 64675 -40921 64917 -40919
rect 64773 -41075 64819 -40921
rect 64969 -41075 65015 -40919
rect 62969 -41974 63015 -41674
rect 62616 -42169 62813 -42115
rect 60638 -42646 60930 -42347
rect 62871 -42510 62917 -42211
rect 62870 -42547 62917 -42510
rect 62969 -42511 63015 -42211
rect 63067 -42547 63113 -42211
rect 63165 -42511 63211 -41674
rect 63578 -41829 63624 -41673
rect 63774 -41827 63820 -41673
rect 63676 -41829 63918 -41827
rect 63970 -41829 64016 -41673
rect 63578 -41875 64215 -41829
rect 63578 -42004 63624 -41904
rect 63676 -42004 63722 -41875
rect 63774 -42004 63820 -41904
rect 63872 -42004 63918 -41875
rect 64416 -42185 64462 -41585
rect 64627 -42185 64673 -41585
rect 64725 -42185 64771 -41585
rect 64823 -42185 64869 -41585
rect 65035 -42185 65081 -41585
rect 63263 -42547 63309 -42211
rect 65266 -42316 65371 -42244
rect 65272 -42399 65337 -42316
rect 64317 -42464 65337 -42399
rect 62870 -42594 63309 -42547
rect 64416 -42797 64462 -42497
rect 64514 -42797 64560 -42497
rect 64612 -42797 64658 -42497
rect 64854 -42797 64900 -42497
rect 64952 -42797 64998 -42497
rect 65559 -42905 65672 -40709
rect 66377 -40742 66507 -40592
rect 66663 -40646 66709 -40446
rect 66761 -40674 66807 -40446
rect 66859 -40646 66905 -40446
rect 66957 -40674 67003 -40446
rect 67194 -40592 67248 -40302
rect 67538 -40568 67584 -40269
rect 67636 -40568 67682 -40268
rect 67734 -40568 67780 -40232
rect 67194 -40646 67522 -40592
rect 66663 -40720 67300 -40674
rect 67468 -40701 67522 -40646
rect 66427 -42146 66481 -40742
rect 66663 -40976 66709 -40720
rect 66761 -40722 67003 -40720
rect 66859 -40976 66905 -40722
rect 67055 -40976 67101 -40720
rect 67442 -40759 67601 -40701
rect 67636 -41105 67682 -40805
rect 67832 -41105 67878 -40268
rect 67930 -40568 67976 -40232
rect 68632 -40740 69340 -40627
rect 68245 -40875 68291 -40775
rect 68343 -40904 68389 -40775
rect 68441 -40875 68487 -40775
rect 68539 -40904 68585 -40775
rect 68245 -40950 68882 -40904
rect 68245 -41106 68291 -40950
rect 68343 -40952 68585 -40950
rect 68441 -41106 68487 -40952
rect 68637 -41106 68683 -40950
rect 66637 -42005 66683 -41705
rect 66284 -42200 66481 -42146
rect 66539 -42541 66585 -42242
rect 66538 -42578 66585 -42541
rect 66637 -42542 66683 -42242
rect 66735 -42578 66781 -42242
rect 66833 -42542 66879 -41705
rect 67246 -41860 67292 -41704
rect 67442 -41858 67488 -41704
rect 67344 -41860 67586 -41858
rect 67638 -41860 67684 -41704
rect 67246 -41906 67883 -41860
rect 67246 -42035 67292 -41935
rect 67344 -42035 67390 -41906
rect 67442 -42035 67488 -41935
rect 67540 -42035 67586 -41906
rect 68084 -42216 68130 -41616
rect 68295 -42216 68341 -41616
rect 68393 -42216 68439 -41616
rect 68491 -42216 68537 -41616
rect 68703 -42216 68749 -41616
rect 66931 -42578 66977 -42242
rect 68934 -42347 69039 -42275
rect 68940 -42430 69005 -42347
rect 67985 -42495 69005 -42430
rect 66538 -42625 66977 -42578
rect 68084 -42828 68130 -42528
rect 68182 -42828 68228 -42528
rect 68280 -42828 68326 -42528
rect 68522 -42828 68568 -42528
rect 68620 -42828 68666 -42528
rect 56241 -43084 60586 -43002
rect 64995 -42936 65672 -42905
rect 69227 -42936 69340 -40740
rect 69445 -42289 69622 -36892
rect 69930 -40017 70230 -36567
rect 71353 -36747 71621 -36656
rect 73030 -36731 73469 -36684
rect 71353 -36801 72741 -36747
rect 73030 -36768 73077 -36731
rect 71353 -36896 71621 -36801
rect 71870 -37241 72000 -37091
rect 72156 -37145 72202 -36945
rect 72254 -37173 72300 -36945
rect 72352 -37145 72398 -36945
rect 72450 -37173 72496 -36945
rect 72687 -37091 72741 -36801
rect 73031 -37067 73077 -36768
rect 73129 -37067 73175 -36767
rect 73227 -37067 73273 -36731
rect 72687 -37145 73015 -37091
rect 72156 -37219 72793 -37173
rect 72961 -37200 73015 -37145
rect 71920 -38645 71974 -37241
rect 72156 -37475 72202 -37219
rect 72254 -37221 72496 -37219
rect 72352 -37475 72398 -37221
rect 72548 -37475 72594 -37219
rect 72935 -37258 73094 -37200
rect 73129 -37604 73175 -37304
rect 73325 -37604 73371 -36767
rect 73423 -37067 73469 -36731
rect 74125 -37239 74833 -37126
rect 73738 -37374 73784 -37274
rect 73836 -37403 73882 -37274
rect 73934 -37374 73980 -37274
rect 74032 -37403 74078 -37274
rect 73738 -37449 74375 -37403
rect 73738 -37605 73784 -37449
rect 73836 -37451 74078 -37449
rect 73934 -37605 73980 -37451
rect 74130 -37605 74176 -37449
rect 72130 -38504 72176 -38204
rect 71777 -38699 71974 -38645
rect 72032 -39040 72078 -38741
rect 72031 -39077 72078 -39040
rect 72130 -39041 72176 -38741
rect 72228 -39077 72274 -38741
rect 72326 -39041 72372 -38204
rect 72739 -38359 72785 -38203
rect 72935 -38357 72981 -38203
rect 72837 -38359 73079 -38357
rect 73131 -38359 73177 -38203
rect 72739 -38405 73376 -38359
rect 72739 -38534 72785 -38434
rect 72837 -38534 72883 -38405
rect 72935 -38534 72981 -38434
rect 73033 -38534 73079 -38405
rect 73577 -38715 73623 -38115
rect 73788 -38715 73834 -38115
rect 73886 -38715 73932 -38115
rect 73984 -38715 74030 -38115
rect 74196 -38715 74242 -38115
rect 72424 -39077 72470 -38741
rect 74427 -38846 74532 -38774
rect 74433 -38929 74498 -38846
rect 73478 -38994 74498 -38929
rect 72031 -39124 72470 -39077
rect 73577 -39327 73623 -39027
rect 73675 -39327 73721 -39027
rect 73773 -39327 73819 -39027
rect 74015 -39327 74061 -39027
rect 74113 -39327 74159 -39027
rect 74346 -39435 74459 -39434
rect 74720 -39435 74833 -37239
rect 75569 -38473 75615 -37973
rect 75838 -38473 75884 -37973
rect 75936 -38473 75982 -37973
rect 76034 -38473 76080 -37973
rect 76164 -38473 76210 -37973
rect 76490 -38473 76536 -37973
rect 76718 -38273 76764 -37973
rect 75338 -38633 75476 -38629
rect 76144 -38633 76282 -38629
rect 76529 -38633 76583 -38560
rect 75338 -38677 76583 -38633
rect 75338 -38683 75476 -38677
rect 76144 -38683 76282 -38677
rect 76529 -38698 76583 -38677
rect 76701 -38713 76767 -38701
rect 78011 -38713 78318 -36567
rect 75177 -39020 75280 -38929
rect 74156 -39548 74833 -39435
rect 69930 -40200 71420 -40017
rect 73022 -40184 73461 -40137
rect 69930 -40254 72733 -40200
rect 73022 -40221 73069 -40184
rect 69930 -40317 71420 -40254
rect 71862 -40694 71992 -40544
rect 72148 -40598 72194 -40398
rect 72246 -40626 72292 -40398
rect 72344 -40598 72390 -40398
rect 72442 -40626 72488 -40398
rect 72679 -40544 72733 -40254
rect 73023 -40520 73069 -40221
rect 73121 -40520 73167 -40220
rect 73219 -40520 73265 -40184
rect 72679 -40598 73007 -40544
rect 72148 -40672 72785 -40626
rect 72953 -40653 73007 -40598
rect 71912 -42098 71966 -40694
rect 72148 -40928 72194 -40672
rect 72246 -40674 72488 -40672
rect 72344 -40928 72390 -40674
rect 72540 -40928 72586 -40672
rect 72927 -40711 73086 -40653
rect 73121 -41057 73167 -40757
rect 73317 -41057 73363 -40220
rect 73415 -40520 73461 -40184
rect 74346 -40579 74459 -39548
rect 75189 -39653 75268 -39020
rect 75471 -39269 75517 -38969
rect 75569 -39269 75615 -38969
rect 75941 -39269 75987 -38769
rect 76039 -39269 76085 -38769
rect 76164 -39269 76210 -38769
rect 76262 -39269 76308 -38769
rect 76392 -39269 76438 -38769
rect 76490 -39269 76536 -38769
rect 76588 -39269 76634 -38769
rect 76701 -38775 78323 -38713
rect 76701 -38784 76767 -38775
rect 76718 -39269 76764 -38969
rect 76816 -39269 76862 -38969
rect 74689 -39732 75268 -39653
rect 74689 -40087 74768 -39732
rect 74663 -40184 74779 -40087
rect 76690 -40215 77129 -40168
rect 75292 -40231 75389 -40225
rect 75292 -40285 76401 -40231
rect 76690 -40252 76737 -40215
rect 75292 -40291 75389 -40285
rect 74117 -40692 74825 -40579
rect 73730 -40827 73776 -40727
rect 73828 -40856 73874 -40727
rect 73926 -40827 73972 -40727
rect 74024 -40856 74070 -40727
rect 73730 -40902 74367 -40856
rect 73730 -41058 73776 -40902
rect 73828 -40904 74070 -40902
rect 73926 -41058 73972 -40904
rect 74122 -41058 74168 -40902
rect 72122 -41957 72168 -41657
rect 71769 -42152 71966 -42098
rect 69403 -42593 69664 -42289
rect 72024 -42493 72070 -42194
rect 72023 -42530 72070 -42493
rect 72122 -42494 72168 -42194
rect 72220 -42530 72266 -42194
rect 72318 -42494 72364 -41657
rect 72731 -41812 72777 -41656
rect 72927 -41810 72973 -41656
rect 72829 -41812 73071 -41810
rect 73123 -41812 73169 -41656
rect 72731 -41858 73368 -41812
rect 72731 -41987 72777 -41887
rect 72829 -41987 72875 -41858
rect 72927 -41987 72973 -41887
rect 73025 -41987 73071 -41858
rect 73569 -42168 73615 -41568
rect 73780 -42168 73826 -41568
rect 73878 -42168 73924 -41568
rect 73976 -42168 74022 -41568
rect 74188 -42168 74234 -41568
rect 72416 -42530 72462 -42194
rect 74419 -42299 74524 -42227
rect 74425 -42382 74490 -42299
rect 73470 -42447 74490 -42382
rect 72023 -42577 72462 -42530
rect 73569 -42780 73615 -42480
rect 73667 -42780 73713 -42480
rect 73765 -42780 73811 -42480
rect 74007 -42780 74053 -42480
rect 74105 -42780 74151 -42480
rect 74712 -42888 74825 -40692
rect 75530 -40725 75660 -40575
rect 75816 -40629 75862 -40429
rect 75914 -40657 75960 -40429
rect 76012 -40629 76058 -40429
rect 76110 -40657 76156 -40429
rect 76347 -40575 76401 -40285
rect 76691 -40551 76737 -40252
rect 76789 -40551 76835 -40251
rect 76887 -40551 76933 -40215
rect 76347 -40629 76675 -40575
rect 75816 -40703 76453 -40657
rect 76621 -40684 76675 -40629
rect 75580 -42129 75634 -40725
rect 75816 -40959 75862 -40703
rect 75914 -40705 76156 -40703
rect 76012 -40959 76058 -40705
rect 76208 -40959 76254 -40703
rect 76595 -40742 76754 -40684
rect 76789 -41088 76835 -40788
rect 76985 -41088 77031 -40251
rect 77083 -40551 77129 -40215
rect 77785 -40723 78493 -40610
rect 77398 -40858 77444 -40758
rect 77496 -40887 77542 -40758
rect 77594 -40858 77640 -40758
rect 77692 -40887 77738 -40758
rect 77398 -40933 78035 -40887
rect 77398 -41089 77444 -40933
rect 77496 -40935 77738 -40933
rect 77594 -41089 77640 -40935
rect 77790 -41089 77836 -40933
rect 75790 -41988 75836 -41688
rect 75437 -42183 75634 -42129
rect 75692 -42524 75738 -42225
rect 75691 -42561 75738 -42524
rect 75790 -42525 75836 -42225
rect 75888 -42561 75934 -42225
rect 75986 -42525 76032 -41688
rect 76399 -41843 76445 -41687
rect 76595 -41841 76641 -41687
rect 76497 -41843 76739 -41841
rect 76791 -41843 76837 -41687
rect 76399 -41889 77036 -41843
rect 76399 -42018 76445 -41918
rect 76497 -42018 76543 -41889
rect 76595 -42018 76641 -41918
rect 76693 -42018 76739 -41889
rect 77237 -42199 77283 -41599
rect 77448 -42199 77494 -41599
rect 77546 -42199 77592 -41599
rect 77644 -42199 77690 -41599
rect 77856 -42199 77902 -41599
rect 76084 -42561 76130 -42225
rect 78087 -42330 78192 -42258
rect 78093 -42413 78158 -42330
rect 77138 -42478 78158 -42413
rect 75691 -42608 76130 -42561
rect 77237 -42811 77283 -42511
rect 77335 -42811 77381 -42511
rect 77433 -42811 77479 -42511
rect 77675 -42811 77721 -42511
rect 77773 -42811 77819 -42511
rect 64995 -43018 69340 -42936
rect 74148 -42919 74825 -42888
rect 78380 -42919 78493 -40723
rect 78579 -42613 78890 -32969
rect 79155 -36485 87674 -36266
rect 79155 -40123 79374 -36485
rect 80608 -36709 80903 -36594
rect 82394 -36693 82833 -36646
rect 80608 -36763 82105 -36709
rect 82394 -36730 82441 -36693
rect 80608 -36867 80903 -36763
rect 81234 -37203 81364 -37053
rect 81520 -37107 81566 -36907
rect 81618 -37135 81664 -36907
rect 81716 -37107 81762 -36907
rect 81814 -37135 81860 -36907
rect 82051 -37053 82105 -36763
rect 82395 -37029 82441 -36730
rect 82493 -37029 82539 -36729
rect 82591 -37029 82637 -36693
rect 82051 -37107 82379 -37053
rect 81520 -37181 82157 -37135
rect 82325 -37162 82379 -37107
rect 81284 -38607 81338 -37203
rect 81520 -37437 81566 -37181
rect 81618 -37183 81860 -37181
rect 81716 -37437 81762 -37183
rect 81912 -37437 81958 -37181
rect 82299 -37220 82458 -37162
rect 82493 -37566 82539 -37266
rect 82689 -37566 82735 -36729
rect 82787 -37029 82833 -36693
rect 83489 -37201 84197 -37088
rect 83102 -37336 83148 -37236
rect 83200 -37365 83246 -37236
rect 83298 -37336 83344 -37236
rect 83396 -37365 83442 -37236
rect 83102 -37411 83739 -37365
rect 83102 -37567 83148 -37411
rect 83200 -37413 83442 -37411
rect 83298 -37567 83344 -37413
rect 83494 -37567 83540 -37411
rect 81494 -38466 81540 -38166
rect 81141 -38661 81338 -38607
rect 81396 -39002 81442 -38703
rect 81395 -39039 81442 -39002
rect 81494 -39003 81540 -38703
rect 81592 -39039 81638 -38703
rect 81690 -39003 81736 -38166
rect 82103 -38321 82149 -38165
rect 82299 -38319 82345 -38165
rect 82201 -38321 82443 -38319
rect 82495 -38321 82541 -38165
rect 82103 -38367 82740 -38321
rect 82103 -38496 82149 -38396
rect 82201 -38496 82247 -38367
rect 82299 -38496 82345 -38396
rect 82397 -38496 82443 -38367
rect 82941 -38677 82987 -38077
rect 83152 -38677 83198 -38077
rect 83250 -38677 83296 -38077
rect 83348 -38677 83394 -38077
rect 83560 -38677 83606 -38077
rect 81788 -39039 81834 -38703
rect 83791 -38808 83896 -38736
rect 83797 -38891 83862 -38808
rect 82842 -38956 83862 -38891
rect 81395 -39086 81834 -39039
rect 82941 -39289 82987 -38989
rect 83039 -39289 83085 -38989
rect 83137 -39289 83183 -38989
rect 83379 -39289 83425 -38989
rect 83477 -39289 83523 -38989
rect 83710 -39397 83823 -39396
rect 84084 -39397 84197 -37201
rect 84933 -38435 84979 -37935
rect 85202 -38435 85248 -37935
rect 85300 -38435 85346 -37935
rect 85398 -38435 85444 -37935
rect 85528 -38435 85574 -37935
rect 85854 -38435 85900 -37935
rect 86082 -38235 86128 -37935
rect 84702 -38595 84840 -38591
rect 85508 -38595 85646 -38591
rect 85893 -38595 85947 -38522
rect 84702 -38639 85947 -38595
rect 84702 -38645 84840 -38639
rect 85508 -38645 85646 -38639
rect 85893 -38660 85947 -38639
rect 86065 -38675 86131 -38663
rect 87455 -38675 87674 -36485
rect 84541 -38982 84644 -38891
rect 83520 -39510 84197 -39397
rect 79155 -40162 80934 -40123
rect 82386 -40146 82825 -40099
rect 79155 -40216 82097 -40162
rect 82386 -40183 82433 -40146
rect 79155 -40342 80934 -40216
rect 81226 -40656 81356 -40506
rect 81512 -40560 81558 -40360
rect 81610 -40588 81656 -40360
rect 81708 -40560 81754 -40360
rect 81806 -40588 81852 -40360
rect 82043 -40506 82097 -40216
rect 82387 -40482 82433 -40183
rect 82485 -40482 82531 -40182
rect 82583 -40482 82629 -40146
rect 82043 -40560 82371 -40506
rect 81512 -40634 82149 -40588
rect 82317 -40615 82371 -40560
rect 81276 -42060 81330 -40656
rect 81512 -40890 81558 -40634
rect 81610 -40636 81852 -40634
rect 81708 -40890 81754 -40636
rect 81904 -40890 81950 -40634
rect 82291 -40673 82450 -40615
rect 82485 -41019 82531 -40719
rect 82681 -41019 82727 -40182
rect 82779 -40482 82825 -40146
rect 83710 -40541 83823 -39510
rect 84553 -39615 84632 -38982
rect 84835 -39231 84881 -38931
rect 84933 -39231 84979 -38931
rect 85305 -39231 85351 -38731
rect 85403 -39231 85449 -38731
rect 85528 -39231 85574 -38731
rect 85626 -39231 85672 -38731
rect 85756 -39231 85802 -38731
rect 85854 -39231 85900 -38731
rect 85952 -39231 85998 -38731
rect 86065 -38737 87687 -38675
rect 86065 -38746 86131 -38737
rect 86082 -39231 86128 -38931
rect 86180 -39231 86226 -38931
rect 84053 -39694 84632 -39615
rect 84053 -40049 84132 -39694
rect 84027 -40146 84143 -40049
rect 86054 -40177 86493 -40130
rect 84656 -40193 84753 -40187
rect 84656 -40247 85765 -40193
rect 86054 -40214 86101 -40177
rect 84656 -40253 84753 -40247
rect 83481 -40654 84189 -40541
rect 83094 -40789 83140 -40689
rect 83192 -40818 83238 -40689
rect 83290 -40789 83336 -40689
rect 83388 -40818 83434 -40689
rect 83094 -40864 83731 -40818
rect 83094 -41020 83140 -40864
rect 83192 -40866 83434 -40864
rect 83290 -41020 83336 -40866
rect 83486 -41020 83532 -40864
rect 81486 -41919 81532 -41619
rect 81133 -42114 81330 -42060
rect 81388 -42455 81434 -42156
rect 81387 -42492 81434 -42455
rect 81486 -42456 81532 -42156
rect 81584 -42492 81630 -42156
rect 81682 -42456 81728 -41619
rect 82095 -41774 82141 -41618
rect 82291 -41772 82337 -41618
rect 82193 -41774 82435 -41772
rect 82487 -41774 82533 -41618
rect 82095 -41820 82732 -41774
rect 82095 -41949 82141 -41849
rect 82193 -41949 82239 -41820
rect 82291 -41949 82337 -41849
rect 82389 -41949 82435 -41820
rect 82933 -42130 82979 -41530
rect 83144 -42130 83190 -41530
rect 83242 -42130 83288 -41530
rect 83340 -42130 83386 -41530
rect 83552 -42130 83598 -41530
rect 81780 -42492 81826 -42156
rect 83783 -42261 83888 -42189
rect 83789 -42344 83854 -42261
rect 82834 -42409 83854 -42344
rect 81387 -42539 81826 -42492
rect 82933 -42742 82979 -42442
rect 83031 -42742 83077 -42442
rect 83129 -42742 83175 -42442
rect 83371 -42742 83417 -42442
rect 83469 -42742 83515 -42442
rect 84076 -42850 84189 -40654
rect 84894 -40687 85024 -40537
rect 85180 -40591 85226 -40391
rect 85278 -40619 85324 -40391
rect 85376 -40591 85422 -40391
rect 85474 -40619 85520 -40391
rect 85711 -40537 85765 -40247
rect 86055 -40513 86101 -40214
rect 86153 -40513 86199 -40213
rect 86251 -40513 86297 -40177
rect 85711 -40591 86039 -40537
rect 85180 -40665 85817 -40619
rect 85985 -40646 86039 -40591
rect 84944 -42091 84998 -40687
rect 85180 -40921 85226 -40665
rect 85278 -40667 85520 -40665
rect 85376 -40921 85422 -40667
rect 85572 -40921 85618 -40665
rect 85959 -40704 86118 -40646
rect 86153 -41050 86199 -40750
rect 86349 -41050 86395 -40213
rect 86447 -40513 86493 -40177
rect 87149 -40685 87857 -40572
rect 86762 -40820 86808 -40720
rect 86860 -40849 86906 -40720
rect 86958 -40820 87004 -40720
rect 87056 -40849 87102 -40720
rect 86762 -40895 87399 -40849
rect 86762 -41051 86808 -40895
rect 86860 -40897 87102 -40895
rect 86958 -41051 87004 -40897
rect 87154 -41051 87200 -40895
rect 85154 -41950 85200 -41650
rect 84801 -42145 84998 -42091
rect 85056 -42486 85102 -42187
rect 85055 -42523 85102 -42486
rect 85154 -42487 85200 -42187
rect 85252 -42523 85298 -42187
rect 85350 -42487 85396 -41650
rect 85763 -41805 85809 -41649
rect 85959 -41803 86005 -41649
rect 85861 -41805 86103 -41803
rect 86155 -41805 86201 -41649
rect 85763 -41851 86400 -41805
rect 85763 -41980 85809 -41880
rect 85861 -41980 85907 -41851
rect 85959 -41980 86005 -41880
rect 86057 -41980 86103 -41851
rect 86601 -42161 86647 -41561
rect 86812 -42161 86858 -41561
rect 86910 -42161 86956 -41561
rect 87008 -42161 87054 -41561
rect 87220 -42161 87266 -41561
rect 85448 -42523 85494 -42187
rect 87451 -42292 87556 -42220
rect 87457 -42375 87522 -42292
rect 86502 -42440 87522 -42375
rect 85055 -42570 85494 -42523
rect 86601 -42773 86647 -42473
rect 86699 -42773 86745 -42473
rect 86797 -42773 86843 -42473
rect 87039 -42773 87085 -42473
rect 87137 -42773 87183 -42473
rect 74148 -43001 78493 -42919
rect 83512 -42881 84189 -42850
rect 87744 -42881 87857 -40685
rect 88110 -42245 88394 -32036
rect 88080 -42588 88439 -42245
rect 83512 -42963 87857 -42881
rect 83516 -42994 87857 -42963
rect 64999 -43049 69340 -43018
rect 74152 -43032 78493 -43001
rect 56245 -43115 60586 -43084
rect 47047 -43149 51388 -43118
rect 42275 -43723 42592 -43640
rect 26575 -43904 35375 -43723
rect 42275 -43904 82025 -43723
rect 42275 -43931 42592 -43904
rect 42232 -44823 42601 -44446
rect 43552 -44744 82025 -44459
rect 42241 -46611 42541 -44823
rect 24763 -46911 42541 -46611
rect 43552 -47154 43837 -44744
rect 24558 -47213 43837 -47154
rect 24295 -47334 43837 -47213
rect 24558 -47439 43837 -47334
rect 13476 -50147 89097 -49863
rect -28640 -52302 -28240 -52256
rect -28640 -52420 -28240 -52374
rect -28640 -52538 -28240 -52492
rect -29536 -60594 -29081 -52616
rect -28640 -52656 -28240 -52610
rect -28640 -52774 -28240 -52728
rect -28640 -52892 -28240 -52846
rect -15203 -52837 9205 -52647
rect -28640 -53010 -28240 -52964
rect -28640 -53128 -28240 -53082
rect -28640 -53246 -28240 -53200
rect -28640 -53364 -28240 -53318
rect -28640 -53482 -28240 -53436
rect -28640 -53600 -28240 -53554
rect -28640 -53718 -28240 -53672
rect -28640 -53836 -28240 -53790
rect -28640 -53954 -28240 -53908
rect -28640 -54072 -28240 -54026
rect -28640 -54190 -28240 -54144
rect -28640 -54308 -28240 -54262
rect -28640 -54426 -28240 -54380
rect -28640 -54544 -28240 -54498
rect -28640 -54662 -28240 -54616
rect -28640 -54780 -28240 -54734
rect -28640 -54898 -28240 -54852
rect -28640 -55016 -28240 -54970
rect -28640 -55134 -28240 -55088
rect -28640 -55252 -28240 -55206
rect -28640 -55370 -28240 -55324
rect -28640 -55488 -28240 -55442
rect -28640 -55606 -28240 -55560
rect -28640 -55724 -28240 -55678
rect -28640 -55842 -28240 -55796
rect -28640 -56078 -28240 -56032
rect -28640 -56314 -28240 -56268
rect -28640 -56550 -28240 -56504
rect -28640 -56786 -28240 -56740
rect -28640 -57022 -28240 -56976
rect -28640 -57258 -28240 -57212
rect -28640 -57494 -28240 -57448
rect -27977 -56182 -27903 -56067
rect -27977 -56228 -27432 -56182
rect -27977 -56418 -27903 -56228
rect -27977 -56464 -27432 -56418
rect -27977 -56654 -27903 -56464
rect -27977 -56700 -27432 -56654
rect -27977 -56890 -27903 -56700
rect -27977 -56936 -27432 -56890
rect -27977 -57126 -27903 -56936
rect -27977 -57172 -27432 -57126
rect -27977 -57362 -27903 -57172
rect -27977 -57408 -27432 -57362
rect -27977 -57598 -27903 -57408
rect -27977 -57644 -27432 -57598
rect -28640 -57730 -28240 -57684
rect -28640 -57841 -28105 -57802
rect -27977 -57834 -27903 -57644
rect -27977 -57841 -27432 -57834
rect -28640 -57848 -27432 -57841
rect -28151 -57880 -27432 -57848
rect -28151 -57887 -27903 -57880
rect -28640 -57966 -28240 -57920
rect -28151 -58038 -28105 -57887
rect -27977 -58012 -27903 -57887
rect -28640 -58084 -28105 -58038
rect -28640 -58202 -28240 -58156
rect -28151 -58274 -28105 -58084
rect -28640 -58320 -28105 -58274
rect -28640 -58438 -28240 -58392
rect -28151 -58510 -28105 -58320
rect -28640 -58556 -28105 -58510
rect -27977 -58200 -27903 -58073
rect -27977 -58246 -27432 -58200
rect -27977 -58436 -27903 -58246
rect -27977 -58482 -27432 -58436
rect -28640 -58674 -28240 -58628
rect -27977 -58672 -27903 -58482
rect -27977 -58718 -27432 -58672
rect -28640 -58792 -28117 -58746
rect -28163 -58823 -28117 -58792
rect -27977 -58823 -27903 -58718
rect -28640 -58910 -28240 -58864
rect -28163 -58869 -27903 -58823
rect -28163 -58982 -28117 -58869
rect -28640 -59028 -28117 -58982
rect -27977 -58908 -27903 -58869
rect -27977 -58954 -27432 -58908
rect -27977 -59083 -27903 -58954
rect -28640 -59146 -28240 -59100
rect -27977 -59218 -27903 -59144
rect -28640 -59264 -27903 -59218
rect -27977 -59274 -27903 -59264
rect -27977 -59320 -27432 -59274
rect -28640 -59382 -28240 -59336
rect -27977 -59510 -27903 -59320
rect -27977 -59556 -27432 -59510
rect -27977 -59561 -27903 -59556
rect -27322 -60594 -26810 -60453
rect -29536 -61049 -26810 -60594
rect -27322 -61078 -26810 -61049
rect -21245 -54086 -21199 -53886
rect -21049 -54086 -21003 -53886
rect -20853 -54086 -20807 -53886
rect -20115 -54086 -20069 -53886
rect -15203 -53926 -15013 -52837
rect -13646 -53299 -13600 -53099
rect -13450 -53299 -13404 -53099
rect -13254 -53299 -13208 -53099
rect -13024 -53352 -12967 -53117
rect -12809 -53299 -12763 -53099
rect -12613 -53299 -12567 -53099
rect -12417 -53299 -12371 -53099
rect -12198 -53214 -12152 -53114
rect -12100 -53214 -12054 -53114
rect -12002 -53214 -11956 -53114
rect -11904 -53214 -11858 -53114
rect -11806 -53214 -11760 -53114
rect -11708 -53214 -11662 -53114
rect -11610 -53214 -11564 -53114
rect -11512 -53214 -11466 -53114
rect -10946 -53299 -10900 -53099
rect -10750 -53299 -10704 -53099
rect -10554 -53299 -10508 -53099
rect -12195 -53352 -12026 -53342
rect -13024 -53409 -12026 -53352
rect -10324 -53352 -10267 -53117
rect -10109 -53299 -10063 -53099
rect -9913 -53299 -9867 -53099
rect -9717 -53299 -9671 -53099
rect -9498 -53214 -9452 -53114
rect -9400 -53214 -9354 -53114
rect -9302 -53214 -9256 -53114
rect -9204 -53214 -9158 -53114
rect -9106 -53214 -9060 -53114
rect -9008 -53214 -8962 -53114
rect -8910 -53214 -8864 -53114
rect -8812 -53214 -8766 -53114
rect -9495 -53352 -9326 -53342
rect -11183 -53374 -11123 -53368
rect -11418 -53395 -11377 -53394
rect -12195 -53416 -12026 -53409
rect -13744 -53579 -13698 -53479
rect -13646 -53579 -13600 -53479
rect -13548 -53579 -13502 -53479
rect -13450 -53579 -13404 -53479
rect -13352 -53579 -13306 -53479
rect -13254 -53579 -13208 -53479
rect -13510 -53802 -13373 -53742
rect -13858 -53860 -13798 -53813
rect -14120 -53924 -13798 -53860
rect -19246 -54308 -19200 -54008
rect -19653 -54363 -19516 -54346
rect -19681 -54404 -19516 -54363
rect -21343 -54793 -21297 -54493
rect -21245 -54793 -21199 -54493
rect -21147 -54793 -21101 -54493
rect -21033 -54794 -20987 -54494
rect -20935 -54794 -20889 -54494
rect -20837 -54794 -20791 -54494
rect -20724 -54794 -20678 -54494
rect -20626 -54794 -20580 -54494
rect -20528 -54794 -20482 -54494
rect -20213 -54794 -20167 -54594
rect -20115 -54710 -20069 -54594
rect -20115 -54745 -19756 -54710
rect -20115 -54794 -20069 -54745
rect -21971 -63599 -21910 -55032
rect -22040 -63600 -21910 -63599
rect -22040 -63633 -21909 -63600
rect -22039 -63718 -21909 -63633
rect -21857 -63727 -21793 -56504
rect -21859 -63899 -21793 -63727
rect -21880 -63900 -21793 -63899
rect -21712 -60975 -21652 -56073
rect -21188 -56217 -21142 -55917
rect -21286 -56753 -21240 -56454
rect -21287 -56790 -21240 -56753
rect -21188 -56754 -21142 -56454
rect -21090 -56790 -21044 -56454
rect -20992 -56754 -20946 -55917
rect -20579 -56072 -20533 -55916
rect -20383 -56070 -20337 -55916
rect -20481 -56072 -20239 -56070
rect -20187 -56072 -20141 -55916
rect -20579 -56118 -19942 -56072
rect -20579 -56247 -20533 -56147
rect -20481 -56247 -20435 -56118
rect -20383 -56247 -20337 -56147
rect -20285 -56247 -20239 -56118
rect -19791 -56279 -19756 -54745
rect -19681 -55114 -19645 -54404
rect -19683 -55246 -19630 -55114
rect -19344 -54844 -19298 -54545
rect -19345 -54881 -19298 -54844
rect -19246 -54845 -19200 -54545
rect -19148 -54881 -19102 -54545
rect -19050 -54845 -19004 -54008
rect -18637 -54163 -18591 -54007
rect -18441 -54161 -18395 -54007
rect -18539 -54163 -18297 -54161
rect -18245 -54163 -18199 -54007
rect -15584 -54039 -14907 -53926
rect -18637 -54209 -18000 -54163
rect -18637 -54338 -18591 -54238
rect -18539 -54338 -18493 -54209
rect -18441 -54338 -18395 -54238
rect -18343 -54338 -18297 -54209
rect -17917 -54234 -17771 -54176
rect -17917 -54260 -17836 -54234
rect -18229 -54295 -17836 -54260
rect -18952 -54881 -18906 -54545
rect -19345 -54928 -18906 -54881
rect -18229 -55365 -18194 -54295
rect -17709 -54397 -17270 -54350
rect -17709 -54434 -17662 -54397
rect -17708 -54733 -17662 -54434
rect -17610 -54733 -17564 -54433
rect -17512 -54733 -17466 -54397
rect -17963 -54829 -17766 -54775
rect -19725 -55400 -18194 -55365
rect -19725 -56148 -19690 -55400
rect -19415 -56022 -19369 -55822
rect -19219 -56022 -19173 -55822
rect -19023 -56022 -18977 -55822
rect -18285 -56022 -18239 -55822
rect -19725 -56194 -19641 -56148
rect -20894 -56790 -20848 -56454
rect -20010 -56513 -19952 -56376
rect -19796 -56416 -19738 -56279
rect -19699 -56285 -19641 -56194
rect -17820 -56233 -17766 -54829
rect -17610 -55270 -17564 -54970
rect -17414 -55270 -17368 -54433
rect -17316 -54733 -17270 -54397
rect -16163 -54447 -16117 -54147
rect -16065 -54447 -16019 -54147
rect -15967 -54447 -15921 -54147
rect -15725 -54447 -15679 -54147
rect -15627 -54447 -15581 -54147
rect -16262 -54545 -15242 -54480
rect -15307 -54628 -15242 -54545
rect -15313 -54700 -15208 -54628
rect -17001 -55040 -16955 -54940
rect -16903 -55069 -16857 -54940
rect -16805 -55040 -16759 -54940
rect -16707 -55069 -16661 -54940
rect -17001 -55115 -16364 -55069
rect -17001 -55271 -16955 -55115
rect -16903 -55117 -16661 -55115
rect -16805 -55271 -16759 -55117
rect -16609 -55271 -16563 -55115
rect -16163 -55359 -16117 -54759
rect -15952 -55359 -15906 -54759
rect -15854 -55359 -15808 -54759
rect -15756 -55359 -15710 -54759
rect -15544 -55359 -15498 -54759
rect -17870 -56383 -17740 -56233
rect -17584 -56255 -17538 -55999
rect -17388 -56253 -17342 -55999
rect -17486 -56255 -17244 -56253
rect -17192 -56255 -17146 -55999
rect -16611 -56170 -16565 -55870
rect -17584 -56301 -16947 -56255
rect -16805 -56274 -16646 -56216
rect -19513 -56729 -19467 -56429
rect -19415 -56729 -19369 -56429
rect -19317 -56729 -19271 -56429
rect -19203 -56730 -19157 -56430
rect -19105 -56730 -19059 -56430
rect -19007 -56730 -18961 -56430
rect -18894 -56730 -18848 -56430
rect -18796 -56730 -18750 -56430
rect -18698 -56730 -18652 -56430
rect -17584 -56529 -17538 -56329
rect -17486 -56529 -17440 -56301
rect -17388 -56529 -17342 -56329
rect -17290 -56529 -17244 -56301
rect -16779 -56329 -16725 -56274
rect -17053 -56383 -16725 -56329
rect -18383 -56730 -18337 -56530
rect -18285 -56730 -18239 -56530
rect -17053 -56673 -16999 -56383
rect -18096 -56727 -16999 -56673
rect -16709 -56706 -16663 -56407
rect -21287 -56837 -20848 -56790
rect -18084 -57441 -17844 -56727
rect -16710 -56743 -16663 -56706
rect -16611 -56707 -16565 -56407
rect -16513 -56743 -16467 -56407
rect -16415 -56707 -16369 -55870
rect -16002 -56025 -15956 -55869
rect -15806 -56023 -15760 -55869
rect -15904 -56025 -15662 -56023
rect -15610 -56025 -15564 -55869
rect -16002 -56071 -15365 -56025
rect -16002 -56200 -15956 -56100
rect -15904 -56200 -15858 -56071
rect -15806 -56200 -15760 -56100
rect -15708 -56200 -15662 -56071
rect -15020 -56235 -14907 -54039
rect -14120 -55840 -14056 -53924
rect -13858 -53950 -13798 -53924
rect -13495 -54020 -13400 -53802
rect -13085 -53920 -13025 -53453
rect -11513 -53455 -11376 -53395
rect -11183 -53434 -11040 -53374
rect -10324 -53409 -9326 -53352
rect -9495 -53416 -9326 -53409
rect -12907 -53579 -12861 -53479
rect -12809 -53579 -12763 -53479
rect -12711 -53579 -12665 -53479
rect -12613 -53579 -12567 -53479
rect -12515 -53579 -12469 -53479
rect -12417 -53579 -12371 -53479
rect -12198 -53629 -12152 -53529
rect -12100 -53629 -12054 -53529
rect -12002 -53629 -11956 -53529
rect -11904 -53629 -11858 -53529
rect -11806 -53629 -11760 -53529
rect -11708 -53629 -11662 -53529
rect -11610 -53629 -11564 -53529
rect -11512 -53629 -11466 -53529
rect -13121 -53980 -12989 -53920
rect -11418 -53940 -11377 -53455
rect -11348 -53891 -11211 -53831
rect -12908 -53988 -11377 -53940
rect -13519 -54080 -13387 -54020
rect -13744 -54237 -13698 -54137
rect -13646 -54237 -13600 -54137
rect -13548 -54237 -13502 -54137
rect -13450 -54237 -13404 -54137
rect -13352 -54237 -13306 -54137
rect -13254 -54237 -13208 -54137
rect -12908 -54142 -12860 -53988
rect -12906 -54187 -12860 -54142
rect -12808 -54187 -12762 -54087
rect -12716 -54106 -12655 -53988
rect -12710 -54187 -12664 -54106
rect -12612 -54187 -12566 -54087
rect -12520 -54108 -12459 -53988
rect -12514 -54187 -12468 -54108
rect -12416 -54187 -12370 -54087
rect -12329 -54106 -12268 -53988
rect -12318 -54187 -12272 -54106
rect -12220 -54187 -12174 -54087
rect -12001 -54237 -11955 -54137
rect -11903 -54237 -11857 -54137
rect -11805 -54237 -11759 -54137
rect -11707 -54237 -11661 -54137
rect -11609 -54237 -11563 -54137
rect -11511 -54237 -11465 -54137
rect -12346 -54307 -12177 -54300
rect -12346 -54364 -11348 -54307
rect -11299 -54339 -11239 -53891
rect -11183 -54182 -11123 -53434
rect -8824 -53457 -8670 -53397
rect -11044 -53579 -10998 -53479
rect -10946 -53579 -10900 -53479
rect -10848 -53579 -10802 -53479
rect -10750 -53579 -10704 -53479
rect -10652 -53579 -10606 -53479
rect -10554 -53579 -10508 -53479
rect -10913 -53808 -10776 -53748
rect -10902 -54016 -10807 -53808
rect -10373 -53832 -10313 -53468
rect -10207 -53579 -10161 -53479
rect -10109 -53579 -10063 -53479
rect -10011 -53579 -9965 -53479
rect -9913 -53579 -9867 -53479
rect -9815 -53579 -9769 -53479
rect -9717 -53579 -9671 -53479
rect -9498 -53629 -9452 -53529
rect -9400 -53629 -9354 -53529
rect -9302 -53629 -9256 -53529
rect -9204 -53629 -9158 -53529
rect -9106 -53629 -9060 -53529
rect -9008 -53629 -8962 -53529
rect -8910 -53629 -8864 -53529
rect -8812 -53629 -8766 -53529
rect -8716 -53732 -8670 -53457
rect -9489 -53777 -8670 -53732
rect -9489 -53778 -8678 -53777
rect -10402 -53892 -10270 -53832
rect -9489 -53944 -9443 -53778
rect -8275 -53808 -8143 -53748
rect -8258 -53873 -8163 -53808
rect -7723 -53873 -7628 -52837
rect -7480 -53709 -7434 -53109
rect -7268 -53709 -7222 -53109
rect -7170 -53709 -7124 -53109
rect -7072 -53709 -7026 -53109
rect -6861 -53709 -6815 -53109
rect -6050 -53505 -6004 -53305
rect -5952 -53505 -5906 -53305
rect -5854 -53505 -5808 -53305
rect -5734 -53505 -5688 -53305
rect -5636 -53505 -5590 -53305
rect -5538 -53505 -5492 -53305
rect -5176 -53505 -5130 -53305
rect -4980 -53505 -4934 -53305
rect -4670 -53505 -4624 -53305
rect -4361 -53505 -4315 -53305
rect -3550 -53505 -3504 -53305
rect -3452 -53505 -3406 -53305
rect -3354 -53505 -3308 -53305
rect -3234 -53505 -3188 -53305
rect -3136 -53505 -3090 -53305
rect -3038 -53505 -2992 -53305
rect -2676 -53505 -2630 -53305
rect -2480 -53505 -2434 -53305
rect -2170 -53505 -2124 -53305
rect -1861 -53505 -1815 -53305
rect -1050 -53505 -1004 -53305
rect -952 -53505 -906 -53305
rect -854 -53505 -808 -53305
rect -734 -53505 -688 -53305
rect -636 -53505 -590 -53305
rect -538 -53505 -492 -53305
rect -176 -53505 -130 -53305
rect 20 -53505 66 -53305
rect 330 -53505 376 -53305
rect 639 -53505 685 -53305
rect 1450 -53505 1496 -53305
rect 1548 -53505 1594 -53305
rect 1646 -53505 1692 -53305
rect 1766 -53505 1812 -53305
rect 1864 -53505 1910 -53305
rect 1962 -53505 2008 -53305
rect 2324 -53505 2370 -53305
rect 2520 -53505 2566 -53305
rect 2830 -53505 2876 -53305
rect 3139 -53505 3185 -53305
rect 3950 -53505 3996 -53305
rect 4048 -53505 4094 -53305
rect 4146 -53505 4192 -53305
rect 4266 -53505 4312 -53305
rect 4364 -53505 4410 -53305
rect 4462 -53505 4508 -53305
rect 4824 -53505 4870 -53305
rect 5020 -53505 5066 -53305
rect 5330 -53505 5376 -53305
rect 5639 -53505 5685 -53305
rect 6950 -53505 6996 -53305
rect 7048 -53505 7094 -53305
rect 7146 -53505 7192 -53305
rect 7266 -53505 7312 -53305
rect 7364 -53505 7410 -53305
rect 7462 -53505 7508 -53305
rect 7824 -53505 7870 -53305
rect 8020 -53505 8066 -53305
rect 8330 -53505 8376 -53305
rect 8639 -53505 8685 -53305
rect -4887 -53633 -4748 -53615
rect -4272 -53633 -4133 -53621
rect -2387 -53633 -2248 -53615
rect -1772 -53633 -1633 -53621
rect 113 -53633 252 -53615
rect 728 -53633 867 -53621
rect 2613 -53633 2752 -53615
rect 3228 -53633 3367 -53621
rect 5113 -53633 5252 -53615
rect 5728 -53633 5867 -53621
rect 8113 -53633 8252 -53615
rect 8728 -53633 8867 -53621
rect 9429 -53633 9629 -53281
rect -6045 -53672 -5906 -53659
rect -4887 -53661 -3982 -53633
rect -4887 -53669 -4748 -53661
rect -6045 -53700 -5691 -53672
rect -4272 -53675 -4133 -53661
rect -6045 -53713 -5906 -53700
rect -10203 -53990 -9443 -53944
rect -8598 -53978 -8466 -53918
rect -8258 -53968 -7628 -53873
rect -10920 -54076 -10783 -54016
rect -10203 -54087 -10157 -53990
rect -10008 -54087 -9966 -53990
rect -9813 -54087 -9771 -53990
rect -9617 -54087 -9575 -53990
rect -11184 -54227 -11123 -54182
rect -11184 -54314 -11124 -54227
rect -11044 -54237 -10998 -54137
rect -10946 -54237 -10900 -54137
rect -10848 -54237 -10802 -54137
rect -10750 -54237 -10704 -54137
rect -10652 -54237 -10606 -54137
rect -10554 -54237 -10508 -54137
rect -10206 -54187 -10157 -54087
rect -10108 -54187 -10062 -54087
rect -10010 -54187 -9964 -54087
rect -9912 -54187 -9866 -54087
rect -9814 -54187 -9768 -54087
rect -9716 -54187 -9670 -54087
rect -9618 -54187 -9572 -54087
rect -9520 -54187 -9474 -54087
rect -9301 -54237 -9255 -54137
rect -9203 -54237 -9157 -54137
rect -9105 -54237 -9059 -54137
rect -9007 -54237 -8961 -54137
rect -8909 -54237 -8863 -54137
rect -8811 -54237 -8765 -54137
rect -8565 -54206 -8507 -53978
rect -8258 -54017 -8163 -53968
rect -8293 -54077 -8156 -54017
rect -9646 -54307 -9477 -54300
rect -12346 -54374 -12177 -54364
rect -13744 -54617 -13698 -54417
rect -13548 -54617 -13502 -54417
rect -13352 -54617 -13306 -54417
rect -12906 -54570 -12860 -54502
rect -12906 -54602 -12855 -54570
rect -12808 -54602 -12762 -54502
rect -12710 -54545 -12664 -54502
rect -12905 -54685 -12855 -54602
rect -12714 -54685 -12663 -54545
rect -12612 -54602 -12566 -54502
rect -12514 -54564 -12468 -54502
rect -12514 -54685 -12463 -54564
rect -12416 -54602 -12370 -54502
rect -12318 -54564 -12272 -54502
rect -12320 -54685 -12269 -54564
rect -12220 -54602 -12174 -54502
rect -12001 -54617 -11955 -54417
rect -11805 -54617 -11759 -54417
rect -11609 -54617 -11563 -54417
rect -11405 -54599 -11348 -54364
rect -9646 -54364 -8648 -54307
rect -8567 -54338 -8507 -54206
rect -8419 -54237 -8373 -54137
rect -8321 -54237 -8275 -54137
rect -8223 -54237 -8177 -54137
rect -8125 -54237 -8079 -54137
rect -8027 -54237 -7981 -54137
rect -7929 -54237 -7883 -54137
rect -9646 -54374 -9477 -54364
rect -11044 -54617 -10998 -54417
rect -10848 -54617 -10802 -54417
rect -10652 -54617 -10606 -54417
rect -10206 -54602 -10160 -54502
rect -10108 -54602 -10062 -54502
rect -10010 -54602 -9964 -54502
rect -9912 -54602 -9866 -54502
rect -9814 -54602 -9768 -54502
rect -9716 -54602 -9670 -54502
rect -9618 -54602 -9572 -54502
rect -9520 -54602 -9474 -54502
rect -9301 -54617 -9255 -54417
rect -9105 -54617 -9059 -54417
rect -8909 -54617 -8863 -54417
rect -8705 -54685 -8648 -54364
rect -8419 -54617 -8373 -54417
rect -8223 -54617 -8177 -54417
rect -8027 -54617 -7981 -54417
rect -12905 -54742 -8648 -54685
rect -7723 -54902 -7628 -53968
rect -7397 -54321 -7351 -54021
rect -7299 -54321 -7253 -54021
rect -7057 -54321 -7011 -54021
rect -6959 -54321 -6913 -54021
rect -6861 -54321 -6815 -54021
rect -10595 -55015 -7627 -54902
rect -12720 -55373 -12281 -55326
rect -12720 -55410 -12673 -55373
rect -12719 -55709 -12673 -55410
rect -12621 -55709 -12575 -55409
rect -12523 -55709 -12477 -55373
rect -13258 -55840 -13072 -55798
rect -14120 -55904 -13072 -55840
rect -13258 -55952 -13072 -55904
rect -15615 -56348 -14907 -56235
rect -16317 -56743 -16271 -56407
rect -16710 -56790 -16271 -56743
rect -15698 -57099 -15430 -56834
rect -15649 -57654 -15461 -57099
rect -15693 -57919 -15425 -57654
rect -21123 -59711 -21077 -59111
rect -20911 -59711 -20865 -59111
rect -20813 -59711 -20767 -59111
rect -20715 -59711 -20669 -59111
rect -20602 -59711 -20556 -59111
rect -20504 -59711 -20458 -59111
rect -20406 -59711 -20360 -59111
rect -19917 -59440 -19871 -59040
rect -19706 -59440 -19660 -59040
rect -19608 -59440 -19562 -59040
rect -19510 -59440 -19464 -59040
rect -19012 -59441 -18966 -59041
rect -18801 -59441 -18755 -59041
rect -18703 -59441 -18657 -59041
rect -18605 -59441 -18559 -59041
rect -20385 -60037 -20248 -59979
rect -21123 -60275 -21077 -60075
rect -21025 -60275 -20979 -60075
rect -20927 -60275 -20881 -60075
rect -20829 -60275 -20783 -60075
rect -21257 -60521 -20453 -60371
rect -21245 -60933 -21158 -60521
rect -21065 -60933 -20978 -60521
rect -20892 -60933 -20805 -60521
rect -20708 -60933 -20621 -60521
rect -20583 -60933 -20496 -60521
rect -21470 -60975 -20487 -60933
rect -21712 -61035 -20487 -60975
rect -21880 -64023 -21757 -63900
rect -21712 -64267 -21652 -61035
rect -21470 -61048 -20487 -61035
rect -20373 -61035 -20283 -60037
rect -19273 -59603 -19215 -59466
rect -20114 -59640 -20056 -59636
rect -20115 -59773 -20056 -59640
rect -19498 -59688 -19361 -59630
rect -20115 -60590 -20072 -59773
rect -19917 -59932 -19871 -59732
rect -19819 -59932 -19773 -59732
rect -19721 -59932 -19675 -59732
rect -20116 -60727 -20058 -60590
rect -20373 -61125 -20056 -61035
rect -21460 -61421 -21414 -61221
rect -21362 -61421 -21316 -61221
rect -21047 -61521 -21001 -61221
rect -20949 -61521 -20903 -61221
rect -20851 -61521 -20805 -61221
rect -20738 -61521 -20692 -61221
rect -20640 -61521 -20594 -61221
rect -20542 -61521 -20496 -61221
rect -20428 -61522 -20382 -61222
rect -20330 -61522 -20284 -61222
rect -20232 -61522 -20186 -61222
rect -20146 -61713 -20056 -61125
rect -19407 -61658 -19372 -59688
rect -19273 -60669 -19238 -59603
rect -19196 -59775 -19138 -59638
rect -18567 -59689 -18430 -59631
rect -19295 -60806 -19237 -60669
rect -19196 -60746 -19161 -59775
rect -19012 -59933 -18966 -59733
rect -18914 -59933 -18868 -59733
rect -18816 -59933 -18770 -59733
rect -19202 -60883 -19144 -60746
rect -19415 -61795 -19357 -61658
rect -21460 -62129 -21414 -61929
rect -20722 -62129 -20676 -61929
rect -20526 -62129 -20480 -61929
rect -20330 -62129 -20284 -61929
rect -21459 -62400 -21416 -62129
rect -18482 -61744 -18447 -59689
rect -18306 -59987 -18189 -59864
rect -18405 -61392 -18347 -61255
rect -18490 -61881 -18432 -61744
rect -21509 -62516 -21351 -62400
rect -18404 -62428 -18365 -61392
rect -18303 -62251 -18211 -59987
rect -15020 -58926 -14907 -56348
rect -12621 -56246 -12575 -55946
rect -12425 -56246 -12379 -55409
rect -12327 -55709 -12281 -55373
rect -11174 -55423 -11128 -55123
rect -11076 -55423 -11030 -55123
rect -10978 -55423 -10932 -55123
rect -10736 -55423 -10690 -55123
rect -10638 -55423 -10592 -55123
rect -11273 -55521 -10253 -55456
rect -10318 -55604 -10253 -55521
rect -10324 -55676 -10219 -55604
rect -12012 -56016 -11966 -55916
rect -11914 -56045 -11868 -55916
rect -11816 -56016 -11770 -55916
rect -11718 -56045 -11672 -55916
rect -12012 -56091 -11375 -56045
rect -12012 -56247 -11966 -56091
rect -11914 -56093 -11672 -56091
rect -11816 -56247 -11770 -56093
rect -11620 -56247 -11574 -56091
rect -11174 -56335 -11128 -55735
rect -10963 -56335 -10917 -55735
rect -10865 -56335 -10819 -55735
rect -10767 -56335 -10721 -55735
rect -10555 -56335 -10509 -55735
rect -15584 -59039 -14907 -58926
rect -17709 -59397 -17270 -59350
rect -17709 -59434 -17662 -59397
rect -17708 -59733 -17662 -59434
rect -17610 -59733 -17564 -59433
rect -17512 -59733 -17466 -59397
rect -17963 -59829 -17766 -59775
rect -17820 -61233 -17766 -59829
rect -17610 -60270 -17564 -59970
rect -17414 -60270 -17368 -59433
rect -17316 -59733 -17270 -59397
rect -16163 -59447 -16117 -59147
rect -16065 -59447 -16019 -59147
rect -15967 -59447 -15921 -59147
rect -15725 -59447 -15679 -59147
rect -15627 -59447 -15581 -59147
rect -16262 -59545 -15242 -59480
rect -15307 -59628 -15242 -59545
rect -15313 -59700 -15208 -59628
rect -17001 -60040 -16955 -59940
rect -16903 -60069 -16857 -59940
rect -16805 -60040 -16759 -59940
rect -16707 -60069 -16661 -59940
rect -17001 -60115 -16364 -60069
rect -17001 -60271 -16955 -60115
rect -16903 -60117 -16661 -60115
rect -16805 -60271 -16759 -60117
rect -16609 -60271 -16563 -60115
rect -16163 -60359 -16117 -59759
rect -15952 -60359 -15906 -59759
rect -15854 -60359 -15808 -59759
rect -15756 -60359 -15710 -59759
rect -15544 -60359 -15498 -59759
rect -17870 -61383 -17740 -61233
rect -17584 -61255 -17538 -60999
rect -17388 -61253 -17342 -60999
rect -17486 -61255 -17244 -61253
rect -17192 -61255 -17146 -60999
rect -16611 -61170 -16565 -60870
rect -17584 -61301 -16947 -61255
rect -16805 -61274 -16646 -61216
rect -17584 -61529 -17538 -61329
rect -17486 -61529 -17440 -61301
rect -17388 -61529 -17342 -61329
rect -17290 -61529 -17244 -61301
rect -16779 -61329 -16725 -61274
rect -17053 -61383 -16725 -61329
rect -17053 -61673 -16999 -61383
rect -18096 -61727 -16999 -61673
rect -16709 -61706 -16663 -61407
rect -18096 -61997 -18042 -61727
rect -16710 -61743 -16663 -61706
rect -16611 -61707 -16565 -61407
rect -16513 -61743 -16467 -61407
rect -16415 -61707 -16369 -60870
rect -16002 -61025 -15956 -60869
rect -15806 -61023 -15760 -60869
rect -15904 -61025 -15662 -61023
rect -15610 -61025 -15564 -60869
rect -16002 -61071 -15365 -61025
rect -16002 -61200 -15956 -61100
rect -15904 -61200 -15858 -61071
rect -15806 -61200 -15760 -61100
rect -15708 -61200 -15662 -61071
rect -15020 -61235 -14907 -59039
rect -14754 -59631 -14546 -57235
rect -15615 -61348 -14907 -61235
rect -16317 -61743 -16271 -61407
rect -16710 -61790 -16271 -61743
rect -18126 -62133 -17982 -61997
rect -18303 -62388 -18165 -62251
rect -18441 -62486 -18304 -62428
rect -12595 -57231 -12549 -56975
rect -12399 -57229 -12353 -56975
rect -12497 -57231 -12255 -57229
rect -12203 -57231 -12157 -56975
rect -11622 -57146 -11576 -56846
rect -12595 -57277 -11958 -57231
rect -11816 -57250 -11657 -57192
rect -12595 -57505 -12549 -57305
rect -12497 -57505 -12451 -57277
rect -12399 -57505 -12353 -57305
rect -12301 -57505 -12255 -57277
rect -11790 -57305 -11736 -57250
rect -12064 -57359 -11736 -57305
rect -12064 -57649 -12010 -57359
rect -14178 -57703 -12010 -57649
rect -11720 -57682 -11674 -57383
rect -14178 -58787 -14124 -57703
rect -11721 -57719 -11674 -57682
rect -11622 -57683 -11576 -57383
rect -11524 -57719 -11478 -57383
rect -11426 -57683 -11380 -56846
rect -11013 -57001 -10967 -56845
rect -10817 -56999 -10771 -56845
rect -10915 -57001 -10673 -56999
rect -10621 -57001 -10575 -56845
rect -11013 -57047 -10376 -57001
rect -11013 -57176 -10967 -57076
rect -10915 -57176 -10869 -57047
rect -10817 -57176 -10771 -57076
rect -10719 -57176 -10673 -57047
rect -10031 -57211 -9918 -55015
rect -10626 -57324 -9918 -57211
rect -11328 -57719 -11282 -57383
rect -11721 -57766 -11282 -57719
rect -13646 -58226 -13600 -58026
rect -13450 -58226 -13404 -58026
rect -13254 -58226 -13208 -58026
rect -13024 -58279 -12967 -58044
rect -12809 -58226 -12763 -58026
rect -12613 -58226 -12567 -58026
rect -12417 -58226 -12371 -58026
rect -12198 -58141 -12152 -58041
rect -12100 -58141 -12054 -58041
rect -12002 -58141 -11956 -58041
rect -11904 -58141 -11858 -58041
rect -11806 -58141 -11760 -58041
rect -11708 -58141 -11662 -58041
rect -11610 -58141 -11564 -58041
rect -11512 -58141 -11466 -58041
rect -10946 -58226 -10900 -58026
rect -10750 -58226 -10704 -58026
rect -10554 -58226 -10508 -58026
rect -12195 -58279 -12026 -58269
rect -13024 -58336 -12026 -58279
rect -10324 -58279 -10267 -58044
rect -10109 -58226 -10063 -58026
rect -9913 -58226 -9867 -58026
rect -9717 -58226 -9671 -58026
rect -9498 -58141 -9452 -58041
rect -9400 -58141 -9354 -58041
rect -9302 -58141 -9256 -58041
rect -9204 -58141 -9158 -58041
rect -9106 -58141 -9060 -58041
rect -9008 -58141 -8962 -58041
rect -8910 -58141 -8864 -58041
rect -8812 -58141 -8766 -58041
rect -9495 -58279 -9326 -58269
rect -11183 -58301 -11123 -58295
rect -11418 -58322 -11377 -58321
rect -12195 -58343 -12026 -58336
rect -13744 -58506 -13698 -58406
rect -13646 -58506 -13600 -58406
rect -13548 -58506 -13502 -58406
rect -13450 -58506 -13404 -58406
rect -13352 -58506 -13306 -58406
rect -13254 -58506 -13208 -58406
rect -13510 -58729 -13373 -58669
rect -13858 -58787 -13798 -58740
rect -14178 -58851 -13798 -58787
rect -13858 -58877 -13798 -58851
rect -13495 -58947 -13400 -58729
rect -13085 -58847 -13025 -58380
rect -11513 -58382 -11376 -58322
rect -11183 -58361 -11040 -58301
rect -10324 -58336 -9326 -58279
rect -9495 -58343 -9326 -58336
rect -12907 -58506 -12861 -58406
rect -12809 -58506 -12763 -58406
rect -12711 -58506 -12665 -58406
rect -12613 -58506 -12567 -58406
rect -12515 -58506 -12469 -58406
rect -12417 -58506 -12371 -58406
rect -12198 -58556 -12152 -58456
rect -12100 -58556 -12054 -58456
rect -12002 -58556 -11956 -58456
rect -11904 -58556 -11858 -58456
rect -11806 -58556 -11760 -58456
rect -11708 -58556 -11662 -58456
rect -11610 -58556 -11564 -58456
rect -11512 -58556 -11466 -58456
rect -13121 -58907 -12989 -58847
rect -11418 -58867 -11377 -58382
rect -11348 -58818 -11211 -58758
rect -12908 -58915 -11377 -58867
rect -13519 -59007 -13387 -58947
rect -13744 -59164 -13698 -59064
rect -13646 -59164 -13600 -59064
rect -13548 -59164 -13502 -59064
rect -13450 -59164 -13404 -59064
rect -13352 -59164 -13306 -59064
rect -13254 -59164 -13208 -59064
rect -12908 -59069 -12860 -58915
rect -12906 -59114 -12860 -59069
rect -12808 -59114 -12762 -59014
rect -12716 -59033 -12655 -58915
rect -12710 -59114 -12664 -59033
rect -12612 -59114 -12566 -59014
rect -12520 -59035 -12459 -58915
rect -12514 -59114 -12468 -59035
rect -12416 -59114 -12370 -59014
rect -12329 -59033 -12268 -58915
rect -12318 -59114 -12272 -59033
rect -12220 -59114 -12174 -59014
rect -12001 -59164 -11955 -59064
rect -11903 -59164 -11857 -59064
rect -11805 -59164 -11759 -59064
rect -11707 -59164 -11661 -59064
rect -11609 -59164 -11563 -59064
rect -11511 -59164 -11465 -59064
rect -12346 -59234 -12177 -59227
rect -12346 -59291 -11348 -59234
rect -11299 -59266 -11239 -58818
rect -11183 -59109 -11123 -58361
rect -8824 -58384 -8670 -58324
rect -11044 -58506 -10998 -58406
rect -10946 -58506 -10900 -58406
rect -10848 -58506 -10802 -58406
rect -10750 -58506 -10704 -58406
rect -10652 -58506 -10606 -58406
rect -10554 -58506 -10508 -58406
rect -10913 -58735 -10776 -58675
rect -10902 -58943 -10807 -58735
rect -10373 -58759 -10313 -58395
rect -10207 -58506 -10161 -58406
rect -10109 -58506 -10063 -58406
rect -10011 -58506 -9965 -58406
rect -9913 -58506 -9867 -58406
rect -9815 -58506 -9769 -58406
rect -9717 -58506 -9671 -58406
rect -9498 -58556 -9452 -58456
rect -9400 -58556 -9354 -58456
rect -9302 -58556 -9256 -58456
rect -9204 -58556 -9158 -58456
rect -9106 -58556 -9060 -58456
rect -9008 -58556 -8962 -58456
rect -8910 -58556 -8864 -58456
rect -8812 -58556 -8766 -58456
rect -8716 -58659 -8670 -58384
rect -9489 -58704 -8670 -58659
rect -8258 -58675 -8163 -55015
rect -9489 -58705 -8678 -58704
rect -10402 -58819 -10270 -58759
rect -9489 -58871 -9443 -58705
rect -8275 -58735 -8143 -58675
rect -10203 -58917 -9443 -58871
rect -8598 -58905 -8466 -58845
rect -10920 -59003 -10783 -58943
rect -10203 -59014 -10157 -58917
rect -10008 -59014 -9966 -58917
rect -9813 -59014 -9771 -58917
rect -9617 -59014 -9575 -58917
rect -11184 -59154 -11123 -59109
rect -11184 -59241 -11124 -59154
rect -11044 -59164 -10998 -59064
rect -10946 -59164 -10900 -59064
rect -10848 -59164 -10802 -59064
rect -10750 -59164 -10704 -59064
rect -10652 -59164 -10606 -59064
rect -10554 -59164 -10508 -59064
rect -10206 -59114 -10157 -59014
rect -10108 -59114 -10062 -59014
rect -10010 -59114 -9964 -59014
rect -9912 -59114 -9866 -59014
rect -9814 -59114 -9768 -59014
rect -9716 -59114 -9670 -59014
rect -9618 -59114 -9572 -59014
rect -9520 -59114 -9474 -59014
rect -9301 -59164 -9255 -59064
rect -9203 -59164 -9157 -59064
rect -9105 -59164 -9059 -59064
rect -9007 -59164 -8961 -59064
rect -8909 -59164 -8863 -59064
rect -8811 -59164 -8765 -59064
rect -8565 -59133 -8507 -58905
rect -8258 -58944 -8163 -58735
rect -8293 -59004 -8156 -58944
rect -9646 -59234 -9477 -59227
rect -12346 -59301 -12177 -59291
rect -13744 -59544 -13698 -59344
rect -13548 -59544 -13502 -59344
rect -13352 -59544 -13306 -59344
rect -12906 -59497 -12860 -59429
rect -12906 -59529 -12855 -59497
rect -12808 -59529 -12762 -59429
rect -12710 -59472 -12664 -59429
rect -12905 -59612 -12855 -59529
rect -12714 -59612 -12663 -59472
rect -12612 -59529 -12566 -59429
rect -12514 -59491 -12468 -59429
rect -12514 -59612 -12463 -59491
rect -12416 -59529 -12370 -59429
rect -12318 -59491 -12272 -59429
rect -12320 -59612 -12269 -59491
rect -12220 -59529 -12174 -59429
rect -12001 -59544 -11955 -59344
rect -11805 -59544 -11759 -59344
rect -11609 -59544 -11563 -59344
rect -11405 -59526 -11348 -59291
rect -9646 -59291 -8648 -59234
rect -8567 -59265 -8507 -59133
rect -8419 -59164 -8373 -59064
rect -8321 -59164 -8275 -59064
rect -8223 -59164 -8177 -59064
rect -8125 -59164 -8079 -59064
rect -8027 -59164 -7981 -59064
rect -7929 -59164 -7883 -59064
rect -9646 -59301 -9477 -59291
rect -11044 -59544 -10998 -59344
rect -10848 -59544 -10802 -59344
rect -10652 -59544 -10606 -59344
rect -10206 -59529 -10160 -59429
rect -10108 -59529 -10062 -59429
rect -10010 -59529 -9964 -59429
rect -9912 -59529 -9866 -59429
rect -9814 -59529 -9768 -59429
rect -9716 -59529 -9670 -59429
rect -9618 -59529 -9572 -59429
rect -9520 -59529 -9474 -59429
rect -9301 -59544 -9255 -59344
rect -9105 -59544 -9059 -59344
rect -8909 -59544 -8863 -59344
rect -8705 -59612 -8648 -59291
rect -8419 -59544 -8373 -59344
rect -8223 -59544 -8177 -59344
rect -8027 -59544 -7981 -59344
rect -12905 -59669 -8648 -59612
rect -7732 -61973 -7556 -55458
rect -7453 -58643 -7407 -58043
rect -7241 -58643 -7195 -58043
rect -7143 -58643 -7097 -58043
rect -7045 -58643 -6999 -58043
rect -6834 -58643 -6788 -58043
rect -7370 -59255 -7324 -58955
rect -7272 -59255 -7226 -58955
rect -7030 -59255 -6984 -58955
rect -6932 -59255 -6886 -58955
rect -6834 -59255 -6788 -58955
rect -7745 -62144 -7545 -61973
rect -6597 -62231 -6465 -53759
rect -5719 -53845 -5691 -53700
rect -5296 -53698 -5157 -53689
rect -4459 -53698 -4323 -53689
rect -5296 -53726 -4323 -53698
rect -5296 -53743 -5157 -53726
rect -4459 -53735 -4323 -53726
rect -5663 -53772 -5524 -53763
rect -4585 -53770 -4446 -53769
rect -4585 -53772 -4054 -53770
rect -5663 -53798 -4054 -53772
rect -5663 -53800 -4446 -53798
rect -5663 -53817 -5524 -53800
rect -4585 -53823 -4446 -53800
rect -4765 -53845 -4634 -53833
rect -5719 -53873 -4634 -53845
rect -4765 -53879 -4634 -53873
rect -6050 -54111 -6004 -53911
rect -5952 -54111 -5906 -53911
rect -5636 -54111 -5590 -53911
rect -5538 -54111 -5492 -53911
rect -5274 -54111 -5228 -53911
rect -5176 -54111 -5130 -53911
rect -4980 -54111 -4934 -53911
rect -4882 -54111 -4836 -53911
rect -4670 -54111 -4624 -53911
rect -4572 -54111 -4526 -53911
rect -4361 -54111 -4315 -53911
rect -4263 -54111 -4217 -53911
rect -5613 -54454 -5567 -54354
rect -5515 -54454 -5469 -54354
rect -5417 -54454 -5371 -54354
rect -5319 -54454 -5273 -54354
rect -5221 -54454 -5175 -54354
rect -5123 -54454 -5077 -54354
rect -4082 -54437 -4054 -53798
rect -4100 -54573 -4054 -54437
rect -5515 -54834 -5469 -54634
rect -5319 -54834 -5273 -54634
rect -5123 -54834 -5077 -54634
rect -4010 -54869 -3982 -53661
rect -3545 -53672 -3406 -53659
rect -2387 -53661 -1411 -53633
rect -2387 -53669 -2248 -53661
rect -3545 -53700 -3191 -53672
rect -1772 -53675 -1633 -53661
rect -3545 -53713 -3406 -53700
rect -3219 -53845 -3191 -53700
rect -2796 -53698 -2657 -53689
rect -1959 -53698 -1823 -53689
rect -2796 -53726 -1823 -53698
rect -2796 -53743 -2657 -53726
rect -1959 -53735 -1823 -53726
rect -3163 -53772 -3024 -53763
rect -2085 -53770 -1946 -53769
rect -2085 -53772 -1497 -53770
rect -3163 -53798 -1497 -53772
rect -3163 -53800 -1946 -53798
rect -3163 -53817 -3024 -53800
rect -2085 -53823 -1946 -53800
rect -2265 -53845 -2134 -53833
rect -3219 -53873 -2134 -53845
rect -2265 -53879 -2134 -53873
rect -3718 -54078 -3672 -53942
rect -3717 -54648 -3673 -54078
rect -3550 -54111 -3504 -53911
rect -3452 -54111 -3406 -53911
rect -3136 -54111 -3090 -53911
rect -3038 -54111 -2992 -53911
rect -2774 -54111 -2728 -53911
rect -2676 -54111 -2630 -53911
rect -2480 -54111 -2434 -53911
rect -2382 -54111 -2336 -53911
rect -2170 -54111 -2124 -53911
rect -2072 -54111 -2026 -53911
rect -1861 -54111 -1815 -53911
rect -1763 -54111 -1717 -53911
rect -3718 -54784 -3672 -54648
rect -1525 -54802 -1497 -53798
rect -1439 -54719 -1411 -53661
rect -1045 -53672 -906 -53659
rect 113 -53661 1061 -53633
rect 113 -53669 252 -53661
rect -1045 -53700 -691 -53672
rect 728 -53675 867 -53661
rect -1045 -53713 -906 -53700
rect -719 -53845 -691 -53700
rect -296 -53698 -157 -53689
rect 541 -53698 677 -53689
rect -296 -53726 677 -53698
rect -296 -53743 -157 -53726
rect 541 -53735 677 -53726
rect -663 -53772 -524 -53763
rect 415 -53770 554 -53769
rect 415 -53772 987 -53770
rect -663 -53798 987 -53772
rect -663 -53800 554 -53798
rect -663 -53817 -524 -53800
rect 415 -53823 554 -53800
rect 235 -53845 366 -53833
rect -719 -53873 366 -53845
rect 235 -53879 366 -53873
rect -1170 -54082 -1124 -53946
rect -1169 -54319 -1125 -54082
rect -1050 -54111 -1004 -53911
rect -952 -54111 -906 -53911
rect -636 -54111 -590 -53911
rect -538 -54111 -492 -53911
rect -274 -54111 -228 -53911
rect -176 -54111 -130 -53911
rect 20 -54111 66 -53911
rect 118 -54111 164 -53911
rect 330 -54111 376 -53911
rect 428 -54111 474 -53911
rect 639 -54111 685 -53911
rect 737 -54111 783 -53911
rect -1005 -54319 -869 -54318
rect -1170 -54363 -869 -54319
rect -1005 -54364 -869 -54363
rect 959 -54663 987 -53798
rect 1033 -54606 1061 -53661
rect 1455 -53672 1594 -53659
rect 2613 -53661 3536 -53633
rect 2613 -53669 2752 -53661
rect 1455 -53700 1809 -53672
rect 3228 -53675 3367 -53661
rect 1455 -53713 1594 -53700
rect 1781 -53845 1809 -53700
rect 2204 -53698 2343 -53689
rect 3041 -53698 3177 -53689
rect 2204 -53726 3177 -53698
rect 2204 -53743 2343 -53726
rect 3041 -53735 3177 -53726
rect 1837 -53772 1976 -53763
rect 2915 -53770 3054 -53769
rect 2915 -53772 3453 -53770
rect 1837 -53798 3453 -53772
rect 1837 -53800 3054 -53798
rect 1837 -53817 1976 -53800
rect 2915 -53823 3054 -53800
rect 2735 -53845 2866 -53833
rect 1781 -53873 2866 -53845
rect 2735 -53879 2866 -53873
rect 1310 -54082 1356 -53946
rect 1311 -54332 1355 -54082
rect 1450 -54111 1496 -53911
rect 1548 -54111 1594 -53911
rect 1864 -54111 1910 -53911
rect 1962 -54111 2008 -53911
rect 2226 -54111 2272 -53911
rect 2324 -54111 2370 -53911
rect 2520 -54111 2566 -53911
rect 2618 -54111 2664 -53911
rect 2830 -54111 2876 -53911
rect 2928 -54111 2974 -53911
rect 3139 -54111 3185 -53911
rect 3237 -54111 3283 -53911
rect 1492 -54332 1628 -54331
rect 1311 -54376 1628 -54332
rect 1492 -54377 1628 -54376
rect 3425 -54543 3453 -53798
rect 3508 -54469 3536 -53661
rect 3955 -53672 4094 -53659
rect 5113 -53661 6841 -53633
rect 5113 -53669 5252 -53661
rect 3955 -53700 4309 -53672
rect 5728 -53675 5867 -53661
rect 3955 -53713 4094 -53700
rect 4281 -53845 4309 -53700
rect 4704 -53698 4843 -53689
rect 5541 -53698 5677 -53689
rect 4704 -53726 5677 -53698
rect 4704 -53743 4843 -53726
rect 5541 -53735 5677 -53726
rect 5235 -53845 5366 -53833
rect 4281 -53873 5366 -53845
rect 5235 -53879 5366 -53873
rect 3727 -54082 3773 -53946
rect 3728 -54394 3772 -54082
rect 3950 -54111 3996 -53911
rect 4048 -54111 4094 -53911
rect 4364 -54111 4410 -53911
rect 4462 -54111 4508 -53911
rect 4726 -54111 4772 -53911
rect 4824 -54111 4870 -53911
rect 5020 -54111 5066 -53911
rect 5118 -54111 5164 -53911
rect 5330 -54111 5376 -53911
rect 5428 -54111 5474 -53911
rect 5639 -54111 5685 -53911
rect 5737 -54111 5783 -53911
rect 6632 -54082 6678 -53946
rect 6633 -54378 6677 -54082
rect 3675 -54440 3811 -54394
rect 6580 -54424 6716 -54378
rect 6813 -54336 6841 -53661
rect 6955 -53672 7094 -53659
rect 8113 -53661 10998 -53633
rect 8113 -53669 8252 -53661
rect 6955 -53700 7309 -53672
rect 8728 -53675 8867 -53661
rect 6955 -53713 7094 -53700
rect 7281 -53845 7309 -53700
rect 7704 -53698 7843 -53689
rect 8541 -53698 8677 -53689
rect 7704 -53726 8677 -53698
rect 7704 -53743 7843 -53726
rect 8541 -53735 8677 -53726
rect 8235 -53845 8366 -53833
rect 7281 -53873 8366 -53845
rect 8235 -53879 8366 -53873
rect 6950 -54111 6996 -53911
rect 7048 -54111 7094 -53911
rect 7364 -54111 7410 -53911
rect 7462 -54111 7508 -53911
rect 7726 -54111 7772 -53911
rect 7824 -54111 7870 -53911
rect 8020 -54111 8066 -53911
rect 8118 -54111 8164 -53911
rect 8330 -54111 8376 -53911
rect 8428 -54111 8474 -53911
rect 8639 -54111 8685 -53911
rect 8737 -54111 8783 -53911
rect 9641 -54336 10833 -54219
rect 6813 -54364 10842 -54336
rect 3508 -54507 10689 -54469
rect 3425 -54571 10614 -54543
rect 1033 -54634 10537 -54606
rect 959 -54691 10452 -54663
rect -1439 -54770 10378 -54719
rect -1525 -54838 10293 -54802
rect -4010 -54920 10222 -54869
rect -3715 -55039 -3579 -55037
rect 3334 -55039 3470 -55035
rect -3715 -55081 3470 -55039
rect -3715 -55083 -3579 -55081
rect -6195 -55121 -6059 -55119
rect 3230 -55121 3385 -55119
rect -6195 -55163 3385 -55121
rect -6195 -55165 -6059 -55163
rect 3230 -55165 3385 -55163
rect -5870 -55737 -5824 -55537
rect -5674 -55737 -5628 -55537
rect -5478 -55737 -5432 -55537
rect -5032 -55652 -4986 -55552
rect -4934 -55652 -4888 -55552
rect -4836 -55652 -4790 -55552
rect -4738 -55652 -4692 -55552
rect -4640 -55652 -4594 -55552
rect -4542 -55652 -4496 -55552
rect -4444 -55652 -4398 -55552
rect -4346 -55652 -4300 -55552
rect -4127 -55737 -4081 -55537
rect -3931 -55737 -3885 -55537
rect -3735 -55737 -3689 -55537
rect -4472 -55790 -4303 -55780
rect -3531 -55790 -3474 -55555
rect -3170 -55737 -3124 -55537
rect -2974 -55737 -2928 -55537
rect -2778 -55737 -2732 -55537
rect -2332 -55652 -2286 -55552
rect -2234 -55652 -2188 -55552
rect -2136 -55652 -2090 -55552
rect -2038 -55652 -1992 -55552
rect -1940 -55652 -1894 -55552
rect -1842 -55652 -1796 -55552
rect -1744 -55652 -1698 -55552
rect -1646 -55652 -1600 -55552
rect -1427 -55737 -1381 -55537
rect -1231 -55737 -1185 -55537
rect -1035 -55737 -989 -55537
rect -4472 -55847 -3474 -55790
rect -1772 -55790 -1603 -55780
rect -831 -55790 -774 -55555
rect -545 -55737 -499 -55537
rect -349 -55737 -303 -55537
rect -153 -55737 -107 -55537
rect 385 -55754 431 -55554
rect 1123 -55754 1169 -55554
rect 1319 -55754 1365 -55554
rect 1515 -55754 1561 -55554
rect 1741 -55715 1787 -55713
rect -4472 -55854 -4303 -55847
rect -5870 -56017 -5824 -55917
rect -5772 -56017 -5726 -55917
rect -5674 -56017 -5628 -55917
rect -5576 -56017 -5530 -55917
rect -5478 -56017 -5432 -55917
rect -5380 -56017 -5334 -55917
rect -5032 -56012 -4986 -55967
rect -5645 -56134 -5513 -56074
rect -5984 -56230 -5924 -56204
rect -6339 -56293 -5924 -56230
rect -6322 -56294 -5924 -56293
rect -5984 -56341 -5924 -56294
rect -5621 -56352 -5526 -56134
rect -5034 -56166 -4986 -56012
rect -4934 -56067 -4888 -55967
rect -4836 -56048 -4790 -55967
rect -4842 -56166 -4781 -56048
rect -4738 -56067 -4692 -55967
rect -4640 -56046 -4594 -55967
rect -4646 -56166 -4585 -56046
rect -4542 -56067 -4496 -55967
rect -4444 -56048 -4398 -55967
rect -4455 -56166 -4394 -56048
rect -4346 -56067 -4300 -55967
rect -4127 -56017 -4081 -55917
rect -4029 -56017 -3983 -55917
rect -3931 -56017 -3885 -55917
rect -3833 -56017 -3787 -55917
rect -3735 -56017 -3689 -55917
rect -3637 -56017 -3591 -55917
rect -5034 -56214 -3503 -56166
rect -5636 -56412 -5499 -56352
rect -5870 -56675 -5824 -56575
rect -5772 -56675 -5726 -56575
rect -5674 -56675 -5628 -56575
rect -5576 -56675 -5530 -56575
rect -5478 -56675 -5432 -56575
rect -5380 -56675 -5334 -56575
rect -5033 -56675 -4987 -56575
rect -4935 -56675 -4889 -56575
rect -4837 -56675 -4791 -56575
rect -4739 -56675 -4693 -56575
rect -4641 -56675 -4595 -56575
rect -4543 -56675 -4497 -56575
rect -4324 -56625 -4278 -56525
rect -4226 -56625 -4180 -56525
rect -4128 -56625 -4082 -56525
rect -4030 -56625 -3984 -56525
rect -3932 -56625 -3886 -56525
rect -3834 -56625 -3788 -56525
rect -3736 -56625 -3690 -56525
rect -3638 -56625 -3592 -56525
rect -3544 -56699 -3503 -56214
rect -3425 -56263 -3365 -55815
rect -3310 -55927 -3250 -55840
rect -1772 -55847 -774 -55790
rect -1772 -55854 -1603 -55847
rect -3310 -55972 -3249 -55927
rect -3474 -56323 -3337 -56263
rect -4321 -56745 -4152 -56738
rect -5150 -56802 -4152 -56745
rect -3639 -56759 -3502 -56699
rect -3309 -56720 -3249 -55972
rect -3170 -56017 -3124 -55917
rect -3072 -56017 -3026 -55917
rect -2974 -56017 -2928 -55917
rect -2876 -56017 -2830 -55917
rect -2778 -56017 -2732 -55917
rect -2680 -56017 -2634 -55917
rect -2332 -56067 -2283 -55967
rect -2234 -56067 -2188 -55967
rect -2136 -56067 -2090 -55967
rect -2038 -56067 -1992 -55967
rect -1940 -56067 -1894 -55967
rect -1842 -56067 -1796 -55967
rect -1744 -56067 -1698 -55967
rect -1646 -56067 -1600 -55967
rect -1427 -56017 -1381 -55917
rect -1329 -56017 -1283 -55917
rect -1231 -56017 -1185 -55917
rect -1133 -56017 -1087 -55917
rect -1035 -56017 -989 -55917
rect -937 -56017 -891 -55917
rect -3046 -56138 -2909 -56078
rect -3028 -56346 -2933 -56138
rect -2329 -56164 -2283 -56067
rect -2134 -56164 -2092 -56067
rect -1939 -56164 -1897 -56067
rect -1743 -56164 -1701 -56067
rect -2329 -56210 -1569 -56164
rect -2528 -56322 -2396 -56262
rect -3039 -56406 -2902 -56346
rect -3170 -56675 -3124 -56575
rect -3072 -56675 -3026 -56575
rect -2974 -56675 -2928 -56575
rect -2876 -56675 -2830 -56575
rect -2778 -56675 -2732 -56575
rect -2680 -56675 -2634 -56575
rect -2499 -56686 -2439 -56322
rect -1615 -56376 -1569 -56210
rect -831 -56284 -774 -55847
rect -693 -55948 -633 -55816
rect 1733 -55849 1787 -55715
rect 2118 -55723 2164 -55567
rect 2314 -55721 2360 -55567
rect 2216 -55723 2458 -55721
rect 2510 -55723 2556 -55567
rect 2093 -55769 2556 -55723
rect -691 -56176 -633 -55948
rect -545 -56017 -499 -55917
rect -447 -56017 -401 -55917
rect -349 -56017 -303 -55917
rect -251 -56017 -205 -55917
rect -153 -56017 -107 -55917
rect -55 -56017 -9 -55917
rect 240 -56013 381 -55960
rect -289 -56137 -152 -56077
rect -691 -56234 -452 -56176
rect -510 -56263 -452 -56234
rect -831 -56341 -565 -56284
rect -514 -56323 -382 -56263
rect -1615 -56377 -804 -56376
rect -1615 -56422 -796 -56377
rect -2333 -56675 -2287 -56575
rect -2235 -56675 -2189 -56575
rect -2137 -56675 -2091 -56575
rect -2039 -56675 -1993 -56575
rect -1941 -56675 -1895 -56575
rect -1843 -56675 -1797 -56575
rect -1624 -56625 -1578 -56525
rect -1526 -56625 -1480 -56525
rect -1428 -56625 -1382 -56525
rect -1330 -56625 -1284 -56525
rect -1232 -56625 -1186 -56525
rect -1134 -56625 -1088 -56525
rect -1036 -56625 -990 -56525
rect -938 -56625 -892 -56525
rect -842 -56697 -796 -56422
rect -622 -56462 -565 -56341
rect -254 -56346 -159 -56137
rect -271 -56406 -139 -56346
rect 240 -56462 297 -56013
rect 385 -56462 431 -56262
rect 483 -56462 529 -56262
rect 798 -56462 844 -56162
rect 896 -56462 942 -56162
rect 994 -56462 1040 -56162
rect 1107 -56462 1153 -56162
rect 1205 -56462 1251 -56162
rect 1303 -56462 1349 -56162
rect 1417 -56461 1463 -56161
rect 1515 -56461 1561 -56161
rect 1613 -56461 1659 -56161
rect -622 -56519 297 -56462
rect -3544 -56760 -3503 -56759
rect -3309 -56780 -3166 -56720
rect -1621 -56745 -1452 -56738
rect -3309 -56786 -3249 -56780
rect -5772 -57055 -5726 -56855
rect -5576 -57055 -5530 -56855
rect -5380 -57055 -5334 -56855
rect -5150 -57037 -5093 -56802
rect -4321 -56812 -4152 -56802
rect -2450 -56802 -1452 -56745
rect -950 -56757 -796 -56697
rect 1733 -56654 1779 -55849
rect 1822 -55933 1958 -55887
rect 2216 -55898 2262 -55769
rect 2314 -55898 2360 -55798
rect 2412 -55898 2458 -55769
rect 2510 -55898 2556 -55798
rect 1886 -56542 1932 -55933
rect 2825 -56441 2871 -56105
rect 2923 -56405 2969 -55568
rect 3119 -55868 3165 -55568
rect 3723 -55725 3769 -55569
rect 3919 -55723 3965 -55569
rect 3821 -55725 4063 -55723
rect 4115 -55725 4161 -55569
rect 3698 -55771 4161 -55725
rect 3821 -55900 3867 -55771
rect 3919 -55900 3965 -55800
rect 4017 -55900 4063 -55771
rect 4115 -55900 4161 -55800
rect 3021 -56441 3067 -56105
rect 3119 -56405 3165 -56105
rect 3217 -56404 3263 -56105
rect 3217 -56441 3264 -56404
rect 2825 -56488 3264 -56441
rect 4430 -56443 4476 -56107
rect 4528 -56407 4574 -55570
rect 4724 -55870 4770 -55570
rect 5347 -55745 5393 -55545
rect 6085 -55745 6131 -55545
rect 6281 -55745 6327 -55545
rect 6477 -55745 6523 -55545
rect 6960 -55756 7006 -55556
rect 7058 -55787 7104 -55556
rect 7156 -55756 7202 -55556
rect 7276 -55756 7322 -55556
rect 7374 -55756 7420 -55556
rect 7472 -55756 7518 -55556
rect 7834 -55756 7880 -55556
rect 8030 -55756 8076 -55556
rect 8340 -55756 8386 -55556
rect 8649 -55756 8695 -55556
rect 6552 -55833 7104 -55787
rect 6556 -55842 6692 -55833
rect 8123 -55884 8262 -55866
rect 8738 -55877 8877 -55872
rect 9669 -55877 9887 -55818
rect 8738 -55884 9887 -55877
rect 8123 -55905 9887 -55884
rect 6965 -55923 7104 -55910
rect 8123 -55912 8978 -55905
rect 9669 -55907 9887 -55905
rect 8123 -55920 8262 -55912
rect 6965 -55951 7319 -55923
rect 8738 -55926 8877 -55912
rect 6965 -55964 7104 -55951
rect 7291 -56096 7319 -55951
rect 7714 -55949 7853 -55940
rect 8551 -55949 8687 -55940
rect 7714 -55977 8687 -55949
rect 7714 -55994 7853 -55977
rect 8551 -55986 8687 -55977
rect 8245 -56096 8376 -56084
rect 4626 -56443 4672 -56107
rect 4724 -56407 4770 -56107
rect 4822 -56406 4868 -56107
rect 7291 -56124 8376 -56096
rect 8245 -56130 8376 -56124
rect 4822 -56443 4869 -56406
rect 4430 -56490 4869 -56443
rect 5347 -56453 5393 -56253
rect 5445 -56453 5491 -56253
rect 5760 -56453 5806 -56153
rect 5858 -56453 5904 -56153
rect 5956 -56453 6002 -56153
rect 6069 -56453 6115 -56153
rect 6167 -56453 6213 -56153
rect 6265 -56453 6311 -56153
rect 6379 -56452 6425 -56152
rect 6477 -56452 6523 -56152
rect 6575 -56452 6621 -56152
rect 6960 -56362 7006 -56162
rect 7058 -56362 7104 -56162
rect 7374 -56362 7420 -56162
rect 7472 -56362 7518 -56162
rect 7736 -56362 7782 -56162
rect 7834 -56362 7880 -56162
rect 8030 -56362 8076 -56162
rect 8128 -56362 8174 -56162
rect 8340 -56362 8386 -56162
rect 8438 -56362 8484 -56162
rect 8649 -56362 8695 -56162
rect 8747 -56362 8793 -56162
rect 1886 -56588 3635 -56542
rect 1733 -56700 5203 -56654
rect -4935 -57055 -4889 -56855
rect -4739 -57055 -4693 -56855
rect -4543 -57055 -4497 -56855
rect -4324 -57040 -4278 -56940
rect -4226 -57040 -4180 -56940
rect -4128 -57040 -4082 -56940
rect -4030 -57040 -3984 -56940
rect -3932 -57040 -3886 -56940
rect -3834 -57040 -3788 -56940
rect -3736 -57040 -3690 -56940
rect -3638 -57040 -3592 -56940
rect -3072 -57055 -3026 -56855
rect -2876 -57055 -2830 -56855
rect -2680 -57055 -2634 -56855
rect -2450 -57037 -2393 -56802
rect -1621 -56812 -1452 -56802
rect -2235 -57055 -2189 -56855
rect -2039 -57055 -1993 -56855
rect -1843 -57055 -1797 -56855
rect -1624 -57040 -1578 -56940
rect -1526 -57040 -1480 -56940
rect -1428 -57040 -1382 -56940
rect -1330 -57040 -1284 -56940
rect -1232 -57040 -1186 -56940
rect -1134 -57040 -1088 -56940
rect -1036 -57040 -990 -56940
rect -938 -57040 -892 -56940
rect -5772 -58493 -5726 -58293
rect -5576 -58493 -5530 -58293
rect -5380 -58493 -5334 -58293
rect -5150 -58546 -5093 -58311
rect -4935 -58493 -4889 -58293
rect -4739 -58493 -4693 -58293
rect -4543 -58493 -4497 -58293
rect -4324 -58408 -4278 -58308
rect -4226 -58408 -4180 -58308
rect -4128 -58408 -4082 -58308
rect -4030 -58408 -3984 -58308
rect -3932 -58408 -3886 -58308
rect -3834 -58408 -3788 -58308
rect -3736 -58408 -3690 -58308
rect -3638 -58408 -3592 -58308
rect -3072 -58493 -3026 -58293
rect -2876 -58493 -2830 -58293
rect -2680 -58493 -2634 -58293
rect -4321 -58546 -4152 -58536
rect -5150 -58603 -4152 -58546
rect -2450 -58546 -2393 -58311
rect -2235 -58493 -2189 -58293
rect -2039 -58493 -1993 -58293
rect -1843 -58493 -1797 -58293
rect -1624 -58408 -1578 -58308
rect -1526 -58408 -1480 -58308
rect -1428 -58408 -1382 -58308
rect -1330 -58408 -1284 -58308
rect -1232 -58408 -1186 -58308
rect -1134 -58408 -1088 -58308
rect -1036 -58408 -990 -58308
rect -938 -58408 -892 -58308
rect -1621 -58546 -1452 -58536
rect -3309 -58568 -3249 -58562
rect -3544 -58589 -3503 -58588
rect -4321 -58610 -4152 -58603
rect -5870 -58773 -5824 -58673
rect -5772 -58773 -5726 -58673
rect -5674 -58773 -5628 -58673
rect -5576 -58773 -5530 -58673
rect -5478 -58773 -5432 -58673
rect -5380 -58773 -5334 -58673
rect -6330 -59054 -6155 -58835
rect -5636 -58996 -5499 -58936
rect -5984 -59054 -5924 -59007
rect -6330 -59118 -5924 -59054
rect -6330 -59149 -6155 -59118
rect -5984 -59144 -5924 -59118
rect -5621 -59184 -5526 -58996
rect -5211 -59114 -5151 -58647
rect -3639 -58649 -3502 -58589
rect -3309 -58628 -3166 -58568
rect -2450 -58603 -1452 -58546
rect -1621 -58610 -1452 -58603
rect -5033 -58773 -4987 -58673
rect -4935 -58773 -4889 -58673
rect -4837 -58773 -4791 -58673
rect -4739 -58773 -4693 -58673
rect -4641 -58773 -4595 -58673
rect -4543 -58773 -4497 -58673
rect -4324 -58823 -4278 -58723
rect -4226 -58823 -4180 -58723
rect -4128 -58823 -4082 -58723
rect -4030 -58823 -3984 -58723
rect -3932 -58823 -3886 -58723
rect -3834 -58823 -3788 -58723
rect -3736 -58823 -3690 -58723
rect -3638 -58823 -3592 -58723
rect -5247 -59174 -5115 -59114
rect -3544 -59134 -3503 -58649
rect -6108 -59214 -5526 -59184
rect -5034 -59182 -3503 -59134
rect -6108 -59274 -5513 -59214
rect -6108 -59279 -5526 -59274
rect -6108 -59358 -6013 -59279
rect -6323 -59453 -6013 -59358
rect -5870 -59431 -5824 -59331
rect -5772 -59431 -5726 -59331
rect -5674 -59431 -5628 -59331
rect -5576 -59431 -5530 -59331
rect -5478 -59431 -5432 -59331
rect -5380 -59431 -5334 -59331
rect -5034 -59336 -4986 -59182
rect -5032 -59381 -4986 -59336
rect -4934 -59381 -4888 -59281
rect -4842 -59300 -4781 -59182
rect -4836 -59381 -4790 -59300
rect -4738 -59381 -4692 -59281
rect -4646 -59302 -4585 -59182
rect -4640 -59381 -4594 -59302
rect -4542 -59381 -4496 -59281
rect -4455 -59300 -4394 -59182
rect -4444 -59381 -4398 -59300
rect -4346 -59381 -4300 -59281
rect -4127 -59431 -4081 -59331
rect -4029 -59431 -3983 -59331
rect -3931 -59431 -3885 -59331
rect -3833 -59431 -3787 -59331
rect -3735 -59431 -3689 -59331
rect -3637 -59431 -3591 -59331
rect -4472 -59501 -4303 -59494
rect -4472 -59558 -3474 -59501
rect -3309 -59376 -3249 -58628
rect -950 -58651 -796 -58591
rect -3170 -58773 -3124 -58673
rect -3072 -58773 -3026 -58673
rect -2974 -58773 -2928 -58673
rect -2876 -58773 -2830 -58673
rect -2778 -58773 -2732 -58673
rect -2680 -58773 -2634 -58673
rect -3039 -59002 -2902 -58942
rect -3028 -59210 -2933 -59002
rect -2333 -58773 -2287 -58673
rect -2235 -58773 -2189 -58673
rect -2137 -58773 -2091 -58673
rect -2039 -58773 -1993 -58673
rect -1941 -58773 -1895 -58673
rect -1843 -58773 -1797 -58673
rect -1624 -58823 -1578 -58723
rect -1526 -58823 -1480 -58723
rect -1428 -58823 -1382 -58723
rect -1330 -58823 -1284 -58723
rect -1232 -58823 -1186 -58723
rect -1134 -58823 -1088 -58723
rect -1036 -58823 -990 -58723
rect -938 -58823 -892 -58723
rect -842 -58926 -796 -58651
rect 1733 -58694 5203 -58648
rect -1615 -58971 -796 -58926
rect -622 -58886 297 -58829
rect -1615 -58972 -804 -58971
rect -1615 -59138 -1569 -58972
rect -622 -59007 -565 -58886
rect -401 -59002 -269 -58942
rect -2329 -59184 -1569 -59138
rect -831 -59064 -565 -59007
rect -3046 -59270 -2909 -59210
rect -2329 -59281 -2283 -59184
rect -2134 -59281 -2092 -59184
rect -1939 -59281 -1897 -59184
rect -1743 -59281 -1701 -59184
rect -3310 -59421 -3249 -59376
rect -3310 -59508 -3250 -59421
rect -3170 -59431 -3124 -59331
rect -3072 -59431 -3026 -59331
rect -2974 -59431 -2928 -59331
rect -2876 -59431 -2830 -59331
rect -2778 -59431 -2732 -59331
rect -2680 -59431 -2634 -59331
rect -2332 -59381 -2283 -59281
rect -2234 -59381 -2188 -59281
rect -2136 -59381 -2090 -59281
rect -2038 -59381 -1992 -59281
rect -1940 -59381 -1894 -59281
rect -1842 -59381 -1796 -59281
rect -1744 -59381 -1698 -59281
rect -1646 -59381 -1600 -59281
rect -1427 -59431 -1381 -59331
rect -1329 -59431 -1283 -59331
rect -1231 -59431 -1185 -59331
rect -1133 -59431 -1087 -59331
rect -1035 -59431 -989 -59331
rect -937 -59431 -891 -59331
rect -1772 -59501 -1603 -59494
rect -831 -59501 -774 -59064
rect -724 -59172 -592 -59112
rect -691 -59400 -633 -59172
rect -384 -59211 -289 -59002
rect -419 -59271 -282 -59211
rect -4472 -59568 -4303 -59558
rect -5870 -59811 -5824 -59611
rect -5674 -59811 -5628 -59611
rect -5478 -59811 -5432 -59611
rect -5032 -59796 -4986 -59696
rect -4934 -59796 -4888 -59696
rect -4836 -59796 -4790 -59696
rect -4738 -59796 -4692 -59696
rect -4640 -59796 -4594 -59696
rect -4542 -59796 -4496 -59696
rect -4444 -59796 -4398 -59696
rect -4346 -59796 -4300 -59696
rect -4127 -59811 -4081 -59611
rect -3931 -59811 -3885 -59611
rect -3735 -59811 -3689 -59611
rect -3531 -59793 -3474 -59558
rect -1772 -59558 -774 -59501
rect -693 -59532 -633 -59400
rect -545 -59431 -499 -59331
rect -447 -59431 -401 -59331
rect -349 -59431 -303 -59331
rect -251 -59431 -205 -59331
rect -153 -59431 -107 -59331
rect -55 -59431 -9 -59331
rect 240 -59335 297 -58886
rect 385 -59086 431 -58886
rect 483 -59086 529 -58886
rect 798 -59186 844 -58886
rect 896 -59186 942 -58886
rect 994 -59186 1040 -58886
rect 1107 -59186 1153 -58886
rect 1205 -59186 1251 -58886
rect 1303 -59186 1349 -58886
rect 1417 -59187 1463 -58887
rect 1515 -59187 1561 -58887
rect 1613 -59187 1659 -58887
rect 240 -59388 381 -59335
rect 1733 -59499 1779 -58694
rect 1886 -58806 3635 -58760
rect 1886 -59415 1932 -58806
rect 2825 -58907 3264 -58860
rect 2825 -59243 2871 -58907
rect 1822 -59461 1958 -59415
rect -1772 -59568 -1603 -59558
rect -3170 -59811 -3124 -59611
rect -2974 -59811 -2928 -59611
rect -2778 -59811 -2732 -59611
rect -2332 -59796 -2286 -59696
rect -2234 -59796 -2188 -59696
rect -2136 -59796 -2090 -59696
rect -2038 -59796 -1992 -59696
rect -1940 -59796 -1894 -59696
rect -1842 -59796 -1796 -59696
rect -1744 -59796 -1698 -59696
rect -1646 -59796 -1600 -59696
rect -1427 -59811 -1381 -59611
rect -1231 -59811 -1185 -59611
rect -1035 -59811 -989 -59611
rect -831 -59793 -774 -59558
rect -545 -59811 -499 -59611
rect -349 -59811 -303 -59611
rect -153 -59811 -107 -59611
rect 385 -59794 431 -59594
rect 1123 -59794 1169 -59594
rect 1319 -59794 1365 -59594
rect 1515 -59794 1561 -59594
rect 1733 -59633 1787 -59499
rect 2216 -59579 2262 -59450
rect 2314 -59550 2360 -59450
rect 2412 -59579 2458 -59450
rect 2510 -59550 2556 -59450
rect 2093 -59625 2556 -59579
rect 1741 -59635 1787 -59633
rect 2118 -59781 2164 -59625
rect 2216 -59627 2458 -59625
rect 2314 -59781 2360 -59627
rect 2510 -59781 2556 -59625
rect 2923 -59780 2969 -58943
rect 3021 -59243 3067 -58907
rect 3119 -59243 3165 -58943
rect 3217 -58944 3264 -58907
rect 4430 -58905 4869 -58858
rect 3217 -59243 3263 -58944
rect 4430 -59241 4476 -58905
rect 3119 -59780 3165 -59480
rect 3821 -59577 3867 -59448
rect 3919 -59548 3965 -59448
rect 4017 -59577 4063 -59448
rect 4115 -59548 4161 -59448
rect 3698 -59623 4161 -59577
rect 3723 -59779 3769 -59623
rect 3821 -59625 4063 -59623
rect 3919 -59779 3965 -59625
rect 4115 -59779 4161 -59623
rect 4528 -59778 4574 -58941
rect 4626 -59241 4672 -58905
rect 4724 -59241 4770 -58941
rect 4822 -58942 4869 -58905
rect 4822 -59241 4868 -58942
rect 5347 -59095 5393 -58895
rect 5445 -59095 5491 -58895
rect 5760 -59195 5806 -58895
rect 5858 -59195 5904 -58895
rect 5956 -59195 6002 -58895
rect 6069 -59195 6115 -58895
rect 6167 -59195 6213 -58895
rect 6265 -59195 6311 -58895
rect 6379 -59196 6425 -58896
rect 6477 -59196 6523 -58896
rect 6575 -59196 6621 -58896
rect 6960 -59186 7006 -58986
rect 7058 -59186 7104 -58986
rect 7374 -59186 7420 -58986
rect 7472 -59186 7518 -58986
rect 7736 -59186 7782 -58986
rect 7834 -59186 7880 -58986
rect 8030 -59186 8076 -58986
rect 8128 -59186 8174 -58986
rect 8340 -59186 8386 -58986
rect 8438 -59186 8484 -58986
rect 8649 -59186 8695 -58986
rect 8747 -59186 8793 -58986
rect 8245 -59224 8376 -59218
rect 7291 -59252 8376 -59224
rect 6965 -59397 7104 -59384
rect 7291 -59397 7319 -59252
rect 8245 -59264 8376 -59252
rect 6965 -59425 7319 -59397
rect 7714 -59371 7853 -59354
rect 8551 -59371 8687 -59362
rect 7714 -59399 8687 -59371
rect 7714 -59408 7853 -59399
rect 8551 -59408 8687 -59399
rect 6965 -59438 7104 -59425
rect 8123 -59436 8262 -59428
rect 8738 -59436 8877 -59422
rect 8123 -59443 8978 -59436
rect 9836 -59443 9864 -55907
rect 8123 -59464 9864 -59443
rect 4724 -59778 4770 -59478
rect 8123 -59482 8262 -59464
rect 8738 -59471 9864 -59464
rect 8738 -59476 8877 -59471
rect 6556 -59515 6692 -59506
rect 6552 -59561 7104 -59515
rect 5347 -59803 5393 -59603
rect 6085 -59803 6131 -59603
rect 6281 -59803 6327 -59603
rect 6477 -59803 6523 -59603
rect 6960 -59792 7006 -59592
rect 7058 -59792 7104 -59561
rect 7156 -59792 7202 -59592
rect 7276 -59792 7322 -59592
rect 7374 -59792 7420 -59592
rect 7472 -59792 7518 -59592
rect 7834 -59792 7880 -59592
rect 8030 -59792 8076 -59592
rect 8340 -59792 8386 -59592
rect 8649 -59792 8695 -59592
rect 3230 -60185 3385 -60183
rect -6071 -60192 3385 -60185
rect -6195 -60227 3385 -60192
rect -6195 -60238 -6059 -60227
rect 3230 -60229 3385 -60227
rect -3715 -60267 -3579 -60265
rect -3715 -60309 3470 -60267
rect -3715 -60311 -3579 -60309
rect 3334 -60313 3470 -60309
rect 10171 -58598 10222 -54920
rect 10168 -58693 10227 -58598
rect -6050 -61437 -6004 -61237
rect -5952 -61437 -5906 -61237
rect -5636 -61437 -5590 -61237
rect -5538 -61437 -5492 -61237
rect -5274 -61437 -5228 -61237
rect -5176 -61437 -5130 -61237
rect -4980 -61437 -4934 -61237
rect -4882 -61437 -4836 -61237
rect -4670 -61437 -4624 -61237
rect -4572 -61437 -4526 -61237
rect -4361 -61437 -4315 -61237
rect -4263 -61437 -4217 -61237
rect -4765 -61475 -4634 -61469
rect -5719 -61503 -4634 -61475
rect -6045 -61648 -5906 -61635
rect -5719 -61648 -5691 -61503
rect -4765 -61515 -4634 -61503
rect 10171 -60428 10222 -58693
rect -4010 -60474 10222 -60428
rect -4010 -60479 9798 -60474
rect -6045 -61676 -5691 -61648
rect -5296 -61622 -5157 -61605
rect -4459 -61622 -4323 -61613
rect -5296 -61650 -4323 -61622
rect -5296 -61659 -5157 -61650
rect -4459 -61659 -4323 -61650
rect -6045 -61689 -5906 -61676
rect -4887 -61687 -4748 -61679
rect -4272 -61687 -4133 -61673
rect -4010 -61687 -3982 -60479
rect 9986 -60510 10134 -60502
rect 10257 -60510 10293 -54838
rect 10327 -59390 10378 -54770
rect 10321 -59529 10390 -59390
rect -1525 -60546 10293 -60510
rect -3718 -60700 -3672 -60564
rect -3717 -61270 -3673 -60700
rect -3718 -61406 -3672 -61270
rect -3550 -61437 -3504 -61237
rect -3452 -61437 -3406 -61237
rect -3136 -61437 -3090 -61237
rect -3038 -61437 -2992 -61237
rect -2774 -61437 -2728 -61237
rect -2676 -61437 -2630 -61237
rect -2480 -61437 -2434 -61237
rect -2382 -61437 -2336 -61237
rect -2170 -61437 -2124 -61237
rect -2072 -61437 -2026 -61237
rect -1861 -61437 -1815 -61237
rect -1763 -61437 -1717 -61237
rect -2265 -61475 -2134 -61469
rect -3219 -61503 -2134 -61475
rect -4887 -61715 -3982 -61687
rect -3545 -61648 -3406 -61635
rect -3219 -61648 -3191 -61503
rect -2265 -61515 -2134 -61503
rect -3163 -61548 -3024 -61531
rect -2085 -61548 -1946 -61525
rect -3163 -61550 -1946 -61548
rect -1525 -61550 -1497 -60546
rect 9986 -60550 10134 -60546
rect 10327 -60578 10378 -59529
rect -3163 -61576 -1497 -61550
rect -3163 -61585 -3024 -61576
rect -2085 -61578 -1497 -61576
rect -1439 -60609 10378 -60578
rect -1439 -60629 9798 -60609
rect 9991 -60616 10378 -60609
rect -2085 -61579 -1946 -61578
rect -3545 -61676 -3191 -61648
rect -2796 -61622 -2657 -61605
rect -1959 -61622 -1823 -61613
rect -2796 -61650 -1823 -61622
rect -2796 -61659 -2657 -61650
rect -1959 -61659 -1823 -61650
rect -3545 -61689 -3406 -61676
rect -2387 -61687 -2248 -61679
rect -1772 -61687 -1633 -61673
rect -1439 -61687 -1411 -60629
rect 9826 -60657 9969 -60639
rect 10424 -60657 10452 -54691
rect 10509 -58278 10537 -54634
rect 10489 -58396 10553 -58278
rect 959 -60685 10452 -60657
rect -1005 -60985 -869 -60984
rect -1170 -61029 -869 -60985
rect -1169 -61266 -1125 -61029
rect -1005 -61030 -869 -61029
rect -1170 -61402 -1124 -61266
rect -1050 -61437 -1004 -61237
rect -952 -61437 -906 -61237
rect -636 -61437 -590 -61237
rect -538 -61437 -492 -61237
rect -274 -61437 -228 -61237
rect -176 -61437 -130 -61237
rect 20 -61437 66 -61237
rect 118 -61437 164 -61237
rect 330 -61437 376 -61237
rect 428 -61437 474 -61237
rect 639 -61437 685 -61237
rect 737 -61437 783 -61237
rect 235 -61475 366 -61469
rect -719 -61503 366 -61475
rect -2387 -61715 -1411 -61687
rect -1045 -61648 -906 -61635
rect -719 -61648 -691 -61503
rect 235 -61515 366 -61503
rect -663 -61548 -524 -61531
rect 415 -61548 554 -61525
rect -663 -61550 554 -61548
rect 959 -61550 987 -60685
rect 9826 -60686 9969 -60685
rect 10509 -60714 10537 -58396
rect -663 -61576 987 -61550
rect -663 -61585 -524 -61576
rect 415 -61578 987 -61576
rect 1033 -60742 10537 -60714
rect 415 -61579 554 -61578
rect -1045 -61676 -691 -61648
rect -296 -61622 -157 -61605
rect 541 -61622 677 -61613
rect -296 -61650 677 -61622
rect -296 -61659 -157 -61650
rect 541 -61659 677 -61650
rect -1045 -61689 -906 -61676
rect 113 -61687 252 -61679
rect 728 -61687 867 -61673
rect 1033 -61687 1061 -60742
rect 9700 -60777 9844 -60770
rect 10586 -60777 10614 -54571
rect 3425 -60805 10614 -60777
rect 10651 -56041 10689 -54507
rect 10651 -56174 10701 -56041
rect 1492 -60972 1628 -60971
rect 1311 -61016 1628 -60972
rect 1311 -61266 1355 -61016
rect 1492 -61017 1628 -61016
rect 1310 -61402 1356 -61266
rect 1450 -61437 1496 -61237
rect 1548 -61437 1594 -61237
rect 1864 -61437 1910 -61237
rect 1962 -61437 2008 -61237
rect 2226 -61437 2272 -61237
rect 2324 -61437 2370 -61237
rect 2520 -61437 2566 -61237
rect 2618 -61437 2664 -61237
rect 2830 -61437 2876 -61237
rect 2928 -61437 2974 -61237
rect 3139 -61437 3185 -61237
rect 3237 -61437 3283 -61237
rect 2735 -61475 2866 -61469
rect 1781 -61503 2866 -61475
rect 113 -61715 1061 -61687
rect 1455 -61648 1594 -61635
rect 1781 -61648 1809 -61503
rect 2735 -61515 2866 -61503
rect 1837 -61548 1976 -61531
rect 2915 -61548 3054 -61525
rect 1837 -61550 3054 -61548
rect 3425 -61550 3453 -60805
rect 9700 -60817 9844 -60805
rect 10651 -60841 10689 -56174
rect 1837 -61576 3453 -61550
rect 1837 -61585 1976 -61576
rect 2915 -61578 3453 -61576
rect 3508 -60851 9206 -60841
rect 9886 -60851 10689 -60841
rect 3508 -60879 10689 -60851
rect 2915 -61579 3054 -61578
rect 1455 -61676 1809 -61648
rect 2204 -61622 2343 -61605
rect 3041 -61622 3177 -61613
rect 2204 -61650 3177 -61622
rect 2204 -61659 2343 -61650
rect 3041 -61659 3177 -61650
rect 1455 -61689 1594 -61676
rect 2613 -61687 2752 -61679
rect 3228 -61687 3367 -61673
rect 3508 -61687 3536 -60879
rect 3675 -60954 3811 -60908
rect 3728 -61266 3772 -60954
rect 6580 -60970 6716 -60924
rect 3727 -61402 3773 -61266
rect 3950 -61437 3996 -61237
rect 4048 -61437 4094 -61237
rect 4364 -61437 4410 -61237
rect 4462 -61437 4508 -61237
rect 4726 -61437 4772 -61237
rect 4824 -61437 4870 -61237
rect 5020 -61437 5066 -61237
rect 5118 -61437 5164 -61237
rect 5330 -61437 5376 -61237
rect 5428 -61437 5474 -61237
rect 5639 -61437 5685 -61237
rect 5737 -61437 5783 -61237
rect 6633 -61266 6677 -60970
rect 6632 -61402 6678 -61266
rect 5235 -61475 5366 -61469
rect 4281 -61503 5366 -61475
rect 2613 -61715 3536 -61687
rect 3955 -61648 4094 -61635
rect 4281 -61648 4309 -61503
rect 5235 -61515 5366 -61503
rect 10814 -60984 10842 -54364
rect 6813 -61012 10842 -60984
rect 3955 -61676 4309 -61648
rect 4704 -61622 4843 -61605
rect 5541 -61622 5677 -61613
rect 4704 -61650 5677 -61622
rect 4704 -61659 4843 -61650
rect 5541 -61659 5677 -61650
rect 3955 -61689 4094 -61676
rect 5113 -61687 5252 -61679
rect 5728 -61687 5867 -61673
rect 6813 -61687 6841 -61012
rect 6950 -61437 6996 -61237
rect 7048 -61437 7094 -61237
rect 7364 -61437 7410 -61237
rect 7462 -61437 7508 -61237
rect 7726 -61437 7772 -61237
rect 7824 -61437 7870 -61237
rect 8020 -61437 8066 -61237
rect 8118 -61437 8164 -61237
rect 8330 -61437 8376 -61237
rect 8428 -61437 8474 -61237
rect 8639 -61437 8685 -61237
rect 8737 -61437 8783 -61237
rect 8235 -61475 8366 -61469
rect 7281 -61503 8366 -61475
rect 5113 -61715 6841 -61687
rect 6955 -61648 7094 -61635
rect 7281 -61648 7309 -61503
rect 8235 -61515 8366 -61503
rect 6955 -61676 7309 -61648
rect 7704 -61622 7843 -61605
rect 8541 -61622 8677 -61613
rect 7704 -61650 8677 -61622
rect 7704 -61659 7843 -61650
rect 8541 -61659 8677 -61650
rect 6955 -61689 7094 -61676
rect 8113 -61687 8252 -61679
rect 8728 -61687 8867 -61673
rect 10970 -61687 10998 -53661
rect 8113 -61715 10998 -61687
rect -4887 -61733 -4748 -61715
rect -4272 -61727 -4133 -61715
rect -2387 -61733 -2248 -61715
rect -1772 -61727 -1633 -61715
rect 113 -61733 252 -61715
rect 728 -61727 867 -61715
rect 2613 -61733 2752 -61715
rect 3228 -61727 3367 -61715
rect 5113 -61733 5252 -61715
rect 5728 -61727 5867 -61715
rect 8113 -61733 8252 -61715
rect 8728 -61727 8867 -61715
rect -6050 -62043 -6004 -61843
rect -5952 -62043 -5906 -61843
rect -5854 -62043 -5808 -61843
rect -5734 -62043 -5688 -61843
rect -5636 -62043 -5590 -61843
rect -5538 -62043 -5492 -61843
rect -5176 -62043 -5130 -61843
rect -4980 -62043 -4934 -61843
rect -4670 -62043 -4624 -61843
rect -4361 -62043 -4315 -61843
rect -3550 -62043 -3504 -61843
rect -3452 -62043 -3406 -61843
rect -3354 -62043 -3308 -61843
rect -3234 -62043 -3188 -61843
rect -3136 -62043 -3090 -61843
rect -3038 -62043 -2992 -61843
rect -2676 -62043 -2630 -61843
rect -2480 -62043 -2434 -61843
rect -2170 -62043 -2124 -61843
rect -1861 -62043 -1815 -61843
rect -1050 -62043 -1004 -61843
rect -952 -62043 -906 -61843
rect -854 -62043 -808 -61843
rect -734 -62043 -688 -61843
rect -636 -62043 -590 -61843
rect -538 -62043 -492 -61843
rect -176 -62043 -130 -61843
rect 20 -62043 66 -61843
rect 330 -62043 376 -61843
rect 639 -62043 685 -61843
rect 1450 -62043 1496 -61843
rect 1548 -62043 1594 -61843
rect 1646 -62043 1692 -61843
rect 1766 -62043 1812 -61843
rect 1864 -62043 1910 -61843
rect 1962 -62043 2008 -61843
rect 2324 -62043 2370 -61843
rect 2520 -62043 2566 -61843
rect 2830 -62043 2876 -61843
rect 3139 -62043 3185 -61843
rect 3950 -62043 3996 -61843
rect 4048 -62043 4094 -61843
rect 4146 -62043 4192 -61843
rect 4266 -62043 4312 -61843
rect 4364 -62043 4410 -61843
rect 4462 -62043 4508 -61843
rect 4824 -62043 4870 -61843
rect 5020 -62043 5066 -61843
rect 5330 -62043 5376 -61843
rect 5639 -62043 5685 -61843
rect 6950 -62043 6996 -61843
rect 7048 -62043 7094 -61843
rect 7146 -62043 7192 -61843
rect 7266 -62043 7312 -61843
rect 7364 -62043 7410 -61843
rect 7462 -62043 7508 -61843
rect 7824 -62043 7870 -61843
rect 8020 -62043 8066 -61843
rect 8330 -62043 8376 -61843
rect 8639 -62043 8685 -61843
rect -6608 -62406 -6445 -62231
rect -21729 -64390 -21606 -64267
rect -6597 -64761 -6465 -62406
rect 9668 -63594 9729 -62217
rect 9599 -63595 9729 -63594
rect 9599 -63628 9730 -63595
rect 9600 -63713 9730 -63628
rect 9782 -63722 9846 -62213
rect 9780 -63894 9846 -63722
rect 9759 -63895 9846 -63894
rect 9759 -64018 9882 -63895
rect 9927 -64262 9987 -62177
rect 9910 -64385 10033 -64262
rect 11612 -61287 11812 -55231
rect 13476 -58773 13745 -50147
rect 14468 -51080 79593 -50769
rect 13415 -59114 13801 -58773
rect 14468 -59063 14719 -51080
rect 15055 -51530 70325 -51353
rect 15055 -57813 15386 -51530
rect 16167 -52089 61616 -51868
rect 16167 -56033 16257 -52089
rect 17548 -52646 52427 -52420
rect 17156 -53126 43602 -52861
rect 16874 -53532 35121 -53283
rect 16900 -54212 17465 -54211
rect 16615 -54352 17465 -54212
rect 27300 -54644 33765 -54475
rect 16582 -55274 16849 -55196
rect 16582 -55429 26496 -55274
rect 16582 -55494 16849 -55429
rect 16845 -55938 17672 -55787
rect 20978 -55921 21024 -55821
rect 21076 -55921 21122 -55821
rect 21174 -55921 21220 -55821
rect 21272 -55921 21318 -55821
rect 21370 -55921 21416 -55821
rect 21468 -55921 21514 -55821
rect 21566 -55921 21612 -55821
rect 21664 -55921 21710 -55821
rect 16163 -56197 16261 -56033
rect 14951 -58238 15465 -57813
rect 16167 -58362 16257 -56197
rect 18872 -56240 18918 -56040
rect 18970 -56240 19016 -56040
rect 19068 -56240 19114 -56040
rect 19166 -56240 19212 -56040
rect 21883 -56006 21929 -55806
rect 22079 -56006 22125 -55806
rect 22275 -56006 22321 -55806
rect 21538 -56059 21707 -56049
rect 22479 -56059 22536 -55824
rect 22720 -56006 22766 -55806
rect 22916 -56006 22962 -55806
rect 23112 -56006 23158 -55806
rect 23678 -55921 23724 -55821
rect 23776 -55921 23822 -55821
rect 23874 -55921 23920 -55821
rect 23972 -55921 24018 -55821
rect 24070 -55921 24116 -55821
rect 24168 -55921 24214 -55821
rect 24266 -55921 24312 -55821
rect 24364 -55921 24410 -55821
rect 24583 -56006 24629 -55806
rect 24779 -56006 24825 -55806
rect 24975 -56006 25021 -55806
rect 20882 -56164 21036 -56104
rect 21538 -56116 22536 -56059
rect 24238 -56059 24407 -56049
rect 25179 -56059 25236 -55824
rect 25420 -56006 25466 -55806
rect 25616 -56006 25662 -55806
rect 25812 -56006 25858 -55806
rect 23335 -56081 23395 -56075
rect 21538 -56123 21707 -56116
rect 23252 -56141 23395 -56081
rect 23589 -56102 23630 -56101
rect 19708 -56278 19750 -56274
rect 19626 -56338 19758 -56278
rect 18872 -57204 18918 -56604
rect 19084 -57204 19130 -56604
rect 19182 -57204 19228 -56604
rect 19280 -57204 19326 -56604
rect 19393 -57204 19439 -56604
rect 19491 -57204 19537 -56604
rect 19589 -57204 19635 -56604
rect 16707 -58141 18817 -57945
rect 18621 -58147 18817 -58141
rect 18621 -58301 18819 -58147
rect 18614 -58343 19651 -58301
rect 16167 -58375 18150 -58362
rect 16167 -58417 19561 -58375
rect 16167 -58452 18150 -58417
rect 18867 -58858 18913 -58658
rect 18965 -58858 19011 -58658
rect 19063 -58858 19109 -58658
rect 19277 -58963 19409 -58903
rect 14452 -59293 14740 -59063
rect 19364 -59076 19406 -58963
rect 19519 -58988 19561 -58417
rect 19609 -58904 19651 -58343
rect 19708 -58372 19750 -56338
rect 19798 -56399 20708 -56342
rect 19798 -57750 19855 -56399
rect 20355 -56515 20487 -56455
rect 20375 -56724 20470 -56515
rect 20651 -56520 20708 -56399
rect 20882 -56439 20928 -56164
rect 20978 -56336 21024 -56236
rect 21076 -56336 21122 -56236
rect 21174 -56336 21220 -56236
rect 21272 -56336 21318 -56236
rect 21370 -56336 21416 -56236
rect 21468 -56336 21514 -56236
rect 21566 -56336 21612 -56236
rect 21664 -56336 21710 -56236
rect 21883 -56286 21929 -56186
rect 21981 -56286 22027 -56186
rect 22079 -56286 22125 -56186
rect 22177 -56286 22223 -56186
rect 22275 -56286 22321 -56186
rect 22373 -56286 22419 -56186
rect 20882 -56484 21701 -56439
rect 20890 -56485 21701 -56484
rect 20651 -56577 20917 -56520
rect 20678 -56685 20810 -56625
rect 20368 -56784 20505 -56724
rect 20095 -56944 20141 -56844
rect 20193 -56944 20239 -56844
rect 20291 -56944 20337 -56844
rect 20389 -56944 20435 -56844
rect 20487 -56944 20533 -56844
rect 20585 -56944 20631 -56844
rect 20719 -56913 20777 -56685
rect 20719 -57045 20779 -56913
rect 20860 -57014 20917 -56577
rect 21655 -56651 21701 -56485
rect 22720 -56286 22766 -56186
rect 22818 -56286 22864 -56186
rect 22916 -56286 22962 -56186
rect 23014 -56286 23060 -56186
rect 23112 -56286 23158 -56186
rect 23210 -56286 23256 -56186
rect 22988 -56515 23125 -56455
rect 21655 -56697 22415 -56651
rect 21787 -56794 21829 -56697
rect 21983 -56794 22025 -56697
rect 22178 -56794 22220 -56697
rect 22369 -56794 22415 -56697
rect 23019 -56723 23114 -56515
rect 22995 -56783 23132 -56723
rect 20977 -56944 21023 -56844
rect 21075 -56944 21121 -56844
rect 21173 -56944 21219 -56844
rect 21271 -56944 21317 -56844
rect 21369 -56944 21415 -56844
rect 21467 -56944 21513 -56844
rect 21686 -56894 21732 -56794
rect 21784 -56894 21830 -56794
rect 21882 -56894 21928 -56794
rect 21980 -56894 22026 -56794
rect 22078 -56894 22124 -56794
rect 22176 -56894 22222 -56794
rect 22274 -56894 22320 -56794
rect 22369 -56894 22418 -56794
rect 22720 -56944 22766 -56844
rect 22818 -56944 22864 -56844
rect 22916 -56944 22962 -56844
rect 23014 -56944 23060 -56844
rect 23112 -56944 23158 -56844
rect 23210 -56944 23256 -56844
rect 23335 -56889 23395 -56141
rect 23588 -56162 23725 -56102
rect 24238 -56116 25236 -56059
rect 24238 -56123 24407 -56116
rect 23335 -56934 23396 -56889
rect 21689 -57014 21858 -57007
rect 20860 -57071 21858 -57014
rect 23336 -57021 23396 -56934
rect 23589 -56647 23630 -56162
rect 23678 -56336 23724 -56236
rect 23776 -56336 23822 -56236
rect 23874 -56336 23920 -56236
rect 23972 -56336 24018 -56236
rect 24070 -56336 24116 -56236
rect 24168 -56336 24214 -56236
rect 24266 -56336 24312 -56236
rect 24364 -56336 24410 -56236
rect 24583 -56286 24629 -56186
rect 24681 -56286 24727 -56186
rect 24779 -56286 24825 -56186
rect 24877 -56286 24923 -56186
rect 24975 -56286 25021 -56186
rect 25073 -56286 25119 -56186
rect 25237 -56627 25297 -56160
rect 25420 -56286 25466 -56186
rect 25518 -56286 25564 -56186
rect 25616 -56286 25662 -56186
rect 25714 -56286 25760 -56186
rect 25812 -56286 25858 -56186
rect 25910 -56286 25956 -56186
rect 25585 -56509 25722 -56449
rect 23589 -56695 25120 -56647
rect 25201 -56687 25333 -56627
rect 23677 -56944 23723 -56844
rect 23775 -56944 23821 -56844
rect 23873 -56944 23919 -56844
rect 23971 -56944 24017 -56844
rect 24069 -56944 24115 -56844
rect 24167 -56944 24213 -56844
rect 24386 -56894 24432 -56794
rect 24480 -56813 24541 -56695
rect 24484 -56894 24530 -56813
rect 24582 -56894 24628 -56794
rect 24671 -56815 24732 -56695
rect 24680 -56894 24726 -56815
rect 24778 -56894 24824 -56794
rect 24867 -56813 24928 -56695
rect 24876 -56894 24922 -56813
rect 24974 -56894 25020 -56794
rect 25072 -56849 25120 -56695
rect 25612 -56727 25707 -56509
rect 26010 -56567 26070 -56520
rect 26010 -56631 26279 -56567
rect 26010 -56657 26156 -56631
rect 25599 -56787 25731 -56727
rect 25072 -56894 25118 -56849
rect 25420 -56944 25466 -56844
rect 25518 -56944 25564 -56844
rect 25616 -56944 25662 -56844
rect 25714 -56944 25760 -56844
rect 25812 -56944 25858 -56844
rect 25910 -56944 25956 -56844
rect 24389 -57014 24558 -57007
rect 20193 -57324 20239 -57124
rect 20389 -57324 20435 -57124
rect 20585 -57324 20631 -57124
rect 20860 -57306 20917 -57071
rect 21689 -57081 21858 -57071
rect 23560 -57071 24558 -57014
rect 21075 -57324 21121 -57124
rect 21271 -57324 21317 -57124
rect 21467 -57324 21513 -57124
rect 21686 -57309 21732 -57209
rect 21784 -57309 21830 -57209
rect 21882 -57309 21928 -57209
rect 21980 -57309 22026 -57209
rect 22078 -57309 22124 -57209
rect 22176 -57309 22222 -57209
rect 22274 -57309 22320 -57209
rect 22372 -57309 22418 -57209
rect 22818 -57324 22864 -57124
rect 23014 -57324 23060 -57124
rect 23210 -57324 23256 -57124
rect 23560 -57306 23617 -57071
rect 24389 -57081 24558 -57071
rect 23775 -57324 23821 -57124
rect 23971 -57324 24017 -57124
rect 24167 -57324 24213 -57124
rect 24386 -57309 24432 -57209
rect 24484 -57309 24530 -57209
rect 24582 -57309 24628 -57209
rect 24680 -57309 24726 -57209
rect 24778 -57309 24824 -57209
rect 24876 -57309 24922 -57209
rect 24974 -57309 25020 -57209
rect 25072 -57309 25118 -57209
rect 25518 -57324 25564 -57124
rect 25714 -57324 25760 -57124
rect 25910 -57324 25956 -57124
rect 26066 -57501 26156 -56657
rect 22124 -57591 26156 -57501
rect 22124 -57682 22284 -57591
rect 19798 -57807 23070 -57750
rect 22121 -57997 22281 -57865
rect 19708 -58414 20478 -58372
rect 22018 -58380 22150 -58320
rect 19813 -58858 19859 -58658
rect 19911 -58858 19957 -58658
rect 20009 -58858 20055 -58658
rect 19725 -58904 19857 -58897
rect 19609 -58946 19857 -58904
rect 19725 -58957 19857 -58946
rect 19948 -58988 20080 -58977
rect 19519 -59030 20080 -58988
rect 19948 -59037 20080 -59030
rect 20313 -59076 20373 -59046
rect 19364 -59118 20373 -59076
rect 18867 -59550 18913 -59150
rect 19078 -59550 19124 -59150
rect 19176 -59550 19222 -59150
rect 19274 -59550 19320 -59150
rect 19813 -59550 19859 -59150
rect 20024 -59550 20070 -59150
rect 20122 -59550 20168 -59150
rect 20220 -59550 20266 -59150
rect 20313 -59178 20373 -59118
rect 20436 -59296 20478 -58414
rect 20631 -58977 20677 -58677
rect 20729 -58977 20775 -58677
rect 20827 -58977 20873 -58677
rect 20941 -58976 20987 -58676
rect 21039 -58976 21085 -58676
rect 21137 -58976 21183 -58676
rect 21250 -58976 21296 -58676
rect 21348 -58976 21394 -58676
rect 21446 -58976 21492 -58676
rect 21761 -58876 21807 -58676
rect 21859 -58876 21905 -58676
rect 22050 -59065 22110 -58380
rect 22189 -58421 22249 -57997
rect 22638 -58276 22684 -57876
rect 22834 -58276 22880 -57876
rect 23013 -58329 23070 -57807
rect 26341 -57818 26496 -55429
rect 23209 -57888 26496 -57818
rect 23209 -58067 23279 -57888
rect 22189 -58422 22530 -58421
rect 22189 -58480 22531 -58422
rect 22984 -58463 23070 -58329
rect 22189 -58481 22530 -58480
rect 22011 -59125 22142 -59065
rect 22189 -59235 22249 -58481
rect 22540 -58730 22586 -58530
rect 22638 -58730 22684 -58530
rect 22750 -58730 22796 -58530
rect 22848 -58730 22894 -58530
rect 23370 -58621 23416 -57921
rect 23468 -58621 23514 -57921
rect 23770 -58621 23816 -57921
rect 23868 -58621 23914 -57921
rect 24253 -58618 24323 -57888
rect 24370 -58621 24416 -57921
rect 24468 -58621 24514 -57921
rect 24770 -58621 24816 -57921
rect 24868 -58621 24914 -57921
rect 25244 -58619 25314 -57888
rect 25370 -58621 25416 -57921
rect 25468 -58621 25514 -57921
rect 25770 -58621 25816 -57921
rect 25868 -58621 25914 -57921
rect 23982 -58671 24100 -58659
rect 23982 -58705 24189 -58671
rect 25955 -58678 26073 -58674
rect 26506 -58678 26627 -58655
rect 23982 -58717 24100 -58705
rect 22490 -59197 22536 -59097
rect 22588 -59197 22634 -59097
rect 22686 -59197 22732 -59097
rect 22784 -59197 22830 -59097
rect 22882 -59197 22928 -59097
rect 22980 -59197 23026 -59097
rect 22189 -59295 22516 -59235
rect 20428 -59428 20488 -59296
rect 20729 -59584 20775 -59384
rect 20925 -59584 20971 -59384
rect 21121 -59584 21167 -59384
rect 21859 -59584 21905 -59384
rect 22588 -59577 22634 -59377
rect 22784 -59577 22830 -59377
rect 22980 -59577 23026 -59377
rect 23468 -59506 23514 -58806
rect 23868 -59506 23914 -58806
rect 24155 -59606 24189 -58705
rect 25059 -58744 25177 -58686
rect 25955 -58723 26627 -58678
rect 25955 -58732 26073 -58723
rect 24468 -59506 24514 -58806
rect 24868 -59506 24914 -58806
rect 25065 -59541 25099 -58744
rect 25468 -59506 25514 -58806
rect 25868 -59506 25914 -58806
rect 25065 -59575 26373 -59541
rect 24155 -59640 26285 -59606
rect 12065 -60562 12111 -60362
rect 12261 -60562 12307 -60362
rect 12457 -60562 12503 -60362
rect 12732 -60615 12789 -60380
rect 12947 -60562 12993 -60362
rect 13143 -60562 13189 -60362
rect 13339 -60562 13385 -60362
rect 13558 -60477 13604 -60377
rect 13656 -60477 13702 -60377
rect 13754 -60477 13800 -60377
rect 13852 -60477 13898 -60377
rect 13950 -60477 13996 -60377
rect 14048 -60477 14094 -60377
rect 14146 -60477 14192 -60377
rect 14244 -60477 14290 -60377
rect 14690 -60562 14736 -60362
rect 14886 -60562 14932 -60362
rect 15082 -60562 15128 -60362
rect 13561 -60615 13730 -60605
rect 11967 -60842 12013 -60742
rect 12065 -60842 12111 -60742
rect 12163 -60842 12209 -60742
rect 12261 -60842 12307 -60742
rect 12359 -60842 12405 -60742
rect 12457 -60842 12503 -60742
rect 12591 -60773 12651 -60641
rect 12732 -60672 13730 -60615
rect 15432 -60615 15489 -60380
rect 15647 -60562 15693 -60362
rect 15843 -60562 15889 -60362
rect 16039 -60562 16085 -60362
rect 16258 -60477 16304 -60377
rect 16356 -60477 16402 -60377
rect 16454 -60477 16500 -60377
rect 16552 -60477 16598 -60377
rect 16650 -60477 16696 -60377
rect 16748 -60477 16794 -60377
rect 16846 -60477 16892 -60377
rect 16944 -60477 16990 -60377
rect 17390 -60562 17436 -60362
rect 17586 -60562 17632 -60362
rect 17782 -60562 17828 -60362
rect 16261 -60615 16430 -60605
rect 12240 -60962 12377 -60902
rect 12247 -61171 12342 -60962
rect 12591 -61001 12649 -60773
rect 12550 -61061 12682 -61001
rect 12732 -61109 12789 -60672
rect 13561 -60679 13730 -60672
rect 12849 -60842 12895 -60742
rect 12947 -60842 12993 -60742
rect 13045 -60842 13091 -60742
rect 13143 -60842 13189 -60742
rect 13241 -60842 13287 -60742
rect 13339 -60842 13385 -60742
rect 13558 -60892 13604 -60792
rect 13656 -60892 13702 -60792
rect 13754 -60892 13800 -60792
rect 13852 -60892 13898 -60792
rect 13950 -60892 13996 -60792
rect 14048 -60892 14094 -60792
rect 14146 -60892 14192 -60792
rect 14241 -60892 14290 -60792
rect 14592 -60842 14638 -60742
rect 14690 -60842 14736 -60742
rect 14788 -60842 14834 -60742
rect 14886 -60842 14932 -60742
rect 14984 -60842 15030 -60742
rect 15082 -60842 15128 -60742
rect 15208 -60752 15268 -60665
rect 15207 -60797 15268 -60752
rect 13659 -60989 13701 -60892
rect 13855 -60989 13897 -60892
rect 14050 -60989 14092 -60892
rect 14241 -60989 14287 -60892
rect 14867 -60963 15004 -60903
rect 12523 -61166 12789 -61109
rect 13527 -61035 14287 -60989
rect 12227 -61231 12359 -61171
rect 12523 -61287 12580 -61166
rect 13527 -61201 13573 -61035
rect 12762 -61202 13573 -61201
rect 11612 -61344 12580 -61287
rect 12754 -61247 13573 -61202
rect -6597 -64897 -6461 -64761
rect 11612 -65134 11812 -61344
rect 12754 -61522 12800 -61247
rect 12850 -61450 12896 -61350
rect 12948 -61450 12994 -61350
rect 13046 -61450 13092 -61350
rect 13144 -61450 13190 -61350
rect 13242 -61450 13288 -61350
rect 13340 -61450 13386 -61350
rect 13438 -61450 13484 -61350
rect 13536 -61450 13582 -61350
rect 13755 -61500 13801 -61400
rect 13853 -61500 13899 -61400
rect 13951 -61500 13997 -61400
rect 14049 -61500 14095 -61400
rect 14147 -61500 14193 -61400
rect 14245 -61500 14291 -61400
rect 14891 -61171 14986 -60963
rect 14860 -61231 14997 -61171
rect 14592 -61500 14638 -61400
rect 14690 -61500 14736 -61400
rect 14788 -61500 14834 -61400
rect 14886 -61500 14932 -61400
rect 14984 -61500 15030 -61400
rect 15082 -61500 15128 -61400
rect 12754 -61582 12908 -61522
rect 15207 -61545 15267 -60797
rect 15432 -60672 16430 -60615
rect 16261 -60679 16430 -60672
rect 15549 -60842 15595 -60742
rect 15647 -60842 15693 -60742
rect 15745 -60842 15791 -60742
rect 15843 -60842 15889 -60742
rect 15941 -60842 15987 -60742
rect 16039 -60842 16085 -60742
rect 16258 -60892 16304 -60792
rect 16356 -60873 16402 -60792
rect 16352 -60991 16413 -60873
rect 16454 -60892 16500 -60792
rect 16552 -60871 16598 -60792
rect 16543 -60991 16604 -60871
rect 16650 -60892 16696 -60792
rect 16748 -60873 16794 -60792
rect 16739 -60991 16800 -60873
rect 16846 -60892 16892 -60792
rect 16944 -60837 16990 -60792
rect 16944 -60991 16992 -60837
rect 17292 -60842 17338 -60742
rect 17390 -60842 17436 -60742
rect 17488 -60842 17534 -60742
rect 17586 -60842 17632 -60742
rect 17684 -60842 17730 -60742
rect 17782 -60842 17828 -60742
rect 17471 -60959 17603 -60899
rect 15461 -61039 16992 -60991
rect 15461 -61524 15502 -61039
rect 17073 -61059 17205 -60999
rect 15550 -61450 15596 -61350
rect 15648 -61450 15694 -61350
rect 15746 -61450 15792 -61350
rect 15844 -61450 15890 -61350
rect 15942 -61450 15988 -61350
rect 16040 -61450 16086 -61350
rect 16138 -61450 16184 -61350
rect 16236 -61450 16282 -61350
rect 16455 -61500 16501 -61400
rect 16553 -61500 16599 -61400
rect 16651 -61500 16697 -61400
rect 16749 -61500 16795 -61400
rect 16847 -61500 16893 -61400
rect 16945 -61500 16991 -61400
rect 13410 -61570 13579 -61563
rect 13410 -61627 14408 -61570
rect 15124 -61605 15267 -61545
rect 15460 -61584 15597 -61524
rect 17109 -61526 17169 -61059
rect 17484 -61177 17579 -60959
rect 17882 -61055 17942 -61029
rect 17882 -61119 18338 -61055
rect 17882 -61166 17942 -61119
rect 17457 -61237 17594 -61177
rect 17292 -61500 17338 -61400
rect 17390 -61500 17436 -61400
rect 17488 -61500 17534 -61400
rect 17586 -61500 17632 -61400
rect 17684 -61500 17730 -61400
rect 17782 -61500 17828 -61400
rect 16110 -61570 16279 -61563
rect 15461 -61585 15502 -61584
rect 15207 -61611 15267 -61605
rect 13410 -61637 13579 -61627
rect 12850 -61865 12896 -61765
rect 12948 -61865 12994 -61765
rect 13046 -61865 13092 -61765
rect 13144 -61865 13190 -61765
rect 13242 -61865 13288 -61765
rect 13340 -61865 13386 -61765
rect 13438 -61865 13484 -61765
rect 13536 -61865 13582 -61765
rect 13755 -61880 13801 -61680
rect 13951 -61880 13997 -61680
rect 14147 -61880 14193 -61680
rect 14351 -61862 14408 -61627
rect 16110 -61627 17108 -61570
rect 16110 -61637 16279 -61627
rect 14592 -61880 14638 -61680
rect 14788 -61880 14834 -61680
rect 14984 -61880 15030 -61680
rect 15550 -61865 15596 -61765
rect 15648 -61865 15694 -61765
rect 15746 -61865 15792 -61765
rect 15844 -61865 15890 -61765
rect 15942 -61865 15988 -61765
rect 16040 -61865 16086 -61765
rect 16138 -61865 16184 -61765
rect 16236 -61865 16282 -61765
rect 16455 -61880 16501 -61680
rect 16651 -61880 16697 -61680
rect 16847 -61880 16893 -61680
rect 17051 -61862 17108 -61627
rect 17292 -61880 17338 -61680
rect 17488 -61880 17534 -61680
rect 17684 -61880 17730 -61680
rect 18210 -64761 18338 -61119
rect 25712 -61811 25782 -59640
rect 26339 -59703 26373 -59575
rect 25593 -62031 25964 -61811
rect 26278 -62360 26399 -59703
rect 18205 -64897 18338 -64761
rect 24998 -62481 26399 -62360
rect 24998 -65324 25119 -62481
rect 26506 -64722 26627 -58723
rect 27300 -58292 27469 -54644
rect 29325 -54909 29764 -54862
rect 29325 -54946 29372 -54909
rect 28165 -55419 28295 -55269
rect 28451 -55323 28497 -55123
rect 28549 -55351 28595 -55123
rect 28647 -55323 28693 -55123
rect 28745 -55351 28791 -55123
rect 29326 -55245 29372 -54946
rect 29424 -55245 29470 -54945
rect 29522 -55245 29568 -54909
rect 28451 -55397 29088 -55351
rect 28215 -56823 28269 -55419
rect 28451 -55653 28497 -55397
rect 28549 -55399 28791 -55397
rect 28647 -55653 28693 -55399
rect 28843 -55653 28889 -55397
rect 29424 -55782 29470 -55482
rect 29620 -55782 29666 -54945
rect 29718 -55245 29764 -54909
rect 30420 -55417 31128 -55304
rect 30033 -55552 30079 -55452
rect 30131 -55581 30177 -55452
rect 30229 -55552 30275 -55452
rect 30327 -55581 30373 -55452
rect 30033 -55627 30670 -55581
rect 30033 -55783 30079 -55627
rect 30131 -55629 30373 -55627
rect 30229 -55783 30275 -55629
rect 30425 -55783 30471 -55627
rect 28425 -56682 28471 -56382
rect 28072 -56877 28269 -56823
rect 28327 -57218 28373 -56919
rect 28326 -57255 28373 -57218
rect 28425 -57219 28471 -56919
rect 28523 -57255 28569 -56919
rect 28621 -57219 28667 -56382
rect 29034 -56537 29080 -56381
rect 29230 -56535 29276 -56381
rect 29132 -56537 29374 -56535
rect 29426 -56537 29472 -56381
rect 29034 -56583 29671 -56537
rect 29034 -56712 29080 -56612
rect 29132 -56712 29178 -56583
rect 29230 -56712 29276 -56612
rect 29328 -56712 29374 -56583
rect 29872 -56893 29918 -56293
rect 30083 -56893 30129 -56293
rect 30181 -56893 30227 -56293
rect 30279 -56893 30325 -56293
rect 30491 -56893 30537 -56293
rect 28719 -57255 28765 -56919
rect 30722 -57024 30827 -56952
rect 30728 -57107 30793 -57024
rect 29773 -57172 30793 -57107
rect 28326 -57302 28765 -57255
rect 29872 -57505 29918 -57205
rect 29970 -57505 30016 -57205
rect 30068 -57505 30114 -57205
rect 30310 -57505 30356 -57205
rect 30408 -57505 30454 -57205
rect 30641 -57613 30754 -57612
rect 31015 -57613 31128 -55417
rect 31864 -56651 31910 -56151
rect 32133 -56651 32179 -56151
rect 32231 -56651 32277 -56151
rect 32329 -56651 32375 -56151
rect 32459 -56651 32505 -56151
rect 32785 -56651 32831 -56151
rect 33013 -56451 33059 -56151
rect 31633 -56811 31771 -56807
rect 32439 -56811 32577 -56807
rect 32824 -56811 32878 -56738
rect 31633 -56855 32878 -56811
rect 31633 -56861 31771 -56855
rect 32439 -56861 32577 -56855
rect 32824 -56876 32878 -56855
rect 32996 -56891 33062 -56879
rect 33596 -56891 33765 -54644
rect 34872 -54766 35121 -53532
rect 35283 -54592 42365 -54401
rect 34781 -54902 35138 -54766
rect 34781 -54956 35144 -54902
rect 34781 -55033 35138 -54956
rect 31472 -57198 31575 -57107
rect 30451 -57726 31128 -57613
rect 27300 -58378 27650 -58292
rect 29317 -58362 29756 -58315
rect 27300 -58432 29028 -58378
rect 29317 -58399 29364 -58362
rect 27300 -58461 27650 -58432
rect 28157 -58872 28287 -58722
rect 28443 -58776 28489 -58576
rect 28541 -58804 28587 -58576
rect 28639 -58776 28685 -58576
rect 28737 -58804 28783 -58576
rect 28974 -58722 29028 -58432
rect 29318 -58698 29364 -58399
rect 29416 -58698 29462 -58398
rect 29514 -58698 29560 -58362
rect 28974 -58776 29302 -58722
rect 28443 -58850 29080 -58804
rect 29248 -58831 29302 -58776
rect 28207 -60276 28261 -58872
rect 28443 -59106 28489 -58850
rect 28541 -58852 28783 -58850
rect 28639 -59106 28685 -58852
rect 28835 -59106 28881 -58850
rect 29222 -58889 29381 -58831
rect 29416 -59235 29462 -58935
rect 29612 -59235 29658 -58398
rect 29710 -58698 29756 -58362
rect 30641 -58757 30754 -57726
rect 31484 -57831 31563 -57198
rect 31766 -57447 31812 -57147
rect 31864 -57447 31910 -57147
rect 32236 -57447 32282 -56947
rect 32334 -57447 32380 -56947
rect 32459 -57447 32505 -56947
rect 32557 -57447 32603 -56947
rect 32687 -57447 32733 -56947
rect 32785 -57447 32831 -56947
rect 32883 -57447 32929 -56947
rect 32996 -56953 34618 -56891
rect 32996 -56962 33062 -56953
rect 33013 -57447 33059 -57147
rect 33111 -57447 33157 -57147
rect 30984 -57910 31563 -57831
rect 30984 -58265 31063 -57910
rect 30958 -58362 31074 -58265
rect 32985 -58393 33424 -58346
rect 31587 -58409 31684 -58403
rect 31587 -58463 32696 -58409
rect 32985 -58430 33032 -58393
rect 31587 -58469 31684 -58463
rect 30412 -58870 31120 -58757
rect 30025 -59005 30071 -58905
rect 30123 -59034 30169 -58905
rect 30221 -59005 30267 -58905
rect 30319 -59034 30365 -58905
rect 30025 -59080 30662 -59034
rect 30025 -59236 30071 -59080
rect 30123 -59082 30365 -59080
rect 30221 -59236 30267 -59082
rect 30417 -59236 30463 -59080
rect 28417 -60135 28463 -59835
rect 28064 -60330 28261 -60276
rect 28319 -60671 28365 -60372
rect 28318 -60708 28365 -60671
rect 28417 -60672 28463 -60372
rect 28515 -60708 28561 -60372
rect 28613 -60672 28659 -59835
rect 29026 -59990 29072 -59834
rect 29222 -59988 29268 -59834
rect 29124 -59990 29366 -59988
rect 29418 -59990 29464 -59834
rect 29026 -60036 29663 -59990
rect 29026 -60165 29072 -60065
rect 29124 -60165 29170 -60036
rect 29222 -60165 29268 -60065
rect 29320 -60165 29366 -60036
rect 29864 -60346 29910 -59746
rect 30075 -60346 30121 -59746
rect 30173 -60346 30219 -59746
rect 30271 -60346 30317 -59746
rect 30483 -60346 30529 -59746
rect 28711 -60708 28757 -60372
rect 30714 -60477 30819 -60405
rect 30720 -60560 30785 -60477
rect 29765 -60625 30785 -60560
rect 28318 -60755 28757 -60708
rect 29864 -60958 29910 -60658
rect 29962 -60958 30008 -60658
rect 30060 -60958 30106 -60658
rect 30302 -60958 30348 -60658
rect 30400 -60958 30446 -60658
rect 31007 -61066 31120 -58870
rect 31825 -58903 31955 -58753
rect 32111 -58807 32157 -58607
rect 32209 -58835 32255 -58607
rect 32307 -58807 32353 -58607
rect 32405 -58835 32451 -58607
rect 32642 -58753 32696 -58463
rect 32986 -58729 33032 -58430
rect 33084 -58729 33130 -58429
rect 33182 -58729 33228 -58393
rect 32642 -58807 32970 -58753
rect 32111 -58881 32748 -58835
rect 32916 -58862 32970 -58807
rect 31875 -60307 31929 -58903
rect 32111 -59137 32157 -58881
rect 32209 -58883 32451 -58881
rect 32307 -59137 32353 -58883
rect 32503 -59137 32549 -58881
rect 32890 -58920 33049 -58862
rect 33084 -59266 33130 -58966
rect 33280 -59266 33326 -58429
rect 33378 -58729 33424 -58393
rect 34080 -58901 34788 -58788
rect 33693 -59036 33739 -58936
rect 33791 -59065 33837 -58936
rect 33889 -59036 33935 -58936
rect 33987 -59065 34033 -58936
rect 33693 -59111 34330 -59065
rect 33693 -59267 33739 -59111
rect 33791 -59113 34033 -59111
rect 33889 -59267 33935 -59113
rect 34085 -59267 34131 -59111
rect 32085 -60166 32131 -59866
rect 31732 -60361 31929 -60307
rect 31987 -60702 32033 -60403
rect 31986 -60739 32033 -60702
rect 32085 -60703 32131 -60403
rect 32183 -60739 32229 -60403
rect 32281 -60703 32327 -59866
rect 32694 -60021 32740 -59865
rect 32890 -60019 32936 -59865
rect 32792 -60021 33034 -60019
rect 33086 -60021 33132 -59865
rect 32694 -60067 33331 -60021
rect 32694 -60196 32740 -60096
rect 32792 -60196 32838 -60067
rect 32890 -60196 32936 -60096
rect 32988 -60196 33034 -60067
rect 33532 -60377 33578 -59777
rect 33743 -60377 33789 -59777
rect 33841 -60377 33887 -59777
rect 33939 -60377 33985 -59777
rect 34151 -60377 34197 -59777
rect 32379 -60739 32425 -60403
rect 34382 -60508 34487 -60436
rect 34388 -60591 34453 -60508
rect 33433 -60656 34453 -60591
rect 31986 -60786 32425 -60739
rect 33532 -60989 33578 -60689
rect 33630 -60989 33676 -60689
rect 33728 -60989 33774 -60689
rect 33970 -60989 34016 -60689
rect 34068 -60989 34114 -60689
rect 30443 -61097 31120 -61066
rect 34675 -61097 34788 -58901
rect 34872 -60522 35121 -55033
rect 35283 -58306 35474 -54592
rect 35959 -54936 36316 -54800
rect 37765 -54920 38204 -54873
rect 35959 -54990 37476 -54936
rect 37765 -54957 37812 -54920
rect 35959 -55067 36316 -54990
rect 36605 -55430 36735 -55280
rect 36891 -55334 36937 -55134
rect 36989 -55362 37035 -55134
rect 37087 -55334 37133 -55134
rect 37185 -55362 37231 -55134
rect 37422 -55280 37476 -54990
rect 37766 -55256 37812 -54957
rect 37864 -55256 37910 -54956
rect 37962 -55256 38008 -54920
rect 37422 -55334 37750 -55280
rect 36891 -55408 37528 -55362
rect 37696 -55389 37750 -55334
rect 36655 -56834 36709 -55430
rect 36891 -55664 36937 -55408
rect 36989 -55410 37231 -55408
rect 37087 -55664 37133 -55410
rect 37283 -55664 37329 -55408
rect 37670 -55447 37829 -55389
rect 37864 -55793 37910 -55493
rect 38060 -55793 38106 -54956
rect 38158 -55256 38204 -54920
rect 38860 -55428 39568 -55315
rect 38473 -55563 38519 -55463
rect 38571 -55592 38617 -55463
rect 38669 -55563 38715 -55463
rect 38767 -55592 38813 -55463
rect 38473 -55638 39110 -55592
rect 38473 -55794 38519 -55638
rect 38571 -55640 38813 -55638
rect 38669 -55794 38715 -55640
rect 38865 -55794 38911 -55638
rect 36865 -56693 36911 -56393
rect 36512 -56888 36709 -56834
rect 36767 -57229 36813 -56930
rect 36766 -57266 36813 -57229
rect 36865 -57230 36911 -56930
rect 36963 -57266 37009 -56930
rect 37061 -57230 37107 -56393
rect 37474 -56548 37520 -56392
rect 37670 -56546 37716 -56392
rect 37572 -56548 37814 -56546
rect 37866 -56548 37912 -56392
rect 37474 -56594 38111 -56548
rect 37474 -56723 37520 -56623
rect 37572 -56723 37618 -56594
rect 37670 -56723 37716 -56623
rect 37768 -56723 37814 -56594
rect 38312 -56904 38358 -56304
rect 38523 -56904 38569 -56304
rect 38621 -56904 38667 -56304
rect 38719 -56904 38765 -56304
rect 38931 -56904 38977 -56304
rect 37159 -57266 37205 -56930
rect 39162 -57035 39267 -56963
rect 39168 -57118 39233 -57035
rect 38213 -57183 39233 -57118
rect 36766 -57313 37205 -57266
rect 38312 -57516 38358 -57216
rect 38410 -57516 38456 -57216
rect 38508 -57516 38554 -57216
rect 38750 -57516 38796 -57216
rect 38848 -57516 38894 -57216
rect 39081 -57624 39194 -57623
rect 39455 -57624 39568 -55428
rect 40304 -56662 40350 -56162
rect 40573 -56662 40619 -56162
rect 40671 -56662 40717 -56162
rect 40769 -56662 40815 -56162
rect 40899 -56662 40945 -56162
rect 41225 -56662 41271 -56162
rect 41453 -56462 41499 -56162
rect 40073 -56822 40211 -56818
rect 40879 -56822 41017 -56818
rect 41264 -56822 41318 -56749
rect 40073 -56866 41318 -56822
rect 40073 -56872 40211 -56866
rect 40879 -56872 41017 -56866
rect 41264 -56887 41318 -56866
rect 41436 -56902 41502 -56890
rect 42149 -56902 42365 -54592
rect 39912 -57209 40015 -57118
rect 38891 -57737 39568 -57624
rect 35283 -58389 36133 -58306
rect 37757 -58373 38196 -58326
rect 35283 -58443 37468 -58389
rect 37757 -58410 37804 -58373
rect 35283 -58497 36133 -58443
rect 36597 -58883 36727 -58733
rect 36883 -58787 36929 -58587
rect 36981 -58815 37027 -58587
rect 37079 -58787 37125 -58587
rect 37177 -58815 37223 -58587
rect 37414 -58733 37468 -58443
rect 37758 -58709 37804 -58410
rect 37856 -58709 37902 -58409
rect 37954 -58709 38000 -58373
rect 37414 -58787 37742 -58733
rect 36883 -58861 37520 -58815
rect 37688 -58842 37742 -58787
rect 36647 -60287 36701 -58883
rect 36883 -59117 36929 -58861
rect 36981 -58863 37223 -58861
rect 37079 -59117 37125 -58863
rect 37275 -59117 37321 -58861
rect 37662 -58900 37821 -58842
rect 37856 -59246 37902 -58946
rect 38052 -59246 38098 -58409
rect 38150 -58709 38196 -58373
rect 39081 -58768 39194 -57737
rect 39924 -57842 40003 -57209
rect 40206 -57458 40252 -57158
rect 40304 -57458 40350 -57158
rect 40676 -57458 40722 -56958
rect 40774 -57458 40820 -56958
rect 40899 -57458 40945 -56958
rect 40997 -57458 41043 -56958
rect 41127 -57458 41173 -56958
rect 41225 -57458 41271 -56958
rect 41323 -57458 41369 -56958
rect 41436 -56964 43058 -56902
rect 41436 -56973 41502 -56964
rect 41453 -57458 41499 -57158
rect 41551 -57458 41597 -57158
rect 39424 -57921 40003 -57842
rect 39424 -58276 39503 -57921
rect 39398 -58373 39514 -58276
rect 41425 -58404 41864 -58357
rect 40027 -58420 40124 -58414
rect 40027 -58474 41136 -58420
rect 41425 -58441 41472 -58404
rect 40027 -58480 40124 -58474
rect 38852 -58881 39560 -58768
rect 38465 -59016 38511 -58916
rect 38563 -59045 38609 -58916
rect 38661 -59016 38707 -58916
rect 38759 -59045 38805 -58916
rect 38465 -59091 39102 -59045
rect 38465 -59247 38511 -59091
rect 38563 -59093 38805 -59091
rect 38661 -59247 38707 -59093
rect 38857 -59247 38903 -59091
rect 36857 -60146 36903 -59846
rect 36504 -60341 36701 -60287
rect 34888 -60691 35111 -60522
rect 36759 -60682 36805 -60383
rect 36758 -60719 36805 -60682
rect 36857 -60683 36903 -60383
rect 36955 -60719 37001 -60383
rect 37053 -60683 37099 -59846
rect 37466 -60001 37512 -59845
rect 37662 -59999 37708 -59845
rect 37564 -60001 37806 -59999
rect 37858 -60001 37904 -59845
rect 37466 -60047 38103 -60001
rect 37466 -60176 37512 -60076
rect 37564 -60176 37610 -60047
rect 37662 -60176 37708 -60076
rect 37760 -60176 37806 -60047
rect 38304 -60357 38350 -59757
rect 38515 -60357 38561 -59757
rect 38613 -60357 38659 -59757
rect 38711 -60357 38757 -59757
rect 38923 -60357 38969 -59757
rect 37151 -60719 37197 -60383
rect 39154 -60488 39259 -60416
rect 39160 -60571 39225 -60488
rect 38205 -60636 39225 -60571
rect 36758 -60766 37197 -60719
rect 38304 -60969 38350 -60669
rect 38402 -60969 38448 -60669
rect 38500 -60969 38546 -60669
rect 38742 -60969 38788 -60669
rect 38840 -60969 38886 -60669
rect 39447 -61077 39560 -58881
rect 40265 -58914 40395 -58764
rect 40551 -58818 40597 -58618
rect 40649 -58846 40695 -58618
rect 40747 -58818 40793 -58618
rect 40845 -58846 40891 -58618
rect 41082 -58764 41136 -58474
rect 41426 -58740 41472 -58441
rect 41524 -58740 41570 -58440
rect 41622 -58740 41668 -58404
rect 41082 -58818 41410 -58764
rect 40551 -58892 41188 -58846
rect 41356 -58873 41410 -58818
rect 40315 -60318 40369 -58914
rect 40551 -59148 40597 -58892
rect 40649 -58894 40891 -58892
rect 40747 -59148 40793 -58894
rect 40943 -59148 40989 -58892
rect 41330 -58931 41489 -58873
rect 41524 -59277 41570 -58977
rect 41720 -59277 41766 -58440
rect 41818 -58740 41864 -58404
rect 42520 -58912 43228 -58799
rect 42133 -59047 42179 -58947
rect 42231 -59076 42277 -58947
rect 42329 -59047 42375 -58947
rect 42427 -59076 42473 -58947
rect 42133 -59122 42770 -59076
rect 42133 -59278 42179 -59122
rect 42231 -59124 42473 -59122
rect 42329 -59278 42375 -59124
rect 42525 -59278 42571 -59122
rect 40525 -60177 40571 -59877
rect 40172 -60372 40369 -60318
rect 40427 -60713 40473 -60414
rect 40426 -60750 40473 -60713
rect 40525 -60714 40571 -60414
rect 40623 -60750 40669 -60414
rect 40721 -60714 40767 -59877
rect 41134 -60032 41180 -59876
rect 41330 -60030 41376 -59876
rect 41232 -60032 41474 -60030
rect 41526 -60032 41572 -59876
rect 41134 -60078 41771 -60032
rect 41134 -60207 41180 -60107
rect 41232 -60207 41278 -60078
rect 41330 -60207 41376 -60107
rect 41428 -60207 41474 -60078
rect 41972 -60388 42018 -59788
rect 42183 -60388 42229 -59788
rect 42281 -60388 42327 -59788
rect 42379 -60388 42425 -59788
rect 42591 -60388 42637 -59788
rect 40819 -60750 40865 -60414
rect 42822 -60519 42927 -60447
rect 42828 -60602 42893 -60519
rect 41873 -60667 42893 -60602
rect 40426 -60797 40865 -60750
rect 41972 -61000 42018 -60700
rect 42070 -61000 42116 -60700
rect 42168 -61000 42214 -60700
rect 42410 -61000 42456 -60700
rect 42508 -61000 42554 -60700
rect 30443 -61179 34788 -61097
rect 30447 -61210 34788 -61179
rect 38883 -61108 39560 -61077
rect 43115 -61108 43228 -58912
rect 43337 -60459 43602 -53126
rect 43779 -54585 51740 -54383
rect 43779 -58375 43981 -54585
rect 44863 -54975 45160 -54889
rect 46628 -54959 47067 -54912
rect 44863 -55029 46339 -54975
rect 46628 -54996 46675 -54959
rect 44863 -55111 45160 -55029
rect 45468 -55469 45598 -55319
rect 45754 -55373 45800 -55173
rect 45852 -55401 45898 -55173
rect 45950 -55373 45996 -55173
rect 46048 -55401 46094 -55173
rect 46285 -55319 46339 -55029
rect 46629 -55295 46675 -54996
rect 46727 -55295 46773 -54995
rect 46825 -55295 46871 -54959
rect 46285 -55373 46613 -55319
rect 45754 -55447 46391 -55401
rect 46559 -55428 46613 -55373
rect 45518 -56873 45572 -55469
rect 45754 -55703 45800 -55447
rect 45852 -55449 46094 -55447
rect 45950 -55703 45996 -55449
rect 46146 -55703 46192 -55447
rect 46533 -55486 46692 -55428
rect 46727 -55832 46773 -55532
rect 46923 -55832 46969 -54995
rect 47021 -55295 47067 -54959
rect 47723 -55467 48431 -55354
rect 47336 -55602 47382 -55502
rect 47434 -55631 47480 -55502
rect 47532 -55602 47578 -55502
rect 47630 -55631 47676 -55502
rect 47336 -55677 47973 -55631
rect 47336 -55833 47382 -55677
rect 47434 -55679 47676 -55677
rect 47532 -55833 47578 -55679
rect 47728 -55833 47774 -55677
rect 45728 -56732 45774 -56432
rect 45375 -56927 45572 -56873
rect 45630 -57268 45676 -56969
rect 45629 -57305 45676 -57268
rect 45728 -57269 45774 -56969
rect 45826 -57305 45872 -56969
rect 45924 -57269 45970 -56432
rect 46337 -56587 46383 -56431
rect 46533 -56585 46579 -56431
rect 46435 -56587 46677 -56585
rect 46729 -56587 46775 -56431
rect 46337 -56633 46974 -56587
rect 46337 -56762 46383 -56662
rect 46435 -56762 46481 -56633
rect 46533 -56762 46579 -56662
rect 46631 -56762 46677 -56633
rect 47175 -56943 47221 -56343
rect 47386 -56943 47432 -56343
rect 47484 -56943 47530 -56343
rect 47582 -56943 47628 -56343
rect 47794 -56943 47840 -56343
rect 46022 -57305 46068 -56969
rect 48025 -57074 48130 -57002
rect 48031 -57157 48096 -57074
rect 47076 -57222 48096 -57157
rect 45629 -57352 46068 -57305
rect 47175 -57555 47221 -57255
rect 47273 -57555 47319 -57255
rect 47371 -57555 47417 -57255
rect 47613 -57555 47659 -57255
rect 47711 -57555 47757 -57255
rect 47944 -57663 48057 -57662
rect 48318 -57663 48431 -55467
rect 49167 -56701 49213 -56201
rect 49436 -56701 49482 -56201
rect 49534 -56701 49580 -56201
rect 49632 -56701 49678 -56201
rect 49762 -56701 49808 -56201
rect 50088 -56701 50134 -56201
rect 50316 -56501 50362 -56201
rect 48936 -56861 49074 -56857
rect 49742 -56861 49880 -56857
rect 50127 -56861 50181 -56788
rect 48936 -56905 50181 -56861
rect 48936 -56911 49074 -56905
rect 49742 -56911 49880 -56905
rect 50127 -56926 50181 -56905
rect 50299 -56941 50365 -56929
rect 51538 -56941 51740 -54585
rect 48775 -57248 48878 -57157
rect 47754 -57776 48431 -57663
rect 43779 -58428 45109 -58375
rect 46620 -58412 47059 -58365
rect 43779 -58482 46331 -58428
rect 46620 -58449 46667 -58412
rect 43779 -58577 45109 -58482
rect 45460 -58922 45590 -58772
rect 45746 -58826 45792 -58626
rect 45844 -58854 45890 -58626
rect 45942 -58826 45988 -58626
rect 46040 -58854 46086 -58626
rect 46277 -58772 46331 -58482
rect 46621 -58748 46667 -58449
rect 46719 -58748 46765 -58448
rect 46817 -58748 46863 -58412
rect 46277 -58826 46605 -58772
rect 45746 -58900 46383 -58854
rect 46551 -58881 46605 -58826
rect 45510 -60326 45564 -58922
rect 45746 -59156 45792 -58900
rect 45844 -58902 46086 -58900
rect 45942 -59156 45988 -58902
rect 46138 -59156 46184 -58900
rect 46525 -58939 46684 -58881
rect 46719 -59285 46765 -58985
rect 46915 -59285 46961 -58448
rect 47013 -58748 47059 -58412
rect 47944 -58807 48057 -57776
rect 48787 -57881 48866 -57248
rect 49069 -57497 49115 -57197
rect 49167 -57497 49213 -57197
rect 49539 -57497 49585 -56997
rect 49637 -57497 49683 -56997
rect 49762 -57497 49808 -56997
rect 49860 -57497 49906 -56997
rect 49990 -57497 50036 -56997
rect 50088 -57497 50134 -56997
rect 50186 -57497 50232 -56997
rect 50299 -57003 51921 -56941
rect 50299 -57012 50365 -57003
rect 50316 -57497 50362 -57197
rect 50414 -57497 50460 -57197
rect 48287 -57960 48866 -57881
rect 48287 -58315 48366 -57960
rect 48261 -58412 48377 -58315
rect 50288 -58443 50727 -58396
rect 48890 -58459 48987 -58453
rect 48890 -58513 49999 -58459
rect 50288 -58480 50335 -58443
rect 48890 -58519 48987 -58513
rect 47715 -58920 48423 -58807
rect 47328 -59055 47374 -58955
rect 47426 -59084 47472 -58955
rect 47524 -59055 47570 -58955
rect 47622 -59084 47668 -58955
rect 47328 -59130 47965 -59084
rect 47328 -59286 47374 -59130
rect 47426 -59132 47668 -59130
rect 47524 -59286 47570 -59132
rect 47720 -59286 47766 -59130
rect 45720 -60185 45766 -59885
rect 45367 -60380 45564 -60326
rect 43337 -60790 43674 -60459
rect 45622 -60721 45668 -60422
rect 45621 -60758 45668 -60721
rect 45720 -60722 45766 -60422
rect 45818 -60758 45864 -60422
rect 45916 -60722 45962 -59885
rect 46329 -60040 46375 -59884
rect 46525 -60038 46571 -59884
rect 46427 -60040 46669 -60038
rect 46721 -60040 46767 -59884
rect 46329 -60086 46966 -60040
rect 46329 -60215 46375 -60115
rect 46427 -60215 46473 -60086
rect 46525 -60215 46571 -60115
rect 46623 -60215 46669 -60086
rect 47167 -60396 47213 -59796
rect 47378 -60396 47424 -59796
rect 47476 -60396 47522 -59796
rect 47574 -60396 47620 -59796
rect 47786 -60396 47832 -59796
rect 46014 -60758 46060 -60422
rect 48017 -60527 48122 -60455
rect 48023 -60610 48088 -60527
rect 47068 -60675 48088 -60610
rect 45621 -60805 46060 -60758
rect 47167 -61008 47213 -60708
rect 47265 -61008 47311 -60708
rect 47363 -61008 47409 -60708
rect 47605 -61008 47651 -60708
rect 47703 -61008 47749 -60708
rect 38883 -61190 43228 -61108
rect 48310 -61116 48423 -58920
rect 49128 -58953 49258 -58803
rect 49414 -58857 49460 -58657
rect 49512 -58885 49558 -58657
rect 49610 -58857 49656 -58657
rect 49708 -58885 49754 -58657
rect 49945 -58803 49999 -58513
rect 50289 -58779 50335 -58480
rect 50387 -58779 50433 -58479
rect 50485 -58779 50531 -58443
rect 49945 -58857 50273 -58803
rect 49414 -58931 50051 -58885
rect 50219 -58912 50273 -58857
rect 49178 -60357 49232 -58953
rect 49414 -59187 49460 -58931
rect 49512 -58933 49754 -58931
rect 49610 -59187 49656 -58933
rect 49806 -59187 49852 -58931
rect 50193 -58970 50352 -58912
rect 50387 -59316 50433 -59016
rect 50583 -59316 50629 -58479
rect 50681 -58779 50727 -58443
rect 51383 -58951 52091 -58838
rect 50996 -59086 51042 -58986
rect 51094 -59115 51140 -58986
rect 51192 -59086 51238 -58986
rect 51290 -59115 51336 -58986
rect 50996 -59161 51633 -59115
rect 50996 -59317 51042 -59161
rect 51094 -59163 51336 -59161
rect 51192 -59317 51238 -59163
rect 51388 -59317 51434 -59161
rect 49388 -60216 49434 -59916
rect 49035 -60411 49232 -60357
rect 49290 -60752 49336 -60453
rect 49289 -60789 49336 -60752
rect 49388 -60753 49434 -60453
rect 49486 -60789 49532 -60453
rect 49584 -60753 49630 -59916
rect 49997 -60071 50043 -59915
rect 50193 -60069 50239 -59915
rect 50095 -60071 50337 -60069
rect 50389 -60071 50435 -59915
rect 49997 -60117 50634 -60071
rect 49997 -60246 50043 -60146
rect 50095 -60246 50141 -60117
rect 50193 -60246 50239 -60146
rect 50291 -60246 50337 -60117
rect 50835 -60427 50881 -59827
rect 51046 -60427 51092 -59827
rect 51144 -60427 51190 -59827
rect 51242 -60427 51288 -59827
rect 51454 -60427 51500 -59827
rect 49682 -60789 49728 -60453
rect 51685 -60558 51790 -60486
rect 51691 -60641 51756 -60558
rect 50736 -60706 51756 -60641
rect 49289 -60836 49728 -60789
rect 50835 -61039 50881 -60739
rect 50933 -61039 50979 -60739
rect 51031 -61039 51077 -60739
rect 51273 -61039 51319 -60739
rect 51371 -61039 51417 -60739
rect 38887 -61221 43228 -61190
rect 47746 -61147 48423 -61116
rect 51978 -61147 52091 -58951
rect 52201 -60320 52427 -52646
rect 53058 -54650 61044 -54391
rect 53058 -58254 53317 -54650
rect 53854 -54941 54100 -54845
rect 55826 -54925 56265 -54878
rect 53854 -54995 55537 -54941
rect 55826 -54962 55873 -54925
rect 53854 -55065 54100 -54995
rect 54666 -55435 54796 -55285
rect 54952 -55339 54998 -55139
rect 55050 -55367 55096 -55139
rect 55148 -55339 55194 -55139
rect 55246 -55367 55292 -55139
rect 55483 -55285 55537 -54995
rect 55827 -55261 55873 -54962
rect 55925 -55261 55971 -54961
rect 56023 -55261 56069 -54925
rect 55483 -55339 55811 -55285
rect 54952 -55413 55589 -55367
rect 55757 -55394 55811 -55339
rect 54716 -56839 54770 -55435
rect 54952 -55669 54998 -55413
rect 55050 -55415 55292 -55413
rect 55148 -55669 55194 -55415
rect 55344 -55669 55390 -55413
rect 55731 -55452 55890 -55394
rect 55925 -55798 55971 -55498
rect 56121 -55798 56167 -54961
rect 56219 -55261 56265 -54925
rect 56921 -55433 57629 -55320
rect 56534 -55568 56580 -55468
rect 56632 -55597 56678 -55468
rect 56730 -55568 56776 -55468
rect 56828 -55597 56874 -55468
rect 56534 -55643 57171 -55597
rect 56534 -55799 56580 -55643
rect 56632 -55645 56874 -55643
rect 56730 -55799 56776 -55645
rect 56926 -55799 56972 -55643
rect 54926 -56698 54972 -56398
rect 54573 -56893 54770 -56839
rect 54828 -57234 54874 -56935
rect 54827 -57271 54874 -57234
rect 54926 -57235 54972 -56935
rect 55024 -57271 55070 -56935
rect 55122 -57235 55168 -56398
rect 55535 -56553 55581 -56397
rect 55731 -56551 55777 -56397
rect 55633 -56553 55875 -56551
rect 55927 -56553 55973 -56397
rect 55535 -56599 56172 -56553
rect 55535 -56728 55581 -56628
rect 55633 -56728 55679 -56599
rect 55731 -56728 55777 -56628
rect 55829 -56728 55875 -56599
rect 56373 -56909 56419 -56309
rect 56584 -56909 56630 -56309
rect 56682 -56909 56728 -56309
rect 56780 -56909 56826 -56309
rect 56992 -56909 57038 -56309
rect 55220 -57271 55266 -56935
rect 57223 -57040 57328 -56968
rect 57229 -57123 57294 -57040
rect 56274 -57188 57294 -57123
rect 54827 -57318 55266 -57271
rect 56373 -57521 56419 -57221
rect 56471 -57521 56517 -57221
rect 56569 -57521 56615 -57221
rect 56811 -57521 56857 -57221
rect 56909 -57521 56955 -57221
rect 57142 -57629 57255 -57628
rect 57516 -57629 57629 -55433
rect 58365 -56667 58411 -56167
rect 58634 -56667 58680 -56167
rect 58732 -56667 58778 -56167
rect 58830 -56667 58876 -56167
rect 58960 -56667 59006 -56167
rect 59286 -56667 59332 -56167
rect 59514 -56467 59560 -56167
rect 58134 -56827 58272 -56823
rect 58940 -56827 59078 -56823
rect 59325 -56827 59379 -56754
rect 58134 -56871 59379 -56827
rect 58134 -56877 58272 -56871
rect 58940 -56877 59078 -56871
rect 59325 -56892 59379 -56871
rect 59497 -56907 59563 -56895
rect 60785 -56907 61044 -54650
rect 61395 -54707 61616 -52089
rect 61847 -54670 69831 -54432
rect 61292 -55021 61668 -54707
rect 57973 -57214 58076 -57123
rect 56952 -57742 57629 -57629
rect 53058 -58394 54266 -58254
rect 55818 -58378 56257 -58331
rect 53058 -58448 55529 -58394
rect 55818 -58415 55865 -58378
rect 53058 -58513 54266 -58448
rect 54658 -58888 54788 -58738
rect 54944 -58792 54990 -58592
rect 55042 -58820 55088 -58592
rect 55140 -58792 55186 -58592
rect 55238 -58820 55284 -58592
rect 55475 -58738 55529 -58448
rect 55819 -58714 55865 -58415
rect 55917 -58714 55963 -58414
rect 56015 -58714 56061 -58378
rect 55475 -58792 55803 -58738
rect 54944 -58866 55581 -58820
rect 55749 -58847 55803 -58792
rect 54708 -60292 54762 -58888
rect 54944 -59122 54990 -58866
rect 55042 -58868 55284 -58866
rect 55140 -59122 55186 -58868
rect 55336 -59122 55382 -58866
rect 55723 -58905 55882 -58847
rect 55917 -59251 55963 -58951
rect 56113 -59251 56159 -58414
rect 56211 -58714 56257 -58378
rect 57142 -58773 57255 -57742
rect 57985 -57847 58064 -57214
rect 58267 -57463 58313 -57163
rect 58365 -57463 58411 -57163
rect 58737 -57463 58783 -56963
rect 58835 -57463 58881 -56963
rect 58960 -57463 59006 -56963
rect 59058 -57463 59104 -56963
rect 59188 -57463 59234 -56963
rect 59286 -57463 59332 -56963
rect 59384 -57463 59430 -56963
rect 59497 -56969 61119 -56907
rect 59497 -56978 59563 -56969
rect 59514 -57463 59560 -57163
rect 59612 -57463 59658 -57163
rect 57485 -57926 58064 -57847
rect 57485 -58281 57564 -57926
rect 57459 -58378 57575 -58281
rect 59486 -58409 59925 -58362
rect 58088 -58425 58185 -58419
rect 58088 -58479 59197 -58425
rect 59486 -58446 59533 -58409
rect 58088 -58485 58185 -58479
rect 56913 -58886 57621 -58773
rect 56526 -59021 56572 -58921
rect 56624 -59050 56670 -58921
rect 56722 -59021 56768 -58921
rect 56820 -59050 56866 -58921
rect 56526 -59096 57163 -59050
rect 56526 -59252 56572 -59096
rect 56624 -59098 56866 -59096
rect 56722 -59252 56768 -59098
rect 56918 -59252 56964 -59096
rect 54918 -60151 54964 -59851
rect 52179 -60820 52477 -60320
rect 54565 -60346 54762 -60292
rect 54820 -60687 54866 -60388
rect 54819 -60724 54866 -60687
rect 54918 -60688 54964 -60388
rect 55016 -60724 55062 -60388
rect 55114 -60688 55160 -59851
rect 55527 -60006 55573 -59850
rect 55723 -60004 55769 -59850
rect 55625 -60006 55867 -60004
rect 55919 -60006 55965 -59850
rect 55527 -60052 56164 -60006
rect 55527 -60181 55573 -60081
rect 55625 -60181 55671 -60052
rect 55723 -60181 55769 -60081
rect 55821 -60181 55867 -60052
rect 56365 -60362 56411 -59762
rect 56576 -60362 56622 -59762
rect 56674 -60362 56720 -59762
rect 56772 -60362 56818 -59762
rect 56984 -60362 57030 -59762
rect 55212 -60724 55258 -60388
rect 57215 -60493 57320 -60421
rect 57221 -60576 57286 -60493
rect 56266 -60641 57286 -60576
rect 54819 -60771 55258 -60724
rect 56365 -60974 56411 -60674
rect 56463 -60974 56509 -60674
rect 56561 -60974 56607 -60674
rect 56803 -60974 56849 -60674
rect 56901 -60974 56947 -60674
rect 57508 -61082 57621 -58886
rect 58326 -58919 58456 -58769
rect 58612 -58823 58658 -58623
rect 58710 -58851 58756 -58623
rect 58808 -58823 58854 -58623
rect 58906 -58851 58952 -58623
rect 59143 -58769 59197 -58479
rect 59487 -58745 59533 -58446
rect 59585 -58745 59631 -58445
rect 59683 -58745 59729 -58409
rect 59143 -58823 59471 -58769
rect 58612 -58897 59249 -58851
rect 59417 -58878 59471 -58823
rect 58376 -60323 58430 -58919
rect 58612 -59153 58658 -58897
rect 58710 -58899 58952 -58897
rect 58808 -59153 58854 -58899
rect 59004 -59153 59050 -58897
rect 59391 -58936 59550 -58878
rect 59585 -59282 59631 -58982
rect 59781 -59282 59827 -58445
rect 59879 -58745 59925 -58409
rect 60581 -58917 61289 -58804
rect 60194 -59052 60240 -58952
rect 60292 -59081 60338 -58952
rect 60390 -59052 60436 -58952
rect 60488 -59081 60534 -58952
rect 60194 -59127 60831 -59081
rect 60194 -59283 60240 -59127
rect 60292 -59129 60534 -59127
rect 60390 -59283 60436 -59129
rect 60586 -59283 60632 -59127
rect 58586 -60182 58632 -59882
rect 58233 -60377 58430 -60323
rect 58488 -60718 58534 -60419
rect 58487 -60755 58534 -60718
rect 58586 -60719 58632 -60419
rect 58684 -60755 58730 -60419
rect 58782 -60719 58828 -59882
rect 59195 -60037 59241 -59881
rect 59391 -60035 59437 -59881
rect 59293 -60037 59535 -60035
rect 59587 -60037 59633 -59881
rect 59195 -60083 59832 -60037
rect 59195 -60212 59241 -60112
rect 59293 -60212 59339 -60083
rect 59391 -60212 59437 -60112
rect 59489 -60212 59535 -60083
rect 60033 -60393 60079 -59793
rect 60244 -60393 60290 -59793
rect 60342 -60393 60388 -59793
rect 60440 -60393 60486 -59793
rect 60652 -60393 60698 -59793
rect 58880 -60755 58926 -60419
rect 60883 -60524 60988 -60452
rect 60889 -60607 60954 -60524
rect 59934 -60672 60954 -60607
rect 58487 -60802 58926 -60755
rect 60033 -61005 60079 -60705
rect 60131 -61005 60177 -60705
rect 60229 -61005 60275 -60705
rect 60471 -61005 60517 -60705
rect 60569 -61005 60615 -60705
rect 47746 -61229 52091 -61147
rect 56944 -61113 57621 -61082
rect 61176 -61113 61289 -58917
rect 61395 -60458 61616 -55021
rect 61847 -58194 62085 -54670
rect 62893 -54875 63143 -54775
rect 64580 -54859 65019 -54812
rect 62893 -54929 64291 -54875
rect 64580 -54896 64627 -54859
rect 62893 -55004 63143 -54929
rect 63420 -55369 63550 -55219
rect 63706 -55273 63752 -55073
rect 63804 -55301 63850 -55073
rect 63902 -55273 63948 -55073
rect 64000 -55301 64046 -55073
rect 64237 -55219 64291 -54929
rect 64581 -55195 64627 -54896
rect 64679 -55195 64725 -54895
rect 64777 -55195 64823 -54859
rect 64237 -55273 64565 -55219
rect 63706 -55347 64343 -55301
rect 64511 -55328 64565 -55273
rect 63470 -56773 63524 -55369
rect 63706 -55603 63752 -55347
rect 63804 -55349 64046 -55347
rect 63902 -55603 63948 -55349
rect 64098 -55603 64144 -55347
rect 64485 -55386 64644 -55328
rect 64679 -55732 64725 -55432
rect 64875 -55732 64921 -54895
rect 64973 -55195 65019 -54859
rect 65675 -55367 66383 -55254
rect 65288 -55502 65334 -55402
rect 65386 -55531 65432 -55402
rect 65484 -55502 65530 -55402
rect 65582 -55531 65628 -55402
rect 65288 -55577 65925 -55531
rect 65288 -55733 65334 -55577
rect 65386 -55579 65628 -55577
rect 65484 -55733 65530 -55579
rect 65680 -55733 65726 -55577
rect 63680 -56632 63726 -56332
rect 63327 -56827 63524 -56773
rect 63582 -57168 63628 -56869
rect 63581 -57205 63628 -57168
rect 63680 -57169 63726 -56869
rect 63778 -57205 63824 -56869
rect 63876 -57169 63922 -56332
rect 64289 -56487 64335 -56331
rect 64485 -56485 64531 -56331
rect 64387 -56487 64629 -56485
rect 64681 -56487 64727 -56331
rect 64289 -56533 64926 -56487
rect 64289 -56662 64335 -56562
rect 64387 -56662 64433 -56533
rect 64485 -56662 64531 -56562
rect 64583 -56662 64629 -56533
rect 65127 -56843 65173 -56243
rect 65338 -56843 65384 -56243
rect 65436 -56843 65482 -56243
rect 65534 -56843 65580 -56243
rect 65746 -56843 65792 -56243
rect 63974 -57205 64020 -56869
rect 65977 -56974 66082 -56902
rect 65983 -57057 66048 -56974
rect 65028 -57122 66048 -57057
rect 63581 -57252 64020 -57205
rect 65127 -57455 65173 -57155
rect 65225 -57455 65271 -57155
rect 65323 -57455 65369 -57155
rect 65565 -57455 65611 -57155
rect 65663 -57455 65709 -57155
rect 65896 -57563 66009 -57562
rect 66270 -57563 66383 -55367
rect 67119 -56601 67165 -56101
rect 67388 -56601 67434 -56101
rect 67486 -56601 67532 -56101
rect 67584 -56601 67630 -56101
rect 67714 -56601 67760 -56101
rect 68040 -56601 68086 -56101
rect 68268 -56401 68314 -56101
rect 66888 -56761 67026 -56757
rect 67694 -56761 67832 -56757
rect 68079 -56761 68133 -56688
rect 66888 -56805 68133 -56761
rect 66888 -56811 67026 -56805
rect 67694 -56811 67832 -56805
rect 68079 -56826 68133 -56805
rect 68251 -56841 68317 -56829
rect 69593 -56841 69831 -54670
rect 70148 -54712 70325 -51530
rect 70633 -54678 79021 -54378
rect 70068 -55003 70406 -54712
rect 66727 -57148 66830 -57057
rect 65706 -57676 66383 -57563
rect 61847 -58328 62983 -58194
rect 64572 -58312 65011 -58265
rect 61847 -58382 64283 -58328
rect 64572 -58349 64619 -58312
rect 61847 -58432 62983 -58382
rect 63412 -58822 63542 -58672
rect 63698 -58726 63744 -58526
rect 63796 -58754 63842 -58526
rect 63894 -58726 63940 -58526
rect 63992 -58754 64038 -58526
rect 64229 -58672 64283 -58382
rect 64573 -58648 64619 -58349
rect 64671 -58648 64717 -58348
rect 64769 -58648 64815 -58312
rect 64229 -58726 64557 -58672
rect 63698 -58800 64335 -58754
rect 64503 -58781 64557 -58726
rect 63462 -60226 63516 -58822
rect 63698 -59056 63744 -58800
rect 63796 -58802 64038 -58800
rect 63894 -59056 63940 -58802
rect 64090 -59056 64136 -58800
rect 64477 -58839 64636 -58781
rect 64671 -59185 64717 -58885
rect 64867 -59185 64913 -58348
rect 64965 -58648 65011 -58312
rect 65896 -58707 66009 -57676
rect 66739 -57781 66818 -57148
rect 67021 -57397 67067 -57097
rect 67119 -57397 67165 -57097
rect 67491 -57397 67537 -56897
rect 67589 -57397 67635 -56897
rect 67714 -57397 67760 -56897
rect 67812 -57397 67858 -56897
rect 67942 -57397 67988 -56897
rect 68040 -57397 68086 -56897
rect 68138 -57397 68184 -56897
rect 68251 -56903 69873 -56841
rect 68251 -56912 68317 -56903
rect 68268 -57397 68314 -57097
rect 68366 -57397 68412 -57097
rect 66239 -57860 66818 -57781
rect 66239 -58215 66318 -57860
rect 66213 -58312 66329 -58215
rect 68240 -58343 68679 -58296
rect 66842 -58359 66939 -58353
rect 66842 -58413 67951 -58359
rect 68240 -58380 68287 -58343
rect 66842 -58419 66939 -58413
rect 65667 -58820 66375 -58707
rect 65280 -58955 65326 -58855
rect 65378 -58984 65424 -58855
rect 65476 -58955 65522 -58855
rect 65574 -58984 65620 -58855
rect 65280 -59030 65917 -58984
rect 65280 -59186 65326 -59030
rect 65378 -59032 65620 -59030
rect 65476 -59186 65522 -59032
rect 65672 -59186 65718 -59030
rect 63672 -60085 63718 -59785
rect 63319 -60280 63516 -60226
rect 61341 -60757 61633 -60458
rect 63574 -60621 63620 -60322
rect 63573 -60658 63620 -60621
rect 63672 -60622 63718 -60322
rect 63770 -60658 63816 -60322
rect 63868 -60622 63914 -59785
rect 64281 -59940 64327 -59784
rect 64477 -59938 64523 -59784
rect 64379 -59940 64621 -59938
rect 64673 -59940 64719 -59784
rect 64281 -59986 64918 -59940
rect 64281 -60115 64327 -60015
rect 64379 -60115 64425 -59986
rect 64477 -60115 64523 -60015
rect 64575 -60115 64621 -59986
rect 65119 -60296 65165 -59696
rect 65330 -60296 65376 -59696
rect 65428 -60296 65474 -59696
rect 65526 -60296 65572 -59696
rect 65738 -60296 65784 -59696
rect 63966 -60658 64012 -60322
rect 65969 -60427 66074 -60355
rect 65975 -60510 66040 -60427
rect 65020 -60575 66040 -60510
rect 63573 -60705 64012 -60658
rect 65119 -60908 65165 -60608
rect 65217 -60908 65263 -60608
rect 65315 -60908 65361 -60608
rect 65557 -60908 65603 -60608
rect 65655 -60908 65701 -60608
rect 66262 -61016 66375 -58820
rect 67080 -58853 67210 -58703
rect 67366 -58757 67412 -58557
rect 67464 -58785 67510 -58557
rect 67562 -58757 67608 -58557
rect 67660 -58785 67706 -58557
rect 67897 -58703 67951 -58413
rect 68241 -58679 68287 -58380
rect 68339 -58679 68385 -58379
rect 68437 -58679 68483 -58343
rect 67897 -58757 68225 -58703
rect 67366 -58831 68003 -58785
rect 68171 -58812 68225 -58757
rect 67130 -60257 67184 -58853
rect 67366 -59087 67412 -58831
rect 67464 -58833 67706 -58831
rect 67562 -59087 67608 -58833
rect 67758 -59087 67804 -58831
rect 68145 -58870 68304 -58812
rect 68339 -59216 68385 -58916
rect 68535 -59216 68581 -58379
rect 68633 -58679 68679 -58343
rect 69335 -58851 70043 -58738
rect 68948 -58986 68994 -58886
rect 69046 -59015 69092 -58886
rect 69144 -58986 69190 -58886
rect 69242 -59015 69288 -58886
rect 68948 -59061 69585 -59015
rect 68948 -59217 68994 -59061
rect 69046 -59063 69288 -59061
rect 69144 -59217 69190 -59063
rect 69340 -59217 69386 -59061
rect 67340 -60116 67386 -59816
rect 66987 -60311 67184 -60257
rect 67242 -60652 67288 -60353
rect 67241 -60689 67288 -60652
rect 67340 -60653 67386 -60353
rect 67438 -60689 67484 -60353
rect 67536 -60653 67582 -59816
rect 67949 -59971 67995 -59815
rect 68145 -59969 68191 -59815
rect 68047 -59971 68289 -59969
rect 68341 -59971 68387 -59815
rect 67949 -60017 68586 -59971
rect 67949 -60146 67995 -60046
rect 68047 -60146 68093 -60017
rect 68145 -60146 68191 -60046
rect 68243 -60146 68289 -60017
rect 68787 -60327 68833 -59727
rect 68998 -60327 69044 -59727
rect 69096 -60327 69142 -59727
rect 69194 -60327 69240 -59727
rect 69406 -60327 69452 -59727
rect 67634 -60689 67680 -60353
rect 69637 -60458 69742 -60386
rect 69643 -60541 69708 -60458
rect 68688 -60606 69708 -60541
rect 67241 -60736 67680 -60689
rect 68787 -60939 68833 -60639
rect 68885 -60939 68931 -60639
rect 68983 -60939 69029 -60639
rect 69225 -60939 69271 -60639
rect 69323 -60939 69369 -60639
rect 56944 -61195 61289 -61113
rect 65698 -61047 66375 -61016
rect 69930 -61047 70043 -58851
rect 70148 -60400 70325 -55003
rect 70633 -58128 70933 -54678
rect 72056 -54858 72324 -54767
rect 73733 -54842 74172 -54795
rect 72056 -54912 73444 -54858
rect 73733 -54879 73780 -54842
rect 72056 -55007 72324 -54912
rect 72573 -55352 72703 -55202
rect 72859 -55256 72905 -55056
rect 72957 -55284 73003 -55056
rect 73055 -55256 73101 -55056
rect 73153 -55284 73199 -55056
rect 73390 -55202 73444 -54912
rect 73734 -55178 73780 -54879
rect 73832 -55178 73878 -54878
rect 73930 -55178 73976 -54842
rect 73390 -55256 73718 -55202
rect 72859 -55330 73496 -55284
rect 73664 -55311 73718 -55256
rect 72623 -56756 72677 -55352
rect 72859 -55586 72905 -55330
rect 72957 -55332 73199 -55330
rect 73055 -55586 73101 -55332
rect 73251 -55586 73297 -55330
rect 73638 -55369 73797 -55311
rect 73832 -55715 73878 -55415
rect 74028 -55715 74074 -54878
rect 74126 -55178 74172 -54842
rect 74828 -55350 75536 -55237
rect 74441 -55485 74487 -55385
rect 74539 -55514 74585 -55385
rect 74637 -55485 74683 -55385
rect 74735 -55514 74781 -55385
rect 74441 -55560 75078 -55514
rect 74441 -55716 74487 -55560
rect 74539 -55562 74781 -55560
rect 74637 -55716 74683 -55562
rect 74833 -55716 74879 -55560
rect 72833 -56615 72879 -56315
rect 72480 -56810 72677 -56756
rect 72735 -57151 72781 -56852
rect 72734 -57188 72781 -57151
rect 72833 -57152 72879 -56852
rect 72931 -57188 72977 -56852
rect 73029 -57152 73075 -56315
rect 73442 -56470 73488 -56314
rect 73638 -56468 73684 -56314
rect 73540 -56470 73782 -56468
rect 73834 -56470 73880 -56314
rect 73442 -56516 74079 -56470
rect 73442 -56645 73488 -56545
rect 73540 -56645 73586 -56516
rect 73638 -56645 73684 -56545
rect 73736 -56645 73782 -56516
rect 74280 -56826 74326 -56226
rect 74491 -56826 74537 -56226
rect 74589 -56826 74635 -56226
rect 74687 -56826 74733 -56226
rect 74899 -56826 74945 -56226
rect 73127 -57188 73173 -56852
rect 75130 -56957 75235 -56885
rect 75136 -57040 75201 -56957
rect 74181 -57105 75201 -57040
rect 72734 -57235 73173 -57188
rect 74280 -57438 74326 -57138
rect 74378 -57438 74424 -57138
rect 74476 -57438 74522 -57138
rect 74718 -57438 74764 -57138
rect 74816 -57438 74862 -57138
rect 75049 -57546 75162 -57545
rect 75423 -57546 75536 -55350
rect 76272 -56584 76318 -56084
rect 76541 -56584 76587 -56084
rect 76639 -56584 76685 -56084
rect 76737 -56584 76783 -56084
rect 76867 -56584 76913 -56084
rect 77193 -56584 77239 -56084
rect 77421 -56384 77467 -56084
rect 76041 -56744 76179 -56740
rect 76847 -56744 76985 -56740
rect 77232 -56744 77286 -56671
rect 76041 -56788 77286 -56744
rect 76041 -56794 76179 -56788
rect 76847 -56794 76985 -56788
rect 77232 -56809 77286 -56788
rect 77404 -56824 77470 -56812
rect 78714 -56824 79021 -54678
rect 75880 -57131 75983 -57040
rect 74859 -57659 75536 -57546
rect 70633 -58311 72123 -58128
rect 73725 -58295 74164 -58248
rect 70633 -58365 73436 -58311
rect 73725 -58332 73772 -58295
rect 70633 -58428 72123 -58365
rect 72565 -58805 72695 -58655
rect 72851 -58709 72897 -58509
rect 72949 -58737 72995 -58509
rect 73047 -58709 73093 -58509
rect 73145 -58737 73191 -58509
rect 73382 -58655 73436 -58365
rect 73726 -58631 73772 -58332
rect 73824 -58631 73870 -58331
rect 73922 -58631 73968 -58295
rect 73382 -58709 73710 -58655
rect 72851 -58783 73488 -58737
rect 73656 -58764 73710 -58709
rect 72615 -60209 72669 -58805
rect 72851 -59039 72897 -58783
rect 72949 -58785 73191 -58783
rect 73047 -59039 73093 -58785
rect 73243 -59039 73289 -58783
rect 73630 -58822 73789 -58764
rect 73824 -59168 73870 -58868
rect 74020 -59168 74066 -58331
rect 74118 -58631 74164 -58295
rect 75049 -58690 75162 -57659
rect 75892 -57764 75971 -57131
rect 76174 -57380 76220 -57080
rect 76272 -57380 76318 -57080
rect 76644 -57380 76690 -56880
rect 76742 -57380 76788 -56880
rect 76867 -57380 76913 -56880
rect 76965 -57380 77011 -56880
rect 77095 -57380 77141 -56880
rect 77193 -57380 77239 -56880
rect 77291 -57380 77337 -56880
rect 77404 -56886 79026 -56824
rect 77404 -56895 77470 -56886
rect 77421 -57380 77467 -57080
rect 77519 -57380 77565 -57080
rect 75392 -57843 75971 -57764
rect 75392 -58198 75471 -57843
rect 75366 -58295 75482 -58198
rect 77393 -58326 77832 -58279
rect 75995 -58342 76092 -58336
rect 75995 -58396 77104 -58342
rect 77393 -58363 77440 -58326
rect 75995 -58402 76092 -58396
rect 74820 -58803 75528 -58690
rect 74433 -58938 74479 -58838
rect 74531 -58967 74577 -58838
rect 74629 -58938 74675 -58838
rect 74727 -58967 74773 -58838
rect 74433 -59013 75070 -58967
rect 74433 -59169 74479 -59013
rect 74531 -59015 74773 -59013
rect 74629 -59169 74675 -59015
rect 74825 -59169 74871 -59013
rect 72825 -60068 72871 -59768
rect 72472 -60263 72669 -60209
rect 70106 -60704 70367 -60400
rect 72727 -60604 72773 -60305
rect 72726 -60641 72773 -60604
rect 72825 -60605 72871 -60305
rect 72923 -60641 72969 -60305
rect 73021 -60605 73067 -59768
rect 73434 -59923 73480 -59767
rect 73630 -59921 73676 -59767
rect 73532 -59923 73774 -59921
rect 73826 -59923 73872 -59767
rect 73434 -59969 74071 -59923
rect 73434 -60098 73480 -59998
rect 73532 -60098 73578 -59969
rect 73630 -60098 73676 -59998
rect 73728 -60098 73774 -59969
rect 74272 -60279 74318 -59679
rect 74483 -60279 74529 -59679
rect 74581 -60279 74627 -59679
rect 74679 -60279 74725 -59679
rect 74891 -60279 74937 -59679
rect 73119 -60641 73165 -60305
rect 75122 -60410 75227 -60338
rect 75128 -60493 75193 -60410
rect 74173 -60558 75193 -60493
rect 72726 -60688 73165 -60641
rect 74272 -60891 74318 -60591
rect 74370 -60891 74416 -60591
rect 74468 -60891 74514 -60591
rect 74710 -60891 74756 -60591
rect 74808 -60891 74854 -60591
rect 75415 -60999 75528 -58803
rect 76233 -58836 76363 -58686
rect 76519 -58740 76565 -58540
rect 76617 -58768 76663 -58540
rect 76715 -58740 76761 -58540
rect 76813 -58768 76859 -58540
rect 77050 -58686 77104 -58396
rect 77394 -58662 77440 -58363
rect 77492 -58662 77538 -58362
rect 77590 -58662 77636 -58326
rect 77050 -58740 77378 -58686
rect 76519 -58814 77156 -58768
rect 77324 -58795 77378 -58740
rect 76283 -60240 76337 -58836
rect 76519 -59070 76565 -58814
rect 76617 -58816 76859 -58814
rect 76715 -59070 76761 -58816
rect 76911 -59070 76957 -58814
rect 77298 -58853 77457 -58795
rect 77492 -59199 77538 -58899
rect 77688 -59199 77734 -58362
rect 77786 -58662 77832 -58326
rect 78488 -58834 79196 -58721
rect 78101 -58969 78147 -58869
rect 78199 -58998 78245 -58869
rect 78297 -58969 78343 -58869
rect 78395 -58998 78441 -58869
rect 78101 -59044 78738 -58998
rect 78101 -59200 78147 -59044
rect 78199 -59046 78441 -59044
rect 78297 -59200 78343 -59046
rect 78493 -59200 78539 -59044
rect 76493 -60099 76539 -59799
rect 76140 -60294 76337 -60240
rect 76395 -60635 76441 -60336
rect 76394 -60672 76441 -60635
rect 76493 -60636 76539 -60336
rect 76591 -60672 76637 -60336
rect 76689 -60636 76735 -59799
rect 77102 -59954 77148 -59798
rect 77298 -59952 77344 -59798
rect 77200 -59954 77442 -59952
rect 77494 -59954 77540 -59798
rect 77102 -60000 77739 -59954
rect 77102 -60129 77148 -60029
rect 77200 -60129 77246 -60000
rect 77298 -60129 77344 -60029
rect 77396 -60129 77442 -60000
rect 77940 -60310 77986 -59710
rect 78151 -60310 78197 -59710
rect 78249 -60310 78295 -59710
rect 78347 -60310 78393 -59710
rect 78559 -60310 78605 -59710
rect 76787 -60672 76833 -60336
rect 78790 -60441 78895 -60369
rect 78796 -60524 78861 -60441
rect 77841 -60589 78861 -60524
rect 76394 -60719 76833 -60672
rect 77940 -60922 77986 -60622
rect 78038 -60922 78084 -60622
rect 78136 -60922 78182 -60622
rect 78378 -60922 78424 -60622
rect 78476 -60922 78522 -60622
rect 65698 -61129 70043 -61047
rect 74851 -61030 75528 -60999
rect 79083 -61030 79196 -58834
rect 79282 -60724 79593 -51080
rect 79858 -54596 88377 -54377
rect 79858 -58234 80077 -54596
rect 81311 -54820 81606 -54705
rect 83097 -54804 83536 -54757
rect 81311 -54874 82808 -54820
rect 83097 -54841 83144 -54804
rect 81311 -54978 81606 -54874
rect 81937 -55314 82067 -55164
rect 82223 -55218 82269 -55018
rect 82321 -55246 82367 -55018
rect 82419 -55218 82465 -55018
rect 82517 -55246 82563 -55018
rect 82754 -55164 82808 -54874
rect 83098 -55140 83144 -54841
rect 83196 -55140 83242 -54840
rect 83294 -55140 83340 -54804
rect 82754 -55218 83082 -55164
rect 82223 -55292 82860 -55246
rect 83028 -55273 83082 -55218
rect 81987 -56718 82041 -55314
rect 82223 -55548 82269 -55292
rect 82321 -55294 82563 -55292
rect 82419 -55548 82465 -55294
rect 82615 -55548 82661 -55292
rect 83002 -55331 83161 -55273
rect 83196 -55677 83242 -55377
rect 83392 -55677 83438 -54840
rect 83490 -55140 83536 -54804
rect 84192 -55312 84900 -55199
rect 83805 -55447 83851 -55347
rect 83903 -55476 83949 -55347
rect 84001 -55447 84047 -55347
rect 84099 -55476 84145 -55347
rect 83805 -55522 84442 -55476
rect 83805 -55678 83851 -55522
rect 83903 -55524 84145 -55522
rect 84001 -55678 84047 -55524
rect 84197 -55678 84243 -55522
rect 82197 -56577 82243 -56277
rect 81844 -56772 82041 -56718
rect 82099 -57113 82145 -56814
rect 82098 -57150 82145 -57113
rect 82197 -57114 82243 -56814
rect 82295 -57150 82341 -56814
rect 82393 -57114 82439 -56277
rect 82806 -56432 82852 -56276
rect 83002 -56430 83048 -56276
rect 82904 -56432 83146 -56430
rect 83198 -56432 83244 -56276
rect 82806 -56478 83443 -56432
rect 82806 -56607 82852 -56507
rect 82904 -56607 82950 -56478
rect 83002 -56607 83048 -56507
rect 83100 -56607 83146 -56478
rect 83644 -56788 83690 -56188
rect 83855 -56788 83901 -56188
rect 83953 -56788 83999 -56188
rect 84051 -56788 84097 -56188
rect 84263 -56788 84309 -56188
rect 82491 -57150 82537 -56814
rect 84494 -56919 84599 -56847
rect 84500 -57002 84565 -56919
rect 83545 -57067 84565 -57002
rect 82098 -57197 82537 -57150
rect 83644 -57400 83690 -57100
rect 83742 -57400 83788 -57100
rect 83840 -57400 83886 -57100
rect 84082 -57400 84128 -57100
rect 84180 -57400 84226 -57100
rect 84413 -57508 84526 -57507
rect 84787 -57508 84900 -55312
rect 85636 -56546 85682 -56046
rect 85905 -56546 85951 -56046
rect 86003 -56546 86049 -56046
rect 86101 -56546 86147 -56046
rect 86231 -56546 86277 -56046
rect 86557 -56546 86603 -56046
rect 86785 -56346 86831 -56046
rect 85405 -56706 85543 -56702
rect 86211 -56706 86349 -56702
rect 86596 -56706 86650 -56633
rect 85405 -56750 86650 -56706
rect 85405 -56756 85543 -56750
rect 86211 -56756 86349 -56750
rect 86596 -56771 86650 -56750
rect 86768 -56786 86834 -56774
rect 88158 -56786 88377 -54596
rect 85244 -57093 85347 -57002
rect 84223 -57621 84900 -57508
rect 79858 -58273 81637 -58234
rect 83089 -58257 83528 -58210
rect 79858 -58327 82800 -58273
rect 83089 -58294 83136 -58257
rect 79858 -58453 81637 -58327
rect 81929 -58767 82059 -58617
rect 82215 -58671 82261 -58471
rect 82313 -58699 82359 -58471
rect 82411 -58671 82457 -58471
rect 82509 -58699 82555 -58471
rect 82746 -58617 82800 -58327
rect 83090 -58593 83136 -58294
rect 83188 -58593 83234 -58293
rect 83286 -58593 83332 -58257
rect 82746 -58671 83074 -58617
rect 82215 -58745 82852 -58699
rect 83020 -58726 83074 -58671
rect 81979 -60171 82033 -58767
rect 82215 -59001 82261 -58745
rect 82313 -58747 82555 -58745
rect 82411 -59001 82457 -58747
rect 82607 -59001 82653 -58745
rect 82994 -58784 83153 -58726
rect 83188 -59130 83234 -58830
rect 83384 -59130 83430 -58293
rect 83482 -58593 83528 -58257
rect 84413 -58652 84526 -57621
rect 85256 -57726 85335 -57093
rect 85538 -57342 85584 -57042
rect 85636 -57342 85682 -57042
rect 86008 -57342 86054 -56842
rect 86106 -57342 86152 -56842
rect 86231 -57342 86277 -56842
rect 86329 -57342 86375 -56842
rect 86459 -57342 86505 -56842
rect 86557 -57342 86603 -56842
rect 86655 -57342 86701 -56842
rect 86768 -56848 88390 -56786
rect 86768 -56857 86834 -56848
rect 86785 -57342 86831 -57042
rect 86883 -57342 86929 -57042
rect 84756 -57805 85335 -57726
rect 84756 -58160 84835 -57805
rect 84730 -58257 84846 -58160
rect 86757 -58288 87196 -58241
rect 85359 -58304 85456 -58298
rect 85359 -58358 86468 -58304
rect 86757 -58325 86804 -58288
rect 85359 -58364 85456 -58358
rect 84184 -58765 84892 -58652
rect 83797 -58900 83843 -58800
rect 83895 -58929 83941 -58800
rect 83993 -58900 84039 -58800
rect 84091 -58929 84137 -58800
rect 83797 -58975 84434 -58929
rect 83797 -59131 83843 -58975
rect 83895 -58977 84137 -58975
rect 83993 -59131 84039 -58977
rect 84189 -59131 84235 -58975
rect 82189 -60030 82235 -59730
rect 81836 -60225 82033 -60171
rect 82091 -60566 82137 -60267
rect 82090 -60603 82137 -60566
rect 82189 -60567 82235 -60267
rect 82287 -60603 82333 -60267
rect 82385 -60567 82431 -59730
rect 82798 -59885 82844 -59729
rect 82994 -59883 83040 -59729
rect 82896 -59885 83138 -59883
rect 83190 -59885 83236 -59729
rect 82798 -59931 83435 -59885
rect 82798 -60060 82844 -59960
rect 82896 -60060 82942 -59931
rect 82994 -60060 83040 -59960
rect 83092 -60060 83138 -59931
rect 83636 -60241 83682 -59641
rect 83847 -60241 83893 -59641
rect 83945 -60241 83991 -59641
rect 84043 -60241 84089 -59641
rect 84255 -60241 84301 -59641
rect 82483 -60603 82529 -60267
rect 84486 -60372 84591 -60300
rect 84492 -60455 84557 -60372
rect 83537 -60520 84557 -60455
rect 82090 -60650 82529 -60603
rect 83636 -60853 83682 -60553
rect 83734 -60853 83780 -60553
rect 83832 -60853 83878 -60553
rect 84074 -60853 84120 -60553
rect 84172 -60853 84218 -60553
rect 84779 -60961 84892 -58765
rect 85597 -58798 85727 -58648
rect 85883 -58702 85929 -58502
rect 85981 -58730 86027 -58502
rect 86079 -58702 86125 -58502
rect 86177 -58730 86223 -58502
rect 86414 -58648 86468 -58358
rect 86758 -58624 86804 -58325
rect 86856 -58624 86902 -58324
rect 86954 -58624 87000 -58288
rect 86414 -58702 86742 -58648
rect 85883 -58776 86520 -58730
rect 86688 -58757 86742 -58702
rect 85647 -60202 85701 -58798
rect 85883 -59032 85929 -58776
rect 85981 -58778 86223 -58776
rect 86079 -59032 86125 -58778
rect 86275 -59032 86321 -58776
rect 86662 -58815 86821 -58757
rect 86856 -59161 86902 -58861
rect 87052 -59161 87098 -58324
rect 87150 -58624 87196 -58288
rect 87852 -58796 88560 -58683
rect 87465 -58931 87511 -58831
rect 87563 -58960 87609 -58831
rect 87661 -58931 87707 -58831
rect 87759 -58960 87805 -58831
rect 87465 -59006 88102 -58960
rect 87465 -59162 87511 -59006
rect 87563 -59008 87805 -59006
rect 87661 -59162 87707 -59008
rect 87857 -59162 87903 -59006
rect 85857 -60061 85903 -59761
rect 85504 -60256 85701 -60202
rect 85759 -60597 85805 -60298
rect 85758 -60634 85805 -60597
rect 85857 -60598 85903 -60298
rect 85955 -60634 86001 -60298
rect 86053 -60598 86099 -59761
rect 86466 -59916 86512 -59760
rect 86662 -59914 86708 -59760
rect 86564 -59916 86806 -59914
rect 86858 -59916 86904 -59760
rect 86466 -59962 87103 -59916
rect 86466 -60091 86512 -59991
rect 86564 -60091 86610 -59962
rect 86662 -60091 86708 -59991
rect 86760 -60091 86806 -59962
rect 87304 -60272 87350 -59672
rect 87515 -60272 87561 -59672
rect 87613 -60272 87659 -59672
rect 87711 -60272 87757 -59672
rect 87923 -60272 87969 -59672
rect 86151 -60634 86197 -60298
rect 88154 -60403 88259 -60331
rect 88160 -60486 88225 -60403
rect 87205 -60551 88225 -60486
rect 85758 -60681 86197 -60634
rect 87304 -60884 87350 -60584
rect 87402 -60884 87448 -60584
rect 87500 -60884 87546 -60584
rect 87742 -60884 87788 -60584
rect 87840 -60884 87886 -60584
rect 74851 -61112 79196 -61030
rect 84215 -60992 84892 -60961
rect 88447 -60992 88560 -58796
rect 88813 -60356 89097 -50147
rect 88783 -60699 89142 -60356
rect 84215 -61074 88560 -60992
rect 84219 -61105 88560 -61074
rect 65702 -61160 70043 -61129
rect 74855 -61143 79196 -61112
rect 56948 -61226 61289 -61195
rect 47750 -61260 52091 -61229
rect 42978 -61834 43295 -61751
rect 27278 -62015 36078 -61834
rect 42978 -62015 82728 -61834
rect 42978 -62042 43295 -62015
rect 42935 -62934 43304 -62557
rect 44255 -62855 82728 -62570
rect 42944 -64722 43244 -62934
rect 25466 -65022 43244 -64722
rect 44255 -65265 44540 -62855
rect 25261 -65324 44540 -65265
rect 24998 -65445 44540 -65324
rect 25261 -65550 44540 -65445
<< metal2 >>
rect 16949 11350 17282 16839
<< obsm2 >>
rect -157 10922 87 12457
rect 93931 12460 95152 38495
rect 1499 1854 1718 1933
rect 1635 931 1718 1854
<< metal3 >>
rect 18260 83864 23340 89236
rect 23580 83864 28660 89236
rect 28900 83864 33980 89236
rect 34220 83864 39300 89236
rect 39540 83864 44620 89236
rect 44860 83864 49940 89236
rect 50180 83864 55260 89236
rect 55500 83864 60580 89236
rect 60820 83864 65900 89236
rect 66140 83864 71220 89236
rect 71460 83864 76540 89236
rect 76780 83864 81860 89236
rect 82100 83864 87180 89236
rect 87420 83864 92500 89236
rect 18260 78252 23340 83624
rect 23580 78252 28660 83624
rect 28900 78252 33980 83624
rect 34220 78252 39300 83624
rect 39540 78252 44620 83624
rect 44860 78252 49940 83624
rect 50180 78252 55260 83624
rect 55500 78252 60580 83624
rect 60820 78252 65900 83624
rect 66140 78252 71220 83624
rect 71460 78252 76540 83624
rect 76780 78252 81860 83624
rect 82100 78252 87180 83624
rect 87420 78252 92500 83624
rect 18260 72640 23340 78012
rect 23580 72640 28660 78012
rect 28900 72640 33980 78012
rect 34220 72640 39300 78012
rect 39540 72640 44620 78012
rect 44860 72640 49940 78012
rect 50180 72640 55260 78012
rect 55500 72640 60580 78012
rect 60820 72640 65900 78012
rect 66140 72640 71220 78012
rect 71460 72640 76540 78012
rect 76780 72640 81860 78012
rect 82100 72640 87180 78012
rect 87420 72640 92500 78012
rect 18260 67028 23340 72400
rect 23580 67028 28660 72400
rect 28900 67028 33980 72400
rect 34220 67028 39300 72400
rect 39540 67028 44620 72400
rect 44860 67028 49940 72400
rect 50180 67028 55260 72400
rect 55500 67028 60580 72400
rect 60820 67028 65900 72400
rect 66140 67028 71220 72400
rect 71460 67028 76540 72400
rect 76780 67028 81860 72400
rect 82100 67028 87180 72400
rect 87420 67028 92500 72400
rect 18260 61416 23340 66788
rect 23580 61416 28660 66788
rect 28900 61416 33980 66788
rect 34220 61416 39300 66788
rect 39540 61416 44620 66788
rect 44860 61416 49940 66788
rect 50180 61416 55260 66788
rect 55500 61416 60580 66788
rect 60820 61416 65900 66788
rect 66140 61416 71220 66788
rect 71460 61416 76540 66788
rect 76780 61416 81860 66788
rect 82100 61416 87180 66788
rect 87420 61416 92500 66788
rect 18260 55804 23340 61176
rect 23580 55804 28660 61176
rect 28900 55804 33980 61176
rect 34220 55804 39300 61176
rect 39540 55804 44620 61176
rect 44860 55804 49940 61176
rect 50180 55804 55260 61176
rect 55500 55804 60580 61176
rect 60820 55804 65900 61176
rect 66140 55804 71220 61176
rect 71460 55804 76540 61176
rect 76780 55804 81860 61176
rect 82100 55804 87180 61176
rect 87420 55804 92500 61176
rect 18260 50192 23340 55564
rect 23580 50192 28660 55564
rect 28900 50192 33980 55564
rect 34220 50192 39300 55564
rect 39540 50192 44620 55564
rect 44860 50192 49940 55564
rect 50180 50192 55260 55564
rect 55500 50192 60580 55564
rect 60820 50192 65900 55564
rect 66140 50192 71220 55564
rect 71460 50192 76540 55564
rect 76780 50192 81860 55564
rect 82100 50192 87180 55564
rect 87420 50192 92500 55564
rect 18260 44580 23340 49952
rect 23580 44580 28660 49952
rect 28900 44580 33980 49952
rect 34220 44580 39300 49952
rect 39540 44580 44620 49952
rect 44860 44580 49940 49952
rect 50180 44580 55260 49952
rect 55500 44580 60580 49952
rect 60820 44580 65900 49952
rect 66140 44580 71220 49952
rect 71460 44580 76540 49952
rect 76780 44580 81860 49952
rect 82100 44580 87180 49952
rect 87420 44580 92500 49952
rect 18260 38968 23340 44340
rect 23580 38968 28660 44340
rect 28900 38968 33980 44340
rect 34220 38968 39300 44340
rect 39540 38968 44620 44340
rect 44860 38968 49940 44340
rect 50180 38968 55260 44340
rect 55500 38968 60580 44340
rect 60820 38968 65900 44340
rect 66140 38968 71220 44340
rect 71460 38968 76540 44340
rect 76780 38968 81860 44340
rect 82100 38968 87180 44340
rect 87420 38968 92500 44340
rect 18260 33356 23340 38728
rect 23580 33356 28660 38728
rect 28900 33356 33980 38728
rect 34220 33356 39300 38728
rect 39540 33356 44620 38728
rect 44860 33356 49940 38728
rect 50180 33356 55260 38728
rect 55500 33356 60580 38728
rect 60820 33356 65900 38728
rect 66140 33356 71220 38728
rect 71460 33356 76540 38728
rect 76780 33356 81860 38728
rect 82100 33356 87180 38728
rect 87420 33356 92500 38728
rect 317 26487 2397 28859
rect 2637 26487 4717 28859
rect 4957 26487 7037 28859
rect 7277 26487 9357 28859
rect 9597 26487 11677 28859
rect 11917 26487 13997 28859
rect 14237 26487 16317 28859
rect 18260 27744 23340 33116
rect 23580 27744 28660 33116
rect 28900 27744 33980 33116
rect 34220 27744 39300 33116
rect 39540 27744 44620 33116
rect 44860 27744 49940 33116
rect 50180 27744 55260 33116
rect 55500 27744 60580 33116
rect 60820 27744 65900 33116
rect 66140 27744 71220 33116
rect 71460 27744 76540 33116
rect 76780 27744 81860 33116
rect 82100 27744 87180 33116
rect 87420 27744 92500 33116
rect 317 23875 2397 26247
rect 2637 23875 4717 26247
rect 4957 23875 7037 26247
rect 7277 23875 9357 26247
rect 9597 23875 11677 26247
rect 11917 23875 13997 26247
rect 14237 23875 16317 26247
rect 317 21263 2397 23635
rect 2637 21263 4717 23635
rect 4957 21263 7037 23635
rect 7277 21263 9357 23635
rect 9597 21263 11677 23635
rect 11917 21263 13997 23635
rect 14237 21263 16317 23635
rect 18260 22132 23340 27504
rect 23580 22132 28660 27504
rect 28900 22132 33980 27504
rect 34220 22132 39300 27504
rect 39540 22132 44620 27504
rect 44860 22132 49940 27504
rect 50180 22132 55260 27504
rect 55500 22132 60580 27504
rect 60820 22132 65900 27504
rect 66140 22132 71220 27504
rect 71460 22132 76540 27504
rect 76780 22132 81860 27504
rect 82100 22132 87180 27504
rect 87420 22132 92500 27504
rect 317 18651 2397 21023
rect 2637 18651 4717 21023
rect 4957 18651 7037 21023
rect 7277 18651 9357 21023
rect 9597 18651 11677 21023
rect 11917 18651 13997 21023
rect 14237 18651 16317 21023
rect 317 16039 2397 18411
rect 2637 16039 4717 18411
rect 4957 16039 7037 18411
rect 7277 16039 9357 18411
rect 9597 16039 11677 18411
rect 11917 16039 13997 18411
rect 14237 16039 16317 18411
rect 317 13427 2397 15799
rect 2637 13427 4717 15799
rect 4957 13427 7037 15799
rect 7277 13427 9357 15799
rect 9597 13427 11677 15799
rect 11917 13427 13997 15799
rect 14237 13427 16317 15799
rect 317 10815 2397 13187
rect 2637 10815 4717 13187
rect 4957 10815 7037 13187
rect 7277 10815 9357 13187
rect 9597 10815 11677 13187
rect 11917 10815 13997 13187
rect 14237 10815 16317 13187
rect 16949 11350 17282 16839
rect 18260 16520 23340 21892
rect 23580 16520 28660 21892
rect 28900 16520 33980 21892
rect 34220 16520 39300 21892
rect 39540 16520 44620 21892
rect 44860 16520 49940 21892
rect 50180 16520 55260 21892
rect 55500 16520 60580 21892
rect 60820 16520 65900 21892
rect 66140 16520 71220 21892
rect 71460 16520 76540 21892
rect 76780 16520 81860 21892
rect 82100 16520 87180 21892
rect 87420 16520 92500 21892
rect 18260 10908 23340 16280
rect 23580 10908 28660 16280
rect 28900 10908 33980 16280
rect 34220 10908 39300 16280
rect 39540 10908 44620 16280
rect 44860 10908 49940 16280
rect 50180 10908 55260 16280
rect 55500 10908 60580 16280
rect 60820 10908 65900 16280
rect 66140 10908 71220 16280
rect 71460 10908 76540 16280
rect 76780 10908 81860 16280
rect 82100 10908 87180 16280
rect 87420 10908 92500 16280
<< obsm3 >>
rect -157 10922 87 12457
rect 93931 12460 95152 38495
<< metal4 >>
rect 17174 89236 18030 89308
rect 17174 89132 92620 89236
rect 17174 83624 18030 89132
rect 17174 83520 92620 83624
rect 17174 78012 18030 83520
rect 17174 77908 92620 78012
rect 17174 72400 18030 77908
rect 17174 72296 92620 72400
rect 17174 66788 18030 72296
rect 17174 66684 92620 66788
rect 17174 61176 18030 66684
rect 17174 61072 92620 61176
rect 17174 55564 18030 61072
rect 17174 55460 92620 55564
rect 17174 49952 18030 55460
rect 17174 49848 92620 49952
rect 17174 44340 18030 49848
rect 17174 44236 92620 44340
rect 17174 38728 18030 44236
rect 17174 38624 92620 38728
rect 17174 33116 18030 38624
rect 17174 33012 92620 33116
rect 17174 28859 18030 33012
rect 197 28755 18030 28859
rect 16812 27504 18030 28755
rect 16812 27400 92620 27504
rect 16812 26247 18030 27400
rect 197 26143 18030 26247
rect 16812 23635 18030 26143
rect 197 23531 18030 23635
rect 16812 21892 18030 23531
rect 16812 21788 92620 21892
rect 16812 21023 18030 21788
rect 197 20919 18030 21023
rect 16812 18411 18030 20919
rect 197 18307 18030 18411
rect 16812 16280 18030 18307
rect 16812 16176 92620 16280
rect 16812 15799 18030 16176
rect 197 15695 18030 15799
rect 16812 13187 18030 15695
rect 197 13083 18030 13187
rect 16812 11509 18030 13083
rect 16812 11245 17392 11509
<< obsm4 >>
rect 18339 86456 23261 88865
rect 23659 86456 28581 88865
rect 28979 86456 33901 88865
rect 34299 86456 39221 88865
rect 39619 86456 44541 88865
rect 44939 86456 49861 88865
rect 50259 86456 55181 88865
rect 55579 86456 60501 88865
rect 60899 86456 65821 88865
rect 66219 86456 71141 88865
rect 71539 86456 76461 88865
rect 76859 86456 81781 88865
rect 82179 86456 87101 88865
rect 87499 86456 92421 88865
rect 93577 86456 95600 89068
rect 18140 86352 95600 86456
rect 18339 83943 23261 86352
rect 23659 83943 28581 86352
rect 28979 83943 33901 86352
rect 34299 83943 39221 86352
rect 39619 83943 44541 86352
rect 44939 83943 49861 86352
rect 50259 83943 55181 86352
rect 55579 83943 60501 86352
rect 60899 83943 65821 86352
rect 66219 83943 71141 86352
rect 71539 83943 76461 86352
rect 76859 83943 81781 86352
rect 82179 83943 87101 86352
rect 87499 83943 92421 86352
rect 18339 80844 23261 83253
rect 23659 80844 28581 83253
rect 28979 80844 33901 83253
rect 34299 80844 39221 83253
rect 39619 80844 44541 83253
rect 44939 80844 49861 83253
rect 50259 80844 55181 83253
rect 55579 80844 60501 83253
rect 60899 80844 65821 83253
rect 66219 80844 71141 83253
rect 71539 80844 76461 83253
rect 76859 80844 81781 83253
rect 82179 80844 87101 83253
rect 87499 80844 92421 83253
rect 93577 80844 95600 86352
rect 18140 80740 95600 80844
rect 18339 78331 23261 80740
rect 23659 78331 28581 80740
rect 28979 78331 33901 80740
rect 34299 78331 39221 80740
rect 39619 78331 44541 80740
rect 44939 78331 49861 80740
rect 50259 78331 55181 80740
rect 55579 78331 60501 80740
rect 60899 78331 65821 80740
rect 66219 78331 71141 80740
rect 71539 78331 76461 80740
rect 76859 78331 81781 80740
rect 82179 78331 87101 80740
rect 87499 78331 92421 80740
rect 18339 75232 23261 77641
rect 23659 75232 28581 77641
rect 28979 75232 33901 77641
rect 34299 75232 39221 77641
rect 39619 75232 44541 77641
rect 44939 75232 49861 77641
rect 50259 75232 55181 77641
rect 55579 75232 60501 77641
rect 60899 75232 65821 77641
rect 66219 75232 71141 77641
rect 71539 75232 76461 77641
rect 76859 75232 81781 77641
rect 82179 75232 87101 77641
rect 87499 75232 92421 77641
rect 93577 75232 95600 80740
rect 18140 75128 95600 75232
rect 18339 72719 23261 75128
rect 23659 72719 28581 75128
rect 28979 72719 33901 75128
rect 34299 72719 39221 75128
rect 39619 72719 44541 75128
rect 44939 72719 49861 75128
rect 50259 72719 55181 75128
rect 55579 72719 60501 75128
rect 60899 72719 65821 75128
rect 66219 72719 71141 75128
rect 71539 72719 76461 75128
rect 76859 72719 81781 75128
rect 82179 72719 87101 75128
rect 87499 72719 92421 75128
rect 18339 69620 23261 72029
rect 23659 69620 28581 72029
rect 28979 69620 33901 72029
rect 34299 69620 39221 72029
rect 39619 69620 44541 72029
rect 44939 69620 49861 72029
rect 50259 69620 55181 72029
rect 55579 69620 60501 72029
rect 60899 69620 65821 72029
rect 66219 69620 71141 72029
rect 71539 69620 76461 72029
rect 76859 69620 81781 72029
rect 82179 69620 87101 72029
rect 87499 69620 92421 72029
rect 93577 69620 95600 75128
rect 18140 69516 95600 69620
rect 18339 67107 23261 69516
rect 23659 67107 28581 69516
rect 28979 67107 33901 69516
rect 34299 67107 39221 69516
rect 39619 67107 44541 69516
rect 44939 67107 49861 69516
rect 50259 67107 55181 69516
rect 55579 67107 60501 69516
rect 60899 67107 65821 69516
rect 66219 67107 71141 69516
rect 71539 67107 76461 69516
rect 76859 67107 81781 69516
rect 82179 67107 87101 69516
rect 87499 67107 92421 69516
rect 18339 64008 23261 66417
rect 23659 64008 28581 66417
rect 28979 64008 33901 66417
rect 34299 64008 39221 66417
rect 39619 64008 44541 66417
rect 44939 64008 49861 66417
rect 50259 64008 55181 66417
rect 55579 64008 60501 66417
rect 60899 64008 65821 66417
rect 66219 64008 71141 66417
rect 71539 64008 76461 66417
rect 76859 64008 81781 66417
rect 82179 64008 87101 66417
rect 87499 64008 92421 66417
rect 93577 64008 95600 69516
rect 18140 63904 95600 64008
rect 18339 61495 23261 63904
rect 23659 61495 28581 63904
rect 28979 61495 33901 63904
rect 34299 61495 39221 63904
rect 39619 61495 44541 63904
rect 44939 61495 49861 63904
rect 50259 61495 55181 63904
rect 55579 61495 60501 63904
rect 60899 61495 65821 63904
rect 66219 61495 71141 63904
rect 71539 61495 76461 63904
rect 76859 61495 81781 63904
rect 82179 61495 87101 63904
rect 87499 61495 92421 63904
rect 18339 58396 23261 60805
rect 23659 58396 28581 60805
rect 28979 58396 33901 60805
rect 34299 58396 39221 60805
rect 39619 58396 44541 60805
rect 44939 58396 49861 60805
rect 50259 58396 55181 60805
rect 55579 58396 60501 60805
rect 60899 58396 65821 60805
rect 66219 58396 71141 60805
rect 71539 58396 76461 60805
rect 76859 58396 81781 60805
rect 82179 58396 87101 60805
rect 87499 58396 92421 60805
rect 93577 58396 95600 63904
rect 18140 58292 95600 58396
rect 18339 55883 23261 58292
rect 23659 55883 28581 58292
rect 28979 55883 33901 58292
rect 34299 55883 39221 58292
rect 39619 55883 44541 58292
rect 44939 55883 49861 58292
rect 50259 55883 55181 58292
rect 55579 55883 60501 58292
rect 60899 55883 65821 58292
rect 66219 55883 71141 58292
rect 71539 55883 76461 58292
rect 76859 55883 81781 58292
rect 82179 55883 87101 58292
rect 87499 55883 92421 58292
rect 18339 52784 23261 55193
rect 23659 52784 28581 55193
rect 28979 52784 33901 55193
rect 34299 52784 39221 55193
rect 39619 52784 44541 55193
rect 44939 52784 49861 55193
rect 50259 52784 55181 55193
rect 55579 52784 60501 55193
rect 60899 52784 65821 55193
rect 66219 52784 71141 55193
rect 71539 52784 76461 55193
rect 76859 52784 81781 55193
rect 82179 52784 87101 55193
rect 87499 52784 92421 55193
rect 93577 52784 95600 58292
rect 18140 52680 95600 52784
rect 18339 50271 23261 52680
rect 23659 50271 28581 52680
rect 28979 50271 33901 52680
rect 34299 50271 39221 52680
rect 39619 50271 44541 52680
rect 44939 50271 49861 52680
rect 50259 50271 55181 52680
rect 55579 50271 60501 52680
rect 60899 50271 65821 52680
rect 66219 50271 71141 52680
rect 71539 50271 76461 52680
rect 76859 50271 81781 52680
rect 82179 50271 87101 52680
rect 87499 50271 92421 52680
rect 18339 47172 23261 49581
rect 23659 47172 28581 49581
rect 28979 47172 33901 49581
rect 34299 47172 39221 49581
rect 39619 47172 44541 49581
rect 44939 47172 49861 49581
rect 50259 47172 55181 49581
rect 55579 47172 60501 49581
rect 60899 47172 65821 49581
rect 66219 47172 71141 49581
rect 71539 47172 76461 49581
rect 76859 47172 81781 49581
rect 82179 47172 87101 49581
rect 87499 47172 92421 49581
rect 93577 47172 95600 52680
rect 18140 47068 95600 47172
rect 18339 44659 23261 47068
rect 23659 44659 28581 47068
rect 28979 44659 33901 47068
rect 34299 44659 39221 47068
rect 39619 44659 44541 47068
rect 44939 44659 49861 47068
rect 50259 44659 55181 47068
rect 55579 44659 60501 47068
rect 60899 44659 65821 47068
rect 66219 44659 71141 47068
rect 71539 44659 76461 47068
rect 76859 44659 81781 47068
rect 82179 44659 87101 47068
rect 87499 44659 92421 47068
rect 18339 41560 23261 43969
rect 23659 41560 28581 43969
rect 28979 41560 33901 43969
rect 34299 41560 39221 43969
rect 39619 41560 44541 43969
rect 44939 41560 49861 43969
rect 50259 41560 55181 43969
rect 55579 41560 60501 43969
rect 60899 41560 65821 43969
rect 66219 41560 71141 43969
rect 71539 41560 76461 43969
rect 76859 41560 81781 43969
rect 82179 41560 87101 43969
rect 87499 41560 92421 43969
rect 93577 41560 95600 47068
rect 18140 41456 95600 41560
rect 18339 39047 23261 41456
rect 23659 39047 28581 41456
rect 28979 39047 33901 41456
rect 34299 39047 39221 41456
rect 39619 39047 44541 41456
rect 44939 39047 49861 41456
rect 50259 39047 55181 41456
rect 55579 39047 60501 41456
rect 60899 39047 65821 41456
rect 66219 39047 71141 41456
rect 71539 39047 76461 41456
rect 76859 39047 81781 41456
rect 82179 39047 87101 41456
rect 87499 39047 92421 41456
rect 18339 35948 23261 38357
rect 23659 35948 28581 38357
rect 28979 35948 33901 38357
rect 34299 35948 39221 38357
rect 39619 35948 44541 38357
rect 44939 35948 49861 38357
rect 50259 35948 55181 38357
rect 55579 35948 60501 38357
rect 60899 35948 65821 38357
rect 66219 35948 71141 38357
rect 71539 35948 76461 38357
rect 76859 35948 81781 38357
rect 82179 35948 87101 38357
rect 87499 35948 92421 38357
rect 93577 35948 95600 41456
rect 18140 35844 95600 35948
rect 18339 33435 23261 35844
rect 23659 33435 28581 35844
rect 28979 33435 33901 35844
rect 34299 33435 39221 35844
rect 39619 33435 44541 35844
rect 44939 33435 49861 35844
rect 50259 33435 55181 35844
rect 55579 33435 60501 35844
rect 60899 33435 65821 35844
rect 66219 33435 71141 35844
rect 71539 33435 76461 35844
rect 76859 33435 81781 35844
rect 82179 33435 87101 35844
rect 87499 33435 92421 35844
rect -194 27579 97 28914
rect 18339 30336 23261 32745
rect 23659 30336 28581 32745
rect 28979 30336 33901 32745
rect 34299 30336 39221 32745
rect 39619 30336 44541 32745
rect 44939 30336 49861 32745
rect 50259 30336 55181 32745
rect 55579 30336 60501 32745
rect 60899 30336 65821 32745
rect 66219 30336 71141 32745
rect 71539 30336 76461 32745
rect 76859 30336 81781 32745
rect 82179 30336 87101 32745
rect 87499 30336 92421 32745
rect 93577 30336 95600 35844
rect 18140 30232 95600 30336
rect 396 27579 2318 28488
rect 2716 27579 4638 28488
rect 5036 27579 6958 28488
rect 7356 27579 9278 28488
rect 9676 27579 11598 28488
rect 11996 27579 13918 28488
rect 14316 27579 16238 28488
rect -194 27475 16437 27579
rect 18339 27823 23261 30232
rect 23659 27823 28581 30232
rect 28979 27823 33901 30232
rect 34299 27823 39221 30232
rect 39619 27823 44541 30232
rect 44939 27823 49861 30232
rect 50259 27823 55181 30232
rect 55579 27823 60501 30232
rect 60899 27823 65821 30232
rect 66219 27823 71141 30232
rect 71539 27823 76461 30232
rect 76859 27823 81781 30232
rect 82179 27823 87101 30232
rect 87499 27823 92421 30232
rect -194 24967 97 27475
rect 396 26566 2318 27475
rect 2716 26566 4638 27475
rect 5036 26566 6958 27475
rect 7356 26566 9278 27475
rect 9676 26566 11598 27475
rect 11996 26566 13918 27475
rect 14316 26566 16238 27475
rect 396 24967 2318 25876
rect 2716 24967 4638 25876
rect 5036 24967 6958 25876
rect 7356 24967 9278 25876
rect 9676 24967 11598 25876
rect 11996 24967 13918 25876
rect 14316 24967 16238 25876
rect -194 24863 16437 24967
rect -194 22355 97 24863
rect 396 23954 2318 24863
rect 2716 23954 4638 24863
rect 5036 23954 6958 24863
rect 7356 23954 9278 24863
rect 9676 23954 11598 24863
rect 11996 23954 13918 24863
rect 14316 23954 16238 24863
rect 18339 24724 23261 27133
rect 23659 24724 28581 27133
rect 28979 24724 33901 27133
rect 34299 24724 39221 27133
rect 39619 24724 44541 27133
rect 44939 24724 49861 27133
rect 50259 24724 55181 27133
rect 55579 24724 60501 27133
rect 60899 24724 65821 27133
rect 66219 24724 71141 27133
rect 71539 24724 76461 27133
rect 76859 24724 81781 27133
rect 82179 24724 87101 27133
rect 87499 24724 92421 27133
rect 93577 24724 95600 30232
rect 18140 24620 95600 24724
rect 396 22355 2318 23264
rect 2716 22355 4638 23264
rect 5036 22355 6958 23264
rect 7356 22355 9278 23264
rect 9676 22355 11598 23264
rect 11996 22355 13918 23264
rect 14316 22355 16238 23264
rect -194 22251 16437 22355
rect -194 19743 97 22251
rect 396 21342 2318 22251
rect 2716 21342 4638 22251
rect 5036 21342 6958 22251
rect 7356 21342 9278 22251
rect 9676 21342 11598 22251
rect 11996 21342 13918 22251
rect 14316 21342 16238 22251
rect 18339 22211 23261 24620
rect 23659 22211 28581 24620
rect 28979 22211 33901 24620
rect 34299 22211 39221 24620
rect 39619 22211 44541 24620
rect 44939 22211 49861 24620
rect 50259 22211 55181 24620
rect 55579 22211 60501 24620
rect 60899 22211 65821 24620
rect 66219 22211 71141 24620
rect 71539 22211 76461 24620
rect 76859 22211 81781 24620
rect 82179 22211 87101 24620
rect 87499 22211 92421 24620
rect 396 19743 2318 20652
rect 2716 19743 4638 20652
rect 5036 19743 6958 20652
rect 7356 19743 9278 20652
rect 9676 19743 11598 20652
rect 11996 19743 13918 20652
rect 14316 19743 16238 20652
rect -194 19639 16437 19743
rect -194 17131 97 19639
rect 396 18730 2318 19639
rect 2716 18730 4638 19639
rect 5036 18730 6958 19639
rect 7356 18730 9278 19639
rect 9676 18730 11598 19639
rect 11996 18730 13918 19639
rect 14316 18730 16238 19639
rect 18339 19112 23261 21521
rect 23659 19112 28581 21521
rect 28979 19112 33901 21521
rect 34299 19112 39221 21521
rect 39619 19112 44541 21521
rect 44939 19112 49861 21521
rect 50259 19112 55181 21521
rect 55579 19112 60501 21521
rect 60899 19112 65821 21521
rect 66219 19112 71141 21521
rect 71539 19112 76461 21521
rect 76859 19112 81781 21521
rect 82179 19112 87101 21521
rect 87499 19112 92421 21521
rect 93577 19112 95600 24620
rect 18140 19008 95600 19112
rect 396 17131 2318 18040
rect 2716 17131 4638 18040
rect 5036 17131 6958 18040
rect 7356 17131 9278 18040
rect 9676 17131 11598 18040
rect 11996 17131 13918 18040
rect 14316 17131 16238 18040
rect -194 17027 16437 17131
rect -194 14519 97 17027
rect 396 16118 2318 17027
rect 2716 16118 4638 17027
rect 5036 16118 6958 17027
rect 7356 16118 9278 17027
rect 9676 16118 11598 17027
rect 11996 16118 13918 17027
rect 14316 16118 16238 17027
rect 18339 16599 23261 19008
rect 23659 16599 28581 19008
rect 28979 16599 33901 19008
rect 34299 16599 39221 19008
rect 39619 16599 44541 19008
rect 44939 16599 49861 19008
rect 50259 16599 55181 19008
rect 55579 16599 60501 19008
rect 60899 16599 65821 19008
rect 66219 16599 71141 19008
rect 71539 16599 76461 19008
rect 76859 16599 81781 19008
rect 82179 16599 87101 19008
rect 87499 16599 92421 19008
rect 396 14519 2318 15428
rect 2716 14519 4638 15428
rect 5036 14519 6958 15428
rect 7356 14519 9278 15428
rect 9676 14519 11598 15428
rect 11996 14519 13918 15428
rect 14316 14519 16238 15428
rect -194 14415 16437 14519
rect -194 11907 97 14415
rect 396 13506 2318 14415
rect 2716 13506 4638 14415
rect 5036 13506 6958 14415
rect 7356 13506 9278 14415
rect 9676 13506 11598 14415
rect 11996 13506 13918 14415
rect 14316 13506 16238 14415
rect 18339 13500 23261 15909
rect 23659 13500 28581 15909
rect 28979 13500 33901 15909
rect 34299 13500 39221 15909
rect 39619 13500 44541 15909
rect 44939 13500 49861 15909
rect 50259 13500 55181 15909
rect 55579 13500 60501 15909
rect 60899 13500 65821 15909
rect 66219 13500 71141 15909
rect 71539 13500 76461 15909
rect 76859 13500 81781 15909
rect 82179 13500 87101 15909
rect 87499 13500 92421 15909
rect 93577 13500 95600 19008
rect 18140 13396 95600 13500
rect 396 11907 2318 12816
rect 2716 11907 4638 12816
rect 5036 11907 6958 12816
rect 7356 11907 9278 12816
rect 9676 11907 11598 12816
rect 11996 11907 13918 12816
rect 14316 11907 16238 12816
rect -194 11803 16437 11907
rect -194 10865 97 11803
rect 396 10894 2318 11803
rect 2716 10894 4638 11803
rect 5036 10894 6958 11803
rect 7356 10894 9278 11803
rect 9676 10894 11598 11803
rect 11996 10894 13918 11803
rect 14316 10894 16238 11803
rect 18339 10987 23261 13396
rect 23659 10987 28581 13396
rect 28979 10987 33901 13396
rect 34299 10987 39221 13396
rect 39619 10987 44541 13396
rect 44939 10987 49861 13396
rect 50259 10987 55181 13396
rect 55579 10987 60501 13396
rect 60899 10987 65821 13396
rect 66219 10987 71141 13396
rect 71539 10987 76461 13396
rect 76859 10987 81781 13396
rect 82179 10987 87101 13396
rect 87499 10987 92421 13396
rect 93577 10777 95600 13396
<< labels >>
rlabel locali s -4314 -1342 -4146 -1334 2 S6
port 1 nsew
rlabel locali s -5167 -1334 -4146 -1282 2 S6
port 1 nsew
rlabel locali s -4314 -1282 -4146 -1268 2 S6
port 1 nsew
rlabel locali s -5167 -1282 -5115 -677 2 S6
port 1 nsew
rlabel locali s -22114 -677 -4996 -603 2 S6
port 1 nsew
rlabel metal1 s 3985 76 4186 265 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6789 938 6835 1138 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6593 938 6639 1138 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6397 938 6443 1138 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6201 938 6247 1138 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6005 938 6051 1138 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6789 1284 6835 1484 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6593 1284 6639 1484 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6397 1284 6443 1484 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6201 1284 6247 1484 6 UP_INPUT
port 2 nsew
rlabel metal1 s 6005 1284 6051 1454 6 UP_INPUT
port 2 nsew
rlabel metal1 s 4064 265 4108 1310 6 UP_INPUT
port 2 nsew
rlabel metal1 s 4064 1310 5294 1354 6 UP_INPUT
port 2 nsew
rlabel metal1 s 5250 1354 5294 1454 6 UP_INPUT
port 2 nsew
rlabel metal1 s 5250 1454 6052 1498 6 UP_INPUT
port 2 nsew
rlabel locali s -26391 -2075 -1693 -1962 2 UP_INPUT
port 2 nsew
rlabel locali s 3985 76 4186 100 6 UP_INPUT
port 2 nsew
rlabel locali s -1806 -1962 -1693 100 2 UP_INPUT
port 2 nsew
rlabel locali s -1806 100 4186 213 6 UP_INPUT
port 2 nsew
rlabel locali s 3985 213 4186 265 6 UP_INPUT
port 2 nsew
rlabel locali s 6795 934 6829 1191 6 UP_INPUT
port 2 nsew
rlabel locali s 6599 934 6633 1191 6 UP_INPUT
port 2 nsew
rlabel locali s 6403 934 6437 1191 6 UP_INPUT
port 2 nsew
rlabel locali s 6207 934 6241 1191 6 UP_INPUT
port 2 nsew
rlabel locali s 6011 934 6045 1191 6 UP_INPUT
port 2 nsew
rlabel locali s 6011 1191 6829 1225 6 UP_INPUT
port 2 nsew
rlabel locali s 6795 1225 6829 1488 6 UP_INPUT
port 2 nsew
rlabel locali s 6599 1225 6633 1488 6 UP_INPUT
port 2 nsew
rlabel locali s 6403 1225 6437 1488 6 UP_INPUT
port 2 nsew
rlabel locali s 6207 1225 6241 1488 6 UP_INPUT
port 2 nsew
rlabel locali s 6011 1225 6045 1488 6 UP_INPUT
port 2 nsew
rlabel metal1 s 4310 -2309 4465 -2171 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6804 -1752 6850 -1552 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6608 -1752 6654 -1552 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6412 -1752 6458 -1552 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6216 -1752 6262 -1552 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6020 -1752 6066 -1552 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6804 -1406 6850 -1206 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6608 -1406 6654 -1206 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6412 -1406 6458 -1206 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6216 -1406 6262 -1206 8 DN_INPUT
port 3 nsew
rlabel metal1 s 6020 -1406 6066 -1236 8 DN_INPUT
port 3 nsew
rlabel metal1 s 4353 -2171 4397 -1380 8 DN_INPUT
port 3 nsew
rlabel metal1 s 4333 -1380 5309 -1336 8 DN_INPUT
port 3 nsew
rlabel metal1 s 5265 -1336 5309 -1236 8 DN_INPUT
port 3 nsew
rlabel metal1 s 5265 -1236 6067 -1192 8 DN_INPUT
port 3 nsew
rlabel locali s 4310 -2309 4465 -2300 8 DN_INPUT
port 3 nsew
rlabel locali s -26307 -2300 4465 -2204 2 DN_INPUT
port 3 nsew
rlabel locali s 4310 -2204 4465 -2171 8 DN_INPUT
port 3 nsew
rlabel locali s 6810 -1756 6844 -1499 8 DN_INPUT
port 3 nsew
rlabel locali s 6614 -1756 6648 -1499 8 DN_INPUT
port 3 nsew
rlabel locali s 6418 -1756 6452 -1499 8 DN_INPUT
port 3 nsew
rlabel locali s 6222 -1756 6256 -1499 8 DN_INPUT
port 3 nsew
rlabel locali s 6026 -1756 6060 -1499 8 DN_INPUT
port 3 nsew
rlabel locali s 6026 -1499 6844 -1465 8 DN_INPUT
port 3 nsew
rlabel locali s 6810 -1465 6844 -1202 8 DN_INPUT
port 3 nsew
rlabel locali s 6614 -1465 6648 -1202 8 DN_INPUT
port 3 nsew
rlabel locali s 6418 -1465 6452 -1202 8 DN_INPUT
port 3 nsew
rlabel locali s 6222 -1465 6256 -1202 8 DN_INPUT
port 3 nsew
rlabel locali s 6026 -1465 6060 -1202 8 DN_INPUT
port 3 nsew
rlabel metal1 s -1585 -2584 -1283 -2369 2 S2
port 4 nsew
rlabel metal1 s -1517 -2369 -1361 -342 2 S2
port 4 nsew
rlabel metal1 s 4383 -213 4585 -15 8 S2
port 4 nsew
rlabel metal1 s -1581 -342 -1323 -85 2 S2
port 4 nsew
rlabel metal1 s 4408 -15 4507 1066 6 S2
port 4 nsew
rlabel metal1 s 4388 1066 4549 1243 6 S2
port 4 nsew
rlabel locali s -1585 -2584 -1283 -2533 2 S2
port 4 nsew
rlabel locali s -26253 -2533 -1283 -2393 2 S2
port 4 nsew
rlabel locali s -1585 -2393 -1283 -2369 2 S2
port 4 nsew
rlabel locali s 4383 -213 4585 -175 8 S2
port 4 nsew
rlabel locali s -1581 -342 -1323 -175 2 S2
port 4 nsew
rlabel locali s -1581 -175 4585 -85 8 S2
port 4 nsew
rlabel locali s -1577 -85 4585 -36 8 S2
port 4 nsew
rlabel locali s 4383 -36 4585 -15 8 S2
port 4 nsew
rlabel locali s 5253 1206 5421 1214 6 S2
port 4 nsew
rlabel locali s 4388 1066 4549 1214 6 S2
port 4 nsew
rlabel locali s 4388 1214 5421 1243 6 S2
port 4 nsew
rlabel locali s 4400 1243 5421 1266 6 S2
port 4 nsew
rlabel locali s 5253 1266 5421 1280 6 S2
port 4 nsew
rlabel locali s 4400 1266 4452 1871 6 S2
port 4 nsew
rlabel locali s 4272 1871 4571 1945 6 S2
port 4 nsew
rlabel metal1 s 3196 -2900 3624 -2539 8 S3
port 5 nsew
rlabel metal1 s 3313 -2539 3558 -911 8 S3
port 5 nsew
rlabel metal1 s 3281 -911 3574 -645 8 S3
port 5 nsew
rlabel locali s 3196 -2900 3624 -2873 8 S3
port 5 nsew
rlabel locali s -26211 -2873 3624 -2628 2 S3
port 5 nsew
rlabel locali s 3196 -2628 3624 -2539 8 S3
port 5 nsew
rlabel locali s 5268 -1484 5436 -1476 8 S3
port 5 nsew
rlabel locali s 4415 -1476 5436 -1424 8 S3
port 5 nsew
rlabel locali s 5268 -1424 5436 -1410 8 S3
port 5 nsew
rlabel locali s 4415 -1424 4467 -819 8 S3
port 5 nsew
rlabel locali s 3281 -911 3574 -819 8 S3
port 5 nsew
rlabel locali s 3281 -819 4586 -745 8 S3
port 5 nsew
rlabel locali s 3281 -745 3574 -645 8 S3
port 5 nsew
rlabel metal1 s 15440 -3211 15853 -2842 8 UP_OUT
port 6 nsew
rlabel metal1 s 15547 -2842 15703 1597 8 UP_OUT
port 6 nsew
rlabel metal1 s 11326 1049 11372 1550 6 UP_OUT
port 6 nsew
rlabel metal1 s 11090 1049 11136 1550 6 UP_OUT
port 6 nsew
rlabel metal1 s 10854 1049 10900 1550 6 UP_OUT
port 6 nsew
rlabel metal1 s 10618 1049 10664 1550 6 UP_OUT
port 6 nsew
rlabel metal1 s 10382 1049 10428 1550 6 UP_OUT
port 6 nsew
rlabel metal1 s 10146 1049 10192 1550 6 UP_OUT
port 6 nsew
rlabel metal1 s 9910 1049 9956 1550 6 UP_OUT
port 6 nsew
rlabel metal1 s 9674 1049 9720 1550 6 UP_OUT
port 6 nsew
rlabel metal1 s 9674 1550 11372 1596 6 UP_OUT
port 6 nsew
rlabel metal1 s 15522 1597 15742 1833 6 UP_OUT
port 6 nsew
rlabel metal1 s 11326 1596 11372 1712 6 UP_OUT
port 6 nsew
rlabel metal1 s 11280 1712 15157 1786 6 UP_OUT
port 6 nsew
rlabel metal1 s 15082 1786 15128 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 14846 1786 14892 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 14610 1786 14656 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 14374 1786 14420 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 14138 1786 14184 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 13902 1786 13948 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 13666 1786 13712 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 13430 1786 13476 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 13194 1786 13240 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 12958 1786 13004 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 12722 1786 12768 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 12486 1786 12532 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 12250 1786 12296 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 12014 1786 12060 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 11778 1786 11824 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 11542 1786 11588 2257 6 UP_OUT
port 6 nsew
rlabel metal1 s 11306 1786 11352 2257 6 UP_OUT
port 6 nsew
rlabel locali s 15440 -3211 15853 -3188 8 UP_OUT
port 6 nsew
rlabel locali s -26114 -3188 15853 -2934 2 UP_OUT
port 6 nsew
rlabel locali s 15440 -2934 15853 -2842 8 UP_OUT
port 6 nsew
rlabel locali s 11332 1045 11366 1453 6 UP_OUT
port 6 nsew
rlabel locali s 11096 1045 11130 1453 6 UP_OUT
port 6 nsew
rlabel locali s 10860 1045 10894 1453 6 UP_OUT
port 6 nsew
rlabel locali s 10624 1045 10658 1453 6 UP_OUT
port 6 nsew
rlabel locali s 10388 1045 10422 1453 6 UP_OUT
port 6 nsew
rlabel locali s 10152 1045 10186 1453 6 UP_OUT
port 6 nsew
rlabel locali s 9916 1045 9950 1453 6 UP_OUT
port 6 nsew
rlabel locali s 9680 1045 9714 1453 6 UP_OUT
port 6 nsew
rlabel locali s 15522 1597 15742 1673 6 UP_OUT
port 6 nsew
rlabel locali s 15088 1673 15742 1707 6 UP_OUT
port 6 nsew
rlabel locali s 15522 1707 15742 1833 6 UP_OUT
port 6 nsew
rlabel locali s 15088 1707 15122 2261 6 UP_OUT
port 6 nsew
rlabel locali s 14852 1853 14886 2261 6 UP_OUT
port 6 nsew
rlabel locali s 14616 1853 14650 2261 6 UP_OUT
port 6 nsew
rlabel locali s 14380 1853 14414 2261 6 UP_OUT
port 6 nsew
rlabel locali s 14144 1853 14178 2261 6 UP_OUT
port 6 nsew
rlabel locali s 13908 1853 13942 2261 6 UP_OUT
port 6 nsew
rlabel locali s 13672 1853 13706 2261 6 UP_OUT
port 6 nsew
rlabel locali s 13436 1853 13470 2261 6 UP_OUT
port 6 nsew
rlabel locali s 13200 1853 13234 2261 6 UP_OUT
port 6 nsew
rlabel locali s 12964 1853 12998 2261 6 UP_OUT
port 6 nsew
rlabel locali s 12728 1853 12762 2261 6 UP_OUT
port 6 nsew
rlabel locali s 12492 1853 12526 2261 6 UP_OUT
port 6 nsew
rlabel locali s 12256 1853 12290 2261 6 UP_OUT
port 6 nsew
rlabel locali s 12020 1853 12054 2261 6 UP_OUT
port 6 nsew
rlabel locali s 11784 1853 11818 2261 6 UP_OUT
port 6 nsew
rlabel locali s 11548 1853 11582 2261 6 UP_OUT
port 6 nsew
rlabel locali s 11312 1853 11346 2261 6 UP_OUT
port 6 nsew
rlabel metal1 s 16088 -3623 16483 -3292 8 DN_OUT
port 7 nsew
rlabel metal1 s 16133 -3292 16375 -1228 8 DN_OUT
port 7 nsew
rlabel metal1 s 16101 -1228 16445 -871 8 DN_OUT
port 7 nsew
rlabel metal1 s 11285 -1707 11331 -1206 8 DN_OUT
port 7 nsew
rlabel metal1 s 11049 -1707 11095 -1206 8 DN_OUT
port 7 nsew
rlabel metal1 s 10813 -1707 10859 -1206 8 DN_OUT
port 7 nsew
rlabel metal1 s 10577 -1707 10623 -1206 8 DN_OUT
port 7 nsew
rlabel metal1 s 10341 -1707 10387 -1206 8 DN_OUT
port 7 nsew
rlabel metal1 s 10105 -1707 10151 -1206 8 DN_OUT
port 7 nsew
rlabel metal1 s 9869 -1707 9915 -1206 8 DN_OUT
port 7 nsew
rlabel metal1 s 9633 -1707 9679 -1206 8 DN_OUT
port 7 nsew
rlabel metal1 s 9633 -1206 11331 -1160 8 DN_OUT
port 7 nsew
rlabel metal1 s 11285 -1160 11331 -1044 8 DN_OUT
port 7 nsew
rlabel metal1 s 11239 -1044 15116 -970 8 DN_OUT
port 7 nsew
rlabel metal1 s 15041 -970 15087 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 14805 -970 14851 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 14569 -970 14615 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 14333 -970 14379 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 14097 -970 14143 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 13861 -970 13907 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 13625 -970 13671 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 13389 -970 13435 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 13153 -970 13199 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 12917 -970 12963 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 12681 -970 12727 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 12445 -970 12491 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 12209 -970 12255 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 11973 -970 12019 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 11737 -970 11783 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 11501 -970 11547 -499 8 DN_OUT
port 7 nsew
rlabel metal1 s 11265 -970 11311 -499 8 DN_OUT
port 7 nsew
rlabel locali s 16088 -3623 16483 -3586 8 DN_OUT
port 7 nsew
rlabel locali s -26140 -3586 16483 -3296 2 DN_OUT
port 7 nsew
rlabel locali s 16088 -3296 16483 -3292 8 DN_OUT
port 7 nsew
rlabel locali s 11291 -1711 11325 -1303 8 DN_OUT
port 7 nsew
rlabel locali s 11055 -1711 11089 -1303 8 DN_OUT
port 7 nsew
rlabel locali s 10819 -1711 10853 -1303 8 DN_OUT
port 7 nsew
rlabel locali s 10583 -1711 10617 -1303 8 DN_OUT
port 7 nsew
rlabel locali s 10347 -1711 10381 -1303 8 DN_OUT
port 7 nsew
rlabel locali s 10111 -1711 10145 -1303 8 DN_OUT
port 7 nsew
rlabel locali s 9875 -1711 9909 -1303 8 DN_OUT
port 7 nsew
rlabel locali s 9639 -1711 9673 -1303 8 DN_OUT
port 7 nsew
rlabel locali s 16101 -1228 16445 -1127 8 DN_OUT
port 7 nsew
rlabel locali s 15047 -1127 16445 -1021 8 DN_OUT
port 7 nsew
rlabel locali s 16101 -1021 16445 -871 8 DN_OUT
port 7 nsew
rlabel locali s 15047 -1021 15081 -495 8 DN_OUT
port 7 nsew
rlabel locali s 14811 -903 14845 -495 8 DN_OUT
port 7 nsew
rlabel locali s 14575 -903 14609 -495 8 DN_OUT
port 7 nsew
rlabel locali s 14339 -903 14373 -495 8 DN_OUT
port 7 nsew
rlabel locali s 14103 -903 14137 -495 8 DN_OUT
port 7 nsew
rlabel locali s 13867 -903 13901 -495 8 DN_OUT
port 7 nsew
rlabel locali s 13631 -903 13665 -495 8 DN_OUT
port 7 nsew
rlabel locali s 13395 -903 13429 -495 8 DN_OUT
port 7 nsew
rlabel locali s 13159 -903 13193 -495 8 DN_OUT
port 7 nsew
rlabel locali s 12923 -903 12957 -495 8 DN_OUT
port 7 nsew
rlabel locali s 12687 -903 12721 -495 8 DN_OUT
port 7 nsew
rlabel locali s 12451 -903 12485 -495 8 DN_OUT
port 7 nsew
rlabel locali s 12215 -903 12249 -495 8 DN_OUT
port 7 nsew
rlabel locali s 11979 -903 12013 -495 8 DN_OUT
port 7 nsew
rlabel locali s 11743 -903 11777 -495 8 DN_OUT
port 7 nsew
rlabel locali s 11507 -903 11541 -495 8 DN_OUT
port 7 nsew
rlabel locali s 11271 -903 11305 -495 8 DN_OUT
port 7 nsew
rlabel metal1 s 17293 -4848 17906 296 8 ITAIL
port 8 nsew
rlabel metal1 s 16519 296 17906 909 6 ITAIL
port 8 nsew
rlabel metal1 s 16519 909 17132 8006 6 ITAIL
port 8 nsew
rlabel metal1 s 10748 4643 10794 5443 6 ITAIL
port 8 nsew
rlabel metal1 s 9032 4643 9078 5443 6 ITAIL
port 8 nsew
rlabel metal1 s 14443 6016 14691 6213 6 ITAIL
port 8 nsew
rlabel metal1 s 14484 6213 14653 7642 6 ITAIL
port 8 nsew
rlabel metal1 s 14484 7642 14795 7749 6 ITAIL
port 8 nsew
rlabel metal1 s 14484 7749 14796 7856 6 ITAIL
port 8 nsew
rlabel metal1 s 14484 7856 14591 7858 6 ITAIL
port 8 nsew
rlabel locali s 17293 -4848 17906 -4766 8 ITAIL
port 8 nsew
rlabel locali s -26205 -4766 17906 -4354 2 ITAIL
port 8 nsew
rlabel locali s 16975 -4354 17906 -4336 8 ITAIL
port 8 nsew
rlabel locali s 17293 -4336 17906 -4235 8 ITAIL
port 8 nsew
rlabel locali s 10754 4639 10788 5501 6 ITAIL
port 8 nsew
rlabel locali s 9038 4639 9072 5496 6 ITAIL
port 8 nsew
rlabel locali s 11815 5565 12295 5710 6 ITAIL
port 8 nsew
rlabel locali s 10711 5501 10837 5592 6 ITAIL
port 8 nsew
rlabel locali s 9012 5496 9098 5582 6 ITAIL
port 8 nsew
rlabel locali s 14443 6016 14691 6038 6 ITAIL
port 8 nsew
rlabel locali s 12023 5710 12136 6038 6 ITAIL
port 8 nsew
rlabel locali s 12023 6038 14691 6151 6 ITAIL
port 8 nsew
rlabel locali s 14443 6151 14691 6213 6 ITAIL
port 8 nsew
rlabel locali s 16664 7621 16961 7685 6 ITAIL
port 8 nsew
rlabel locali s 14552 7642 14795 7685 6 ITAIL
port 8 nsew
rlabel locali s 14552 7685 16961 7821 6 ITAIL
port 8 nsew
rlabel locali s 16664 7821 16961 7884 6 ITAIL
port 8 nsew
rlabel locali s 14552 7821 14795 7846 6 ITAIL
port 8 nsew
rlabel metal1 s 17978 -5437 18468 -4849 8 S4
port 9 nsew
rlabel metal1 s 18137 -4849 18324 2985 8 S4
port 9 nsew
rlabel metal1 s 18137 2985 18330 3181 6 S4
port 9 nsew
rlabel metal1 s 18137 3181 18324 3184 6 S4
port 9 nsew
rlabel locali s 17978 -5437 18468 -5399 8 S4
port 9 nsew
rlabel locali s -26311 -5399 18468 -5013 2 S4
port 9 nsew
rlabel locali s 17978 -5013 18468 -4849 8 S4
port 9 nsew
rlabel locali s 20532 2371 20700 2379 6 S4
port 9 nsew
rlabel locali s 19679 2379 20700 2431 6 S4
port 9 nsew
rlabel locali s 20532 2431 20700 2445 6 S4
port 9 nsew
rlabel locali s 19679 2431 19731 3036 6 S4
port 9 nsew
rlabel locali s 18156 2985 18330 3036 6 S4
port 9 nsew
rlabel locali s 18156 3036 19850 3110 6 S4
port 9 nsew
rlabel locali s 18156 3110 18330 3181 6 S4
port 9 nsew
rlabel metal1 s 18424 -6171 19081 -5532 8 VCTRL_IN
port 10 nsew
rlabel metal1 s 22068 2103 22114 2303 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 21872 2103 21918 2303 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 21676 2103 21722 2303 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 21480 2103 21526 2303 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 21284 2103 21330 2303 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 22068 2449 22114 2649 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 21872 2449 21918 2649 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 21676 2449 21722 2649 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 21480 2449 21526 2649 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 21284 2449 21330 2619 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 19341 2444 19481 2475 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 19341 2475 20573 2519 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 20529 2519 20573 2619 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 19341 2519 19481 2579 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 18621 -5532 18758 2557 8 VCTRL_IN
port 10 nsew
rlabel metal1 s 20529 2619 21331 2663 6 VCTRL_IN
port 10 nsew
rlabel locali s -26321 -6098 18704 -6062 2 VCTRL_IN
port 10 nsew
rlabel locali s -26321 -6062 18990 -5664 2 VCTRL_IN
port 10 nsew
rlabel locali s 18534 -5664 18990 -5587 8 VCTRL_IN
port 10 nsew
rlabel locali s 22074 2099 22108 2356 6 VCTRL_IN
port 10 nsew
rlabel locali s 21878 2099 21912 2356 6 VCTRL_IN
port 10 nsew
rlabel locali s 21682 2099 21716 2356 6 VCTRL_IN
port 10 nsew
rlabel locali s 21486 2099 21520 2356 6 VCTRL_IN
port 10 nsew
rlabel locali s 21290 2099 21324 2356 6 VCTRL_IN
port 10 nsew
rlabel locali s 21290 2356 22108 2390 6 VCTRL_IN
port 10 nsew
rlabel locali s 22074 2390 22108 2653 6 VCTRL_IN
port 10 nsew
rlabel locali s 21878 2390 21912 2653 6 VCTRL_IN
port 10 nsew
rlabel locali s 21682 2390 21716 2653 6 VCTRL_IN
port 10 nsew
rlabel locali s 21486 2390 21520 2653 6 VCTRL_IN
port 10 nsew
rlabel locali s 21290 2390 21324 2653 6 VCTRL_IN
port 10 nsew
rlabel locali s 19341 2444 19481 2447 6 VCTRL_IN
port 10 nsew
rlabel locali s 18629 2441 18739 2447 6 VCTRL_IN
port 10 nsew
rlabel locali s 18629 2447 19481 2540 6 VCTRL_IN
port 10 nsew
rlabel locali s 19341 2540 19481 2579 6 VCTRL_IN
port 10 nsew
rlabel locali s 18629 2540 18739 2549 6 VCTRL_IN
port 10 nsew
rlabel metal1 s 18949 -6850 19611 -6293 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 22240 -1247 22286 -1047 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 22044 -1247 22090 -1047 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 21848 -1247 21894 -1047 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 21652 -1247 21698 -1047 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 21456 -1247 21502 -1047 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 22240 -901 22286 -701 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 22044 -901 22090 -701 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 21848 -901 21894 -701 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 21652 -901 21698 -701 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 21456 -901 21502 -731 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 19212 -6293 19542 -875 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 19212 -875 20745 -831 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 20701 -831 20745 -731 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 19212 -831 19359 -829 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 20701 -731 21503 -687 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 18949 -6850 19611 -6787 8 LF_OFFCHIP
port 11 nsew
rlabel locali s -26653 -6787 19611 -6346 2 LF_OFFCHIP
port 11 nsew
rlabel locali s 18949 -6346 19611 -6293 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 22246 -1251 22280 -994 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 22050 -1251 22084 -994 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 21854 -1251 21888 -994 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 21658 -1251 21692 -994 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 21462 -1251 21496 -994 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 21462 -994 22280 -960 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 22246 -960 22280 -697 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 22050 -960 22084 -697 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 21854 -960 21888 -697 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 21658 -960 21692 -697 8 LF_OFFCHIP
port 11 nsew
rlabel locali s 21462 -960 21496 -697 8 LF_OFFCHIP
port 11 nsew
rlabel metal1 s 19665 -7634 20295 -7025 8 S5
port 12 nsew
rlabel metal1 s 19868 -7025 20066 -1279 8 S5
port 12 nsew
rlabel metal1 s 19836 -1279 20093 -990 8 S5
port 12 nsew
rlabel locali s 19665 -7634 20295 -7593 8 S5
port 12 nsew
rlabel locali s -26746 -7593 20295 -7100 2 S5
port 12 nsew
rlabel locali s 19665 -7100 20295 -7025 8 S5
port 12 nsew
rlabel locali s 19836 -1279 20093 -1129 8 S5
port 12 nsew
rlabel locali s 20704 -979 20872 -971 8 S5
port 12 nsew
rlabel locali s 19836 -1129 20098 -971 8 S5
port 12 nsew
rlabel locali s 19836 -971 20872 -919 8 S5
port 12 nsew
rlabel locali s 20704 -919 20872 -905 8 S5
port 12 nsew
rlabel locali s 19836 -919 20098 -916 8 S5
port 12 nsew
rlabel locali s 19851 -916 19903 -314 8 S5
port 12 nsew
rlabel locali s 19723 -314 20022 -240 8 S5
port 12 nsew
rlabel metal1 s -26820 -39467 -26273 -39421 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26319 -39421 -26273 -39231 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26820 -39231 -26273 -39185 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26319 -39185 -26273 -38995 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26820 -38995 -26273 -38949 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26319 -38949 -26273 -38759 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26820 -38759 -26273 -38713 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26319 -38713 -26273 -38523 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26820 -38523 -26273 -38477 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26319 -38477 -26273 -38287 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26820 -38287 -26273 -38241 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26319 -38241 -26273 -38051 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26820 -38051 -26273 -38005 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -37861 -26083 -37835 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -37835 -25612 -37815 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26319 -38005 -26273 -37815 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26820 -37815 -25612 -37789 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26820 -37789 -26083 -37769 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -37769 -26083 -37599 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -37599 -25612 -37553 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -37553 -26083 -37363 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -37363 -25612 -37317 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -37317 -26083 -37127 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -37127 -25612 -37081 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -37081 -26083 -36891 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -36891 -25612 -36845 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -36845 -26083 -36655 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -36655 -25612 -36609 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -36609 -26083 -36419 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -36419 -25612 -36373 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -36373 -26083 -36183 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -36183 -25612 -36137 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -36137 -26083 -35947 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -35947 -25612 -35901 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -35901 -26083 -35711 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -35711 -25612 -35665 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -35665 -26083 -35475 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -35475 -25612 -35429 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -35429 -26083 -35239 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -35239 -25612 -35193 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -35193 -26083 -35003 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -35003 -25612 -34957 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -34957 -26083 -34767 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -34767 -25612 -34721 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -34721 -26083 -34531 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -34531 -25612 -34485 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -34485 -26083 -34295 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -34295 -25612 -34249 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -34249 -26083 -34059 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -34059 -25612 -34013 2 OUT_CORE
port 13 nsew
rlabel metal1 s -26157 -34013 -26083 -33984 2 OUT_CORE
port 13 nsew
rlabel locali s -26824 -39461 -26416 -39427 2 OUT_CORE
port 13 nsew
rlabel locali s -26824 -39225 -26416 -39191 2 OUT_CORE
port 13 nsew
rlabel locali s -26824 -38989 -26416 -38955 2 OUT_CORE
port 13 nsew
rlabel locali s -26824 -38753 -26416 -38719 2 OUT_CORE
port 13 nsew
rlabel locali s -26824 -38517 -26416 -38483 2 OUT_CORE
port 13 nsew
rlabel locali s -26824 -38281 -26416 -38247 2 OUT_CORE
port 13 nsew
rlabel locali s -26824 -38045 -26416 -38011 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -37829 -25608 -37795 2 OUT_CORE
port 13 nsew
rlabel locali s -26824 -37809 -26416 -37775 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -37593 -25608 -37559 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -37357 -25608 -37323 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -37121 -25608 -37087 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -36885 -25608 -36851 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -36649 -25608 -36615 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -36413 -25608 -36379 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -36177 -25608 -36143 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -35941 -25608 -35907 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -35705 -25608 -35671 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -35469 -25608 -35435 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -35233 -25608 -35199 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -34997 -25608 -34963 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -34761 -25608 -34727 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -34525 -25608 -34491 2 OUT_CORE
port 13 nsew
rlabel locali s -26016 -34289 -25608 -34255 2 OUT_CORE
port 13 nsew
rlabel locali s -26196 -34053 -25608 -34019 2 OUT_CORE
port 13 nsew
rlabel locali s -26196 -34019 -26162 -33893 2 OUT_CORE
port 13 nsew
rlabel locali s -26347 -33893 -26140 -33190 2 OUT_CORE
port 13 nsew
rlabel locali s -32225 -33190 -26140 -32972 2 OUT_CORE
port 13 nsew
rlabel metal1 s -28640 -57612 -28093 -57566 2 OUT_USB
port 14 nsew
rlabel metal1 s -28139 -57566 -28093 -57376 2 OUT_USB
port 14 nsew
rlabel metal1 s -28640 -57376 -28093 -57330 2 OUT_USB
port 14 nsew
rlabel metal1 s -28139 -57330 -28093 -57140 2 OUT_USB
port 14 nsew
rlabel metal1 s -28640 -57140 -28093 -57094 2 OUT_USB
port 14 nsew
rlabel metal1 s -28139 -57094 -28093 -56904 2 OUT_USB
port 14 nsew
rlabel metal1 s -28640 -56904 -28093 -56858 2 OUT_USB
port 14 nsew
rlabel metal1 s -28139 -56858 -28093 -56668 2 OUT_USB
port 14 nsew
rlabel metal1 s -28640 -56668 -28093 -56622 2 OUT_USB
port 14 nsew
rlabel metal1 s -28139 -56622 -28093 -56432 2 OUT_USB
port 14 nsew
rlabel metal1 s -28640 -56432 -28093 -56386 2 OUT_USB
port 14 nsew
rlabel metal1 s -28139 -56386 -28093 -56196 2 OUT_USB
port 14 nsew
rlabel metal1 s -28640 -56196 -28093 -56150 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -56006 -27903 -55980 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -55980 -27432 -55960 2 OUT_USB
port 14 nsew
rlabel metal1 s -28139 -56150 -28093 -55960 2 OUT_USB
port 14 nsew
rlabel metal1 s -28640 -55960 -27432 -55934 2 OUT_USB
port 14 nsew
rlabel metal1 s -28640 -55934 -27903 -55914 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -55914 -27903 -55744 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -55744 -27432 -55698 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -55698 -27903 -55508 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -55508 -27432 -55462 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -55462 -27903 -55272 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -55272 -27432 -55226 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -55226 -27903 -55036 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -55036 -27432 -54990 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -54990 -27903 -54800 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -54800 -27432 -54754 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -54754 -27903 -54564 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -54564 -27432 -54518 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -54518 -27903 -54328 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -54328 -27432 -54282 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -54282 -27903 -54092 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -54092 -27432 -54046 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -54046 -27903 -53856 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -53856 -27432 -53810 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -53810 -27903 -53620 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -53620 -27432 -53574 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -53574 -27903 -53384 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -53384 -27432 -53338 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -53338 -27903 -53148 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -53148 -27432 -53102 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -53102 -27903 -52912 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -52912 -27432 -52866 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -52866 -27903 -52676 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -52676 -27432 -52630 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -52630 -27903 -52440 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -52440 -27432 -52394 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -52394 -27903 -52204 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -52204 -27432 -52158 2 OUT_USB
port 14 nsew
rlabel metal1 s -27977 -52158 -27903 -52129 2 OUT_USB
port 14 nsew
rlabel locali s -28644 -57606 -28236 -57572 2 OUT_USB
port 14 nsew
rlabel locali s -28644 -57370 -28236 -57336 2 OUT_USB
port 14 nsew
rlabel locali s -28644 -57134 -28236 -57100 2 OUT_USB
port 14 nsew
rlabel locali s -28644 -56898 -28236 -56864 2 OUT_USB
port 14 nsew
rlabel locali s -28644 -56662 -28236 -56628 2 OUT_USB
port 14 nsew
rlabel locali s -28644 -56426 -28236 -56392 2 OUT_USB
port 14 nsew
rlabel locali s -28644 -56190 -28236 -56156 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -55974 -27428 -55940 2 OUT_USB
port 14 nsew
rlabel locali s -28644 -55954 -28236 -55920 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -55738 -27428 -55704 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -55502 -27428 -55468 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -55266 -27428 -55232 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -55030 -27428 -54996 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -54794 -27428 -54760 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -54558 -27428 -54524 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -54322 -27428 -54288 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -54086 -27428 -54052 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -53850 -27428 -53816 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -53614 -27428 -53580 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -53378 -27428 -53344 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -53142 -27428 -53108 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -52906 -27428 -52872 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -52670 -27428 -52636 2 OUT_USB
port 14 nsew
rlabel locali s -27836 -52434 -27428 -52400 2 OUT_USB
port 14 nsew
rlabel locali s -28016 -52198 -27428 -52164 2 OUT_USB
port 14 nsew
rlabel locali s -28016 -52164 -27982 -52016 2 OUT_USB
port 14 nsew
rlabel locali s -28065 -52016 -27886 -50847 2 OUT_USB
port 14 nsew
rlabel locali s -32776 -50847 -27886 -50668 2 OUT_USB
port 14 nsew
rlabel metal1 s -5288 -43468 -5149 -43467 2 D12
port 15 nsew
rlabel metal1 s -5288 -43467 -4757 -43465 2 D12
port 15 nsew
rlabel metal1 s -6366 -43474 -6227 -43465 2 D12
port 15 nsew
rlabel metal1 s -6366 -43465 -4757 -43439 2 D12
port 15 nsew
rlabel metal1 s -4785 -43439 -4757 -42289 2 D12
port 15 nsew
rlabel metal1 s -6366 -43439 -5149 -43437 2 D12
port 15 nsew
rlabel metal1 s -5288 -43437 -5149 -43414 2 D12
port 15 nsew
rlabel metal1 s -6366 -43437 -6227 -43420 2 D12
port 15 nsew
rlabel metal1 s -4785 -42289 9423 -42238 8 D12
port 15 nsew
rlabel metal1 s 9372 -42238 9423 -36888 8 D12
port 15 nsew
rlabel metal1 s -13584 -39248 -13454 -39098 2 D12
port 15 nsew
rlabel metal1 s -13534 -39098 -13480 -38901 2 D12
port 15 nsew
rlabel metal1 s -15145 -44640 -14969 -38901 2 D12
port 15 nsew
rlabel metal1 s -23239 -44638 -23116 -44515 2 D12
port 15 nsew
rlabel metal1 s -15145 -38901 -13480 -38725 2 D12
port 15 nsew
rlabel metal1 s -13534 -38725 -13480 -37694 2 D12
port 15 nsew
rlabel metal1 s -13677 -37694 -13480 -37640 2 D12
port 15 nsew
rlabel metal1 s -6442 -36888 9423 -36837 8 D12
port 15 nsew
rlabel metal1 s -6442 -36837 -6391 -36455 2 D12
port 15 nsew
rlabel metal1 s -6442 -36455 -6306 -36381 2 D12
port 15 nsew
rlabel metal1 s -23186 -44515 -23125 -35988 2 D12
port 15 nsew
rlabel locali s -32434 -44640 27308 -44504 2 D12
port 15 nsew
rlabel locali s 27172 -44504 27308 -43278 8 D12
port 15 nsew
rlabel locali s 27172 -43278 30907 -43142 8 D12
port 15 nsew
rlabel locali s 31205 -42156 31340 -42148 8 D12
port 15 nsew
rlabel locali s 31185 -42148 31340 -42146 8 D12
port 15 nsew
rlabel locali s 30771 -43142 30907 -42146 8 D12
port 15 nsew
rlabel locali s 30771 -42146 31340 -42110 8 D12
port 15 nsew
rlabel locali s 27537 -42125 27672 -42117 8 D12
port 15 nsew
rlabel locali s 27517 -42117 27672 -42115 8 D12
port 15 nsew
rlabel locali s 27172 -43142 27308 -42115 8 D12
port 15 nsew
rlabel locali s 8550 -44504 8606 -43094 8 D12
port 15 nsew
rlabel locali s -5288 -43468 -5149 -43414 2 D12
port 15 nsew
rlabel locali s -6366 -43474 -6227 -43420 2 D12
port 15 nsew
rlabel locali s 8549 -43094 8607 -42286 8 D12
port 15 nsew
rlabel locali s 8549 -42286 8673 -42243 8 D12
port 15 nsew
rlabel locali s 8550 -42243 8673 -42242 8 D12
port 15 nsew
rlabel locali s 31185 -42110 31340 -42108 8 D12
port 15 nsew
rlabel locali s 31205 -42108 31340 -42102 8 D12
port 15 nsew
rlabel locali s 26989 -42115 27672 -42079 8 D12
port 15 nsew
rlabel locali s 27517 -42079 27672 -42077 8 D12
port 15 nsew
rlabel locali s 27537 -42077 27672 -42071 8 D12
port 15 nsew
rlabel locali s -21357 -41813 -21212 -41757 2 D12
port 15 nsew
rlabel locali s -21357 -41757 -21297 -41752 2 D12
port 15 nsew
rlabel locali s -23186 -41767 -23126 -41752 2 D12
port 15 nsew
rlabel locali s -23186 -41752 -21297 -41711 2 D12
port 15 nsew
rlabel locali s -23186 -41711 -23126 -41530 2 D12
port 15 nsew
rlabel locali s -13410 -39162 -13337 -39156 2 D12
port 15 nsew
rlabel locali s -13584 -39248 -13454 -39156 2 D12
port 15 nsew
rlabel locali s -13584 -39156 -13337 -39115 2 D12
port 15 nsew
rlabel locali s -13410 -39115 -13337 -39102 2 D12
port 15 nsew
rlabel locali s -13584 -39115 -13454 -39098 2 D12
port 15 nsew
rlabel locali s -13036 -37710 -12962 -37684 2 D12
port 15 nsew
rlabel locali s -13674 -37686 -13447 -37684 2 D12
port 15 nsew
rlabel locali s -13674 -37684 -12962 -37646 2 D12
port 15 nsew
rlabel locali s -13448 -37646 -12962 -37645 2 D12
port 15 nsew
rlabel locali s -13036 -37645 -12962 -37639 2 D12
port 15 nsew
rlabel locali s -13448 -37645 -13377 -37644 2 D12
port 15 nsew
rlabel locali s -6442 -36455 -6254 -36381 2 D12
port 15 nsew
rlabel locali s -21593 -36232 -21458 -36225 2 D12
port 15 nsew
rlabel locali s -23186 -36226 -23125 -36225 2 D12
port 15 nsew
rlabel locali s -23186 -36225 -21458 -36191 2 D12
port 15 nsew
rlabel locali s -21593 -36191 -21458 -36178 2 D12
port 15 nsew
rlabel locali s -23186 -36191 -23125 -35988 2 D12
port 15 nsew
rlabel metal1 s 8591 -44832 8714 -44709 8 D13
port 16 nsew
rlabel metal1 s -23048 -44837 -22925 -44714 2 D13
port 16 nsew
rlabel metal1 s 8644 -44709 8705 -44105 8 D13
port 16 nsew
rlabel metal1 s 8649 -43472 8714 -43467 8 D13
port 16 nsew
rlabel metal1 s 7712 -43468 7851 -43467 8 D13
port 16 nsew
rlabel metal1 s 7610 -43467 10221 -43465 8 D13
port 16 nsew
rlabel metal1 s 6634 -43474 6773 -43465 8 D13
port 16 nsew
rlabel metal1 s 6634 -43465 10221 -43439 8 D13
port 16 nsew
rlabel metal1 s 10193 -43439 10221 -35687 8 D13
port 16 nsew
rlabel metal1 s 8649 -43439 8714 -43335 8 D13
port 16 nsew
rlabel metal1 s 6634 -43439 7851 -43437 8 D13
port 16 nsew
rlabel metal1 s 7712 -43437 7851 -43414 8 D13
port 16 nsew
rlabel metal1 s 6634 -43437 6773 -43420 8 D13
port 16 nsew
rlabel metal1 s -22995 -44714 -22934 -35909 2 D13
port 16 nsew
rlabel metal1 s 7712 -35712 7851 -35689 8 D13
port 16 nsew
rlabel metal1 s 6634 -35706 6773 -35689 8 D13
port 16 nsew
rlabel metal1 s 6634 -35689 7851 -35687 8 D13
port 16 nsew
rlabel metal1 s 6634 -35687 10221 -35661 8 D13
port 16 nsew
rlabel metal1 s 7610 -35661 10221 -35659 8 D13
port 16 nsew
rlabel metal1 s 7712 -35659 7851 -35658 8 D13
port 16 nsew
rlabel metal1 s 6634 -35661 6773 -35652 8 D13
port 16 nsew
rlabel locali s -32450 -44839 35748 -44703 8 D13
port 16 nsew
rlabel locali s 35612 -44703 35748 -43289 8 D13
port 16 nsew
rlabel locali s 8652 -44232 8706 -43472 8 D13
port 16 nsew
rlabel locali s 8649 -43472 8714 -43335 8 D13
port 16 nsew
rlabel locali s 7712 -43468 7851 -43414 8 D13
port 16 nsew
rlabel locali s 6634 -43474 6773 -43420 8 D13
port 16 nsew
rlabel locali s 35612 -43289 39347 -43153 8 D13
port 16 nsew
rlabel locali s 39645 -42167 39780 -42159 8 D13
port 16 nsew
rlabel locali s 39625 -42159 39780 -42157 8 D13
port 16 nsew
rlabel locali s 39211 -43153 39347 -42157 8 D13
port 16 nsew
rlabel locali s 39211 -42157 39780 -42121 8 D13
port 16 nsew
rlabel locali s 35977 -42136 36112 -42128 8 D13
port 16 nsew
rlabel locali s 35957 -42128 36112 -42126 8 D13
port 16 nsew
rlabel locali s 35612 -43153 35748 -42126 8 D13
port 16 nsew
rlabel locali s 39625 -42121 39780 -42119 8 D13
port 16 nsew
rlabel locali s 39645 -42119 39780 -42113 8 D13
port 16 nsew
rlabel locali s 35429 -42126 36112 -42090 8 D13
port 16 nsew
rlabel locali s 35957 -42090 36112 -42088 8 D13
port 16 nsew
rlabel locali s 35977 -42088 36112 -42082 8 D13
port 16 nsew
rlabel locali s -21677 -41845 -21532 -41841 2 D13
port 16 nsew
rlabel locali s -22995 -42024 -22935 -41841 2 D13
port 16 nsew
rlabel locali s -22995 -41841 -21532 -41800 2 D13
port 16 nsew
rlabel locali s -21677 -41800 -21532 -41789 2 D13
port 16 nsew
rlabel locali s -22995 -41800 -22935 -41787 2 D13
port 16 nsew
rlabel locali s -21781 -36154 -21646 -36147 2 D13
port 16 nsew
rlabel locali s -22995 -36147 -21646 -36109 2 D13
port 16 nsew
rlabel locali s -21781 -36109 -21646 -36100 2 D13
port 16 nsew
rlabel locali s -22995 -36109 -22934 -35909 2 D13
port 16 nsew
rlabel locali s 7712 -35712 7851 -35658 8 D13
port 16 nsew
rlabel locali s 6634 -35706 6773 -35652 8 D13
port 16 nsew
rlabel metal1 s 8697 -45065 8820 -44942 8 D14
port 17 nsew
rlabel metal1 s -22942 -45070 -22819 -44947 2 D14
port 17 nsew
rlabel metal1 s 8753 -44942 8813 -44109 8 D14
port 17 nsew
rlabel metal1 s 8762 -44109 8806 -44106 8 D14
port 17 nsew
rlabel metal1 s 4712 -43468 4851 -43467 8 D14
port 17 nsew
rlabel metal1 s 4712 -43467 6071 -43465 8 D14
port 17 nsew
rlabel metal1 s 3634 -43474 3773 -43465 8 D14
port 17 nsew
rlabel metal1 s 3634 -43465 6071 -43439 8 D14
port 17 nsew
rlabel metal1 s 8684 -42845 8823 -42841 8 D14
port 17 nsew
rlabel metal1 s 6043 -43439 6071 -42841 8 D14
port 17 nsew
rlabel metal1 s 3634 -43439 4851 -43437 8 D14
port 17 nsew
rlabel metal1 s 4712 -43437 4851 -43414 8 D14
port 17 nsew
rlabel metal1 s 3634 -43437 3773 -43420 8 D14
port 17 nsew
rlabel metal1 s 6043 -42841 10070 -42813 8 D14
port 17 nsew
rlabel metal1 s 10042 -42813 10070 -36313 8 D14
port 17 nsew
rlabel metal1 s 8684 -42813 8823 -42798 8 D14
port 17 nsew
rlabel metal1 s -22886 -44947 -22826 -42127 2 D14
port 17 nsew
rlabel metal1 s -22886 -42127 -22825 -41890 2 D14
port 17 nsew
rlabel metal1 s 6043 -36313 10070 -36285 8 D14
port 17 nsew
rlabel metal1 s 6043 -36285 6071 -35687 8 D14
port 17 nsew
rlabel metal1 s -22886 -41890 -22826 -36061 2 D14
port 17 nsew
rlabel metal1 s -22886 -36061 -22825 -35823 2 D14
port 17 nsew
rlabel metal1 s 4712 -35712 4851 -35689 8 D14
port 17 nsew
rlabel metal1 s 3634 -35706 3773 -35689 8 D14
port 17 nsew
rlabel metal1 s 3634 -35689 4851 -35687 8 D14
port 17 nsew
rlabel metal1 s 3634 -35687 6071 -35661 8 D14
port 17 nsew
rlabel metal1 s 4712 -35661 6071 -35659 8 D14
port 17 nsew
rlabel metal1 s 4712 -35659 4851 -35658 8 D14
port 17 nsew
rlabel metal1 s 3634 -35661 3773 -35652 8 D14
port 17 nsew
rlabel locali s -32458 -45072 44658 -44936 8 D14
port 17 nsew
rlabel locali s 44522 -44936 44658 -43328 8 D14
port 17 nsew
rlabel locali s 44475 -43328 48210 -43192 8 D14
port 17 nsew
rlabel locali s 48508 -42206 48643 -42198 8 D14
port 17 nsew
rlabel locali s 48488 -42198 48643 -42196 8 D14
port 17 nsew
rlabel locali s 48074 -43192 48210 -42196 8 D14
port 17 nsew
rlabel locali s 44475 -43192 44658 -43178 8 D14
port 17 nsew
rlabel locali s 48074 -42196 48643 -42160 8 D14
port 17 nsew
rlabel locali s 44840 -42175 44975 -42167 8 D14
port 17 nsew
rlabel locali s 44820 -42167 44975 -42165 8 D14
port 17 nsew
rlabel locali s 44475 -43178 44611 -42165 8 D14
port 17 nsew
rlabel locali s 8757 -44232 8811 -42844 8 D14
port 17 nsew
rlabel locali s 4712 -43468 4851 -43414 8 D14
port 17 nsew
rlabel locali s 3634 -43474 3773 -43420 8 D14
port 17 nsew
rlabel locali s 8693 -42844 8816 -42800 8 D14
port 17 nsew
rlabel locali s 48488 -42160 48643 -42158 8 D14
port 17 nsew
rlabel locali s 48508 -42158 48643 -42152 8 D14
port 17 nsew
rlabel locali s 44292 -42165 44975 -42129 8 D14
port 17 nsew
rlabel locali s 44820 -42129 44975 -42127 8 D14
port 17 nsew
rlabel locali s 44840 -42127 44975 -42121 8 D14
port 17 nsew
rlabel locali s -22006 -41940 -21861 -41933 2 D14
port 17 nsew
rlabel locali s -22885 -42127 -22825 -41933 2 D14
port 17 nsew
rlabel locali s -22885 -41933 -21861 -41892 2 D14
port 17 nsew
rlabel locali s -22006 -41892 -21861 -41884 2 D14
port 17 nsew
rlabel locali s -22885 -41892 -22825 -41890 2 D14
port 17 nsew
rlabel locali s -22117 -36072 -21982 -36063 2 D14
port 17 nsew
rlabel locali s -22136 -36063 -21982 -36061 2 D14
port 17 nsew
rlabel locali s -22886 -36061 -21982 -36026 2 D14
port 17 nsew
rlabel locali s -22117 -36026 -21982 -36018 2 D14
port 17 nsew
rlabel locali s -22886 -36026 -22825 -35823 2 D14
port 17 nsew
rlabel locali s 4712 -35712 4851 -35658 8 D14
port 17 nsew
rlabel locali s 3634 -35706 3773 -35652 8 D14
port 17 nsew
rlabel metal1 s 8790 -45322 8914 -45199 8 D15
port 18 nsew
rlabel metal1 s -22849 -45327 -22725 -45204 2 D15
port 18 nsew
rlabel metal1 s 8852 -45199 8913 -44252 8 D15
port 18 nsew
rlabel metal1 s -20912 -42537 -20854 -42400 2 D15
port 18 nsew
rlabel metal1 s -20892 -42400 -20857 -41491 2 D15
port 18 nsew
rlabel metal1 s -20892 -41491 -20834 -41354 2 D15
port 18 nsew
rlabel metal1 s 8833 -41228 8978 -41216 8 D15
port 18 nsew
rlabel metal1 s 7722 -41217 7861 -41216 8 D15
port 18 nsew
rlabel metal1 s 7722 -41216 9095 -41214 8 D15
port 18 nsew
rlabel metal1 s 6644 -41223 6783 -41214 8 D15
port 18 nsew
rlabel metal1 s 6644 -41214 9095 -41188 8 D15
port 18 nsew
rlabel metal1 s 9065 -41188 9093 -37953 8 D15
port 18 nsew
rlabel metal1 s 8833 -41188 8978 -41093 8 D15
port 18 nsew
rlabel metal1 s 6644 -41188 7861 -41186 8 D15
port 18 nsew
rlabel metal1 s 7722 -41186 7861 -41163 8 D15
port 18 nsew
rlabel metal1 s 6644 -41186 6783 -41169 8 D15
port 18 nsew
rlabel metal1 s 9052 -37953 9103 -37938 8 D15
port 18 nsew
rlabel metal1 s 7722 -37963 7861 -37940 8 D15
port 18 nsew
rlabel metal1 s 6644 -37957 6783 -37940 8 D15
port 18 nsew
rlabel metal1 s 6644 -37940 7861 -37938 8 D15
port 18 nsew
rlabel metal1 s 6644 -37938 9103 -37912 8 D15
port 18 nsew
rlabel metal1 s 7722 -37912 9103 -37910 8 D15
port 18 nsew
rlabel metal1 s 9052 -37910 9103 -37902 8 D15
port 18 nsew
rlabel metal1 s 7722 -37910 7861 -37909 8 D15
port 18 nsew
rlabel metal1 s 6644 -37912 6783 -37903 8 D15
port 18 nsew
rlabel metal1 s -20370 -37226 -20238 -37222 2 D15
port 18 nsew
rlabel metal1 s -20417 -37222 -20214 -37182 2 D15
port 18 nsew
rlabel metal1 s -20370 -37182 -20214 -37173 2 D15
port 18 nsew
rlabel metal1 s -20254 -37173 -20214 -36400 2 D15
port 18 nsew
rlabel metal1 s -22787 -45204 -22726 -36988 2 D15
port 18 nsew
rlabel metal1 s -20261 -36400 -20124 -36342 2 D15
port 18 nsew
rlabel locali s -32482 -45327 53809 -45191 8 D15
port 18 nsew
rlabel locali s 53673 -45191 53809 -43294 8 D15
port 18 nsew
rlabel locali s 53673 -43294 57408 -43158 8 D15
port 18 nsew
rlabel locali s 57706 -42172 57841 -42164 8 D15
port 18 nsew
rlabel locali s 57686 -42164 57841 -42162 8 D15
port 18 nsew
rlabel locali s 57272 -43158 57408 -42162 8 D15
port 18 nsew
rlabel locali s 57272 -42162 57841 -42126 8 D15
port 18 nsew
rlabel locali s 54038 -42141 54173 -42133 8 D15
port 18 nsew
rlabel locali s 54018 -42133 54173 -42131 8 D15
port 18 nsew
rlabel locali s 53673 -43158 53809 -42131 8 D15
port 18 nsew
rlabel locali s 57686 -42126 57841 -42124 8 D15
port 18 nsew
rlabel locali s 57706 -42124 57841 -42118 8 D15
port 18 nsew
rlabel locali s 53490 -42131 54173 -42095 8 D15
port 18 nsew
rlabel locali s 54018 -42095 54173 -42093 8 D15
port 18 nsew
rlabel locali s 54038 -42093 54173 -42087 8 D15
port 18 nsew
rlabel locali s 8856 -44449 8912 -41228 8 D15
port 18 nsew
rlabel locali s -22787 -42537 -20854 -42496 2 D15
port 18 nsew
rlabel locali s -20912 -42496 -20854 -42400 2 D15
port 18 nsew
rlabel locali s -22787 -42496 -22729 -42400 2 D15
port 18 nsew
rlabel locali s -20485 -41502 -20342 -41485 2 D15
port 18 nsew
rlabel locali s -20892 -41491 -20834 -41485 2 D15
port 18 nsew
rlabel locali s -20892 -41485 -20342 -41449 2 D15
port 18 nsew
rlabel locali s -20485 -41449 -20342 -41442 2 D15
port 18 nsew
rlabel locali s -20892 -41449 -20834 -41354 2 D15
port 18 nsew
rlabel locali s 8833 -41228 8978 -41093 8 D15
port 18 nsew
rlabel locali s 7722 -41217 7861 -41163 8 D15
port 18 nsew
rlabel locali s 6644 -41223 6783 -41169 8 D15
port 18 nsew
rlabel locali s 7722 -37963 7861 -37909 8 D15
port 18 nsew
rlabel locali s 6644 -37957 6783 -37903 8 D15
port 18 nsew
rlabel locali s -20370 -37226 -20238 -37222 2 D15
port 18 nsew
rlabel locali s -22787 -37226 -22727 -37222 2 D15
port 18 nsew
rlabel locali s -22787 -37222 -20238 -37182 2 D15
port 18 nsew
rlabel locali s -20370 -37182 -20238 -37173 2 D15
port 18 nsew
rlabel locali s -22787 -37182 -22727 -37105 2 D15
port 18 nsew
rlabel locali s -22787 -37105 -22719 -37065 2 D15
port 18 nsew
rlabel locali s -22787 -37065 -22727 -36989 2 D15
port 18 nsew
rlabel locali s -19661 -36393 -19587 -36387 2 D15
port 18 nsew
rlabel locali s -20073 -36388 -20002 -36387 2 D15
port 18 nsew
rlabel locali s -20073 -36387 -19587 -36386 2 D15
port 18 nsew
rlabel locali s -20261 -36400 -20124 -36386 2 D15
port 18 nsew
rlabel locali s -20299 -36386 -19587 -36348 2 D15
port 18 nsew
rlabel locali s -19661 -36348 -19587 -36322 2 D15
port 18 nsew
rlabel locali s -20299 -36348 -20072 -36346 2 D15
port 18 nsew
rlabel locali s -20261 -36346 -20124 -36342 2 D15
port 18 nsew
rlabel metal1 s 61366 -11971 62272 -11116 8 F_IN
port 19 nsew
rlabel metal1 s -6611 -11894 -5937 -11153 2 F_IN
port 19 nsew
rlabel metal1 s 64667 -4113 64713 -3913 8 F_IN
port 19 nsew
rlabel metal1 s 64471 -4113 64517 -3913 8 F_IN
port 19 nsew
rlabel metal1 s 64275 -4113 64321 -3913 8 F_IN
port 19 nsew
rlabel metal1 s 64079 -4113 64125 -3913 8 F_IN
port 19 nsew
rlabel metal1 s 63883 -4113 63929 -3913 8 F_IN
port 19 nsew
rlabel metal1 s 64667 -3767 64713 -3567 8 F_IN
port 19 nsew
rlabel metal1 s 64471 -3767 64517 -3567 8 F_IN
port 19 nsew
rlabel metal1 s 64275 -3767 64321 -3567 8 F_IN
port 19 nsew
rlabel metal1 s 64079 -3767 64125 -3567 8 F_IN
port 19 nsew
rlabel metal1 s 63883 -3767 63929 -3597 8 F_IN
port 19 nsew
rlabel metal1 s 61655 -11116 62108 -3741 8 F_IN
port 19 nsew
rlabel metal1 s 61655 -3741 63172 -3697 8 F_IN
port 19 nsew
rlabel metal1 s 63128 -3697 63172 -3597 8 F_IN
port 19 nsew
rlabel metal1 s 63128 -3597 63930 -3553 8 F_IN
port 19 nsew
rlabel metal1 s -6601 -11153 -6294 224 2 F_IN
port 19 nsew
rlabel metal1 s -6601 224 -5078 257 4 F_IN
port 19 nsew
rlabel metal1 s -6600 257 -5078 308 4 F_IN
port 19 nsew
rlabel metal1 s -6600 308 -5077 389 4 F_IN
port 19 nsew
rlabel metal1 s -6599 389 -5077 473 4 F_IN
port 19 nsew
rlabel metal1 s -1310 762 -1264 962 4 F_IN
port 19 nsew
rlabel metal1 s -1506 762 -1460 962 4 F_IN
port 19 nsew
rlabel metal1 s -1702 762 -1656 962 4 F_IN
port 19 nsew
rlabel metal1 s -1898 762 -1852 962 4 F_IN
port 19 nsew
rlabel metal1 s -2094 762 -2048 962 4 F_IN
port 19 nsew
rlabel metal1 s -5243 473 -5078 1073 4 F_IN
port 19 nsew
rlabel metal1 s -18039 321 -17604 565 4 F_IN
port 19 nsew
rlabel metal1 s -1310 1108 -1264 1308 4 F_IN
port 19 nsew
rlabel metal1 s -1506 1108 -1460 1308 4 F_IN
port 19 nsew
rlabel metal1 s -1702 1108 -1656 1308 4 F_IN
port 19 nsew
rlabel metal1 s -1898 1108 -1852 1308 4 F_IN
port 19 nsew
rlabel metal1 s -2094 1108 -2048 1278 4 F_IN
port 19 nsew
rlabel metal1 s -5243 1073 -3681 1134 4 F_IN
port 19 nsew
rlabel metal1 s -5243 1134 -2805 1178 4 F_IN
port 19 nsew
rlabel metal1 s -2849 1178 -2805 1278 4 F_IN
port 19 nsew
rlabel metal1 s -5243 1178 -3681 1219 4 F_IN
port 19 nsew
rlabel metal1 s -2849 1278 -2047 1322 4 F_IN
port 19 nsew
rlabel metal1 s -16414 9112 -16236 9129 4 F_IN
port 19 nsew
rlabel metal1 s -17836 565 -17700 9129 4 F_IN
port 19 nsew
rlabel metal1 s -17836 9129 -7080 9265 4 F_IN
port 19 nsew
rlabel metal1 s -7311 9265 -7080 9281 4 F_IN
port 19 nsew
rlabel metal1 s -7311 9281 -7025 9369 4 F_IN
port 19 nsew
rlabel metal1 s -16414 9265 -16236 9325 4 F_IN
port 19 nsew
rlabel metal1 s -7268 9369 -7025 9382 4 F_IN
port 19 nsew
rlabel metal1 s -8001 26665 -7941 26701 4 F_IN
port 19 nsew
rlabel metal1 s -8468 26701 -7941 26761 4 F_IN
port 19 nsew
rlabel metal1 s -8001 26761 -7941 26797 4 F_IN
port 19 nsew
rlabel metal1 s -10852 28438 -10792 28487 4 F_IN
port 19 nsew
rlabel metal1 s -11300 28487 -10792 28547 4 F_IN
port 19 nsew
rlabel metal1 s -10852 28547 -10792 28575 4 F_IN
port 19 nsew
rlabel metal1 s -10853 29384 -10793 29413 4 F_IN
port 19 nsew
rlabel metal1 s -10853 29413 -10429 29473 4 F_IN
port 19 nsew
rlabel metal1 s -10853 29473 -10793 29516 4 F_IN
port 19 nsew
rlabel metal1 s -7023 31950 -6972 41862 4 F_IN
port 19 nsew
rlabel metal1 s -11910 31950 -11859 41862 4 F_IN
port 19 nsew
rlabel metal1 s -12088 41742 -11981 41862 4 F_IN
port 19 nsew
rlabel metal1 s -12088 41862 -6972 41913 4 F_IN
port 19 nsew
rlabel metal1 s -12088 41913 -11981 41933 4 F_IN
port 19 nsew
rlabel metal1 s -14142 42120 -13873 43172 4 F_IN
port 19 nsew
rlabel metal1 s -16404 43172 -6583 43467 4 F_IN
port 19 nsew
rlabel metal1 s -12914 46266 -12854 46309 4 F_IN
port 19 nsew
rlabel metal1 s -13278 46309 -12854 46369 4 F_IN
port 19 nsew
rlabel metal1 s -12914 46369 -12854 46398 4 F_IN
port 19 nsew
rlabel metal1 s -12915 47207 -12855 47235 4 F_IN
port 19 nsew
rlabel metal1 s -12915 47235 -12407 47295 4 F_IN
port 19 nsew
rlabel metal1 s -12915 47295 -12855 47344 4 F_IN
port 19 nsew
rlabel metal1 s -6852 48509 -6500 58642 4 F_IN
port 19 nsew
rlabel metal1 s -7809 50353 -7620 50532 4 F_IN
port 19 nsew
rlabel metal1 s -7771 50532 -7696 51948 4 F_IN
port 19 nsew
rlabel metal1 s -7981 51921 -7846 51948 4 F_IN
port 19 nsew
rlabel metal1 s -7981 51948 -7696 52023 4 F_IN
port 19 nsew
rlabel metal1 s -7981 52023 -7846 52053 4 F_IN
port 19 nsew
rlabel metal1 s -8366 54394 -8306 54437 4 F_IN
port 19 nsew
rlabel metal1 s -8366 54437 -7942 54497 4 F_IN
port 19 nsew
rlabel metal1 s -8366 54497 -8306 54526 4 F_IN
port 19 nsew
rlabel metal1 s -8365 55335 -8305 55363 4 F_IN
port 19 nsew
rlabel metal1 s -8813 55363 -8305 55423 4 F_IN
port 19 nsew
rlabel metal1 s -8365 55423 -8305 55472 4 F_IN
port 19 nsew
rlabel metal1 s -14196 58642 -6500 58742 4 F_IN
port 19 nsew
rlabel metal1 s -14196 58742 -6540 58887 4 F_IN
port 19 nsew
rlabel metal1 s -6834 58887 -6540 58922 4 F_IN
port 19 nsew
rlabel metal1 s -6786 59510 -6653 59723 4 F_IN
port 19 nsew
rlabel metal1 s -6746 59723 -6692 60894 4 F_IN
port 19 nsew
rlabel metal1 s -8613 59511 -8350 59770 4 F_IN
port 19 nsew
rlabel metal1 s -7090 60894 -6692 60948 4 F_IN
port 19 nsew
rlabel metal1 s -7090 60948 -7036 61168 4 F_IN
port 19 nsew
rlabel metal1 s -7203 61142 -7145 61168 4 F_IN
port 19 nsew
rlabel metal1 s -7203 61168 -7036 61222 4 F_IN
port 19 nsew
rlabel metal1 s -7203 61222 -7145 61301 4 F_IN
port 19 nsew
rlabel metal1 s -14196 58887 -13951 114640 4 F_IN
port 19 nsew
rlabel locali s 61366 -11971 62272 -11839 8 F_IN
port 19 nsew
rlabel locali s -6611 -11894 -5937 -11839 2 F_IN
port 19 nsew
rlabel locali s -6611 -11839 62272 -11274 8 F_IN
port 19 nsew
rlabel locali s 61366 -11274 62272 -11116 8 F_IN
port 19 nsew
rlabel locali s -6611 -11274 -5937 -11153 2 F_IN
port 19 nsew
rlabel locali s 64673 -4117 64707 -3860 8 F_IN
port 19 nsew
rlabel locali s 64477 -4117 64511 -3860 8 F_IN
port 19 nsew
rlabel locali s 64281 -4117 64315 -3860 8 F_IN
port 19 nsew
rlabel locali s 64085 -4117 64119 -3860 8 F_IN
port 19 nsew
rlabel locali s 63889 -4117 63923 -3860 8 F_IN
port 19 nsew
rlabel locali s 63889 -3860 64707 -3826 8 F_IN
port 19 nsew
rlabel locali s 64673 -3826 64707 -3563 8 F_IN
port 19 nsew
rlabel locali s 64477 -3826 64511 -3563 8 F_IN
port 19 nsew
rlabel locali s 64281 -3826 64315 -3563 8 F_IN
port 19 nsew
rlabel locali s 64085 -3826 64119 -3563 8 F_IN
port 19 nsew
rlabel locali s 63889 -3826 63923 -3563 8 F_IN
port 19 nsew
rlabel locali s -6543 299 -5591 320 4 F_IN
port 19 nsew
rlabel locali s -22512 320 -5591 457 4 F_IN
port 19 nsew
rlabel locali s -6543 457 -5591 465 4 F_IN
port 19 nsew
rlabel locali s -18039 457 -17604 565 4 F_IN
port 19 nsew
rlabel locali s -1304 758 -1270 1015 4 F_IN
port 19 nsew
rlabel locali s -1500 758 -1466 1015 4 F_IN
port 19 nsew
rlabel locali s -1696 758 -1662 1015 4 F_IN
port 19 nsew
rlabel locali s -1892 758 -1858 1015 4 F_IN
port 19 nsew
rlabel locali s -2088 758 -2054 1015 4 F_IN
port 19 nsew
rlabel locali s -2088 1015 -1270 1049 4 F_IN
port 19 nsew
rlabel locali s -1304 1049 -1270 1312 4 F_IN
port 19 nsew
rlabel locali s -1500 1049 -1466 1312 4 F_IN
port 19 nsew
rlabel locali s -1696 1049 -1662 1312 4 F_IN
port 19 nsew
rlabel locali s -1892 1049 -1858 1312 4 F_IN
port 19 nsew
rlabel locali s -2088 1049 -2054 1312 4 F_IN
port 19 nsew
rlabel locali s -16404 8556 -16268 9112 4 F_IN
port 19 nsew
rlabel locali s -7268 9281 -7025 9382 4 F_IN
port 19 nsew
rlabel locali s -16414 9112 -16236 9325 4 F_IN
port 19 nsew
rlabel locali s -6682 13714 -6646 13791 4 F_IN
port 19 nsew
rlabel locali s -7261 9382 -7198 13791 4 F_IN
port 19 nsew
rlabel locali s -7261 13791 -6646 13848 4 F_IN
port 19 nsew
rlabel locali s -6682 13848 -6646 14105 4 F_IN
port 19 nsew
rlabel locali s -6684 14105 -6644 14125 4 F_IN
port 19 nsew
rlabel locali s -6690 14125 -6636 14260 4 F_IN
port 19 nsew
rlabel locali s -7993 26259 -7954 26665 4 F_IN
port 19 nsew
rlabel locali s -8001 26665 -7941 26797 4 F_IN
port 19 nsew
rlabel locali s -8542 26701 -8336 26738 4 F_IN
port 19 nsew
rlabel locali s -8543 26738 -8336 26761 4 F_IN
port 19 nsew
rlabel locali s -8543 26761 -8480 26773 4 F_IN
port 19 nsew
rlabel locali s -7993 26797 -7954 30356 4 F_IN
port 19 nsew
rlabel locali s -8554 26773 -8480 26941 4 F_IN
port 19 nsew
rlabel locali s -10842 26259 -10803 28438 4 F_IN
port 19 nsew
rlabel locali s -11310 28259 -11236 28427 4 F_IN
port 19 nsew
rlabel locali s -10852 28438 -10792 28575 4 F_IN
port 19 nsew
rlabel locali s -11299 28427 -11241 28487 4 F_IN
port 19 nsew
rlabel locali s -11300 28487 -11168 28547 4 F_IN
port 19 nsew
rlabel locali s -10842 28575 -10803 29384 4 F_IN
port 19 nsew
rlabel locali s -10561 29413 -10339 29473 4 F_IN
port 19 nsew
rlabel locali s -10402 29473 -10328 29641 4 F_IN
port 19 nsew
rlabel locali s -10853 29384 -10793 29516 4 F_IN
port 19 nsew
rlabel locali s -7993 30356 -7672 30430 4 F_IN
port 19 nsew
rlabel locali s -7993 30430 -7831 30431 4 F_IN
port 19 nsew
rlabel locali s -7646 30959 -7572 31127 4 F_IN
port 19 nsew
rlabel locali s -7641 31127 -7583 31162 4 F_IN
port 19 nsew
rlabel locali s -7646 31841 -7572 31950 4 F_IN
port 19 nsew
rlabel locali s -7993 30431 -7954 31950 4 F_IN
port 19 nsew
rlabel locali s -7993 31950 -6972 31989 4 F_IN
port 19 nsew
rlabel locali s -10842 29516 -10803 31950 4 F_IN
port 19 nsew
rlabel locali s -11310 31841 -11236 31950 4 F_IN
port 19 nsew
rlabel locali s -11910 31950 -10803 31989 4 F_IN
port 19 nsew
rlabel locali s -7023 31989 -6972 32087 4 F_IN
port 19 nsew
rlabel locali s -7646 31989 -7572 32009 4 F_IN
port 19 nsew
rlabel locali s -11310 31989 -11236 32009 4 F_IN
port 19 nsew
rlabel locali s -11910 31989 -11859 32087 4 F_IN
port 19 nsew
rlabel locali s -12088 41742 -11981 41933 4 F_IN
port 19 nsew
rlabel locali s -12070 41933 -11987 42222 4 F_IN
port 19 nsew
rlabel locali s -14114 42198 -13935 42222 4 F_IN
port 19 nsew
rlabel locali s -14114 42222 -11987 42305 4 F_IN
port 19 nsew
rlabel locali s -14114 42305 -13935 42326 4 F_IN
port 19 nsew
rlabel locali s -6830 43172 -6583 48580 4 F_IN
port 19 nsew
rlabel locali s -12970 43172 -12767 43467 4 F_IN
port 19 nsew
rlabel locali s -16404 9325 -16268 43467 4 F_IN
port 19 nsew
rlabel locali s -12471 43773 -12397 43793 4 F_IN
port 19 nsew
rlabel locali s -12904 43467 -12865 43793 4 F_IN
port 19 nsew
rlabel locali s -12904 43793 -12397 43832 4 F_IN
port 19 nsew
rlabel locali s -12471 43832 -12397 43941 4 F_IN
port 19 nsew
rlabel locali s -12904 43832 -12865 46266 4 F_IN
port 19 nsew
rlabel locali s -12914 46266 -12854 46398 4 F_IN
port 19 nsew
rlabel locali s -13379 46141 -13305 46309 4 F_IN
port 19 nsew
rlabel locali s -13368 46309 -13146 46369 4 F_IN
port 19 nsew
rlabel locali s -12904 46398 -12865 47207 4 F_IN
port 19 nsew
rlabel locali s -12539 47235 -12407 47295 4 F_IN
port 19 nsew
rlabel locali s -12466 47295 -12408 47355 4 F_IN
port 19 nsew
rlabel locali s -12915 47207 -12855 47344 4 F_IN
port 19 nsew
rlabel locali s -12471 47355 -12397 47523 4 F_IN
port 19 nsew
rlabel locali s -6830 48580 -6560 48691 4 F_IN
port 19 nsew
rlabel locali s -6828 48691 -6560 48815 4 F_IN
port 19 nsew
rlabel locali s -12904 47344 -12865 49523 4 F_IN
port 19 nsew
rlabel locali s -6763 50351 -6517 50390 4 F_IN
port 19 nsew
rlabel locali s -7809 50353 -7620 50390 4 F_IN
port 19 nsew
rlabel locali s -7809 50390 -6517 50532 4 F_IN
port 19 nsew
rlabel locali s -6763 50532 -6517 50569 4 F_IN
port 19 nsew
rlabel locali s -8823 51901 -8749 51921 4 F_IN
port 19 nsew
rlabel locali s -8823 51921 -7846 51960 4 F_IN
port 19 nsew
rlabel locali s -8355 51960 -7846 52027 4 F_IN
port 19 nsew
rlabel locali s -7981 52027 -7846 52053 4 F_IN
port 19 nsew
rlabel locali s -7915 54269 -7841 54437 4 F_IN
port 19 nsew
rlabel locali s -8355 52027 -8316 54394 4 F_IN
port 19 nsew
rlabel locali s -8823 51960 -8749 52069 4 F_IN
port 19 nsew
rlabel locali s -8074 54437 -7852 54497 4 F_IN
port 19 nsew
rlabel locali s -8366 54394 -8306 54526 4 F_IN
port 19 nsew
rlabel locali s -8355 54526 -8316 55335 4 F_IN
port 19 nsew
rlabel locali s -8365 55335 -8305 55472 4 F_IN
port 19 nsew
rlabel locali s -8813 55363 -8681 55423 4 F_IN
port 19 nsew
rlabel locali s -8355 55472 -8316 57651 4 F_IN
port 19 nsew
rlabel locali s -8812 55423 -8754 55483 4 F_IN
port 19 nsew
rlabel locali s -8823 55483 -8749 55651 4 F_IN
port 19 nsew
rlabel locali s -6834 58592 -6540 58922 4 F_IN
port 19 nsew
rlabel locali s -6802 58922 -6623 59771 4 F_IN
port 19 nsew
rlabel locali s -8598 58645 -8393 59511 4 F_IN
port 19 nsew
rlabel locali s -14170 59217 -13975 59438 4 F_IN
port 19 nsew
rlabel locali s -8613 59511 -8350 59770 4 F_IN
port 19 nsew
rlabel locali s -8540 59770 -8504 60140 4 F_IN
port 19 nsew
rlabel locali s -8542 60140 -8502 60160 4 F_IN
port 19 nsew
rlabel locali s -8550 60160 -8496 60295 4 F_IN
port 19 nsew
rlabel locali s -7194 60932 -7158 61139 4 F_IN
port 19 nsew
rlabel locali s -7196 61139 -7156 61159 4 F_IN
port 19 nsew
rlabel locali s -7202 61159 -7148 61294 4 F_IN
port 19 nsew
rlabel locali s -14193 67443 -13990 67512 4 F_IN
port 19 nsew
rlabel locali s -14193 67512 -8461 67658 4 F_IN
port 19 nsew
rlabel locali s -8607 67658 -8461 68160 4 F_IN
port 19 nsew
rlabel locali s -14193 67658 -13990 67717 4 F_IN
port 19 nsew
rlabel locali s -8551 68160 -8515 68580 4 F_IN
port 19 nsew
rlabel locali s -8553 68580 -8513 68600 4 F_IN
port 19 nsew
rlabel locali s -8561 68600 -8507 68735 4 F_IN
port 19 nsew
rlabel locali s -14147 76140 -14008 76194 4 F_IN
port 19 nsew
rlabel locali s -14147 76194 -8547 76340 4 F_IN
port 19 nsew
rlabel locali s -8693 76340 -8547 76961 4 F_IN
port 19 nsew
rlabel locali s -14147 76340 -14008 76392 4 F_IN
port 19 nsew
rlabel locali s -8590 76961 -8554 77443 4 F_IN
port 19 nsew
rlabel locali s -8592 77443 -8552 77463 4 F_IN
port 19 nsew
rlabel locali s -8600 77463 -8546 77598 4 F_IN
port 19 nsew
rlabel locali s -14174 85479 -13969 85513 4 F_IN
port 19 nsew
rlabel locali s -14174 85513 -8455 85659 4 F_IN
port 19 nsew
rlabel locali s -8601 85659 -8455 86242 4 F_IN
port 19 nsew
rlabel locali s -14174 85659 -13969 85711 4 F_IN
port 19 nsew
rlabel locali s -8556 86242 -8520 86641 4 F_IN
port 19 nsew
rlabel locali s -8558 86641 -8518 86661 4 F_IN
port 19 nsew
rlabel locali s -8566 86661 -8512 86796 4 F_IN
port 19 nsew
rlabel locali s -14186 93978 -13954 94040 4 F_IN
port 19 nsew
rlabel locali s -14186 94040 -8330 94279 4 F_IN
port 19 nsew
rlabel locali s -8569 94279 -8330 94966 4 F_IN
port 19 nsew
rlabel locali s -14186 94279 -13954 94326 4 F_IN
port 19 nsew
rlabel locali s -8490 94966 -8454 95395 4 F_IN
port 19 nsew
rlabel locali s -8492 95395 -8452 95415 4 F_IN
port 19 nsew
rlabel locali s -8500 95415 -8446 95550 4 F_IN
port 19 nsew
rlabel locali s -14196 103283 -13951 103368 4 F_IN
port 19 nsew
rlabel locali s -14196 103368 -8358 103553 4 F_IN
port 19 nsew
rlabel locali s -8543 103553 -8358 104032 4 F_IN
port 19 nsew
rlabel locali s -14196 103553 -13951 103665 4 F_IN
port 19 nsew
rlabel locali s -8473 104032 -8437 104548 4 F_IN
port 19 nsew
rlabel locali s -8475 104548 -8435 104568 4 F_IN
port 19 nsew
rlabel locali s -8483 104568 -8429 104703 4 F_IN
port 19 nsew
rlabel locali s -14192 112236 -13954 112285 4 F_IN
port 19 nsew
rlabel locali s -14192 112285 -8216 112579 4 F_IN
port 19 nsew
rlabel locali s -8510 112579 -8216 113493 4 F_IN
port 19 nsew
rlabel locali s -14192 112579 -13954 112636 4 F_IN
port 19 nsew
rlabel locali s -8435 113493 -8399 113912 4 F_IN
port 19 nsew
rlabel locali s -8437 113912 -8397 113932 4 F_IN
port 19 nsew
rlabel locali s -8445 113932 -8391 114067 4 F_IN
port 19 nsew
rlabel metal1 s -5986 -26877 -5847 -26876 2 D0
port 20 nsew
rlabel metal1 s -5986 -26876 -5455 -26874 2 D0
port 20 nsew
rlabel metal1 s -7064 -26883 -6925 -26874 2 D0
port 20 nsew
rlabel metal1 s -7064 -26874 -5455 -26848 2 D0
port 20 nsew
rlabel metal1 s -5483 -26848 -5455 -25698 2 D0
port 20 nsew
rlabel metal1 s -7064 -26848 -5847 -26846 2 D0
port 20 nsew
rlabel metal1 s -5986 -26846 -5847 -26823 2 D0
port 20 nsew
rlabel metal1 s -7064 -26846 -6925 -26829 2 D0
port 20 nsew
rlabel metal1 s -5483 -25698 8725 -25647 8 D0
port 20 nsew
rlabel metal1 s 8674 -25647 8725 -20297 8 D0
port 20 nsew
rlabel metal1 s -14282 -22657 -14152 -22507 2 D0
port 20 nsew
rlabel metal1 s -14232 -22507 -14178 -22310 2 D0
port 20 nsew
rlabel metal1 s -15843 -28049 -15667 -22310 2 D0
port 20 nsew
rlabel metal1 s -23937 -28047 -23814 -27924 2 D0
port 20 nsew
rlabel metal1 s -15843 -22310 -14178 -22134 2 D0
port 20 nsew
rlabel metal1 s -14232 -22134 -14178 -21103 2 D0
port 20 nsew
rlabel metal1 s -14375 -21103 -14178 -21049 2 D0
port 20 nsew
rlabel metal1 s -7140 -20297 8725 -20246 8 D0
port 20 nsew
rlabel metal1 s -7140 -20246 -7089 -19864 2 D0
port 20 nsew
rlabel metal1 s -7140 -19864 -7004 -19790 2 D0
port 20 nsew
rlabel metal1 s -23884 -27924 -23823 -19397 2 D0
port 20 nsew
rlabel locali s -32565 -28049 26610 -27913 2 D0
port 20 nsew
rlabel locali s 26474 -27913 26610 -26687 8 D0
port 20 nsew
rlabel locali s 26474 -26687 30209 -26551 8 D0
port 20 nsew
rlabel locali s 30507 -25565 30642 -25557 8 D0
port 20 nsew
rlabel locali s 30487 -25557 30642 -25555 8 D0
port 20 nsew
rlabel locali s 30073 -26551 30209 -25555 8 D0
port 20 nsew
rlabel locali s 30073 -25555 30642 -25519 8 D0
port 20 nsew
rlabel locali s 26839 -25534 26974 -25526 8 D0
port 20 nsew
rlabel locali s 26819 -25526 26974 -25524 8 D0
port 20 nsew
rlabel locali s 26474 -26551 26610 -25524 8 D0
port 20 nsew
rlabel locali s 7852 -27913 7908 -26503 8 D0
port 20 nsew
rlabel locali s -5986 -26877 -5847 -26823 2 D0
port 20 nsew
rlabel locali s -7064 -26883 -6925 -26829 2 D0
port 20 nsew
rlabel locali s 7851 -26503 7909 -25695 8 D0
port 20 nsew
rlabel locali s 7851 -25695 7975 -25652 8 D0
port 20 nsew
rlabel locali s 7852 -25652 7975 -25651 8 D0
port 20 nsew
rlabel locali s 30487 -25519 30642 -25517 8 D0
port 20 nsew
rlabel locali s 30507 -25517 30642 -25511 8 D0
port 20 nsew
rlabel locali s 26291 -25524 26974 -25488 8 D0
port 20 nsew
rlabel locali s 26819 -25488 26974 -25486 8 D0
port 20 nsew
rlabel locali s 26839 -25486 26974 -25480 8 D0
port 20 nsew
rlabel locali s -22055 -25222 -21910 -25166 2 D0
port 20 nsew
rlabel locali s -22055 -25166 -21995 -25161 2 D0
port 20 nsew
rlabel locali s -23884 -25176 -23824 -25161 2 D0
port 20 nsew
rlabel locali s -23884 -25161 -21995 -25120 2 D0
port 20 nsew
rlabel locali s -23884 -25120 -23824 -24939 2 D0
port 20 nsew
rlabel locali s -14108 -22571 -14035 -22565 2 D0
port 20 nsew
rlabel locali s -14282 -22657 -14152 -22565 2 D0
port 20 nsew
rlabel locali s -14282 -22565 -14035 -22524 2 D0
port 20 nsew
rlabel locali s -14108 -22524 -14035 -22511 2 D0
port 20 nsew
rlabel locali s -14282 -22524 -14152 -22507 2 D0
port 20 nsew
rlabel locali s -13734 -21119 -13660 -21093 2 D0
port 20 nsew
rlabel locali s -14372 -21095 -14145 -21093 2 D0
port 20 nsew
rlabel locali s -14372 -21093 -13660 -21055 2 D0
port 20 nsew
rlabel locali s -14146 -21055 -13660 -21054 2 D0
port 20 nsew
rlabel locali s -13734 -21054 -13660 -21048 2 D0
port 20 nsew
rlabel locali s -14146 -21054 -14075 -21053 2 D0
port 20 nsew
rlabel locali s -7140 -19864 -6952 -19790 2 D0
port 20 nsew
rlabel locali s -22291 -19641 -22156 -19634 2 D0
port 20 nsew
rlabel locali s -23884 -19635 -23823 -19634 2 D0
port 20 nsew
rlabel locali s -23884 -19634 -22156 -19600 2 D0
port 20 nsew
rlabel locali s -22291 -19600 -22156 -19587 2 D0
port 20 nsew
rlabel locali s -23884 -19600 -23823 -19397 2 D0
port 20 nsew
rlabel metal1 s 7893 -28241 8016 -28118 8 D1
port 21 nsew
rlabel metal1 s -23746 -28246 -23623 -28123 2 D1
port 21 nsew
rlabel metal1 s 7946 -28118 8007 -27514 8 D1
port 21 nsew
rlabel metal1 s 7951 -26881 8016 -26876 8 D1
port 21 nsew
rlabel metal1 s 7014 -26877 7153 -26876 8 D1
port 21 nsew
rlabel metal1 s 6912 -26876 9523 -26874 8 D1
port 21 nsew
rlabel metal1 s 5936 -26883 6075 -26874 8 D1
port 21 nsew
rlabel metal1 s 5936 -26874 9523 -26848 8 D1
port 21 nsew
rlabel metal1 s 9495 -26848 9523 -19096 8 D1
port 21 nsew
rlabel metal1 s 7951 -26848 8016 -26744 8 D1
port 21 nsew
rlabel metal1 s 5936 -26848 7153 -26846 8 D1
port 21 nsew
rlabel metal1 s 7014 -26846 7153 -26823 8 D1
port 21 nsew
rlabel metal1 s 5936 -26846 6075 -26829 8 D1
port 21 nsew
rlabel metal1 s -23693 -28123 -23632 -19318 2 D1
port 21 nsew
rlabel metal1 s 7014 -19121 7153 -19098 8 D1
port 21 nsew
rlabel metal1 s 5936 -19115 6075 -19098 8 D1
port 21 nsew
rlabel metal1 s 5936 -19098 7153 -19096 8 D1
port 21 nsew
rlabel metal1 s 5936 -19096 9523 -19070 8 D1
port 21 nsew
rlabel metal1 s 6912 -19070 9523 -19068 8 D1
port 21 nsew
rlabel metal1 s 7014 -19068 7153 -19067 8 D1
port 21 nsew
rlabel metal1 s 5936 -19070 6075 -19061 8 D1
port 21 nsew
rlabel locali s -32538 -28248 35050 -28112 8 D1
port 21 nsew
rlabel locali s 34914 -28112 35050 -26698 8 D1
port 21 nsew
rlabel locali s 7954 -27641 8008 -26881 8 D1
port 21 nsew
rlabel locali s 7951 -26881 8016 -26744 8 D1
port 21 nsew
rlabel locali s 7014 -26877 7153 -26823 8 D1
port 21 nsew
rlabel locali s 5936 -26883 6075 -26829 8 D1
port 21 nsew
rlabel locali s 34914 -26698 38649 -26562 8 D1
port 21 nsew
rlabel locali s 38947 -25576 39082 -25568 8 D1
port 21 nsew
rlabel locali s 38927 -25568 39082 -25566 8 D1
port 21 nsew
rlabel locali s 38513 -26562 38649 -25566 8 D1
port 21 nsew
rlabel locali s 38513 -25566 39082 -25530 8 D1
port 21 nsew
rlabel locali s 35279 -25545 35414 -25537 8 D1
port 21 nsew
rlabel locali s 35259 -25537 35414 -25535 8 D1
port 21 nsew
rlabel locali s 34914 -26562 35050 -25535 8 D1
port 21 nsew
rlabel locali s 38927 -25530 39082 -25528 8 D1
port 21 nsew
rlabel locali s 38947 -25528 39082 -25522 8 D1
port 21 nsew
rlabel locali s 34731 -25535 35414 -25499 8 D1
port 21 nsew
rlabel locali s 35259 -25499 35414 -25497 8 D1
port 21 nsew
rlabel locali s 35279 -25497 35414 -25491 8 D1
port 21 nsew
rlabel locali s -22375 -25254 -22230 -25250 2 D1
port 21 nsew
rlabel locali s -23693 -25433 -23633 -25250 2 D1
port 21 nsew
rlabel locali s -23693 -25250 -22230 -25209 2 D1
port 21 nsew
rlabel locali s -22375 -25209 -22230 -25198 2 D1
port 21 nsew
rlabel locali s -23693 -25209 -23633 -25196 2 D1
port 21 nsew
rlabel locali s -22479 -19563 -22344 -19556 2 D1
port 21 nsew
rlabel locali s -23693 -19556 -22344 -19518 2 D1
port 21 nsew
rlabel locali s -22479 -19518 -22344 -19509 2 D1
port 21 nsew
rlabel locali s -23693 -19518 -23632 -19318 2 D1
port 21 nsew
rlabel locali s 7014 -19121 7153 -19067 8 D1
port 21 nsew
rlabel locali s 5936 -19115 6075 -19061 8 D1
port 21 nsew
rlabel metal1 s 7999 -28474 8122 -28351 8 D2
port 22 nsew
rlabel metal1 s -23640 -28479 -23517 -28356 2 D2
port 22 nsew
rlabel metal1 s 8055 -28351 8115 -27518 8 D2
port 22 nsew
rlabel metal1 s 8064 -27518 8108 -27515 8 D2
port 22 nsew
rlabel metal1 s 4014 -26877 4153 -26876 8 D2
port 22 nsew
rlabel metal1 s 4014 -26876 5373 -26874 8 D2
port 22 nsew
rlabel metal1 s 2936 -26883 3075 -26874 8 D2
port 22 nsew
rlabel metal1 s 2936 -26874 5373 -26848 8 D2
port 22 nsew
rlabel metal1 s 7986 -26254 8125 -26250 8 D2
port 22 nsew
rlabel metal1 s 5345 -26848 5373 -26250 8 D2
port 22 nsew
rlabel metal1 s 2936 -26848 4153 -26846 8 D2
port 22 nsew
rlabel metal1 s 4014 -26846 4153 -26823 8 D2
port 22 nsew
rlabel metal1 s 2936 -26846 3075 -26829 8 D2
port 22 nsew
rlabel metal1 s 5345 -26250 9372 -26222 8 D2
port 22 nsew
rlabel metal1 s 9344 -26222 9372 -19722 8 D2
port 22 nsew
rlabel metal1 s 7986 -26222 8125 -26207 8 D2
port 22 nsew
rlabel metal1 s -23584 -28356 -23524 -25536 2 D2
port 22 nsew
rlabel metal1 s -23584 -25536 -23523 -25299 2 D2
port 22 nsew
rlabel metal1 s 5345 -19722 9372 -19694 8 D2
port 22 nsew
rlabel metal1 s 5345 -19694 5373 -19096 8 D2
port 22 nsew
rlabel metal1 s -23584 -25299 -23524 -19470 2 D2
port 22 nsew
rlabel metal1 s -23584 -19470 -23523 -19232 2 D2
port 22 nsew
rlabel metal1 s 4014 -19121 4153 -19098 8 D2
port 22 nsew
rlabel metal1 s 2936 -19115 3075 -19098 8 D2
port 22 nsew
rlabel metal1 s 2936 -19098 4153 -19096 8 D2
port 22 nsew
rlabel metal1 s 2936 -19096 5373 -19070 8 D2
port 22 nsew
rlabel metal1 s 4014 -19070 5373 -19068 8 D2
port 22 nsew
rlabel metal1 s 4014 -19068 4153 -19067 8 D2
port 22 nsew
rlabel metal1 s 2936 -19070 3075 -19061 8 D2
port 22 nsew
rlabel locali s -32538 -28481 43960 -28345 8 D2
port 22 nsew
rlabel locali s 43824 -28345 43960 -26737 8 D2
port 22 nsew
rlabel locali s 43777 -26737 47512 -26601 8 D2
port 22 nsew
rlabel locali s 47810 -25615 47945 -25607 8 D2
port 22 nsew
rlabel locali s 47790 -25607 47945 -25605 8 D2
port 22 nsew
rlabel locali s 47376 -26601 47512 -25605 8 D2
port 22 nsew
rlabel locali s 43777 -26601 43960 -26587 8 D2
port 22 nsew
rlabel locali s 47376 -25605 47945 -25569 8 D2
port 22 nsew
rlabel locali s 44142 -25584 44277 -25576 8 D2
port 22 nsew
rlabel locali s 44122 -25576 44277 -25574 8 D2
port 22 nsew
rlabel locali s 43777 -26587 43913 -25574 8 D2
port 22 nsew
rlabel locali s 8059 -27641 8113 -26253 8 D2
port 22 nsew
rlabel locali s 4014 -26877 4153 -26823 8 D2
port 22 nsew
rlabel locali s 2936 -26883 3075 -26829 8 D2
port 22 nsew
rlabel locali s 7995 -26253 8118 -26209 8 D2
port 22 nsew
rlabel locali s 47790 -25569 47945 -25567 8 D2
port 22 nsew
rlabel locali s 47810 -25567 47945 -25561 8 D2
port 22 nsew
rlabel locali s 43594 -25574 44277 -25538 8 D2
port 22 nsew
rlabel locali s 44122 -25538 44277 -25536 8 D2
port 22 nsew
rlabel locali s 44142 -25536 44277 -25530 8 D2
port 22 nsew
rlabel locali s -22704 -25349 -22559 -25342 2 D2
port 22 nsew
rlabel locali s -23583 -25536 -23523 -25342 2 D2
port 22 nsew
rlabel locali s -23583 -25342 -22559 -25301 2 D2
port 22 nsew
rlabel locali s -22704 -25301 -22559 -25293 2 D2
port 22 nsew
rlabel locali s -23583 -25301 -23523 -25299 2 D2
port 22 nsew
rlabel locali s -22815 -19481 -22680 -19472 2 D2
port 22 nsew
rlabel locali s -22834 -19472 -22680 -19470 2 D2
port 22 nsew
rlabel locali s -23584 -19470 -22680 -19435 2 D2
port 22 nsew
rlabel locali s -22815 -19435 -22680 -19427 2 D2
port 22 nsew
rlabel locali s -23584 -19435 -23523 -19232 2 D2
port 22 nsew
rlabel locali s 4014 -19121 4153 -19067 8 D2
port 22 nsew
rlabel locali s 2936 -19115 3075 -19061 8 D2
port 22 nsew
rlabel metal1 s 8092 -28731 8216 -28608 8 D3
port 23 nsew
rlabel metal1 s -23547 -28736 -23423 -28613 2 D3
port 23 nsew
rlabel metal1 s 8154 -28608 8215 -27661 8 D3
port 23 nsew
rlabel metal1 s -21610 -25946 -21552 -25809 2 D3
port 23 nsew
rlabel metal1 s -21590 -25809 -21555 -24900 2 D3
port 23 nsew
rlabel metal1 s -21590 -24900 -21532 -24763 2 D3
port 23 nsew
rlabel metal1 s 8135 -24637 8280 -24625 8 D3
port 23 nsew
rlabel metal1 s 7024 -24626 7163 -24625 8 D3
port 23 nsew
rlabel metal1 s 7024 -24625 8397 -24623 8 D3
port 23 nsew
rlabel metal1 s 5946 -24632 6085 -24623 8 D3
port 23 nsew
rlabel metal1 s 5946 -24623 8397 -24597 8 D3
port 23 nsew
rlabel metal1 s 8367 -24597 8395 -21362 8 D3
port 23 nsew
rlabel metal1 s 8135 -24597 8280 -24502 8 D3
port 23 nsew
rlabel metal1 s 5946 -24597 7163 -24595 8 D3
port 23 nsew
rlabel metal1 s 7024 -24595 7163 -24572 8 D3
port 23 nsew
rlabel metal1 s 5946 -24595 6085 -24578 8 D3
port 23 nsew
rlabel metal1 s 8354 -21362 8405 -21347 8 D3
port 23 nsew
rlabel metal1 s 7024 -21372 7163 -21349 8 D3
port 23 nsew
rlabel metal1 s 5946 -21366 6085 -21349 8 D3
port 23 nsew
rlabel metal1 s 5946 -21349 7163 -21347 8 D3
port 23 nsew
rlabel metal1 s 5946 -21347 8405 -21321 8 D3
port 23 nsew
rlabel metal1 s 7024 -21321 8405 -21319 8 D3
port 23 nsew
rlabel metal1 s 8354 -21319 8405 -21311 8 D3
port 23 nsew
rlabel metal1 s 7024 -21319 7163 -21318 8 D3
port 23 nsew
rlabel metal1 s 5946 -21321 6085 -21312 8 D3
port 23 nsew
rlabel metal1 s -21068 -20635 -20936 -20631 2 D3
port 23 nsew
rlabel metal1 s -21115 -20631 -20912 -20591 2 D3
port 23 nsew
rlabel metal1 s -21068 -20591 -20912 -20582 2 D3
port 23 nsew
rlabel metal1 s -20952 -20582 -20912 -19809 2 D3
port 23 nsew
rlabel metal1 s -23485 -28613 -23424 -20397 2 D3
port 23 nsew
rlabel metal1 s -20959 -19809 -20822 -19751 2 D3
port 23 nsew
rlabel locali s -32592 -28736 53111 -28600 8 D3
port 23 nsew
rlabel locali s 52975 -28600 53111 -26703 8 D3
port 23 nsew
rlabel locali s 52975 -26703 56710 -26567 8 D3
port 23 nsew
rlabel locali s 57008 -25581 57143 -25573 8 D3
port 23 nsew
rlabel locali s 56988 -25573 57143 -25571 8 D3
port 23 nsew
rlabel locali s 56574 -26567 56710 -25571 8 D3
port 23 nsew
rlabel locali s 56574 -25571 57143 -25535 8 D3
port 23 nsew
rlabel locali s 53340 -25550 53475 -25542 8 D3
port 23 nsew
rlabel locali s 53320 -25542 53475 -25540 8 D3
port 23 nsew
rlabel locali s 52975 -26567 53111 -25540 8 D3
port 23 nsew
rlabel locali s 56988 -25535 57143 -25533 8 D3
port 23 nsew
rlabel locali s 57008 -25533 57143 -25527 8 D3
port 23 nsew
rlabel locali s 52792 -25540 53475 -25504 8 D3
port 23 nsew
rlabel locali s 53320 -25504 53475 -25502 8 D3
port 23 nsew
rlabel locali s 53340 -25502 53475 -25496 8 D3
port 23 nsew
rlabel locali s 8158 -27858 8214 -24637 8 D3
port 23 nsew
rlabel locali s -23485 -25946 -21552 -25905 2 D3
port 23 nsew
rlabel locali s -21610 -25905 -21552 -25809 2 D3
port 23 nsew
rlabel locali s -23485 -25905 -23427 -25809 2 D3
port 23 nsew
rlabel locali s -21183 -24911 -21040 -24894 2 D3
port 23 nsew
rlabel locali s -21590 -24900 -21532 -24894 2 D3
port 23 nsew
rlabel locali s -21590 -24894 -21040 -24858 2 D3
port 23 nsew
rlabel locali s -21183 -24858 -21040 -24851 2 D3
port 23 nsew
rlabel locali s -21590 -24858 -21532 -24763 2 D3
port 23 nsew
rlabel locali s 8135 -24637 8280 -24502 8 D3
port 23 nsew
rlabel locali s 7024 -24626 7163 -24572 8 D3
port 23 nsew
rlabel locali s 5946 -24632 6085 -24578 8 D3
port 23 nsew
rlabel locali s 7024 -21372 7163 -21318 8 D3
port 23 nsew
rlabel locali s 5946 -21366 6085 -21312 8 D3
port 23 nsew
rlabel locali s -21068 -20635 -20936 -20631 2 D3
port 23 nsew
rlabel locali s -23485 -20635 -23425 -20631 2 D3
port 23 nsew
rlabel locali s -23485 -20631 -20936 -20591 2 D3
port 23 nsew
rlabel locali s -21068 -20591 -20936 -20582 2 D3
port 23 nsew
rlabel locali s -23485 -20591 -23425 -20514 2 D3
port 23 nsew
rlabel locali s -23485 -20514 -23417 -20474 2 D3
port 23 nsew
rlabel locali s -23485 -20474 -23425 -20398 2 D3
port 23 nsew
rlabel locali s -20359 -19802 -20285 -19796 2 D3
port 23 nsew
rlabel locali s -20771 -19797 -20700 -19796 2 D3
port 23 nsew
rlabel locali s -20771 -19796 -20285 -19795 2 D3
port 23 nsew
rlabel locali s -20959 -19809 -20822 -19795 2 D3
port 23 nsew
rlabel locali s -20997 -19795 -20285 -19757 2 D3
port 23 nsew
rlabel locali s -20359 -19757 -20285 -19731 2 D3
port 23 nsew
rlabel locali s -20997 -19757 -20770 -19755 2 D3
port 23 nsew
rlabel locali s -20959 -19755 -20822 -19751 2 D3
port 23 nsew
rlabel metal1 s 8199 -29011 8329 -28926 8 D4
port 24 nsew
rlabel metal1 s -23440 -29016 -23310 -28931 2 D4
port 24 nsew
rlabel metal1 s 8198 -28926 8329 -28893 8 D4
port 24 nsew
rlabel metal1 s -23441 -28931 -23310 -28898 2 D4
port 24 nsew
rlabel metal1 s 8198 -28893 8328 -28892 8 D4
port 24 nsew
rlabel metal1 s -23441 -28898 -23311 -28897 2 D4
port 24 nsew
rlabel metal1 s 8267 -28892 8328 -27515 8 D4
port 24 nsew
rlabel metal1 s 1514 -26877 1653 -26876 8 D4
port 24 nsew
rlabel metal1 s 1514 -26876 2052 -26874 8 D4
port 24 nsew
rlabel metal1 s 436 -26883 575 -26874 8 D4
port 24 nsew
rlabel metal1 s 436 -26874 2052 -26848 8 D4
port 24 nsew
rlabel metal1 s 8299 -26115 8443 -26103 8 D4
port 24 nsew
rlabel metal1 s 2024 -26848 2052 -26103 8 D4
port 24 nsew
rlabel metal1 s 436 -26848 1653 -26846 8 D4
port 24 nsew
rlabel metal1 s 1514 -26846 1653 -26823 8 D4
port 24 nsew
rlabel metal1 s 436 -26846 575 -26829 8 D4
port 24 nsew
rlabel metal1 s 2024 -26103 9213 -26075 8 D4
port 24 nsew
rlabel metal1 s 9185 -26075 9213 -19869 8 D4
port 24 nsew
rlabel metal1 s 8299 -26075 8443 -26068 8 D4
port 24 nsew
rlabel metal1 s -21517 -26025 -21459 -25888 2 D4
port 24 nsew
rlabel metal1 s -21516 -25888 -21473 -25071 2 D4
port 24 nsew
rlabel metal1 s -21516 -25071 -21457 -24938 2 D4
port 24 nsew
rlabel metal1 s -21515 -24938 -21457 -24934 2 D4
port 24 nsew
rlabel metal1 s -21084 -20544 -21031 -20412 2 D4
port 24 nsew
rlabel metal1 s 2024 -19869 9213 -19841 8 D4
port 24 nsew
rlabel metal1 s 2024 -19841 2052 -19096 8 D4
port 24 nsew
rlabel metal1 s -21082 -20412 -21046 -19702 2 D4
port 24 nsew
rlabel metal1 s -23372 -28897 -23311 -20330 2 D4
port 24 nsew
rlabel metal1 s -21082 -19702 -20917 -19661 2 D4
port 24 nsew
rlabel metal1 s -21054 -19661 -20917 -19644 2 D4
port 24 nsew
rlabel metal1 s 1514 -19121 1653 -19098 8 D4
port 24 nsew
rlabel metal1 s 436 -19115 575 -19098 8 D4
port 24 nsew
rlabel metal1 s 436 -19098 1653 -19096 8 D4
port 24 nsew
rlabel metal1 s 436 -19096 2052 -19070 8 D4
port 24 nsew
rlabel metal1 s 1514 -19070 2052 -19068 8 D4
port 24 nsew
rlabel metal1 s 1514 -19068 1653 -19067 8 D4
port 24 nsew
rlabel metal1 s 436 -19070 575 -19061 8 D4
port 24 nsew
rlabel locali s -33001 -29027 -22941 -29022 2 D4
port 24 nsew
rlabel locali s -33001 -29022 61865 -28886 8 D4
port 24 nsew
rlabel locali s 61729 -28886 61865 -26637 8 D4
port 24 nsew
rlabel locali s 8289 -28886 8425 -28884 8 D4
port 24 nsew
rlabel locali s 61729 -26637 65464 -26501 8 D4
port 24 nsew
rlabel locali s 65762 -25515 65897 -25507 8 D4
port 24 nsew
rlabel locali s 65742 -25507 65897 -25505 8 D4
port 24 nsew
rlabel locali s 65328 -26501 65464 -25505 8 D4
port 24 nsew
rlabel locali s 65328 -25505 65897 -25469 8 D4
port 24 nsew
rlabel locali s 62094 -25484 62229 -25476 8 D4
port 24 nsew
rlabel locali s 62074 -25476 62229 -25474 8 D4
port 24 nsew
rlabel locali s 61729 -26501 61865 -25474 8 D4
port 24 nsew
rlabel locali s 8270 -27641 8324 -26110 8 D4
port 24 nsew
rlabel locali s 1514 -26877 1653 -26823 8 D4
port 24 nsew
rlabel locali s 436 -26883 575 -26829 8 D4
port 24 nsew
rlabel locali s 8270 -26110 8427 -26070 8 D4
port 24 nsew
rlabel locali s -23372 -26118 -23314 -26025 2 D4
port 24 nsew
rlabel locali s -23372 -26025 -21459 -25984 2 D4
port 24 nsew
rlabel locali s -21517 -25984 -21459 -25888 2 D4
port 24 nsew
rlabel locali s -23372 -25984 -23314 -25981 2 D4
port 24 nsew
rlabel locali s 65742 -25469 65897 -25467 8 D4
port 24 nsew
rlabel locali s 65762 -25467 65897 -25461 8 D4
port 24 nsew
rlabel locali s 61546 -25474 62229 -25438 8 D4
port 24 nsew
rlabel locali s 62074 -25438 62229 -25436 8 D4
port 24 nsew
rlabel locali s 62094 -25436 62229 -25430 8 D4
port 24 nsew
rlabel locali s -21406 -24991 -21260 -24983 2 D4
port 24 nsew
rlabel locali s -21515 -25071 -21457 -24983 2 D4
port 24 nsew
rlabel locali s -21515 -24983 -21260 -24947 2 D4
port 24 nsew
rlabel locali s -21406 -24947 -21260 -24931 2 D4
port 24 nsew
rlabel locali s -21515 -24947 -21457 -24934 2 D4
port 24 nsew
rlabel locali s -23372 -20546 -23311 -20544 2 D4
port 24 nsew
rlabel locali s -23372 -20544 -21031 -20508 2 D4
port 24 nsew
rlabel locali s -21084 -20508 -21031 -20412 2 D4
port 24 nsew
rlabel locali s -23372 -20508 -23311 -20330 2 D4
port 24 nsew
rlabel locali s -20824 -19707 -20689 -19699 2 D4
port 24 nsew
rlabel locali s -20844 -19699 -20689 -19697 2 D4
port 24 nsew
rlabel locali s -21054 -19702 -20917 -19697 2 D4
port 24 nsew
rlabel locali s -21054 -19697 -20689 -19661 2 D4
port 24 nsew
rlabel locali s -20844 -19661 -20689 -19659 2 D4
port 24 nsew
rlabel locali s -20824 -19659 -20689 -19653 2 D4
port 24 nsew
rlabel locali s -21054 -19661 -20917 -19644 2 D4
port 24 nsew
rlabel locali s 1514 -19121 1653 -19067 8 D4
port 24 nsew
rlabel locali s 436 -19115 575 -19061 8 D4
port 24 nsew
rlabel metal1 s 8358 -29316 8481 -29193 8 D5
port 25 nsew
rlabel metal1 s -23281 -29321 -23158 -29198 2 D5
port 25 nsew
rlabel metal1 s 8358 -29193 8445 -29192 8 D5
port 25 nsew
rlabel metal1 s -23281 -29198 -23194 -29197 2 D5
port 25 nsew
rlabel metal1 s 8379 -29192 8445 -29020 8 D5
port 25 nsew
rlabel metal1 s -23260 -29197 -23194 -29025 2 D5
port 25 nsew
rlabel metal1 s 8381 -29020 8445 -27511 8 D5
port 25 nsew
rlabel metal1 s -986 -26877 -847 -26876 2 D5
port 25 nsew
rlabel metal1 s -986 -26876 -414 -26874 2 D5
port 25 nsew
rlabel metal1 s -2064 -26883 -1925 -26874 2 D5
port 25 nsew
rlabel metal1 s -2064 -26874 -414 -26848 2 D5
port 25 nsew
rlabel metal1 s 8425 -25984 8568 -25983 8 D5
port 25 nsew
rlabel metal1 s -442 -26848 -414 -25983 2 D5
port 25 nsew
rlabel metal1 s -2064 -26848 -847 -26846 2 D5
port 25 nsew
rlabel metal1 s -986 -26846 -847 -26823 2 D5
port 25 nsew
rlabel metal1 s -2064 -26846 -1925 -26829 2 D5
port 25 nsew
rlabel metal1 s -442 -25983 9051 -25955 8 D5
port 25 nsew
rlabel metal1 s -20696 -26104 -20638 -25967 2 D5
port 25 nsew
rlabel metal1 s 9023 -25955 9051 -19989 8 D5
port 25 nsew
rlabel metal1 s 8425 -25955 8568 -25937 8 D5
port 25 nsew
rlabel metal1 s -20674 -25967 -20639 -24901 2 D5
port 25 nsew
rlabel metal1 s -20674 -24901 -20616 -24764 2 D5
port 25 nsew
rlabel metal1 s -23258 -29025 -23194 -21802 2 D5
port 25 nsew
rlabel metal1 s -442 -19989 9051 -19961 8 D5
port 25 nsew
rlabel metal1 s -442 -19961 -414 -19096 2 D5
port 25 nsew
rlabel metal1 s -986 -19121 -847 -19098 2 D5
port 25 nsew
rlabel metal1 s -2064 -19115 -1925 -19098 2 D5
port 25 nsew
rlabel metal1 s -2064 -19098 -847 -19096 2 D5
port 25 nsew
rlabel metal1 s -2064 -19096 -414 -19070 2 D5
port 25 nsew
rlabel metal1 s -986 -19070 -414 -19068 2 D5
port 25 nsew
rlabel metal1 s -986 -19068 -847 -19067 2 D5
port 25 nsew
rlabel metal1 s -2064 -19070 -1925 -19061 2 D5
port 25 nsew
rlabel locali s -32755 -29321 71018 -29185 8 D5
port 25 nsew
rlabel locali s 70882 -29185 71018 -26620 8 D5
port 25 nsew
rlabel locali s 70882 -26620 74617 -26484 8 D5
port 25 nsew
rlabel locali s 74915 -25498 75050 -25490 8 D5
port 25 nsew
rlabel locali s 74895 -25490 75050 -25488 8 D5
port 25 nsew
rlabel locali s 74481 -26484 74617 -25488 8 D5
port 25 nsew
rlabel locali s 74481 -25488 75050 -25452 8 D5
port 25 nsew
rlabel locali s 71247 -25467 71382 -25459 8 D5
port 25 nsew
rlabel locali s 71227 -25459 71382 -25457 8 D5
port 25 nsew
rlabel locali s 70882 -26484 71018 -25457 8 D5
port 25 nsew
rlabel locali s 8385 -27641 8439 -26468 8 D5
port 25 nsew
rlabel locali s -986 -26877 -847 -26823 2 D5
port 25 nsew
rlabel locali s -2064 -26883 -1925 -26829 2 D5
port 25 nsew
rlabel locali s 8385 -26468 8538 -26414 8 D5
port 25 nsew
rlabel locali s 8484 -26414 8538 -25983 8 D5
port 25 nsew
rlabel locali s -23258 -26199 -23200 -26104 2 D5
port 25 nsew
rlabel locali s -23258 -26104 -20638 -26063 2 D5
port 25 nsew
rlabel locali s 8429 -25983 8552 -25939 8 D5
port 25 nsew
rlabel locali s -20696 -26063 -20638 -25967 2 D5
port 25 nsew
rlabel locali s -23258 -26063 -23200 -26062 2 D5
port 25 nsew
rlabel locali s 74895 -25452 75050 -25450 8 D5
port 25 nsew
rlabel locali s 74915 -25450 75050 -25444 8 D5
port 25 nsew
rlabel locali s 70699 -25457 71382 -25421 8 D5
port 25 nsew
rlabel locali s 71227 -25421 71382 -25419 8 D5
port 25 nsew
rlabel locali s 71247 -25419 71382 -25413 8 D5
port 25 nsew
rlabel locali s -20278 -24912 -20135 -24895 2 D5
port 25 nsew
rlabel locali s -20674 -24901 -20616 -24895 2 D5
port 25 nsew
rlabel locali s -20674 -24895 -20135 -24859 2 D5
port 25 nsew
rlabel locali s -20278 -24859 -20135 -24852 2 D5
port 25 nsew
rlabel locali s -20674 -24859 -20616 -24764 2 D5
port 25 nsew
rlabel locali s -23256 -22046 -23196 -21809 2 D5
port 25 nsew
rlabel locali s -22301 -21711 -22227 -21705 2 D5
port 25 nsew
rlabel locali s -22713 -21706 -22642 -21705 2 D5
port 25 nsew
rlabel locali s -22713 -21705 -22227 -21704 2 D5
port 25 nsew
rlabel locali s -23239 -21809 -23199 -21704 2 D5
port 25 nsew
rlabel locali s -23239 -21704 -22227 -21666 2 D5
port 25 nsew
rlabel locali s -22301 -21666 -22227 -21640 2 D5
port 25 nsew
rlabel locali s -23239 -21666 -22712 -21664 2 D5
port 25 nsew
rlabel locali s -986 -19121 -847 -19067 2 D5
port 25 nsew
rlabel locali s -2064 -19115 -1925 -19061 2 D5
port 25 nsew
rlabel metal1 s 8509 -29683 8632 -29560 8 D6
port 26 nsew
rlabel metal1 s -23130 -29688 -23007 -29565 2 D6
port 26 nsew
rlabel metal1 s 8526 -29560 8586 -27475 8 D6
port 26 nsew
rlabel metal1 s -3486 -26877 -3347 -26876 2 D6
port 26 nsew
rlabel metal1 s -3486 -26876 -2898 -26874 2 D6
port 26 nsew
rlabel metal1 s -4564 -26883 -4425 -26874 2 D6
port 26 nsew
rlabel metal1 s -4564 -26874 -2898 -26848 2 D6
port 26 nsew
rlabel metal1 s 8585 -25848 8733 -25844 8 D6
port 26 nsew
rlabel metal1 s -2926 -26848 -2898 -25844 2 D6
port 26 nsew
rlabel metal1 s -4564 -26848 -3347 -26846 2 D6
port 26 nsew
rlabel metal1 s -3486 -26846 -3347 -26823 2 D6
port 26 nsew
rlabel metal1 s -4564 -26846 -4425 -26829 2 D6
port 26 nsew
rlabel metal1 s -20603 -26181 -20545 -26044 2 D6
port 26 nsew
rlabel metal1 s -2926 -25844 8892 -25808 8 D6
port 26 nsew
rlabel metal1 s 8856 -25808 8892 -20136 8 D6
port 26 nsew
rlabel metal1 s 8585 -25808 8733 -25800 8 D6
port 26 nsew
rlabel metal1 s -20597 -26044 -20562 -25073 2 D6
port 26 nsew
rlabel metal1 s -20597 -25073 -20539 -24936 2 D6
port 26 nsew
rlabel metal1 s -23113 -29565 -23053 -21371 2 D6
port 26 nsew
rlabel metal1 s -2926 -20136 8892 -20100 8 D6
port 26 nsew
rlabel metal1 s -2926 -20100 -2898 -19096 2 D6
port 26 nsew
rlabel metal1 s -3486 -19121 -3347 -19098 2 D6
port 26 nsew
rlabel metal1 s -4564 -19115 -4425 -19098 2 D6
port 26 nsew
rlabel metal1 s -4564 -19098 -3347 -19096 2 D6
port 26 nsew
rlabel metal1 s -4564 -19096 -2898 -19070 2 D6
port 26 nsew
rlabel metal1 s -3486 -19070 -2898 -19068 2 D6
port 26 nsew
rlabel metal1 s -3486 -19068 -3347 -19067 2 D6
port 26 nsew
rlabel metal1 s -4564 -19070 -4425 -19061 2 D6
port 26 nsew
rlabel locali s -32917 -29691 80406 -29555 8 D6
port 26 nsew
rlabel locali s 80270 -29555 80406 -26582 8 D6
port 26 nsew
rlabel locali s 8529 -27641 8583 -27600 8 D6
port 26 nsew
rlabel locali s 8529 -27600 8681 -27546 8 D6
port 26 nsew
rlabel locali s 80246 -26582 83981 -26446 8 D6
port 26 nsew
rlabel locali s 84279 -25460 84414 -25452 8 D6
port 26 nsew
rlabel locali s 84259 -25452 84414 -25450 8 D6
port 26 nsew
rlabel locali s 83845 -26446 83981 -25450 8 D6
port 26 nsew
rlabel locali s 83845 -25450 84414 -25414 8 D6
port 26 nsew
rlabel locali s 80611 -25429 80746 -25421 8 D6
port 26 nsew
rlabel locali s 80591 -25421 80746 -25419 8 D6
port 26 nsew
rlabel locali s 80246 -26446 80382 -25419 8 D6
port 26 nsew
rlabel locali s 8627 -27546 8681 -25848 8 D6
port 26 nsew
rlabel locali s 8529 -27546 8583 -27516 8 D6
port 26 nsew
rlabel locali s -3486 -26877 -3347 -26823 2 D6
port 26 nsew
rlabel locali s -4564 -26883 -4425 -26829 2 D6
port 26 nsew
rlabel locali s -23113 -26277 -23055 -26181 2 D6
port 26 nsew
rlabel locali s -23113 -26181 -20545 -26140 2 D6
port 26 nsew
rlabel locali s -20603 -26140 -20545 -26044 2 D6
port 26 nsew
rlabel locali s 8585 -25848 8733 -25800 8 D6
port 26 nsew
rlabel locali s 84259 -25414 84414 -25412 8 D6
port 26 nsew
rlabel locali s 84279 -25412 84414 -25406 8 D6
port 26 nsew
rlabel locali s 80063 -25419 80746 -25383 8 D6
port 26 nsew
rlabel locali s 80591 -25383 80746 -25381 8 D6
port 26 nsew
rlabel locali s 80611 -25381 80746 -25375 8 D6
port 26 nsew
rlabel locali s -20501 -24992 -20355 -24984 2 D6
port 26 nsew
rlabel locali s -20597 -25073 -20539 -24984 2 D6
port 26 nsew
rlabel locali s -20597 -24984 -20355 -24948 2 D6
port 26 nsew
rlabel locali s -20501 -24948 -20355 -24932 2 D6
port 26 nsew
rlabel locali s -20597 -24948 -20539 -24936 2 D6
port 26 nsew
rlabel locali s -22766 -21616 -22631 -21608 2 D6
port 26 nsew
rlabel locali s -22786 -21608 -22631 -21606 2 D6
port 26 nsew
rlabel locali s -23113 -21608 -23053 -21606 2 D6
port 26 nsew
rlabel locali s -23113 -21606 -22631 -21570 2 D6
port 26 nsew
rlabel locali s -22786 -21570 -22631 -21568 2 D6
port 26 nsew
rlabel locali s -22766 -21568 -22631 -21562 2 D6
port 26 nsew
rlabel locali s -23113 -21570 -23053 -21371 2 D6
port 26 nsew
rlabel locali s -3486 -19121 -3347 -19067 2 D6
port 26 nsew
rlabel locali s -4564 -19115 -4425 -19061 2 D6
port 26 nsew
rlabel metal1 s -14516 9376 -14393 9429 4 D7
port 27 nsew
rlabel metal1 s -14516 9429 -5866 9490 4 D7
port 27 nsew
rlabel metal1 s -14516 9490 -14393 9499 4 D7
port 27 nsew
rlabel metal1 s -14518 17470 -8603 17646 4 D7
port 27 nsew
rlabel metal1 s -7572 18938 -7518 19081 4 D7
port 27 nsew
rlabel metal1 s -8779 17646 -8603 19081 4 D7
port 27 nsew
rlabel metal1 s -9126 19031 -8976 19081 4 D7
port 27 nsew
rlabel metal1 s -9126 19081 -7518 19135 4 D7
port 27 nsew
rlabel metal1 s -9126 19135 -8976 19161 4 D7
port 27 nsew
rlabel metal1 s -6766 26173 -6259 26224 4 D7
port 27 nsew
rlabel metal1 s -6333 26224 -6259 26309 4 D7
port 27 nsew
rlabel metal1 s -6766 26224 -6715 41987 4 D7
port 27 nsew
rlabel metal1 s -13352 26249 -13298 26388 4 D7
port 27 nsew
rlabel metal1 s -13343 26388 -13315 27327 4 D7
port 27 nsew
rlabel metal1 s -13346 27327 -13292 27466 4 D7
port 27 nsew
rlabel metal1 s -13345 27466 -13317 27830 4 D7
port 27 nsew
rlabel metal1 s -13345 27830 -12116 27858 4 D7
port 27 nsew
rlabel metal1 s -12167 27858 -12116 41987 4 D7
port 27 nsew
rlabel metal1 s -12167 41987 -6715 42038 4 D7
port 27 nsew
rlabel locali s -20516 4336 -14382 4472 4 D7
port 27 nsew
rlabel locali s -6104 9429 -5866 9490 4 D7
port 27 nsew
rlabel locali s -11645 9429 -11408 9489 4 D7
port 27 nsew
rlabel locali s -6103 9490 -6069 11022 4 D7
port 27 nsew
rlabel locali s -6110 11022 -6056 11157 4 D7
port 27 nsew
rlabel locali s -11630 9489 -11589 11258 4 D7
port 27 nsew
rlabel locali s -11691 11258 -11589 11318 4 D7
port 27 nsew
rlabel locali s -11691 11318 -11635 11403 4 D7
port 27 nsew
rlabel locali s -7564 18941 -7524 19167 4 D7
port 27 nsew
rlabel locali s -9126 19031 -8976 19161 4 D7
port 27 nsew
rlabel locali s -7564 19167 -7522 19168 4 D7
port 27 nsew
rlabel locali s -7562 19168 -7522 19238 4 D7
port 27 nsew
rlabel locali s -9034 19161 -8993 19205 4 D7
port 27 nsew
rlabel locali s -7562 19238 -7523 19579 4 D7
port 27 nsew
rlabel locali s -9040 19205 -8980 19278 4 D7
port 27 nsew
rlabel locali s -7588 19579 -7517 19653 4 D7
port 27 nsew
rlabel locali s -6333 26173 -6259 26361 4 D7
port 27 nsew
rlabel locali s -13352 26249 -13298 26388 4 D7
port 27 nsew
rlabel locali s -13346 27327 -13292 27466 4 D7
port 27 nsew
rlabel locali s -12972 41164 -12121 41165 4 D7
port 27 nsew
rlabel locali s -14518 4472 -14382 41165 4 D7
port 27 nsew
rlabel locali s -14518 41165 -12120 41221 4 D7
port 27 nsew
rlabel locali s -12972 41221 -12120 41222 4 D7
port 27 nsew
rlabel locali s -12164 41222 -12120 41288 4 D7
port 27 nsew
rlabel locali s -11993 59604 -11957 59787 4 D7
port 27 nsew
rlabel locali s -14518 41221 -14382 59787 4 D7
port 27 nsew
rlabel locali s -14518 59787 -11957 59923 4 D7
port 27 nsew
rlabel locali s -11993 59923 -11957 60132 4 D7
port 27 nsew
rlabel locali s -11995 60132 -11955 60152 4 D7
port 27 nsew
rlabel locali s -12003 60152 -11949 60287 4 D7
port 27 nsew
rlabel locali s -13156 59923 -13020 63386 4 D7
port 27 nsew
rlabel locali s -13156 63386 -11988 63522 4 D7
port 27 nsew
rlabel locali s -12024 63522 -11988 63800 4 D7
port 27 nsew
rlabel locali s -12026 63800 -11986 63820 4 D7
port 27 nsew
rlabel locali s -12034 63820 -11980 63955 4 D7
port 27 nsew
rlabel metal1 s -14715 9567 -14592 9620 4 D8
port 28 nsew
rlabel metal1 s -14715 9620 -5787 9681 4 D8
port 28 nsew
rlabel metal1 s -14715 9681 -14592 9690 4 D8
port 28 nsew
rlabel metal1 s -5584 39249 -5530 39388 4 D8
port 28 nsew
rlabel metal1 s -13352 39249 -13298 39388 4 D8
port 28 nsew
rlabel metal1 s -5567 39388 -5539 40225 4 D8
port 28 nsew
rlabel metal1 s -5567 40225 -5537 40327 4 D8
port 28 nsew
rlabel metal1 s -13343 39388 -13315 40225 4 D8
port 28 nsew
rlabel metal1 s -13345 40225 -13315 40327 4 D8
port 28 nsew
rlabel metal1 s -5590 40327 -5536 40466 4 D8
port 28 nsew
rlabel metal1 s -13346 40327 -13292 40466 4 D8
port 28 nsew
rlabel metal1 s -5565 40466 -5537 42808 4 D8
port 28 nsew
rlabel metal1 s -13345 40466 -13317 41264 4 D8
port 28 nsew
rlabel metal1 s -14710 41206 -14587 41259 4 D8
port 28 nsew
rlabel metal1 s -13350 41264 -13213 41329 4 D8
port 28 nsew
rlabel metal1 s -14710 41259 -13983 41320 4 D8
port 28 nsew
rlabel metal1 s -14710 41320 -14587 41329 4 D8
port 28 nsew
rlabel metal1 s -13345 41329 -13317 42808 4 D8
port 28 nsew
rlabel metal1 s -13345 42808 -5537 42836 4 D8
port 28 nsew
rlabel locali s -14717 5310 -14581 5353 4 D8
port 28 nsew
rlabel locali s -19980 5353 -14581 5489 4 D8
port 28 nsew
rlabel locali s -6025 9620 -5787 9681 4 D8
port 28 nsew
rlabel locali s -11902 9620 -11665 9680 4 D8
port 28 nsew
rlabel locali s -6025 9681 -5987 10834 4 D8
port 28 nsew
rlabel locali s -6032 10834 -5978 10969 4 D8
port 28 nsew
rlabel locali s -11719 9680 -11678 10938 4 D8
port 28 nsew
rlabel locali s -11723 10938 -11667 11083 4 D8
port 28 nsew
rlabel locali s -5584 39249 -5530 39388 4 D8
port 28 nsew
rlabel locali s -13352 39249 -13298 39388 4 D8
port 28 nsew
rlabel locali s -5590 40327 -5536 40466 4 D8
port 28 nsew
rlabel locali s -13346 40327 -13292 40466 4 D8
port 28 nsew
rlabel locali s -13350 41264 -13213 41267 4 D8
port 28 nsew
rlabel locali s -14110 41267 -13213 41321 4 D8
port 28 nsew
rlabel locali s -13350 41321 -13213 41329 4 D8
port 28 nsew
rlabel locali s -12004 68044 -11968 68227 4 D8
port 28 nsew
rlabel locali s -14717 5489 -14581 68227 4 D8
port 28 nsew
rlabel locali s -14717 68227 -11968 68363 4 D8
port 28 nsew
rlabel locali s -12004 68363 -11968 68572 4 D8
port 28 nsew
rlabel locali s -12006 68572 -11966 68592 4 D8
port 28 nsew
rlabel locali s -12014 68592 -11960 68727 4 D8
port 28 nsew
rlabel locali s -13167 68363 -13031 71826 4 D8
port 28 nsew
rlabel locali s -13167 71826 -11999 71962 4 D8
port 28 nsew
rlabel locali s -12035 71962 -11999 72240 4 D8
port 28 nsew
rlabel locali s -12037 72240 -11997 72260 4 D8
port 28 nsew
rlabel locali s -12045 72260 -11991 72395 4 D8
port 28 nsew
rlabel metal1 s -14948 9673 -14825 9729 4 D9
port 29 nsew
rlabel metal1 s -14948 9729 -5701 9789 4 D9
port 29 nsew
rlabel metal1 s -5939 9789 -5701 9790 4 D9
port 29 nsew
rlabel metal1 s -12005 9789 -11768 9790 4 D9
port 29 nsew
rlabel metal1 s -14948 9789 -14825 9796 4 D9
port 29 nsew
rlabel metal1 s -5584 36249 -5530 36388 4 D9
port 29 nsew
rlabel metal1 s -13352 36249 -13298 36388 4 D9
port 29 nsew
rlabel metal1 s -5567 36388 -5539 37327 4 D9
port 29 nsew
rlabel metal1 s -13343 36388 -13315 37327 4 D9
port 29 nsew
rlabel metal1 s -5590 37327 -5536 37466 4 D9
port 29 nsew
rlabel metal1 s -13346 37327 -13292 37466 4 D9
port 29 nsew
rlabel metal1 s -5565 37466 -5537 38658 4 D9
port 29 nsew
rlabel metal1 s -13345 37466 -13317 38658 4 D9
port 29 nsew
rlabel metal1 s -6191 38658 -5537 38686 4 D9
port 29 nsew
rlabel metal1 s -6191 38686 -6163 42657 4 D9
port 29 nsew
rlabel metal1 s -13345 38658 -12691 38686 4 D9
port 29 nsew
rlabel metal1 s -12719 38686 -12691 41299 4 D9
port 29 nsew
rlabel metal1 s -12723 41299 -12676 41438 4 D9
port 29 nsew
rlabel metal1 s -14943 41312 -14820 41368 4 D9
port 29 nsew
rlabel metal1 s -14943 41368 -13987 41377 4 D9
port 29 nsew
rlabel metal1 s -14943 41377 -13984 41421 4 D9
port 29 nsew
rlabel metal1 s -14943 41421 -13987 41428 4 D9
port 29 nsew
rlabel metal1 s -14943 41428 -14820 41435 4 D9
port 29 nsew
rlabel metal1 s -12719 41438 -12691 42657 4 D9
port 29 nsew
rlabel metal1 s -12719 42657 -6163 42685 4 D9
port 29 nsew
rlabel locali s -19851 7017 -14814 7153 4 D9
port 29 nsew
rlabel locali s -5939 9729 -5701 9790 4 D9
port 29 nsew
rlabel locali s -12005 9730 -11768 9790 4 D9
port 29 nsew
rlabel locali s -5939 9790 -5904 10479 4 D9
port 29 nsew
rlabel locali s -5941 10479 -5904 10498 4 D9
port 29 nsew
rlabel locali s -5950 10498 -5896 10633 4 D9
port 29 nsew
rlabel locali s -11811 9790 -11770 10609 4 D9
port 29 nsew
rlabel locali s -11818 10609 -11762 10754 4 D9
port 29 nsew
rlabel locali s -5584 36249 -5530 36388 4 D9
port 29 nsew
rlabel locali s -13352 36249 -13298 36388 4 D9
port 29 nsew
rlabel locali s -5590 37327 -5536 37466 4 D9
port 29 nsew
rlabel locali s -13346 37327 -13292 37466 4 D9
port 29 nsew
rlabel locali s -12722 41308 -12678 41372 4 D9
port 29 nsew
rlabel locali s -14110 41372 -12678 41426 4 D9
port 29 nsew
rlabel locali s -12722 41426 -12678 41431 4 D9
port 29 nsew
rlabel locali s -12043 76907 -12007 77090 4 D9
port 29 nsew
rlabel locali s -13206 77090 -12007 77137 4 D9
port 29 nsew
rlabel locali s -14950 7153 -14814 77137 4 D9
port 29 nsew
rlabel locali s -14950 77137 -12007 77226 4 D9
port 29 nsew
rlabel locali s -12043 77226 -12007 77435 4 D9
port 29 nsew
rlabel locali s -14950 77226 -13056 77273 4 D9
port 29 nsew
rlabel locali s -12045 77435 -12005 77455 4 D9
port 29 nsew
rlabel locali s -12053 77455 -11999 77590 4 D9
port 29 nsew
rlabel locali s -13206 77273 -13070 80689 4 D9
port 29 nsew
rlabel locali s -13206 80689 -12038 80825 4 D9
port 29 nsew
rlabel locali s -12074 80825 -12038 81103 4 D9
port 29 nsew
rlabel locali s -12076 81103 -12036 81123 4 D9
port 29 nsew
rlabel locali s -12084 81123 -12030 81258 4 D9
port 29 nsew
rlabel metal1 s -15205 9766 -15082 9828 4 D10
port 30 nsew
rlabel metal1 s -15205 9828 -6866 9889 4 D10
port 30 nsew
rlabel metal1 s -15205 9889 -15082 9890 4 D10
port 30 nsew
rlabel metal1 s -12415 11703 -12278 11723 4 D10
port 30 nsew
rlabel metal1 s -12415 11723 -11232 11758 4 D10
port 30 nsew
rlabel metal1 s -11369 11758 -11232 11781 4 D10
port 30 nsew
rlabel metal1 s -12415 11758 -12278 11761 4 D10
port 30 nsew
rlabel metal1 s -7100 12198 -7060 12245 4 D10
port 30 nsew
rlabel metal1 s -6278 12354 -6220 12361 4 D10
port 30 nsew
rlabel metal1 s -7104 12245 -7051 12361 4 D10
port 30 nsew
rlabel metal1 s -7104 12361 -6220 12377 4 D10
port 30 nsew
rlabel metal1 s -7100 12377 -6220 12401 4 D10
port 30 nsew
rlabel metal1 s -6278 12401 -6220 12491 4 D10
port 30 nsew
rlabel metal1 s -7835 39259 -7781 39398 4 D10
port 30 nsew
rlabel metal1 s -11101 39259 -11047 39398 4 D10
port 30 nsew
rlabel metal1 s -7818 39398 -7790 40337 4 D10
port 30 nsew
rlabel metal1 s -11092 39398 -11064 40337 4 D10
port 30 nsew
rlabel metal1 s -7841 40337 -7787 40476 4 D10
port 30 nsew
rlabel metal1 s -11095 40337 -11041 40476 4 D10
port 30 nsew
rlabel metal1 s -7816 40476 -7788 41667 4 D10
port 30 nsew
rlabel metal1 s -11094 40476 -11066 41448 4 D10
port 30 nsew
rlabel metal1 s -11106 41448 -10971 41593 4 D10
port 30 nsew
rlabel metal1 s -15200 41405 -15077 41467 4 D10
port 30 nsew
rlabel metal1 s -15200 41467 -14130 41528 4 D10
port 30 nsew
rlabel metal1 s -15200 41528 -15077 41529 4 D10
port 30 nsew
rlabel metal1 s -7831 41667 -7780 41680 4 D10
port 30 nsew
rlabel metal1 s -11094 41593 -11066 41680 4 D10
port 30 nsew
rlabel metal1 s -11094 41680 -7780 41708 4 D10
port 30 nsew
rlabel metal1 s -7831 41708 -7780 41718 4 D10
port 30 nsew
rlabel metal1 s -11094 41708 -11066 41710 4 D10
port 30 nsew
rlabel locali s -19000 7720 -15069 7856 4 D10
port 30 nsew
rlabel locali s -7104 9828 -6867 9888 4 D10
port 30 nsew
rlabel locali s -12415 9828 -12278 9886 4 D10
port 30 nsew
rlabel locali s -6983 9888 -6943 9896 4 D10
port 30 nsew
rlabel locali s -7100 9888 -7060 12245 4 D10
port 30 nsew
rlabel locali s -12415 9886 -12374 11703 4 D10
port 30 nsew
rlabel locali s -11369 11723 -11232 11781 4 D10
port 30 nsew
rlabel locali s -12415 11703 -12278 11761 4 D10
port 30 nsew
rlabel locali s -11363 11781 -11327 12130 4 D10
port 30 nsew
rlabel locali s -6264 12316 -6224 12354 4 D10
port 30 nsew
rlabel locali s -6278 12354 -6220 12491 4 D10
port 30 nsew
rlabel locali s -7104 12245 -7051 12377 4 D10
port 30 nsew
rlabel locali s -11380 12130 -11320 12273 4 D10
port 30 nsew
rlabel locali s -6264 12491 -6224 12542 4 D10
port 30 nsew
rlabel locali s -6266 12542 -6224 12543 4 D10
port 30 nsew
rlabel locali s -6266 12543 -6226 12613 4 D10
port 30 nsew
rlabel locali s -6265 12613 -6226 12954 4 D10
port 30 nsew
rlabel locali s -6271 12954 -6200 13028 4 D10
port 30 nsew
rlabel locali s -7835 39259 -7781 39398 4 D10
port 30 nsew
rlabel locali s -11101 39259 -11047 39398 4 D10
port 30 nsew
rlabel locali s -7841 40337 -7787 40476 4 D10
port 30 nsew
rlabel locali s -11095 40337 -11041 40476 4 D10
port 30 nsew
rlabel locali s -11106 41448 -10971 41471 4 D10
port 30 nsew
rlabel locali s -14327 41471 -10971 41527 4 D10
port 30 nsew
rlabel locali s -11106 41527 -10971 41593 4 D10
port 30 nsew
rlabel locali s -12009 86105 -11973 86288 4 D10
port 30 nsew
rlabel locali s -15205 7856 -15069 86288 4 D10
port 30 nsew
rlabel locali s -15205 86288 -11973 86424 4 D10
port 30 nsew
rlabel locali s -12009 86424 -11973 86633 4 D10
port 30 nsew
rlabel locali s -12011 86633 -11971 86653 4 D10
port 30 nsew
rlabel locali s -12019 86653 -11965 86788 4 D10
port 30 nsew
rlabel locali s -13172 86424 -13036 89887 4 D10
port 30 nsew
rlabel locali s -13172 89887 -12004 90023 4 D10
port 30 nsew
rlabel locali s -12040 90023 -12004 90301 4 D10
port 30 nsew
rlabel locali s -12042 90301 -12002 90321 4 D10
port 30 nsew
rlabel locali s -12050 90321 -11996 90456 4 D10
port 30 nsew
rlabel metal1 s -4585 -61579 -4446 -61578 2 D16
port 31 nsew
rlabel metal1 s -4585 -61578 -4054 -61576 2 D16
port 31 nsew
rlabel metal1 s -5663 -61585 -5524 -61576 2 D16
port 31 nsew
rlabel metal1 s -5663 -61576 -4054 -61550 2 D16
port 31 nsew
rlabel metal1 s -4082 -61550 -4054 -60400 2 D16
port 31 nsew
rlabel metal1 s -5663 -61550 -4446 -61548 2 D16
port 31 nsew
rlabel metal1 s -4585 -61548 -4446 -61525 2 D16
port 31 nsew
rlabel metal1 s -5663 -61548 -5524 -61531 2 D16
port 31 nsew
rlabel metal1 s -4082 -60400 10126 -60349 8 D16
port 31 nsew
rlabel metal1 s 10075 -60349 10126 -54999 8 D16
port 31 nsew
rlabel metal1 s -12881 -57359 -12751 -57209 2 D16
port 31 nsew
rlabel metal1 s -12831 -57209 -12777 -57012 2 D16
port 31 nsew
rlabel metal1 s -14442 -62751 -14266 -57012 2 D16
port 31 nsew
rlabel metal1 s -22536 -62749 -22413 -62626 2 D16
port 31 nsew
rlabel metal1 s -14442 -57012 -12777 -56836 2 D16
port 31 nsew
rlabel metal1 s -12831 -56836 -12777 -55805 2 D16
port 31 nsew
rlabel metal1 s -12974 -55805 -12777 -55751 2 D16
port 31 nsew
rlabel metal1 s -5739 -54999 10126 -54948 8 D16
port 31 nsew
rlabel metal1 s -5739 -54948 -5688 -54566 2 D16
port 31 nsew
rlabel metal1 s -5739 -54566 -5603 -54492 2 D16
port 31 nsew
rlabel metal1 s -22483 -62626 -22422 -54099 2 D16
port 31 nsew
rlabel locali s -33062 -62751 28011 -62615 2 D16
port 31 nsew
rlabel locali s 27875 -62615 28011 -61389 8 D16
port 31 nsew
rlabel locali s 27875 -61389 31610 -61253 8 D16
port 31 nsew
rlabel locali s 31908 -60267 32043 -60259 8 D16
port 31 nsew
rlabel locali s 31888 -60259 32043 -60257 8 D16
port 31 nsew
rlabel locali s 31474 -61253 31610 -60257 8 D16
port 31 nsew
rlabel locali s 31474 -60257 32043 -60221 8 D16
port 31 nsew
rlabel locali s 28240 -60236 28375 -60228 8 D16
port 31 nsew
rlabel locali s 28220 -60228 28375 -60226 8 D16
port 31 nsew
rlabel locali s 27875 -61253 28011 -60226 8 D16
port 31 nsew
rlabel locali s 9253 -62615 9309 -61205 8 D16
port 31 nsew
rlabel locali s -4585 -61579 -4446 -61525 2 D16
port 31 nsew
rlabel locali s -5663 -61585 -5524 -61531 2 D16
port 31 nsew
rlabel locali s 9252 -61205 9310 -60397 8 D16
port 31 nsew
rlabel locali s 9252 -60397 9376 -60354 8 D16
port 31 nsew
rlabel locali s 9253 -60354 9376 -60353 8 D16
port 31 nsew
rlabel locali s 31888 -60221 32043 -60219 8 D16
port 31 nsew
rlabel locali s 31908 -60219 32043 -60213 8 D16
port 31 nsew
rlabel locali s 27692 -60226 28375 -60190 8 D16
port 31 nsew
rlabel locali s 28220 -60190 28375 -60188 8 D16
port 31 nsew
rlabel locali s 28240 -60188 28375 -60182 8 D16
port 31 nsew
rlabel locali s -20654 -59924 -20509 -59868 2 D16
port 31 nsew
rlabel locali s -20654 -59868 -20594 -59863 2 D16
port 31 nsew
rlabel locali s -22483 -59878 -22423 -59863 2 D16
port 31 nsew
rlabel locali s -22483 -59863 -20594 -59822 2 D16
port 31 nsew
rlabel locali s -22483 -59822 -22423 -59641 2 D16
port 31 nsew
rlabel locali s -12707 -57273 -12634 -57267 2 D16
port 31 nsew
rlabel locali s -12881 -57359 -12751 -57267 2 D16
port 31 nsew
rlabel locali s -12881 -57267 -12634 -57226 2 D16
port 31 nsew
rlabel locali s -12707 -57226 -12634 -57213 2 D16
port 31 nsew
rlabel locali s -12881 -57226 -12751 -57209 2 D16
port 31 nsew
rlabel locali s -12333 -55821 -12259 -55795 2 D16
port 31 nsew
rlabel locali s -12971 -55797 -12744 -55795 2 D16
port 31 nsew
rlabel locali s -12971 -55795 -12259 -55757 2 D16
port 31 nsew
rlabel locali s -12745 -55757 -12259 -55756 2 D16
port 31 nsew
rlabel locali s -12333 -55756 -12259 -55750 2 D16
port 31 nsew
rlabel locali s -12745 -55756 -12674 -55755 2 D16
port 31 nsew
rlabel locali s -5739 -54566 -5551 -54492 2 D16
port 31 nsew
rlabel locali s -20890 -54343 -20755 -54336 2 D16
port 31 nsew
rlabel locali s -22483 -54337 -22422 -54336 2 D16
port 31 nsew
rlabel locali s -22483 -54336 -20755 -54302 2 D16
port 31 nsew
rlabel locali s -20890 -54302 -20755 -54289 2 D16
port 31 nsew
rlabel locali s -22483 -54302 -22422 -54099 2 D16
port 31 nsew
rlabel metal1 s 9294 -62943 9417 -62820 8 D17
port 32 nsew
rlabel metal1 s -22345 -62948 -22222 -62825 2 D17
port 32 nsew
rlabel metal1 s 9347 -62820 9408 -62216 8 D17
port 32 nsew
rlabel metal1 s 9352 -61583 9417 -61578 8 D17
port 32 nsew
rlabel metal1 s 8415 -61579 8554 -61578 8 D17
port 32 nsew
rlabel metal1 s 8313 -61578 10924 -61576 8 D17
port 32 nsew
rlabel metal1 s 7337 -61585 7476 -61576 8 D17
port 32 nsew
rlabel metal1 s 7337 -61576 10924 -61550 8 D17
port 32 nsew
rlabel metal1 s 10896 -61550 10924 -53798 8 D17
port 32 nsew
rlabel metal1 s 9352 -61550 9417 -61446 8 D17
port 32 nsew
rlabel metal1 s 7337 -61550 8554 -61548 8 D17
port 32 nsew
rlabel metal1 s 8415 -61548 8554 -61525 8 D17
port 32 nsew
rlabel metal1 s 7337 -61548 7476 -61531 8 D17
port 32 nsew
rlabel metal1 s -22292 -62825 -22231 -54020 2 D17
port 32 nsew
rlabel metal1 s 8415 -53823 8554 -53800 8 D17
port 32 nsew
rlabel metal1 s 7337 -53817 7476 -53800 8 D17
port 32 nsew
rlabel metal1 s 7337 -53800 8554 -53798 8 D17
port 32 nsew
rlabel metal1 s 7337 -53798 10924 -53772 8 D17
port 32 nsew
rlabel metal1 s 8313 -53772 10924 -53770 8 D17
port 32 nsew
rlabel metal1 s 8415 -53770 8554 -53769 8 D17
port 32 nsew
rlabel metal1 s 7337 -53772 7476 -53763 8 D17
port 32 nsew
rlabel locali s -33463 -62950 36451 -62814 8 D17
port 32 nsew
rlabel locali s 36315 -62814 36451 -61400 8 D17
port 32 nsew
rlabel locali s 9355 -62343 9409 -61583 8 D17
port 32 nsew
rlabel locali s 9352 -61583 9417 -61446 8 D17
port 32 nsew
rlabel locali s 8415 -61579 8554 -61525 8 D17
port 32 nsew
rlabel locali s 7337 -61585 7476 -61531 8 D17
port 32 nsew
rlabel locali s 36315 -61400 40050 -61264 8 D17
port 32 nsew
rlabel locali s 40348 -60278 40483 -60270 8 D17
port 32 nsew
rlabel locali s 40328 -60270 40483 -60268 8 D17
port 32 nsew
rlabel locali s 39914 -61264 40050 -60268 8 D17
port 32 nsew
rlabel locali s 39914 -60268 40483 -60232 8 D17
port 32 nsew
rlabel locali s 36680 -60247 36815 -60239 8 D17
port 32 nsew
rlabel locali s 36660 -60239 36815 -60237 8 D17
port 32 nsew
rlabel locali s 36315 -61264 36451 -60237 8 D17
port 32 nsew
rlabel locali s 40328 -60232 40483 -60230 8 D17
port 32 nsew
rlabel locali s 40348 -60230 40483 -60224 8 D17
port 32 nsew
rlabel locali s 36132 -60237 36815 -60201 8 D17
port 32 nsew
rlabel locali s 36660 -60201 36815 -60199 8 D17
port 32 nsew
rlabel locali s 36680 -60199 36815 -60193 8 D17
port 32 nsew
rlabel locali s -20974 -59956 -20829 -59952 2 D17
port 32 nsew
rlabel locali s -22292 -60135 -22232 -59952 2 D17
port 32 nsew
rlabel locali s -22292 -59952 -20829 -59911 2 D17
port 32 nsew
rlabel locali s -20974 -59911 -20829 -59900 2 D17
port 32 nsew
rlabel locali s -22292 -59911 -22232 -59898 2 D17
port 32 nsew
rlabel locali s -21078 -54265 -20943 -54258 2 D17
port 32 nsew
rlabel locali s -22292 -54258 -20943 -54220 2 D17
port 32 nsew
rlabel locali s -21078 -54220 -20943 -54211 2 D17
port 32 nsew
rlabel locali s -22292 -54220 -22231 -54020 2 D17
port 32 nsew
rlabel locali s 8415 -53823 8554 -53769 8 D17
port 32 nsew
rlabel locali s 7337 -53817 7476 -53763 8 D17
port 32 nsew
rlabel metal1 s 9400 -63176 9523 -63053 8 D18
port 33 nsew
rlabel metal1 s -22239 -63181 -22116 -63058 2 D18
port 33 nsew
rlabel metal1 s 9456 -63053 9516 -62220 8 D18
port 33 nsew
rlabel metal1 s 9465 -62220 9509 -62217 8 D18
port 33 nsew
rlabel metal1 s 5415 -61579 5554 -61578 8 D18
port 33 nsew
rlabel metal1 s 5415 -61578 6774 -61576 8 D18
port 33 nsew
rlabel metal1 s 4337 -61585 4476 -61576 8 D18
port 33 nsew
rlabel metal1 s 4337 -61576 6774 -61550 8 D18
port 33 nsew
rlabel metal1 s 9387 -60956 9526 -60952 8 D18
port 33 nsew
rlabel metal1 s 6746 -61550 6774 -60952 8 D18
port 33 nsew
rlabel metal1 s 4337 -61550 5554 -61548 8 D18
port 33 nsew
rlabel metal1 s 5415 -61548 5554 -61525 8 D18
port 33 nsew
rlabel metal1 s 4337 -61548 4476 -61531 8 D18
port 33 nsew
rlabel metal1 s 6746 -60952 10773 -60924 8 D18
port 33 nsew
rlabel metal1 s 10745 -60924 10773 -54424 8 D18
port 33 nsew
rlabel metal1 s 9387 -60924 9526 -60909 8 D18
port 33 nsew
rlabel metal1 s -22183 -63058 -22123 -60238 2 D18
port 33 nsew
rlabel metal1 s -22183 -60238 -22122 -60001 2 D18
port 33 nsew
rlabel metal1 s 6746 -54424 10773 -54396 8 D18
port 33 nsew
rlabel metal1 s 6746 -54396 6774 -53798 8 D18
port 33 nsew
rlabel metal1 s -22183 -60001 -22123 -54172 2 D18
port 33 nsew
rlabel metal1 s -22183 -54172 -22122 -53934 2 D18
port 33 nsew
rlabel metal1 s 5415 -53823 5554 -53800 8 D18
port 33 nsew
rlabel metal1 s 4337 -53817 4476 -53800 8 D18
port 33 nsew
rlabel metal1 s 4337 -53800 5554 -53798 8 D18
port 33 nsew
rlabel metal1 s 4337 -53798 6774 -53772 8 D18
port 33 nsew
rlabel metal1 s 5415 -53772 6774 -53770 8 D18
port 33 nsew
rlabel metal1 s 5415 -53770 5554 -53769 8 D18
port 33 nsew
rlabel metal1 s 4337 -53772 4476 -53763 8 D18
port 33 nsew
rlabel locali s -32991 -63183 45361 -63047 8 D18
port 33 nsew
rlabel locali s 45225 -63047 45361 -61439 8 D18
port 33 nsew
rlabel locali s 45178 -61439 48913 -61303 8 D18
port 33 nsew
rlabel locali s 49211 -60317 49346 -60309 8 D18
port 33 nsew
rlabel locali s 49191 -60309 49346 -60307 8 D18
port 33 nsew
rlabel locali s 48777 -61303 48913 -60307 8 D18
port 33 nsew
rlabel locali s 45178 -61303 45361 -61289 8 D18
port 33 nsew
rlabel locali s 48777 -60307 49346 -60271 8 D18
port 33 nsew
rlabel locali s 45543 -60286 45678 -60278 8 D18
port 33 nsew
rlabel locali s 45523 -60278 45678 -60276 8 D18
port 33 nsew
rlabel locali s 45178 -61289 45314 -60276 8 D18
port 33 nsew
rlabel locali s 9460 -62343 9514 -60955 8 D18
port 33 nsew
rlabel locali s 5415 -61579 5554 -61525 8 D18
port 33 nsew
rlabel locali s 4337 -61585 4476 -61531 8 D18
port 33 nsew
rlabel locali s 9396 -60955 9519 -60911 8 D18
port 33 nsew
rlabel locali s 49191 -60271 49346 -60269 8 D18
port 33 nsew
rlabel locali s 49211 -60269 49346 -60263 8 D18
port 33 nsew
rlabel locali s 44995 -60276 45678 -60240 8 D18
port 33 nsew
rlabel locali s 45523 -60240 45678 -60238 8 D18
port 33 nsew
rlabel locali s 45543 -60238 45678 -60232 8 D18
port 33 nsew
rlabel locali s -21303 -60051 -21158 -60044 2 D18
port 33 nsew
rlabel locali s -22182 -60238 -22122 -60044 2 D18
port 33 nsew
rlabel locali s -22182 -60044 -21158 -60003 2 D18
port 33 nsew
rlabel locali s -21303 -60003 -21158 -59995 2 D18
port 33 nsew
rlabel locali s -22182 -60003 -22122 -60001 2 D18
port 33 nsew
rlabel locali s -21414 -54183 -21279 -54174 2 D18
port 33 nsew
rlabel locali s -21433 -54174 -21279 -54172 2 D18
port 33 nsew
rlabel locali s -22183 -54172 -21279 -54137 2 D18
port 33 nsew
rlabel locali s -21414 -54137 -21279 -54129 2 D18
port 33 nsew
rlabel locali s -22183 -54137 -22122 -53934 2 D18
port 33 nsew
rlabel locali s 5415 -53823 5554 -53769 8 D18
port 33 nsew
rlabel locali s 4337 -53817 4476 -53763 8 D18
port 33 nsew
rlabel metal1 s 9493 -63433 9617 -63310 8 D19
port 34 nsew
rlabel metal1 s -22146 -63438 -22022 -63315 2 D19
port 34 nsew
rlabel metal1 s 9555 -63310 9616 -62363 8 D19
port 34 nsew
rlabel metal1 s -20209 -60648 -20151 -60511 2 D19
port 34 nsew
rlabel metal1 s -20189 -60511 -20154 -59602 2 D19
port 34 nsew
rlabel metal1 s -20189 -59602 -20131 -59465 2 D19
port 34 nsew
rlabel metal1 s 9536 -59339 9681 -59327 8 D19
port 34 nsew
rlabel metal1 s 8425 -59328 8564 -59327 8 D19
port 34 nsew
rlabel metal1 s 8425 -59327 9798 -59325 8 D19
port 34 nsew
rlabel metal1 s 7347 -59334 7486 -59325 8 D19
port 34 nsew
rlabel metal1 s 7347 -59325 9798 -59299 8 D19
port 34 nsew
rlabel metal1 s 9768 -59299 9796 -56064 8 D19
port 34 nsew
rlabel metal1 s 9536 -59299 9681 -59204 8 D19
port 34 nsew
rlabel metal1 s 7347 -59299 8564 -59297 8 D19
port 34 nsew
rlabel metal1 s 8425 -59297 8564 -59274 8 D19
port 34 nsew
rlabel metal1 s 7347 -59297 7486 -59280 8 D19
port 34 nsew
rlabel metal1 s 9755 -56064 9806 -56049 8 D19
port 34 nsew
rlabel metal1 s 8425 -56074 8564 -56051 8 D19
port 34 nsew
rlabel metal1 s 7347 -56068 7486 -56051 8 D19
port 34 nsew
rlabel metal1 s 7347 -56051 8564 -56049 8 D19
port 34 nsew
rlabel metal1 s 7347 -56049 9806 -56023 8 D19
port 34 nsew
rlabel metal1 s 8425 -56023 9806 -56021 8 D19
port 34 nsew
rlabel metal1 s 9755 -56021 9806 -56013 8 D19
port 34 nsew
rlabel metal1 s 8425 -56021 8564 -56020 8 D19
port 34 nsew
rlabel metal1 s 7347 -56023 7486 -56014 8 D19
port 34 nsew
rlabel metal1 s -19667 -55337 -19535 -55333 2 D19
port 34 nsew
rlabel metal1 s -19714 -55333 -19511 -55293 2 D19
port 34 nsew
rlabel metal1 s -19667 -55293 -19511 -55284 2 D19
port 34 nsew
rlabel metal1 s -19551 -55284 -19511 -54511 2 D19
port 34 nsew
rlabel metal1 s -22084 -63315 -22023 -55099 2 D19
port 34 nsew
rlabel metal1 s -19558 -54511 -19421 -54453 2 D19
port 34 nsew
rlabel locali s -32976 -63438 54512 -63302 8 D19
port 34 nsew
rlabel locali s 54376 -63302 54512 -61405 8 D19
port 34 nsew
rlabel locali s 54376 -61405 58111 -61269 8 D19
port 34 nsew
rlabel locali s 58409 -60283 58544 -60275 8 D19
port 34 nsew
rlabel locali s 58389 -60275 58544 -60273 8 D19
port 34 nsew
rlabel locali s 57975 -61269 58111 -60273 8 D19
port 34 nsew
rlabel locali s 57975 -60273 58544 -60237 8 D19
port 34 nsew
rlabel locali s 54741 -60252 54876 -60244 8 D19
port 34 nsew
rlabel locali s 54721 -60244 54876 -60242 8 D19
port 34 nsew
rlabel locali s 54376 -61269 54512 -60242 8 D19
port 34 nsew
rlabel locali s 58389 -60237 58544 -60235 8 D19
port 34 nsew
rlabel locali s 58409 -60235 58544 -60229 8 D19
port 34 nsew
rlabel locali s 54193 -60242 54876 -60206 8 D19
port 34 nsew
rlabel locali s 54721 -60206 54876 -60204 8 D19
port 34 nsew
rlabel locali s 54741 -60204 54876 -60198 8 D19
port 34 nsew
rlabel locali s 9559 -62560 9615 -59339 8 D19
port 34 nsew
rlabel locali s -22084 -60648 -20151 -60607 2 D19
port 34 nsew
rlabel locali s -20209 -60607 -20151 -60511 2 D19
port 34 nsew
rlabel locali s -22084 -60607 -22026 -60511 2 D19
port 34 nsew
rlabel locali s -19782 -59613 -19639 -59596 2 D19
port 34 nsew
rlabel locali s -20189 -59602 -20131 -59596 2 D19
port 34 nsew
rlabel locali s -20189 -59596 -19639 -59560 2 D19
port 34 nsew
rlabel locali s -19782 -59560 -19639 -59553 2 D19
port 34 nsew
rlabel locali s -20189 -59560 -20131 -59465 2 D19
port 34 nsew
rlabel locali s 9536 -59339 9681 -59204 8 D19
port 34 nsew
rlabel locali s 8425 -59328 8564 -59274 8 D19
port 34 nsew
rlabel locali s 7347 -59334 7486 -59280 8 D19
port 34 nsew
rlabel locali s 8425 -56074 8564 -56020 8 D19
port 34 nsew
rlabel locali s 7347 -56068 7486 -56014 8 D19
port 34 nsew
rlabel locali s -19667 -55337 -19535 -55333 2 D19
port 34 nsew
rlabel locali s -22084 -55337 -22024 -55333 2 D19
port 34 nsew
rlabel locali s -22084 -55333 -19535 -55293 2 D19
port 34 nsew
rlabel locali s -19667 -55293 -19535 -55284 2 D19
port 34 nsew
rlabel locali s -22084 -55293 -22024 -55216 2 D19
port 34 nsew
rlabel locali s -22084 -55216 -22016 -55176 2 D19
port 34 nsew
rlabel locali s -22084 -55176 -22024 -55100 2 D19
port 34 nsew
rlabel locali s -18958 -54504 -18884 -54498 2 D19
port 34 nsew
rlabel locali s -19370 -54499 -19299 -54498 2 D19
port 34 nsew
rlabel locali s -19370 -54498 -18884 -54497 2 D19
port 34 nsew
rlabel locali s -19558 -54511 -19421 -54497 2 D19
port 34 nsew
rlabel locali s -19596 -54497 -18884 -54459 2 D19
port 34 nsew
rlabel locali s -18958 -54459 -18884 -54433 2 D19
port 34 nsew
rlabel locali s -19596 -54459 -19369 -54457 2 D19
port 34 nsew
rlabel locali s -19558 -54457 -19421 -54453 2 D19
port 34 nsew
rlabel metal1 s 26730 -62429 82728 -62184 8 OUTB
port 35 nsew
rlabel metal1 s 27599 -56846 27858 -56583 8 OUTB
port 35 nsew
rlabel metal1 s 29230 -55436 29389 -55378 8 OUTB
port 35 nsew
rlabel metal1 s 29256 -55378 29310 -55323 8 OUTB
port 35 nsew
rlabel metal1 s 28982 -55323 29310 -55269 8 OUTB
port 35 nsew
rlabel metal1 s 28982 -55269 29036 -54979 8 OUTB
port 35 nsew
rlabel metal1 s 26730 -62184 26975 -55085 8 OUTB
port 35 nsew
rlabel metal1 s 11260 -64637 11555 -62375 8 OUTB
port 35 nsew
rlabel metal1 s -22800 -64647 -22587 -64469 2 OUTB
port 35 nsew
rlabel metal1 s 10208 -62375 11555 -62106 8 OUTB
port 35 nsew
rlabel metal1 s 15295 -61148 15432 -61088 8 OUTB
port 35 nsew
rlabel metal1 s 14397 -61511 14457 -61147 8 OUTB
port 35 nsew
rlabel metal1 s 15323 -61088 15383 -60640 8 OUTB
port 35 nsew
rlabel metal1 s 14354 -61147 14486 -61087 8 OUTB
port 35 nsew
rlabel metal1 s 23451 -57046 23511 -56598 8 OUTB
port 35 nsew
rlabel metal1 s 23423 -56598 23560 -56538 8 OUTB
port 35 nsew
rlabel metal1 s 22482 -56599 22614 -56539 8 OUTB
port 35 nsew
rlabel metal1 s 22525 -56539 22585 -56175 8 OUTB
port 35 nsew
rlabel metal1 s 20009 -56214 20141 -56079 8 OUTB
port 35 nsew
rlabel metal1 s 20036 -56079 20111 -56004 8 OUTB
port 35 nsew
rlabel metal1 s 18441 -56042 18620 -56004 8 OUTB
port 35 nsew
rlabel metal1 s 18441 -56004 20111 -55929 8 OUTB
port 35 nsew
rlabel metal1 s 18441 -55929 18620 -55853 8 OUTB
port 35 nsew
rlabel metal1 s 16597 -55085 26975 -55067 8 OUTB
port 35 nsew
rlabel metal1 s 27598 -55019 27811 -54979 8 OUTB
port 35 nsew
rlabel metal1 s 27598 -54979 29036 -54925 8 OUTB
port 35 nsew
rlabel metal1 s 27598 -54925 27811 -54886 8 OUTB
port 35 nsew
rlabel metal1 s 16597 -55067 27010 -54773 8 OUTB
port 35 nsew
rlabel metal1 s 11260 -62106 11555 -54816 8 OUTB
port 35 nsew
rlabel metal1 s 9830 -60321 10021 -60214 8 OUTB
port 35 nsew
rlabel metal1 s 9950 -60214 10001 -60143 8 OUTB
port 35 nsew
rlabel metal1 s 38 -60143 10001 -60092 8 OUTB
port 35 nsew
rlabel metal1 s 9950 -60092 10001 -55256 8 OUTB
port 35 nsew
rlabel metal1 s -2528 -59086 -2396 -59026 2 OUTB
port 35 nsew
rlabel metal1 s -3425 -59533 -3365 -59085 2 OUTB
port 35 nsew
rlabel metal1 s -2499 -59026 -2439 -58662 2 OUTB
port 35 nsew
rlabel metal1 s -3474 -59085 -3337 -59025 2 OUTB
port 35 nsew
rlabel metal1 s -5211 -56701 -5151 -56234 2 OUTB
port 35 nsew
rlabel metal1 s -5247 -56234 -5115 -56174 2 OUTB
port 35 nsew
rlabel metal1 s -22783 -64469 -22647 -55544 2 OUTB
port 35 nsew
rlabel metal1 s -31679 -64865 -30522 -63836 2 OUTB
port 35 nsew
rlabel metal1 s -31679 -63836 -30520 -62597 2 OUTB
port 35 nsew
rlabel metal1 s -22783 -55544 -22543 -55501 2 OUTB
port 35 nsew
rlabel metal1 s -22783 -55501 -22530 -55313 2 OUTB
port 35 nsew
rlabel metal1 s -22631 -55313 -22530 -55258 2 OUTB
port 35 nsew
rlabel metal1 s 38 -55256 10001 -55205 8 OUTB
port 35 nsew
rlabel metal1 s 16597 -54773 26830 -54733 8 OUTB
port 35 nsew
rlabel metal1 s 58913 -9909 59860 -8831 8 OUTB
port 35 nsew
rlabel metal1 s 59172 -8831 59616 2260 8 OUTB
port 35 nsew
rlabel metal1 s -31679 -62597 -30522 -8679 2 OUTB
port 35 nsew
rlabel metal1 s 58706 2260 59616 2704 6 OUTB
port 35 nsew
rlabel metal1 s 54604 1826 54650 2327 6 OUTB
port 35 nsew
rlabel metal1 s 54368 1826 54414 2327 6 OUTB
port 35 nsew
rlabel metal1 s 54132 1826 54178 2327 6 OUTB
port 35 nsew
rlabel metal1 s 53896 1826 53942 2327 6 OUTB
port 35 nsew
rlabel metal1 s 53660 1826 53706 2327 6 OUTB
port 35 nsew
rlabel metal1 s 53424 1826 53470 2327 6 OUTB
port 35 nsew
rlabel metal1 s 53188 1826 53234 2327 6 OUTB
port 35 nsew
rlabel metal1 s 52952 1826 52998 2327 6 OUTB
port 35 nsew
rlabel metal1 s 52952 2327 54650 2373 6 OUTB
port 35 nsew
rlabel metal1 s 54604 2373 54650 2489 6 OUTB
port 35 nsew
rlabel metal1 s 54558 2489 58435 2563 6 OUTB
port 35 nsew
rlabel metal1 s 58360 2563 58406 3034 6 OUTB
port 35 nsew
rlabel metal1 s 58124 2563 58170 3034 6 OUTB
port 35 nsew
rlabel metal1 s 57888 2563 57934 3034 6 OUTB
port 35 nsew
rlabel metal1 s 57652 2563 57698 3034 6 OUTB
port 35 nsew
rlabel metal1 s 57416 2563 57462 3034 6 OUTB
port 35 nsew
rlabel metal1 s 57180 2563 57226 3034 6 OUTB
port 35 nsew
rlabel metal1 s 56944 2563 56990 3034 6 OUTB
port 35 nsew
rlabel metal1 s 56708 2563 56754 3034 6 OUTB
port 35 nsew
rlabel metal1 s 56472 2563 56518 3034 6 OUTB
port 35 nsew
rlabel metal1 s 56236 2563 56282 3034 6 OUTB
port 35 nsew
rlabel metal1 s 56000 2563 56046 3034 6 OUTB
port 35 nsew
rlabel metal1 s 55764 2563 55810 3034 6 OUTB
port 35 nsew
rlabel metal1 s 55528 2563 55574 3034 6 OUTB
port 35 nsew
rlabel metal1 s 55292 2563 55338 3034 6 OUTB
port 35 nsew
rlabel metal1 s 55056 2563 55102 3034 6 OUTB
port 35 nsew
rlabel metal1 s 54820 2563 54866 3034 6 OUTB
port 35 nsew
rlabel metal1 s 54584 2563 54630 3034 6 OUTB
port 35 nsew
rlabel locali s -22800 -64647 -22587 -64637 2 OUTB
port 35 nsew
rlabel locali s -31679 -64865 -30522 -64637 2 OUTB
port 35 nsew
rlabel locali s -31679 -64637 11555 -64501 2 OUTB
port 35 nsew
rlabel locali s -22800 -64501 -22587 -64469 2 OUTB
port 35 nsew
rlabel locali s -31679 -64501 -30522 -63836 2 OUTB
port 35 nsew
rlabel locali s -31679 -63836 -30520 -63625 2 OUTB
port 35 nsew
rlabel locali s 80324 -62425 80724 -62187 8 OUTB
port 35 nsew
rlabel locali s 80373 -62187 80667 -56743 8 OUTB
port 35 nsew
rlabel locali s 71371 -62429 71753 -62184 8 OUTB
port 35 nsew
rlabel locali s 62066 -62419 62414 -62187 8 OUTB
port 35 nsew
rlabel locali s 53567 -62407 53799 -62202 8 OUTB
port 35 nsew
rlabel locali s 44228 -62380 44480 -62241 8 OUTB
port 35 nsew
rlabel locali s 71456 -62184 71641 -56776 8 OUTB
port 35 nsew
rlabel locali s 62128 -62187 62367 -56802 8 OUTB
port 35 nsew
rlabel locali s 53601 -62202 53747 -56834 8 OUTB
port 35 nsew
rlabel locali s 44282 -62241 44428 -56926 8 OUTB
port 35 nsew
rlabel locali s 35531 -62426 35805 -62223 8 OUTB
port 35 nsew
rlabel locali s 82020 -56678 82155 -56670 8 OUTB
port 35 nsew
rlabel locali s 82000 -56670 82155 -56668 8 OUTB
port 35 nsew
rlabel locali s 80373 -56743 81581 -56668 8 OUTB
port 35 nsew
rlabel locali s 80373 -56668 82155 -56632 8 OUTB
port 35 nsew
rlabel locali s 72656 -56716 72791 -56708 8 OUTB
port 35 nsew
rlabel locali s 72636 -56708 72791 -56706 8 OUTB
port 35 nsew
rlabel locali s 71456 -56776 72120 -56706 8 OUTB
port 35 nsew
rlabel locali s 71456 -56706 72791 -56670 8 OUTB
port 35 nsew
rlabel locali s 63503 -56733 63638 -56725 8 OUTB
port 35 nsew
rlabel locali s 63483 -56725 63638 -56723 8 OUTB
port 35 nsew
rlabel locali s 62128 -56802 63054 -56723 8 OUTB
port 35 nsew
rlabel locali s 54749 -56799 54884 -56791 8 OUTB
port 35 nsew
rlabel locali s 54729 -56791 54884 -56789 8 OUTB
port 35 nsew
rlabel locali s 53601 -56834 54330 -56789 8 OUTB
port 35 nsew
rlabel locali s 53601 -56789 54884 -56753 8 OUTB
port 35 nsew
rlabel locali s 45551 -56833 45686 -56825 8 OUTB
port 35 nsew
rlabel locali s 45531 -56825 45686 -56823 8 OUTB
port 35 nsew
rlabel locali s 44282 -56926 45049 -56823 8 OUTB
port 35 nsew
rlabel locali s 35600 -62223 35746 -56840 8 OUTB
port 35 nsew
rlabel locali s 27305 -62403 27526 -62208 8 OUTB
port 35 nsew
rlabel locali s 10286 -62347 10414 -62168 8 OUTB
port 35 nsew
rlabel locali s 14229 -61612 14397 -61601 8 OUTB
port 35 nsew
rlabel locali s 14229 -61601 14457 -61538 8 OUTB
port 35 nsew
rlabel locali s 14397 -61538 14457 -61379 8 OUTB
port 35 nsew
rlabel locali s 15295 -61148 15432 -61137 8 OUTB
port 35 nsew
rlabel locali s 14354 -61147 14486 -61137 8 OUTB
port 35 nsew
rlabel locali s 11260 -61203 11555 -61137 8 OUTB
port 35 nsew
rlabel locali s 11260 -61137 17611 -61098 8 OUTB
port 35 nsew
rlabel locali s 15295 -61098 15432 -61088 8 OUTB
port 35 nsew
rlabel locali s 14354 -61098 14486 -61087 8 OUTB
port 35 nsew
rlabel locali s 15443 -60704 15611 -60699 8 OUTB
port 35 nsew
rlabel locali s 15323 -60772 15383 -60699 8 OUTB
port 35 nsew
rlabel locali s 11881 -61098 11920 -60704 8 OUTB
port 35 nsew
rlabel locali s 11260 -61098 11555 -61000 8 OUTB
port 35 nsew
rlabel locali s 15323 -60699 15611 -60641 8 OUTB
port 35 nsew
rlabel locali s 15443 -60641 15611 -60630 8 OUTB
port 35 nsew
rlabel locali s 15323 -60641 15383 -60640 8 OUTB
port 35 nsew
rlabel locali s 11861 -60704 12029 -60630 8 OUTB
port 35 nsew
rlabel locali s 10310 -62168 10393 -60303 8 OUTB
port 35 nsew
rlabel locali s 9830 -60321 10021 -60303 8 OUTB
port 35 nsew
rlabel locali s 9830 -60303 10393 -60220 8 OUTB
port 35 nsew
rlabel locali s 9830 -60220 10021 -60214 8 OUTB
port 35 nsew
rlabel locali s 38 -60143 175 -60092 8 OUTB
port 35 nsew
rlabel locali s 38 -60092 77 -59543 8 OUTB
port 35 nsew
rlabel locali s -71 -59543 97 -59469 8 OUTB
port 35 nsew
rlabel locali s -3425 -59533 -3365 -59532 2 OUTB
port 35 nsew
rlabel locali s -3653 -59543 -3485 -59532 2 OUTB
port 35 nsew
rlabel locali s -3653 -59532 -3365 -59474 2 OUTB
port 35 nsew
rlabel locali s 38 -59469 77 -59075 8 OUTB
port 35 nsew
rlabel locali s -3425 -59474 -3365 -59401 2 OUTB
port 35 nsew
rlabel locali s -3653 -59474 -3485 -59469 2 OUTB
port 35 nsew
rlabel locali s -2528 -59086 -2396 -59075 2 OUTB
port 35 nsew
rlabel locali s -3474 -59085 -3337 -59075 2 OUTB
port 35 nsew
rlabel locali s -5653 -59075 77 -59036 2 OUTB
port 35 nsew
rlabel locali s -2528 -59036 -2396 -59026 2 OUTB
port 35 nsew
rlabel locali s -3474 -59036 -3337 -59025 2 OUTB
port 35 nsew
rlabel locali s -2499 -58794 -2439 -58635 2 OUTB
port 35 nsew
rlabel locali s -2499 -58635 -2271 -58572 2 OUTB
port 35 nsew
rlabel locali s -2439 -58572 -2271 -58561 2 OUTB
port 35 nsew
rlabel locali s 23571 -57056 23739 -57045 8 OUTB
port 35 nsew
rlabel locali s 23451 -57046 23511 -57045 8 OUTB
port 35 nsew
rlabel locali s 23451 -57045 23739 -56987 8 OUTB
port 35 nsew
rlabel locali s 23571 -56987 23739 -56982 8 OUTB
port 35 nsew
rlabel locali s 23451 -56987 23511 -56914 8 OUTB
port 35 nsew
rlabel locali s 19989 -57056 20157 -56982 8 OUTB
port 35 nsew
rlabel locali s 44282 -56823 45686 -56787 8 OUTB
port 35 nsew
rlabel locali s 45531 -56787 45686 -56785 8 OUTB
port 35 nsew
rlabel locali s 45551 -56785 45686 -56779 8 OUTB
port 35 nsew
rlabel locali s 44282 -56787 45049 -56780 8 OUTB
port 35 nsew
rlabel locali s 36688 -56794 36823 -56786 8 OUTB
port 35 nsew
rlabel locali s 36668 -56786 36823 -56784 8 OUTB
port 35 nsew
rlabel locali s 35600 -56840 36248 -56784 8 OUTB
port 35 nsew
rlabel locali s 54729 -56753 54884 -56751 8 OUTB
port 35 nsew
rlabel locali s 54749 -56751 54884 -56745 8 OUTB
port 35 nsew
rlabel locali s 62128 -56723 63638 -56687 8 OUTB
port 35 nsew
rlabel locali s 53601 -56753 54330 -56688 8 OUTB
port 35 nsew
rlabel locali s 35600 -56784 36823 -56748 8 OUTB
port 35 nsew
rlabel locali s 27599 -56846 27858 -56831 8 OUTB
port 35 nsew
rlabel locali s 36668 -56748 36823 -56746 8 OUTB
port 35 nsew
rlabel locali s 36688 -56746 36823 -56740 8 OUTB
port 35 nsew
rlabel locali s 35600 -56748 36248 -56694 8 OUTB
port 35 nsew
rlabel locali s 28248 -56783 28383 -56775 8 OUTB
port 35 nsew
rlabel locali s 28228 -56775 28383 -56773 8 OUTB
port 35 nsew
rlabel locali s 26733 -56831 27858 -56773 8 OUTB
port 35 nsew
rlabel locali s 26733 -56773 28383 -56737 8 OUTB
port 35 nsew
rlabel locali s 28228 -56737 28383 -56735 8 OUTB
port 35 nsew
rlabel locali s 28248 -56735 28383 -56729 8 OUTB
port 35 nsew
rlabel locali s 63483 -56687 63638 -56685 8 OUTB
port 35 nsew
rlabel locali s 63503 -56685 63638 -56679 8 OUTB
port 35 nsew
rlabel locali s 72636 -56670 72791 -56668 8 OUTB
port 35 nsew
rlabel locali s 72656 -56668 72791 -56662 8 OUTB
port 35 nsew
rlabel locali s 82000 -56632 82155 -56630 8 OUTB
port 35 nsew
rlabel locali s 82020 -56630 82155 -56624 8 OUTB
port 35 nsew
rlabel locali s 80373 -56632 81581 -56449 8 OUTB
port 35 nsew
rlabel locali s 71456 -56670 72120 -56591 8 OUTB
port 35 nsew
rlabel locali s 62128 -56687 63054 -56563 8 OUTB
port 35 nsew
rlabel locali s 26733 -56737 27858 -56626 8 OUTB
port 35 nsew
rlabel locali s 27599 -56626 27858 -56583 8 OUTB
port 35 nsew
rlabel locali s 23423 -56598 23560 -56588 8 OUTB
port 35 nsew
rlabel locali s 22482 -56599 22614 -56588 8 OUTB
port 35 nsew
rlabel locali s 20009 -56982 20048 -56588 8 OUTB
port 35 nsew
rlabel locali s -5139 -56787 -4971 -56776 2 OUTB
port 35 nsew
rlabel locali s -5174 -56776 -4971 -56775 2 OUTB
port 35 nsew
rlabel locali s -5211 -56775 -4971 -56713 2 OUTB
port 35 nsew
rlabel locali s 20009 -56588 25739 -56549 8 OUTB
port 35 nsew
rlabel locali s -5211 -56713 -5151 -56569 2 OUTB
port 35 nsew
rlabel locali s 23423 -56549 23560 -56538 8 OUTB
port 35 nsew
rlabel locali s 22482 -56549 22614 -56539 8 OUTB
port 35 nsew
rlabel locali s 22525 -56307 22585 -56148 8 OUTB
port 35 nsew
rlabel locali s 20009 -56549 20115 -56214 8 OUTB
port 35 nsew
rlabel locali s -5247 -56234 -5115 -56226 2 OUTB
port 35 nsew
rlabel locali s 22357 -56148 22585 -56085 8 OUTB
port 35 nsew
rlabel locali s 22357 -56085 22525 -56074 8 OUTB
port 35 nsew
rlabel locali s 20009 -56214 20141 -56079 8 OUTB
port 35 nsew
rlabel locali s -5653 -56226 77 -56187 2 OUTB
port 35 nsew
rlabel locali s 18441 -56042 18620 -55853 8 OUTB
port 35 nsew
rlabel locali s 38 -56187 77 -55879 8 OUTB
port 35 nsew
rlabel locali s -1556 -56187 -1481 -56064 2 OUTB
port 35 nsew
rlabel locali s -5247 -56187 -5115 -56174 2 OUTB
port 35 nsew
rlabel locali s -1556 -56064 -1482 -55905 2 OUTB
port 35 nsew
rlabel locali s 29247 -55435 29382 -55429 8 OUTB
port 35 nsew
rlabel locali s 29227 -55429 29382 -55427 8 OUTB
port 35 nsew
rlabel locali s 29020 -55427 29382 -55391 8 OUTB
port 35 nsew
rlabel locali s 29227 -55391 29382 -55389 8 OUTB
port 35 nsew
rlabel locali s 29247 -55389 29382 -55381 8 OUTB
port 35 nsew
rlabel locali s 26680 -55067 27010 -55035 8 OUTB
port 35 nsew
rlabel locali s 26680 -55035 27859 -54856 8 OUTB
port 35 nsew
rlabel locali s 18478 -55853 18620 -54996 8 OUTB
port 35 nsew
rlabel locali s -71 -55879 97 -55805 8 OUTB
port 35 nsew
rlabel locali s -953 -55879 -785 -55874 2 OUTB
port 35 nsew
rlabel locali s -953 -55874 -750 -55816 2 OUTB
port 35 nsew
rlabel locali s -953 -55816 -785 -55805 2 OUTB
port 35 nsew
rlabel locali s 38 -55805 77 -55256 8 OUTB
port 35 nsew
rlabel locali s -22631 -55501 -22530 -55494 2 OUTB
port 35 nsew
rlabel locali s 38 -55256 175 -55205 8 OUTB
port 35 nsew
rlabel locali s -22631 -55494 -18064 -55431 2 OUTB
port 35 nsew
rlabel locali s 11260 -55063 16779 -55061 8 OUTB
port 35 nsew
rlabel locali s 26680 -54856 27010 -54773 8 OUTB
port 35 nsew
rlabel locali s 18439 -54996 18657 -54750 8 OUTB
port 35 nsew
rlabel locali s 11260 -55061 16903 -54816 8 OUTB
port 35 nsew
rlabel locali s -17787 -54923 -17652 -54917 2 OUTB
port 35 nsew
rlabel locali s -17807 -54917 -17652 -54915 2 OUTB
port 35 nsew
rlabel locali s -18121 -55431 -18064 -54915 2 OUTB
port 35 nsew
rlabel locali s -22631 -55431 -22530 -55258 2 OUTB
port 35 nsew
rlabel locali s -18198 -54915 -17652 -54879 2 OUTB
port 35 nsew
rlabel locali s -17807 -54879 -17652 -54877 2 OUTB
port 35 nsew
rlabel locali s -17787 -54877 -17652 -54869 2 OUTB
port 35 nsew
rlabel locali s 16668 -54816 16903 -54793 8 OUTB
port 35 nsew
rlabel locali s 58913 -9909 59860 -9713 8 OUTB
port 35 nsew
rlabel locali s -31467 -10014 -30570 -9713 2 OUTB
port 35 nsew
rlabel locali s -34283 -9713 59860 -9060 8 OUTB
port 35 nsew
rlabel locali s 58913 -9060 59860 -8831 8 OUTB
port 35 nsew
rlabel locali s -31467 -9060 -30570 -8797 2 OUTB
port 35 nsew
rlabel locali s 54610 1822 54644 2230 6 OUTB
port 35 nsew
rlabel locali s 54374 1822 54408 2230 6 OUTB
port 35 nsew
rlabel locali s 54138 1822 54172 2230 6 OUTB
port 35 nsew
rlabel locali s 53902 1822 53936 2230 6 OUTB
port 35 nsew
rlabel locali s 53666 1822 53700 2230 6 OUTB
port 35 nsew
rlabel locali s 53430 1822 53464 2230 6 OUTB
port 35 nsew
rlabel locali s 53194 1822 53228 2230 6 OUTB
port 35 nsew
rlabel locali s 52958 1822 52992 2230 6 OUTB
port 35 nsew
rlabel locali s 58711 2334 58930 2450 6 OUTB
port 35 nsew
rlabel locali s 58366 2450 58930 2484 6 OUTB
port 35 nsew
rlabel locali s 58711 2484 58930 2597 6 OUTB
port 35 nsew
rlabel locali s 58366 2484 58400 3038 6 OUTB
port 35 nsew
rlabel locali s 58130 2630 58164 3038 6 OUTB
port 35 nsew
rlabel locali s 57894 2630 57928 3038 6 OUTB
port 35 nsew
rlabel locali s 57658 2630 57692 3038 6 OUTB
port 35 nsew
rlabel locali s 57422 2630 57456 3038 6 OUTB
port 35 nsew
rlabel locali s 57186 2630 57220 3038 6 OUTB
port 35 nsew
rlabel locali s 56950 2630 56984 3038 6 OUTB
port 35 nsew
rlabel locali s 56714 2630 56748 3038 6 OUTB
port 35 nsew
rlabel locali s 56478 2630 56512 3038 6 OUTB
port 35 nsew
rlabel locali s 56242 2630 56276 3038 6 OUTB
port 35 nsew
rlabel locali s 56006 2630 56040 3038 6 OUTB
port 35 nsew
rlabel locali s 55770 2630 55804 3038 6 OUTB
port 35 nsew
rlabel locali s 55534 2630 55568 3038 6 OUTB
port 35 nsew
rlabel locali s 55298 2630 55332 3038 6 OUTB
port 35 nsew
rlabel locali s 55062 2630 55096 3038 6 OUTB
port 35 nsew
rlabel locali s 54826 2630 54860 3038 6 OUTB
port 35 nsew
rlabel locali s 54590 2630 54624 3038 6 OUTB
port 35 nsew
rlabel metal1 s 26027 -44318 82025 -44073 8 OUT
port 36 nsew
rlabel metal1 s 26896 -38735 27155 -38472 8 OUT
port 36 nsew
rlabel metal1 s 28527 -37325 28686 -37267 8 OUT
port 36 nsew
rlabel metal1 s 28553 -37267 28607 -37212 8 OUT
port 36 nsew
rlabel metal1 s 28279 -37212 28607 -37158 8 OUT
port 36 nsew
rlabel metal1 s 28279 -37158 28333 -36868 8 OUT
port 36 nsew
rlabel metal1 s 26027 -44073 26272 -36974 8 OUT
port 36 nsew
rlabel metal1 s 10557 -46526 10852 -44264 8 OUT
port 36 nsew
rlabel metal1 s -23503 -46536 -23290 -46358 2 OUT
port 36 nsew
rlabel metal1 s 9505 -44264 10852 -43995 8 OUT
port 36 nsew
rlabel metal1 s 14592 -43037 14729 -42977 8 OUT
port 36 nsew
rlabel metal1 s 13694 -43400 13754 -43036 8 OUT
port 36 nsew
rlabel metal1 s 14620 -42977 14680 -42529 8 OUT
port 36 nsew
rlabel metal1 s 13651 -43036 13783 -42976 8 OUT
port 36 nsew
rlabel metal1 s 22748 -38935 22808 -38487 8 OUT
port 36 nsew
rlabel metal1 s 22720 -38487 22857 -38427 8 OUT
port 36 nsew
rlabel metal1 s 21779 -38488 21911 -38428 8 OUT
port 36 nsew
rlabel metal1 s 21822 -38428 21882 -38064 8 OUT
port 36 nsew
rlabel metal1 s 19306 -38103 19438 -37968 8 OUT
port 36 nsew
rlabel metal1 s 19333 -37968 19408 -37893 8 OUT
port 36 nsew
rlabel metal1 s 17738 -37931 17917 -37893 8 OUT
port 36 nsew
rlabel metal1 s 17738 -37893 19408 -37818 8 OUT
port 36 nsew
rlabel metal1 s 17738 -37818 17917 -37742 8 OUT
port 36 nsew
rlabel metal1 s 15894 -36974 26272 -36956 8 OUT
port 36 nsew
rlabel metal1 s 26895 -36908 27108 -36868 8 OUT
port 36 nsew
rlabel metal1 s 26895 -36868 28333 -36814 8 OUT
port 36 nsew
rlabel metal1 s 26895 -36814 27108 -36775 8 OUT
port 36 nsew
rlabel metal1 s 15894 -36956 26307 -36662 8 OUT
port 36 nsew
rlabel metal1 s 10557 -43995 10852 -36705 8 OUT
port 36 nsew
rlabel metal1 s 9127 -42210 9318 -42103 8 OUT
port 36 nsew
rlabel metal1 s 9247 -42103 9298 -42032 8 OUT
port 36 nsew
rlabel metal1 s -665 -42032 9298 -41981 8 OUT
port 36 nsew
rlabel metal1 s 9247 -41981 9298 -37145 8 OUT
port 36 nsew
rlabel metal1 s -3231 -40975 -3099 -40915 2 OUT
port 36 nsew
rlabel metal1 s -4128 -41422 -4068 -40974 2 OUT
port 36 nsew
rlabel metal1 s -3202 -40915 -3142 -40551 2 OUT
port 36 nsew
rlabel metal1 s -4177 -40974 -4040 -40914 2 OUT
port 36 nsew
rlabel metal1 s -5914 -38590 -5854 -38123 2 OUT
port 36 nsew
rlabel metal1 s -5950 -38123 -5818 -38063 2 OUT
port 36 nsew
rlabel metal1 s -23486 -46358 -23350 -37433 2 OUT
port 36 nsew
rlabel metal1 s -23486 -37433 -23246 -37390 2 OUT
port 36 nsew
rlabel metal1 s -23486 -37390 -23233 -37202 2 OUT
port 36 nsew
rlabel metal1 s -23334 -37202 -23233 -37147 2 OUT
port 36 nsew
rlabel metal1 s -665 -37145 9298 -37094 8 OUT
port 36 nsew
rlabel metal1 s 15894 -36662 26127 -36622 8 OUT
port 36 nsew
rlabel metal1 s 60423 -10731 61454 -9617 8 OUT
port 36 nsew
rlabel metal1 s -29580 -46472 -28157 -10506 2 OUT
port 36 nsew
rlabel metal1 s 60549 -9617 61159 -228 8 OUT
port 36 nsew
rlabel metal1 s 54401 -1085 54447 -584 8 OUT
port 36 nsew
rlabel metal1 s 54165 -1085 54211 -584 8 OUT
port 36 nsew
rlabel metal1 s 53929 -1085 53975 -584 8 OUT
port 36 nsew
rlabel metal1 s 53693 -1085 53739 -584 8 OUT
port 36 nsew
rlabel metal1 s 53457 -1085 53503 -584 8 OUT
port 36 nsew
rlabel metal1 s 53221 -1085 53267 -584 8 OUT
port 36 nsew
rlabel metal1 s 52985 -1085 53031 -584 8 OUT
port 36 nsew
rlabel metal1 s 52749 -1085 52795 -584 8 OUT
port 36 nsew
rlabel metal1 s 52749 -584 54447 -538 8 OUT
port 36 nsew
rlabel metal1 s 54401 -538 54447 -422 8 OUT
port 36 nsew
rlabel metal1 s 54355 -422 58232 -348 8 OUT
port 36 nsew
rlabel metal1 s 58157 -348 58203 123 8 OUT
port 36 nsew
rlabel metal1 s 57921 -348 57967 123 8 OUT
port 36 nsew
rlabel metal1 s 57685 -348 57731 123 8 OUT
port 36 nsew
rlabel metal1 s 57449 -348 57495 123 8 OUT
port 36 nsew
rlabel metal1 s 57213 -348 57259 123 8 OUT
port 36 nsew
rlabel metal1 s 56977 -348 57023 123 8 OUT
port 36 nsew
rlabel metal1 s 56741 -348 56787 123 8 OUT
port 36 nsew
rlabel metal1 s 56505 -348 56551 123 8 OUT
port 36 nsew
rlabel metal1 s 56269 -348 56315 123 8 OUT
port 36 nsew
rlabel metal1 s 56033 -348 56079 123 8 OUT
port 36 nsew
rlabel metal1 s 55797 -348 55843 123 8 OUT
port 36 nsew
rlabel metal1 s 55561 -348 55607 123 8 OUT
port 36 nsew
rlabel metal1 s 55325 -348 55371 123 8 OUT
port 36 nsew
rlabel metal1 s 55089 -348 55135 123 8 OUT
port 36 nsew
rlabel metal1 s 54853 -348 54899 123 8 OUT
port 36 nsew
rlabel metal1 s 54617 -348 54663 123 8 OUT
port 36 nsew
rlabel metal1 s 54381 -348 54427 123 8 OUT
port 36 nsew
rlabel locali s -23503 -46536 -23290 -46526 2 OUT
port 36 nsew
rlabel locali s -29580 -46526 10852 -46390 2 OUT
port 36 nsew
rlabel locali s -23503 -46390 -23290 -46358 2 OUT
port 36 nsew
rlabel locali s -29580 -46390 -28157 -45411 2 OUT
port 36 nsew
rlabel locali s 79621 -44314 80021 -44076 8 OUT
port 36 nsew
rlabel locali s 79670 -44076 79964 -38632 8 OUT
port 36 nsew
rlabel locali s 70668 -44318 71050 -44073 8 OUT
port 36 nsew
rlabel locali s 61363 -44308 61711 -44076 8 OUT
port 36 nsew
rlabel locali s 52864 -44296 53096 -44091 8 OUT
port 36 nsew
rlabel locali s 43525 -44269 43777 -44130 8 OUT
port 36 nsew
rlabel locali s 70753 -44073 70938 -38665 8 OUT
port 36 nsew
rlabel locali s 61425 -44076 61664 -38691 8 OUT
port 36 nsew
rlabel locali s 52898 -44091 53044 -38723 8 OUT
port 36 nsew
rlabel locali s 43579 -44130 43725 -38815 8 OUT
port 36 nsew
rlabel locali s 34828 -44315 35102 -44112 8 OUT
port 36 nsew
rlabel locali s 81317 -38567 81452 -38559 8 OUT
port 36 nsew
rlabel locali s 81297 -38559 81452 -38557 8 OUT
port 36 nsew
rlabel locali s 79670 -38632 80878 -38557 8 OUT
port 36 nsew
rlabel locali s 79670 -38557 81452 -38521 8 OUT
port 36 nsew
rlabel locali s 71953 -38605 72088 -38597 8 OUT
port 36 nsew
rlabel locali s 71933 -38597 72088 -38595 8 OUT
port 36 nsew
rlabel locali s 70753 -38665 71417 -38595 8 OUT
port 36 nsew
rlabel locali s 70753 -38595 72088 -38559 8 OUT
port 36 nsew
rlabel locali s 62800 -38622 62935 -38614 8 OUT
port 36 nsew
rlabel locali s 62780 -38614 62935 -38612 8 OUT
port 36 nsew
rlabel locali s 61425 -38691 62351 -38612 8 OUT
port 36 nsew
rlabel locali s 54046 -38688 54181 -38680 8 OUT
port 36 nsew
rlabel locali s 54026 -38680 54181 -38678 8 OUT
port 36 nsew
rlabel locali s 52898 -38723 53627 -38678 8 OUT
port 36 nsew
rlabel locali s 52898 -38678 54181 -38642 8 OUT
port 36 nsew
rlabel locali s 44848 -38722 44983 -38714 8 OUT
port 36 nsew
rlabel locali s 44828 -38714 44983 -38712 8 OUT
port 36 nsew
rlabel locali s 43579 -38815 44346 -38712 8 OUT
port 36 nsew
rlabel locali s 34897 -44112 35043 -38729 8 OUT
port 36 nsew
rlabel locali s 26602 -44292 26823 -44097 8 OUT
port 36 nsew
rlabel locali s 9583 -44236 9711 -44057 8 OUT
port 36 nsew
rlabel locali s 13526 -43501 13694 -43490 8 OUT
port 36 nsew
rlabel locali s 13526 -43490 13754 -43427 8 OUT
port 36 nsew
rlabel locali s 13694 -43427 13754 -43268 8 OUT
port 36 nsew
rlabel locali s 14592 -43037 14729 -43026 8 OUT
port 36 nsew
rlabel locali s 13651 -43036 13783 -43026 8 OUT
port 36 nsew
rlabel locali s 10557 -43092 10852 -43026 8 OUT
port 36 nsew
rlabel locali s 10557 -43026 16908 -42987 8 OUT
port 36 nsew
rlabel locali s 14592 -42987 14729 -42977 8 OUT
port 36 nsew
rlabel locali s 13651 -42987 13783 -42976 8 OUT
port 36 nsew
rlabel locali s 14740 -42593 14908 -42588 8 OUT
port 36 nsew
rlabel locali s 14620 -42661 14680 -42588 8 OUT
port 36 nsew
rlabel locali s 11178 -42987 11217 -42593 8 OUT
port 36 nsew
rlabel locali s 10557 -42987 10852 -42889 8 OUT
port 36 nsew
rlabel locali s 14620 -42588 14908 -42530 8 OUT
port 36 nsew
rlabel locali s 14740 -42530 14908 -42519 8 OUT
port 36 nsew
rlabel locali s 14620 -42530 14680 -42529 8 OUT
port 36 nsew
rlabel locali s 11158 -42593 11326 -42519 8 OUT
port 36 nsew
rlabel locali s 9607 -44057 9690 -42192 8 OUT
port 36 nsew
rlabel locali s 9127 -42210 9318 -42192 8 OUT
port 36 nsew
rlabel locali s 9127 -42192 9690 -42109 8 OUT
port 36 nsew
rlabel locali s 9127 -42109 9318 -42103 8 OUT
port 36 nsew
rlabel locali s -665 -42032 -528 -41981 2 OUT
port 36 nsew
rlabel locali s -665 -41981 -626 -41432 2 OUT
port 36 nsew
rlabel locali s -774 -41432 -606 -41358 2 OUT
port 36 nsew
rlabel locali s -4128 -41422 -4068 -41421 2 OUT
port 36 nsew
rlabel locali s -4356 -41432 -4188 -41421 2 OUT
port 36 nsew
rlabel locali s -4356 -41421 -4068 -41363 2 OUT
port 36 nsew
rlabel locali s -665 -41358 -626 -40964 2 OUT
port 36 nsew
rlabel locali s -4128 -41363 -4068 -41290 2 OUT
port 36 nsew
rlabel locali s -4356 -41363 -4188 -41358 2 OUT
port 36 nsew
rlabel locali s -3231 -40975 -3099 -40964 2 OUT
port 36 nsew
rlabel locali s -4177 -40974 -4040 -40964 2 OUT
port 36 nsew
rlabel locali s -6356 -40964 -626 -40925 2 OUT
port 36 nsew
rlabel locali s -3231 -40925 -3099 -40915 2 OUT
port 36 nsew
rlabel locali s -4177 -40925 -4040 -40914 2 OUT
port 36 nsew
rlabel locali s -3202 -40683 -3142 -40524 2 OUT
port 36 nsew
rlabel locali s -3202 -40524 -2974 -40461 2 OUT
port 36 nsew
rlabel locali s -3142 -40461 -2974 -40450 2 OUT
port 36 nsew
rlabel locali s 22868 -38945 23036 -38934 8 OUT
port 36 nsew
rlabel locali s 22748 -38935 22808 -38934 8 OUT
port 36 nsew
rlabel locali s 22748 -38934 23036 -38876 8 OUT
port 36 nsew
rlabel locali s 22868 -38876 23036 -38871 8 OUT
port 36 nsew
rlabel locali s 22748 -38876 22808 -38803 8 OUT
port 36 nsew
rlabel locali s 19286 -38945 19454 -38871 8 OUT
port 36 nsew
rlabel locali s 43579 -38712 44983 -38676 8 OUT
port 36 nsew
rlabel locali s 44828 -38676 44983 -38674 8 OUT
port 36 nsew
rlabel locali s 44848 -38674 44983 -38668 8 OUT
port 36 nsew
rlabel locali s 43579 -38676 44346 -38669 8 OUT
port 36 nsew
rlabel locali s 35985 -38683 36120 -38675 8 OUT
port 36 nsew
rlabel locali s 35965 -38675 36120 -38673 8 OUT
port 36 nsew
rlabel locali s 34897 -38729 35545 -38673 8 OUT
port 36 nsew
rlabel locali s 54026 -38642 54181 -38640 8 OUT
port 36 nsew
rlabel locali s 54046 -38640 54181 -38634 8 OUT
port 36 nsew
rlabel locali s 61425 -38612 62935 -38576 8 OUT
port 36 nsew
rlabel locali s 52898 -38642 53627 -38577 8 OUT
port 36 nsew
rlabel locali s 34897 -38673 36120 -38637 8 OUT
port 36 nsew
rlabel locali s 26896 -38735 27155 -38720 8 OUT
port 36 nsew
rlabel locali s 35965 -38637 36120 -38635 8 OUT
port 36 nsew
rlabel locali s 35985 -38635 36120 -38629 8 OUT
port 36 nsew
rlabel locali s 34897 -38637 35545 -38583 8 OUT
port 36 nsew
rlabel locali s 27545 -38672 27680 -38664 8 OUT
port 36 nsew
rlabel locali s 27525 -38664 27680 -38662 8 OUT
port 36 nsew
rlabel locali s 26030 -38720 27155 -38662 8 OUT
port 36 nsew
rlabel locali s 26030 -38662 27680 -38626 8 OUT
port 36 nsew
rlabel locali s 27525 -38626 27680 -38624 8 OUT
port 36 nsew
rlabel locali s 27545 -38624 27680 -38618 8 OUT
port 36 nsew
rlabel locali s 62780 -38576 62935 -38574 8 OUT
port 36 nsew
rlabel locali s 62800 -38574 62935 -38568 8 OUT
port 36 nsew
rlabel locali s 71933 -38559 72088 -38557 8 OUT
port 36 nsew
rlabel locali s 71953 -38557 72088 -38551 8 OUT
port 36 nsew
rlabel locali s 81297 -38521 81452 -38519 8 OUT
port 36 nsew
rlabel locali s 81317 -38519 81452 -38513 8 OUT
port 36 nsew
rlabel locali s 79670 -38521 80878 -38338 8 OUT
port 36 nsew
rlabel locali s 70753 -38559 71417 -38480 8 OUT
port 36 nsew
rlabel locali s 61425 -38576 62351 -38452 8 OUT
port 36 nsew
rlabel locali s 26030 -38626 27155 -38515 8 OUT
port 36 nsew
rlabel locali s 26896 -38515 27155 -38472 8 OUT
port 36 nsew
rlabel locali s 22720 -38487 22857 -38477 8 OUT
port 36 nsew
rlabel locali s 21779 -38488 21911 -38477 8 OUT
port 36 nsew
rlabel locali s 19306 -38871 19345 -38477 8 OUT
port 36 nsew
rlabel locali s -5842 -38676 -5674 -38665 2 OUT
port 36 nsew
rlabel locali s -5877 -38665 -5674 -38664 2 OUT
port 36 nsew
rlabel locali s -5914 -38664 -5674 -38602 2 OUT
port 36 nsew
rlabel locali s 19306 -38477 25036 -38438 8 OUT
port 36 nsew
rlabel locali s -5914 -38602 -5854 -38458 2 OUT
port 36 nsew
rlabel locali s 22720 -38438 22857 -38427 8 OUT
port 36 nsew
rlabel locali s 21779 -38438 21911 -38428 8 OUT
port 36 nsew
rlabel locali s 21822 -38196 21882 -38037 8 OUT
port 36 nsew
rlabel locali s 19306 -38438 19412 -38103 8 OUT
port 36 nsew
rlabel locali s -5950 -38123 -5818 -38115 2 OUT
port 36 nsew
rlabel locali s 21654 -38037 21882 -37974 8 OUT
port 36 nsew
rlabel locali s 21654 -37974 21822 -37963 8 OUT
port 36 nsew
rlabel locali s 19306 -38103 19438 -37968 8 OUT
port 36 nsew
rlabel locali s -6356 -38115 -626 -38076 2 OUT
port 36 nsew
rlabel locali s 17738 -37931 17917 -37742 8 OUT
port 36 nsew
rlabel locali s -665 -38076 -626 -37768 2 OUT
port 36 nsew
rlabel locali s -2259 -38076 -2184 -37953 2 OUT
port 36 nsew
rlabel locali s -5950 -38076 -5818 -38063 2 OUT
port 36 nsew
rlabel locali s -2259 -37953 -2185 -37794 2 OUT
port 36 nsew
rlabel locali s 28544 -37324 28679 -37318 8 OUT
port 36 nsew
rlabel locali s 28524 -37318 28679 -37316 8 OUT
port 36 nsew
rlabel locali s 28317 -37316 28679 -37280 8 OUT
port 36 nsew
rlabel locali s 28524 -37280 28679 -37278 8 OUT
port 36 nsew
rlabel locali s 28544 -37278 28679 -37270 8 OUT
port 36 nsew
rlabel locali s 25977 -36956 26307 -36924 8 OUT
port 36 nsew
rlabel locali s 25977 -36924 27156 -36745 8 OUT
port 36 nsew
rlabel locali s 17775 -37742 17917 -36885 8 OUT
port 36 nsew
rlabel locali s -774 -37768 -606 -37694 2 OUT
port 36 nsew
rlabel locali s -1656 -37768 -1488 -37763 2 OUT
port 36 nsew
rlabel locali s -1656 -37763 -1453 -37705 2 OUT
port 36 nsew
rlabel locali s -1656 -37705 -1488 -37694 2 OUT
port 36 nsew
rlabel locali s -665 -37694 -626 -37145 2 OUT
port 36 nsew
rlabel locali s -23334 -37390 -23233 -37383 2 OUT
port 36 nsew
rlabel locali s -665 -37145 -528 -37094 2 OUT
port 36 nsew
rlabel locali s -23334 -37383 -18767 -37320 2 OUT
port 36 nsew
rlabel locali s 10557 -36952 16076 -36950 8 OUT
port 36 nsew
rlabel locali s 25977 -36745 26307 -36662 8 OUT
port 36 nsew
rlabel locali s 17736 -36885 17954 -36639 8 OUT
port 36 nsew
rlabel locali s 10557 -36950 16200 -36705 8 OUT
port 36 nsew
rlabel locali s -18490 -36812 -18355 -36806 2 OUT
port 36 nsew
rlabel locali s -18510 -36806 -18355 -36804 2 OUT
port 36 nsew
rlabel locali s -18824 -37320 -18767 -36804 2 OUT
port 36 nsew
rlabel locali s -23334 -37320 -23233 -37147 2 OUT
port 36 nsew
rlabel locali s -18901 -36804 -18355 -36768 2 OUT
port 36 nsew
rlabel locali s -18510 -36768 -18355 -36766 2 OUT
port 36 nsew
rlabel locali s -18490 -36766 -18355 -36758 2 OUT
port 36 nsew
rlabel locali s 15965 -36705 16200 -36682 8 OUT
port 36 nsew
rlabel locali s -34369 -13296 -28472 -12595 2 OUT
port 36 nsew
rlabel locali s -29173 -12595 -28472 -11751 2 OUT
port 36 nsew
rlabel locali s 60423 -10731 61454 -10681 8 OUT
port 36 nsew
rlabel locali s -29564 -11751 -28286 -10681 2 OUT
port 36 nsew
rlabel locali s -29564 -10681 61454 -10522 8 OUT
port 36 nsew
rlabel locali s -29347 -10522 61454 -9983 8 OUT
port 36 nsew
rlabel locali s 60423 -9983 61454 -9617 8 OUT
port 36 nsew
rlabel locali s -29173 -9983 -28472 -9982 2 OUT
port 36 nsew
rlabel locali s 54407 -1089 54441 -681 8 OUT
port 36 nsew
rlabel locali s 54171 -1089 54205 -681 8 OUT
port 36 nsew
rlabel locali s 53935 -1089 53969 -681 8 OUT
port 36 nsew
rlabel locali s 53699 -1089 53733 -681 8 OUT
port 36 nsew
rlabel locali s 53463 -1089 53497 -681 8 OUT
port 36 nsew
rlabel locali s 53227 -1089 53261 -681 8 OUT
port 36 nsew
rlabel locali s 52991 -1089 53025 -681 8 OUT
port 36 nsew
rlabel locali s 52755 -1089 52789 -681 8 OUT
port 36 nsew
rlabel locali s 60613 -669 61078 -618 8 OUT
port 36 nsew
rlabel locali s 58324 -618 61078 -461 8 OUT
port 36 nsew
rlabel locali s 58163 -461 61078 -427 8 OUT
port 36 nsew
rlabel locali s 60613 -427 61078 -338 8 OUT
port 36 nsew
rlabel locali s 58163 -427 58197 127 8 OUT
port 36 nsew
rlabel locali s 57927 -281 57961 127 8 OUT
port 36 nsew
rlabel locali s 57691 -281 57725 127 8 OUT
port 36 nsew
rlabel locali s 57455 -281 57489 127 8 OUT
port 36 nsew
rlabel locali s 57219 -281 57253 127 8 OUT
port 36 nsew
rlabel locali s 56983 -281 57017 127 8 OUT
port 36 nsew
rlabel locali s 56747 -281 56781 127 8 OUT
port 36 nsew
rlabel locali s 56511 -281 56545 127 8 OUT
port 36 nsew
rlabel locali s 56275 -281 56309 127 8 OUT
port 36 nsew
rlabel locali s 56039 -281 56073 127 8 OUT
port 36 nsew
rlabel locali s 55803 -281 55837 127 8 OUT
port 36 nsew
rlabel locali s 55567 -281 55601 127 8 OUT
port 36 nsew
rlabel locali s 55331 -281 55365 127 8 OUT
port 36 nsew
rlabel locali s 55095 -281 55129 127 8 OUT
port 36 nsew
rlabel locali s 54859 -281 54893 127 8 OUT
port 36 nsew
rlabel locali s 54623 -281 54657 127 8 OUT
port 36 nsew
rlabel locali s 54387 -281 54421 127 8 OUT
port 36 nsew
rlabel metal1 s -8007 767 -7961 1268 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -8243 767 -8197 1268 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -8479 767 -8433 1268 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -8715 767 -8669 1268 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -8951 767 -8905 1268 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -9187 767 -9141 1268 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -9423 767 -9377 1268 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -9659 767 -9613 1268 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -9659 1268 -7961 1314 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -9659 1314 -9613 1430 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -13444 1430 -9567 1504 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -9639 1504 -9593 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -9875 1504 -9829 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -10111 1504 -10065 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -10347 1504 -10301 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -10583 1504 -10537 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -10819 1504 -10773 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -11055 1504 -11009 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -11291 1504 -11245 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -11527 1504 -11481 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -11763 1504 -11717 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -11999 1504 -11953 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -12235 1504 -12189 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -12471 1504 -12425 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -12707 1504 -12661 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -12943 1504 -12897 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -13179 1504 -13133 1975 4 PRE_SCALAR
port 37 nsew
rlabel metal1 s -13415 1504 -13369 1975 4 PRE_SCALAR
port 37 nsew
rlabel locali s -8001 763 -7967 1171 4 PRE_SCALAR
port 37 nsew
rlabel locali s -8237 763 -8203 1171 4 PRE_SCALAR
port 37 nsew
rlabel locali s -8473 763 -8439 1171 4 PRE_SCALAR
port 37 nsew
rlabel locali s -8709 763 -8675 1171 4 PRE_SCALAR
port 37 nsew
rlabel locali s -8945 763 -8911 1171 4 PRE_SCALAR
port 37 nsew
rlabel locali s -9181 763 -9147 1171 4 PRE_SCALAR
port 37 nsew
rlabel locali s -9417 763 -9383 1171 4 PRE_SCALAR
port 37 nsew
rlabel locali s -9653 763 -9619 1171 4 PRE_SCALAR
port 37 nsew
rlabel locali s -22664 1391 -13375 1425 4 PRE_SCALAR
port 37 nsew
rlabel locali s -9633 1571 -9599 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -9869 1571 -9835 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -10105 1571 -10071 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -10341 1571 -10307 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -10577 1571 -10543 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -10813 1571 -10779 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -11049 1571 -11015 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -11285 1571 -11251 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -11521 1571 -11487 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -11757 1571 -11723 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -11993 1571 -11959 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -12229 1571 -12195 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -12465 1571 -12431 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -12701 1571 -12667 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -12937 1571 -12903 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -13173 1571 -13139 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -13409 1425 -13375 1979 4 PRE_SCALAR
port 37 nsew
rlabel locali s -22962 160 -3643 212 4 S1
port 38 nsew
rlabel locali s -2846 1030 -2678 1038 4 S1
port 38 nsew
rlabel locali s -3695 212 -3643 1038 4 S1
port 38 nsew
rlabel locali s -3699 1038 -2678 1090 4 S1
port 38 nsew
rlabel locali s -2846 1090 -2678 1104 4 S1
port 38 nsew
rlabel locali s -3699 1090 -3647 1695 4 S1
port 38 nsew
rlabel locali s -3827 1695 -3528 1769 4 S1
port 38 nsew
rlabel metal1 s 62246 -13180 63072 -12441 8 S7
port 39 nsew
rlabel metal1 s 62465 -12441 62732 -4139 8 S7
port 39 nsew
rlabel metal1 s 62432 -4139 62779 -3786 8 S7
port 39 nsew
rlabel locali s -34505 -14566 -26421 -13991 2 S7
port 39 nsew
rlabel locali s 62246 -13180 63072 -13121 8 S7
port 39 nsew
rlabel locali s -26996 -13991 -26421 -13121 2 S7
port 39 nsew
rlabel locali s -26996 -13121 63072 -12546 8 S7
port 39 nsew
rlabel locali s 62246 -12546 63072 -12441 8 S7
port 39 nsew
rlabel locali s 63131 -3845 63299 -3837 8 S7
port 39 nsew
rlabel locali s 62432 -4139 62779 -3837 8 S7
port 39 nsew
rlabel locali s 62278 -3837 63299 -3785 8 S7
port 39 nsew
rlabel locali s 63131 -3785 63299 -3771 8 S7
port 39 nsew
rlabel locali s 62278 -3785 62330 -3180 8 S7
port 39 nsew
rlabel locali s 62150 -3180 62449 -3106 8 S7
port 39 nsew
rlabel metal1 s -11279 -16536 -11233 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -11515 -16536 -11469 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -11751 -16536 -11705 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -11987 -16536 -11941 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -12223 -16536 -12177 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -12459 -16536 -12413 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -12695 -16536 -12649 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -12931 -16536 -12885 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -13167 -16536 -13121 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -13403 -16536 -13357 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -13639 -16536 -13593 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -13875 -16536 -13829 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -14111 -16536 -14065 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -14347 -16536 -14301 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -14583 -16536 -14537 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -14819 -16536 -14773 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -15055 -16536 -15009 -16065 2 DIV_OUT
port 40 nsew
rlabel metal1 s -15084 -16065 -11207 -15991 2 DIV_OUT
port 40 nsew
rlabel metal1 s -11299 -15991 -11253 -15875 2 DIV_OUT
port 40 nsew
rlabel metal1 s -11299 -15875 -9601 -15829 2 DIV_OUT
port 40 nsew
rlabel metal1 s -9647 -15829 -9601 -15328 2 DIV_OUT
port 40 nsew
rlabel metal1 s -9883 -15829 -9837 -15328 2 DIV_OUT
port 40 nsew
rlabel metal1 s -10119 -15829 -10073 -15328 2 DIV_OUT
port 40 nsew
rlabel metal1 s -10355 -15829 -10309 -15328 2 DIV_OUT
port 40 nsew
rlabel metal1 s -10591 -15829 -10545 -15328 2 DIV_OUT
port 40 nsew
rlabel metal1 s -10827 -15829 -10781 -15328 2 DIV_OUT
port 40 nsew
rlabel metal1 s -11063 -15829 -11017 -15328 2 DIV_OUT
port 40 nsew
rlabel metal1 s -11299 -15829 -11253 -15328 2 DIV_OUT
port 40 nsew
rlabel locali s -11273 -16540 -11239 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -11509 -16540 -11475 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -11745 -16540 -11711 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -11981 -16540 -11947 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -12217 -16540 -12183 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -12453 -16540 -12419 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -12689 -16540 -12655 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -12925 -16540 -12891 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -13161 -16540 -13127 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -13397 -16540 -13363 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -13633 -16540 -13599 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -13869 -16540 -13835 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -14105 -16540 -14071 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -14341 -16540 -14307 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -14577 -16540 -14543 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -14813 -16540 -14779 -16132 2 DIV_OUT
port 40 nsew
rlabel locali s -15049 -16540 -15015 -15986 2 DIV_OUT
port 40 nsew
rlabel locali s -34293 -16022 -15114 -15986 2 DIV_OUT
port 40 nsew
rlabel locali s -34293 -15986 -15015 -15952 2 DIV_OUT
port 40 nsew
rlabel locali s -34293 -15952 -15114 -15892 2 DIV_OUT
port 40 nsew
rlabel locali s -9641 -15732 -9607 -15324 2 DIV_OUT
port 40 nsew
rlabel locali s -9877 -15732 -9843 -15324 2 DIV_OUT
port 40 nsew
rlabel locali s -10113 -15732 -10079 -15324 2 DIV_OUT
port 40 nsew
rlabel locali s -10349 -15732 -10315 -15324 2 DIV_OUT
port 40 nsew
rlabel locali s -10585 -15732 -10551 -15324 2 DIV_OUT
port 40 nsew
rlabel locali s -10821 -15732 -10787 -15324 2 DIV_OUT
port 40 nsew
rlabel locali s -11057 -15732 -11023 -15324 2 DIV_OUT
port 40 nsew
rlabel locali s -11293 -15732 -11259 -15324 2 DIV_OUT
port 40 nsew
rlabel metal1 s 17782 -61880 17828 -61680 8 VDD
port 41 nsew
rlabel metal1 s 17586 -61880 17632 -61680 8 VDD
port 41 nsew
rlabel metal1 s 17390 -61880 17436 -61680 8 VDD
port 41 nsew
rlabel metal1 s 16945 -61880 16991 -61680 8 VDD
port 41 nsew
rlabel metal1 s 16749 -61880 16795 -61680 8 VDD
port 41 nsew
rlabel metal1 s 16553 -61880 16599 -61680 8 VDD
port 41 nsew
rlabel metal1 s 15082 -61880 15128 -61680 8 VDD
port 41 nsew
rlabel metal1 s 14886 -61880 14932 -61680 8 VDD
port 41 nsew
rlabel metal1 s 14690 -61880 14736 -61680 8 VDD
port 41 nsew
rlabel metal1 s 14245 -61880 14291 -61680 8 VDD
port 41 nsew
rlabel metal1 s 14049 -61880 14095 -61680 8 VDD
port 41 nsew
rlabel metal1 s 13853 -61880 13899 -61680 8 VDD
port 41 nsew
rlabel metal1 s 8737 -62043 8783 -61843 8 VDD
port 41 nsew
rlabel metal1 s 8541 -62043 8587 -61843 8 VDD
port 41 nsew
rlabel metal1 s 8428 -62043 8474 -61843 8 VDD
port 41 nsew
rlabel metal1 s 8232 -62043 8278 -61843 8 VDD
port 41 nsew
rlabel metal1 s 8118 -62043 8164 -61843 8 VDD
port 41 nsew
rlabel metal1 s 7922 -62043 7968 -61843 8 VDD
port 41 nsew
rlabel metal1 s 7726 -62043 7772 -61843 8 VDD
port 41 nsew
rlabel metal1 s 5737 -62043 5783 -61843 8 VDD
port 41 nsew
rlabel metal1 s 5541 -62043 5587 -61843 8 VDD
port 41 nsew
rlabel metal1 s 5428 -62043 5474 -61843 8 VDD
port 41 nsew
rlabel metal1 s 5232 -62043 5278 -61843 8 VDD
port 41 nsew
rlabel metal1 s 5118 -62043 5164 -61843 8 VDD
port 41 nsew
rlabel metal1 s 4922 -62043 4968 -61843 8 VDD
port 41 nsew
rlabel metal1 s 4726 -62043 4772 -61843 8 VDD
port 41 nsew
rlabel metal1 s 3237 -62043 3283 -61843 8 VDD
port 41 nsew
rlabel metal1 s 3041 -62043 3087 -61843 8 VDD
port 41 nsew
rlabel metal1 s 2928 -62043 2974 -61843 8 VDD
port 41 nsew
rlabel metal1 s 2732 -62043 2778 -61843 8 VDD
port 41 nsew
rlabel metal1 s 2618 -62043 2664 -61843 8 VDD
port 41 nsew
rlabel metal1 s 2422 -62043 2468 -61843 8 VDD
port 41 nsew
rlabel metal1 s 2226 -62043 2272 -61843 8 VDD
port 41 nsew
rlabel metal1 s 737 -62043 783 -61843 8 VDD
port 41 nsew
rlabel metal1 s 541 -62043 587 -61843 8 VDD
port 41 nsew
rlabel metal1 s 428 -62043 474 -61843 8 VDD
port 41 nsew
rlabel metal1 s 232 -62043 278 -61843 8 VDD
port 41 nsew
rlabel metal1 s 118 -62043 164 -61843 8 VDD
port 41 nsew
rlabel metal1 s -78 -62043 -32 -61843 2 VDD
port 41 nsew
rlabel metal1 s -274 -62043 -228 -61843 2 VDD
port 41 nsew
rlabel metal1 s -1763 -62043 -1717 -61843 2 VDD
port 41 nsew
rlabel metal1 s -1959 -62043 -1913 -61843 2 VDD
port 41 nsew
rlabel metal1 s -2072 -62043 -2026 -61843 2 VDD
port 41 nsew
rlabel metal1 s -2268 -62043 -2222 -61843 2 VDD
port 41 nsew
rlabel metal1 s -2382 -62043 -2336 -61843 2 VDD
port 41 nsew
rlabel metal1 s -2578 -62043 -2532 -61843 2 VDD
port 41 nsew
rlabel metal1 s -2774 -62043 -2728 -61843 2 VDD
port 41 nsew
rlabel metal1 s -4263 -62043 -4217 -61843 2 VDD
port 41 nsew
rlabel metal1 s -4459 -62043 -4413 -61843 2 VDD
port 41 nsew
rlabel metal1 s -4572 -62043 -4526 -61843 2 VDD
port 41 nsew
rlabel metal1 s -4768 -62043 -4722 -61843 2 VDD
port 41 nsew
rlabel metal1 s -4882 -62043 -4836 -61843 2 VDD
port 41 nsew
rlabel metal1 s -5078 -62043 -5032 -61843 2 VDD
port 41 nsew
rlabel metal1 s -5274 -62043 -5228 -61843 2 VDD
port 41 nsew
rlabel metal1 s -18948 -62293 -18772 -61662 2 VDD
port 41 nsew
rlabel metal1 s -20232 -62129 -20186 -61929 2 VDD
port 41 nsew
rlabel metal1 s -20428 -62129 -20382 -61929 2 VDD
port 41 nsew
rlabel metal1 s -20624 -62129 -20578 -61929 2 VDD
port 41 nsew
rlabel metal1 s -20820 -62129 -20774 -61929 2 VDD
port 41 nsew
rlabel metal1 s -21362 -62129 -21316 -61929 2 VDD
port 41 nsew
rlabel metal1 s -21558 -62129 -21512 -61929 2 VDD
port 41 nsew
rlabel metal1 s 1104 -61386 1227 -61250 8 VDD
port 41 nsew
rlabel metal1 s -1379 -61386 -1256 -61250 2 VDD
port 41 nsew
rlabel metal1 s -3946 -61421 -3823 -61285 2 VDD
port 41 nsew
rlabel metal1 s 1108 -61250 1222 -60833 8 VDD
port 41 nsew
rlabel metal1 s 1103 -60833 1226 -60832 8 VDD
port 41 nsew
rlabel metal1 s 1103 -60832 1409 -60770 8 VDD
port 41 nsew
rlabel metal1 s -1375 -61250 -1261 -60798 2 VDD
port 41 nsew
rlabel metal1 s -1380 -60798 -1257 -60662 2 VDD
port 41 nsew
rlabel metal1 s -3942 -61285 -3828 -60654 2 VDD
port 41 nsew
rlabel metal1 s -15512 -60969 -15466 -60869 2 VDD
port 41 nsew
rlabel metal1 s -15708 -60969 -15662 -60869 2 VDD
port 41 nsew
rlabel metal1 s -15904 -60969 -15858 -60869 2 VDD
port 41 nsew
rlabel metal1 s -16100 -60969 -16054 -60869 2 VDD
port 41 nsew
rlabel metal1 s -16317 -61170 -16271 -60870 2 VDD
port 41 nsew
rlabel metal1 s -16513 -61170 -16467 -60870 2 VDD
port 41 nsew
rlabel metal1 s -16709 -61170 -16663 -60870 2 VDD
port 41 nsew
rlabel metal1 s -17094 -61199 -17048 -60999 2 VDD
port 41 nsew
rlabel metal1 s -17290 -61199 -17244 -60999 2 VDD
port 41 nsew
rlabel metal1 s -17486 -61199 -17440 -60999 2 VDD
port 41 nsew
rlabel metal1 s -17682 -61199 -17636 -60999 2 VDD
port 41 nsew
rlabel metal1 s 87825 -60272 87871 -59672 8 VDD
port 41 nsew
rlabel metal1 s 87402 -60272 87448 -59672 8 VDD
port 41 nsew
rlabel metal1 s 87206 -60272 87252 -59672 8 VDD
port 41 nsew
rlabel metal1 s 86956 -59860 87002 -59760 8 VDD
port 41 nsew
rlabel metal1 s 86760 -59860 86806 -59760 8 VDD
port 41 nsew
rlabel metal1 s 86564 -59860 86610 -59760 8 VDD
port 41 nsew
rlabel metal1 s 86368 -59860 86414 -59760 8 VDD
port 41 nsew
rlabel metal1 s 86151 -60061 86197 -59761 8 VDD
port 41 nsew
rlabel metal1 s 85955 -60061 86001 -59761 8 VDD
port 41 nsew
rlabel metal1 s 85759 -60061 85805 -59761 8 VDD
port 41 nsew
rlabel metal1 s 84157 -60241 84203 -59641 8 VDD
port 41 nsew
rlabel metal1 s 83734 -60241 83780 -59641 8 VDD
port 41 nsew
rlabel metal1 s 83538 -60241 83584 -59641 8 VDD
port 41 nsew
rlabel metal1 s 83288 -59829 83334 -59729 8 VDD
port 41 nsew
rlabel metal1 s 83092 -59829 83138 -59729 8 VDD
port 41 nsew
rlabel metal1 s 82896 -59829 82942 -59729 8 VDD
port 41 nsew
rlabel metal1 s 82700 -59829 82746 -59729 8 VDD
port 41 nsew
rlabel metal1 s 82483 -60030 82529 -59730 8 VDD
port 41 nsew
rlabel metal1 s 82287 -60030 82333 -59730 8 VDD
port 41 nsew
rlabel metal1 s 82091 -60030 82137 -59730 8 VDD
port 41 nsew
rlabel metal1 s 78461 -60310 78507 -59710 8 VDD
port 41 nsew
rlabel metal1 s 78038 -60310 78084 -59710 8 VDD
port 41 nsew
rlabel metal1 s 77842 -60310 77888 -59710 8 VDD
port 41 nsew
rlabel metal1 s 77592 -59898 77638 -59798 8 VDD
port 41 nsew
rlabel metal1 s 77396 -59898 77442 -59798 8 VDD
port 41 nsew
rlabel metal1 s 77200 -59898 77246 -59798 8 VDD
port 41 nsew
rlabel metal1 s 77004 -59898 77050 -59798 8 VDD
port 41 nsew
rlabel metal1 s 76787 -60099 76833 -59799 8 VDD
port 41 nsew
rlabel metal1 s 76591 -60099 76637 -59799 8 VDD
port 41 nsew
rlabel metal1 s 76395 -60099 76441 -59799 8 VDD
port 41 nsew
rlabel metal1 s 74793 -60279 74839 -59679 8 VDD
port 41 nsew
rlabel metal1 s 74370 -60279 74416 -59679 8 VDD
port 41 nsew
rlabel metal1 s 74174 -60279 74220 -59679 8 VDD
port 41 nsew
rlabel metal1 s 73924 -59867 73970 -59767 8 VDD
port 41 nsew
rlabel metal1 s 73728 -59867 73774 -59767 8 VDD
port 41 nsew
rlabel metal1 s 73532 -59867 73578 -59767 8 VDD
port 41 nsew
rlabel metal1 s 73336 -59867 73382 -59767 8 VDD
port 41 nsew
rlabel metal1 s 73119 -60068 73165 -59768 8 VDD
port 41 nsew
rlabel metal1 s 72923 -60068 72969 -59768 8 VDD
port 41 nsew
rlabel metal1 s 72727 -60068 72773 -59768 8 VDD
port 41 nsew
rlabel metal1 s 69308 -60327 69354 -59727 8 VDD
port 41 nsew
rlabel metal1 s 68885 -60327 68931 -59727 8 VDD
port 41 nsew
rlabel metal1 s 68689 -60327 68735 -59727 8 VDD
port 41 nsew
rlabel metal1 s 68439 -59915 68485 -59815 8 VDD
port 41 nsew
rlabel metal1 s 68243 -59915 68289 -59815 8 VDD
port 41 nsew
rlabel metal1 s 68047 -59915 68093 -59815 8 VDD
port 41 nsew
rlabel metal1 s 67851 -59915 67897 -59815 8 VDD
port 41 nsew
rlabel metal1 s 67634 -60116 67680 -59816 8 VDD
port 41 nsew
rlabel metal1 s 67438 -60116 67484 -59816 8 VDD
port 41 nsew
rlabel metal1 s 67242 -60116 67288 -59816 8 VDD
port 41 nsew
rlabel metal1 s 65640 -60296 65686 -59696 8 VDD
port 41 nsew
rlabel metal1 s 65217 -60296 65263 -59696 8 VDD
port 41 nsew
rlabel metal1 s 65021 -60296 65067 -59696 8 VDD
port 41 nsew
rlabel metal1 s 64771 -59884 64817 -59784 8 VDD
port 41 nsew
rlabel metal1 s 64575 -59884 64621 -59784 8 VDD
port 41 nsew
rlabel metal1 s 64379 -59884 64425 -59784 8 VDD
port 41 nsew
rlabel metal1 s 64183 -59884 64229 -59784 8 VDD
port 41 nsew
rlabel metal1 s 63966 -60085 64012 -59785 8 VDD
port 41 nsew
rlabel metal1 s 63770 -60085 63816 -59785 8 VDD
port 41 nsew
rlabel metal1 s 63574 -60085 63620 -59785 8 VDD
port 41 nsew
rlabel metal1 s 60554 -60393 60600 -59793 8 VDD
port 41 nsew
rlabel metal1 s 60131 -60393 60177 -59793 8 VDD
port 41 nsew
rlabel metal1 s 59935 -60393 59981 -59793 8 VDD
port 41 nsew
rlabel metal1 s 59685 -59981 59731 -59881 8 VDD
port 41 nsew
rlabel metal1 s 59489 -59981 59535 -59881 8 VDD
port 41 nsew
rlabel metal1 s 59293 -59981 59339 -59881 8 VDD
port 41 nsew
rlabel metal1 s 59097 -59981 59143 -59881 8 VDD
port 41 nsew
rlabel metal1 s 58880 -60182 58926 -59882 8 VDD
port 41 nsew
rlabel metal1 s 58684 -60182 58730 -59882 8 VDD
port 41 nsew
rlabel metal1 s 58488 -60182 58534 -59882 8 VDD
port 41 nsew
rlabel metal1 s 56886 -60362 56932 -59762 8 VDD
port 41 nsew
rlabel metal1 s 56463 -60362 56509 -59762 8 VDD
port 41 nsew
rlabel metal1 s 56267 -60362 56313 -59762 8 VDD
port 41 nsew
rlabel metal1 s 56017 -59950 56063 -59850 8 VDD
port 41 nsew
rlabel metal1 s 55821 -59950 55867 -59850 8 VDD
port 41 nsew
rlabel metal1 s 55625 -59950 55671 -59850 8 VDD
port 41 nsew
rlabel metal1 s 55429 -59950 55475 -59850 8 VDD
port 41 nsew
rlabel metal1 s 55212 -60151 55258 -59851 8 VDD
port 41 nsew
rlabel metal1 s 55016 -60151 55062 -59851 8 VDD
port 41 nsew
rlabel metal1 s 54820 -60151 54866 -59851 8 VDD
port 41 nsew
rlabel metal1 s 51356 -60427 51402 -59827 8 VDD
port 41 nsew
rlabel metal1 s 50933 -60427 50979 -59827 8 VDD
port 41 nsew
rlabel metal1 s 50737 -60427 50783 -59827 8 VDD
port 41 nsew
rlabel metal1 s 50487 -60015 50533 -59915 8 VDD
port 41 nsew
rlabel metal1 s 50291 -60015 50337 -59915 8 VDD
port 41 nsew
rlabel metal1 s 50095 -60015 50141 -59915 8 VDD
port 41 nsew
rlabel metal1 s 49899 -60015 49945 -59915 8 VDD
port 41 nsew
rlabel metal1 s 49682 -60216 49728 -59916 8 VDD
port 41 nsew
rlabel metal1 s 49486 -60216 49532 -59916 8 VDD
port 41 nsew
rlabel metal1 s 49290 -60216 49336 -59916 8 VDD
port 41 nsew
rlabel metal1 s 47688 -60396 47734 -59796 8 VDD
port 41 nsew
rlabel metal1 s 47265 -60396 47311 -59796 8 VDD
port 41 nsew
rlabel metal1 s 47069 -60396 47115 -59796 8 VDD
port 41 nsew
rlabel metal1 s 46819 -59984 46865 -59884 8 VDD
port 41 nsew
rlabel metal1 s 46623 -59984 46669 -59884 8 VDD
port 41 nsew
rlabel metal1 s 46427 -59984 46473 -59884 8 VDD
port 41 nsew
rlabel metal1 s 46231 -59984 46277 -59884 8 VDD
port 41 nsew
rlabel metal1 s 46014 -60185 46060 -59885 8 VDD
port 41 nsew
rlabel metal1 s 45818 -60185 45864 -59885 8 VDD
port 41 nsew
rlabel metal1 s 45622 -60185 45668 -59885 8 VDD
port 41 nsew
rlabel metal1 s 42493 -60388 42539 -59788 8 VDD
port 41 nsew
rlabel metal1 s 42070 -60388 42116 -59788 8 VDD
port 41 nsew
rlabel metal1 s 41874 -60388 41920 -59788 8 VDD
port 41 nsew
rlabel metal1 s 41624 -59976 41670 -59876 8 VDD
port 41 nsew
rlabel metal1 s 41428 -59976 41474 -59876 8 VDD
port 41 nsew
rlabel metal1 s 41232 -59976 41278 -59876 8 VDD
port 41 nsew
rlabel metal1 s 41036 -59976 41082 -59876 8 VDD
port 41 nsew
rlabel metal1 s 40819 -60177 40865 -59877 8 VDD
port 41 nsew
rlabel metal1 s 40623 -60177 40669 -59877 8 VDD
port 41 nsew
rlabel metal1 s 40427 -60177 40473 -59877 8 VDD
port 41 nsew
rlabel metal1 s 38825 -60357 38871 -59757 8 VDD
port 41 nsew
rlabel metal1 s 38402 -60357 38448 -59757 8 VDD
port 41 nsew
rlabel metal1 s 38206 -60357 38252 -59757 8 VDD
port 41 nsew
rlabel metal1 s 37956 -59945 38002 -59845 8 VDD
port 41 nsew
rlabel metal1 s 37760 -59945 37806 -59845 8 VDD
port 41 nsew
rlabel metal1 s 37564 -59945 37610 -59845 8 VDD
port 41 nsew
rlabel metal1 s 37368 -59945 37414 -59845 8 VDD
port 41 nsew
rlabel metal1 s 37151 -60146 37197 -59846 8 VDD
port 41 nsew
rlabel metal1 s 36955 -60146 37001 -59846 8 VDD
port 41 nsew
rlabel metal1 s 36759 -60146 36805 -59846 8 VDD
port 41 nsew
rlabel metal1 s 34053 -60377 34099 -59777 8 VDD
port 41 nsew
rlabel metal1 s 33630 -60377 33676 -59777 8 VDD
port 41 nsew
rlabel metal1 s 33434 -60377 33480 -59777 8 VDD
port 41 nsew
rlabel metal1 s 17684 -60562 17730 -60362 8 VDD
port 41 nsew
rlabel metal1 s 17488 -60562 17534 -60362 8 VDD
port 41 nsew
rlabel metal1 s 17292 -60562 17338 -60362 8 VDD
port 41 nsew
rlabel metal1 s 15941 -60562 15987 -60362 8 VDD
port 41 nsew
rlabel metal1 s 15745 -60562 15791 -60362 8 VDD
port 41 nsew
rlabel metal1 s 15549 -60562 15595 -60362 8 VDD
port 41 nsew
rlabel metal1 s 14984 -60562 15030 -60362 8 VDD
port 41 nsew
rlabel metal1 s 14788 -60562 14834 -60362 8 VDD
port 41 nsew
rlabel metal1 s 14592 -60562 14638 -60362 8 VDD
port 41 nsew
rlabel metal1 s 13241 -60562 13287 -60362 8 VDD
port 41 nsew
rlabel metal1 s 13045 -60562 13091 -60362 8 VDD
port 41 nsew
rlabel metal1 s 12849 -60562 12895 -60362 8 VDD
port 41 nsew
rlabel metal1 s 12359 -60562 12405 -60362 8 VDD
port 41 nsew
rlabel metal1 s 12163 -60562 12209 -60362 8 VDD
port 41 nsew
rlabel metal1 s 11967 -60562 12013 -60362 8 VDD
port 41 nsew
rlabel metal1 s -3947 -60654 -3824 -60518 2 VDD
port 41 nsew
rlabel metal1 s -18143 -60667 -17951 -60495 2 VDD
port 41 nsew
rlabel metal1 s 33184 -59965 33230 -59865 8 VDD
port 41 nsew
rlabel metal1 s 32988 -59965 33034 -59865 8 VDD
port 41 nsew
rlabel metal1 s 32792 -59965 32838 -59865 8 VDD
port 41 nsew
rlabel metal1 s 32596 -59965 32642 -59865 8 VDD
port 41 nsew
rlabel metal1 s 32379 -60166 32425 -59866 8 VDD
port 41 nsew
rlabel metal1 s 32183 -60166 32229 -59866 8 VDD
port 41 nsew
rlabel metal1 s 31987 -60166 32033 -59866 8 VDD
port 41 nsew
rlabel metal1 s 30385 -60346 30431 -59746 8 VDD
port 41 nsew
rlabel metal1 s 29962 -60346 30008 -59746 8 VDD
port 41 nsew
rlabel metal1 s 29766 -60346 29812 -59746 8 VDD
port 41 nsew
rlabel metal1 s 29516 -59934 29562 -59834 8 VDD
port 41 nsew
rlabel metal1 s 29320 -59934 29366 -59834 8 VDD
port 41 nsew
rlabel metal1 s 29124 -59934 29170 -59834 8 VDD
port 41 nsew
rlabel metal1 s 28928 -59934 28974 -59834 8 VDD
port 41 nsew
rlabel metal1 s 28711 -60135 28757 -59835 8 VDD
port 41 nsew
rlabel metal1 s 28515 -60135 28561 -59835 8 VDD
port 41 nsew
rlabel metal1 s 28319 -60135 28365 -59835 8 VDD
port 41 nsew
rlabel metal1 s 7741 -59996 7864 -59984 8 VDD
port 41 nsew
rlabel metal1 s 6525 -59997 6648 -59984 8 VDD
port 41 nsew
rlabel metal1 s 6525 -59984 7864 -59879 8 VDD
port 41 nsew
rlabel metal1 s 7741 -59879 7864 -59860 8 VDD
port 41 nsew
rlabel metal1 s 6525 -59879 6648 -59861 8 VDD
port 41 nsew
rlabel metal1 s 5169 -60002 5292 -59991 8 VDD
port 41 nsew
rlabel metal1 s 4768 -60000 4891 -59991 8 VDD
port 41 nsew
rlabel metal1 s 4768 -59991 5292 -59884 8 VDD
port 41 nsew
rlabel metal1 s 5169 -59884 5292 -59866 8 VDD
port 41 nsew
rlabel metal1 s 4768 -59884 4891 -59864 8 VDD
port 41 nsew
rlabel metal1 s 3540 -59977 3663 -59961 8 VDD
port 41 nsew
rlabel metal1 s 173 -59989 296 -59976 8 VDD
port 41 nsew
rlabel metal1 s -121 -59988 2 -59976 2 VDD
port 41 nsew
rlabel metal1 s 3151 -59976 3274 -59961 8 VDD
port 41 nsew
rlabel metal1 s 3151 -59961 3663 -59854 8 VDD
port 41 nsew
rlabel metal1 s 3540 -59854 3663 -59841 8 VDD
port 41 nsew
rlabel metal1 s 3151 -59854 3274 -59840 8 VDD
port 41 nsew
rlabel metal1 s -121 -59976 296 -59861 8 VDD
port 41 nsew
rlabel metal1 s 173 -59861 296 -59853 8 VDD
port 41 nsew
rlabel metal1 s -121 -59861 2 -59852 2 VDD
port 41 nsew
rlabel metal1 s 51796 -59746 51947 -59721 8 VDD
port 41 nsew
rlabel metal1 s 51546 -59733 51637 -59721 8 VDD
port 41 nsew
rlabel metal1 s 60994 -59712 61145 -59687 8 VDD
port 41 nsew
rlabel metal1 s 60744 -59699 60835 -59687 8 VDD
port 41 nsew
rlabel metal1 s 78901 -59629 79052 -59604 8 VDD
port 41 nsew
rlabel metal1 s 69748 -59646 69899 -59621 8 VDD
port 41 nsew
rlabel metal1 s 69498 -59633 69589 -59621 8 VDD
port 41 nsew
rlabel metal1 s 78651 -59616 78742 -59604 8 VDD
port 41 nsew
rlabel metal1 s 88265 -59591 88416 -59566 8 VDD
port 41 nsew
rlabel metal1 s 88015 -59578 88106 -59566 8 VDD
port 41 nsew
rlabel metal1 s 88015 -59566 88416 -59427 8 VDD
port 41 nsew
rlabel metal1 s 88265 -59427 88416 -59400 8 VDD
port 41 nsew
rlabel metal1 s 88015 -59427 88106 -59415 8 VDD
port 41 nsew
rlabel metal1 s 84595 -59513 84691 -59487 8 VDD
port 41 nsew
rlabel metal1 s 83292 -59494 83475 -59487 8 VDD
port 41 nsew
rlabel metal1 s 83292 -59487 84691 -59405 8 VDD
port 41 nsew
rlabel metal1 s 78651 -59604 79052 -59465 8 VDD
port 41 nsew
rlabel metal1 s 78901 -59465 79052 -59438 8 VDD
port 41 nsew
rlabel metal1 s 78651 -59465 78742 -59453 8 VDD
port 41 nsew
rlabel metal1 s 75231 -59551 75327 -59525 8 VDD
port 41 nsew
rlabel metal1 s 73928 -59532 74111 -59525 8 VDD
port 41 nsew
rlabel metal1 s 73928 -59525 75327 -59443 8 VDD
port 41 nsew
rlabel metal1 s 69498 -59621 69899 -59482 8 VDD
port 41 nsew
rlabel metal1 s 69748 -59482 69899 -59455 8 VDD
port 41 nsew
rlabel metal1 s 69498 -59482 69589 -59470 8 VDD
port 41 nsew
rlabel metal1 s 66078 -59568 66174 -59542 8 VDD
port 41 nsew
rlabel metal1 s 64775 -59549 64958 -59542 8 VDD
port 41 nsew
rlabel metal1 s 64775 -59542 66174 -59460 8 VDD
port 41 nsew
rlabel metal1 s 60744 -59687 61145 -59548 8 VDD
port 41 nsew
rlabel metal1 s 60994 -59548 61145 -59521 8 VDD
port 41 nsew
rlabel metal1 s 60744 -59548 60835 -59536 8 VDD
port 41 nsew
rlabel metal1 s 57324 -59634 57420 -59608 8 VDD
port 41 nsew
rlabel metal1 s 56021 -59615 56204 -59608 8 VDD
port 41 nsew
rlabel metal1 s 56021 -59608 57420 -59526 8 VDD
port 41 nsew
rlabel metal1 s 51546 -59721 51947 -59582 8 VDD
port 41 nsew
rlabel metal1 s 42933 -59707 43084 -59682 8 VDD
port 41 nsew
rlabel metal1 s 42683 -59694 42774 -59682 8 VDD
port 41 nsew
rlabel metal1 s 51796 -59582 51947 -59555 8 VDD
port 41 nsew
rlabel metal1 s 51546 -59582 51637 -59570 8 VDD
port 41 nsew
rlabel metal1 s 48126 -59668 48222 -59642 8 VDD
port 41 nsew
rlabel metal1 s 46823 -59649 47006 -59642 8 VDD
port 41 nsew
rlabel metal1 s 46823 -59642 48222 -59560 8 VDD
port 41 nsew
rlabel metal1 s 48126 -59560 48222 -59531 8 VDD
port 41 nsew
rlabel metal1 s 57324 -59526 57420 -59497 8 VDD
port 41 nsew
rlabel metal1 s 56021 -59526 56204 -59485 8 VDD
port 41 nsew
rlabel metal1 s 46823 -59560 47006 -59519 8 VDD
port 41 nsew
rlabel metal1 s 42683 -59682 43084 -59543 8 VDD
port 41 nsew
rlabel metal1 s 34493 -59696 34644 -59671 8 VDD
port 41 nsew
rlabel metal1 s 34243 -59683 34334 -59671 8 VDD
port 41 nsew
rlabel metal1 s 42933 -59543 43084 -59516 8 VDD
port 41 nsew
rlabel metal1 s 42683 -59543 42774 -59531 8 VDD
port 41 nsew
rlabel metal1 s 39263 -59629 39359 -59603 8 VDD
port 41 nsew
rlabel metal1 s 37960 -59610 38143 -59603 8 VDD
port 41 nsew
rlabel metal1 s 37960 -59603 39359 -59521 8 VDD
port 41 nsew
rlabel metal1 s 39263 -59521 39359 -59492 8 VDD
port 41 nsew
rlabel metal1 s 37960 -59521 38143 -59480 8 VDD
port 41 nsew
rlabel metal1 s 34243 -59671 34644 -59532 8 VDD
port 41 nsew
rlabel metal1 s 34493 -59532 34644 -59505 8 VDD
port 41 nsew
rlabel metal1 s 34243 -59532 34334 -59520 8 VDD
port 41 nsew
rlabel metal1 s 30823 -59618 30919 -59592 8 VDD
port 41 nsew
rlabel metal1 s 29520 -59599 29703 -59592 8 VDD
port 41 nsew
rlabel metal1 s 8747 -59792 8793 -59592 8 VDD
port 41 nsew
rlabel metal1 s 8551 -59792 8597 -59592 8 VDD
port 41 nsew
rlabel metal1 s 8438 -59792 8484 -59592 8 VDD
port 41 nsew
rlabel metal1 s 8242 -59792 8288 -59592 8 VDD
port 41 nsew
rlabel metal1 s 8128 -59792 8174 -59592 8 VDD
port 41 nsew
rlabel metal1 s 7932 -59792 7978 -59592 8 VDD
port 41 nsew
rlabel metal1 s 7736 -59792 7782 -59592 8 VDD
port 41 nsew
rlabel metal1 s 6575 -59803 6621 -59603 8 VDD
port 41 nsew
rlabel metal1 s 6379 -59803 6425 -59603 8 VDD
port 41 nsew
rlabel metal1 s 6183 -59803 6229 -59603 8 VDD
port 41 nsew
rlabel metal1 s 5987 -59803 6033 -59603 8 VDD
port 41 nsew
rlabel metal1 s 5445 -59803 5491 -59603 8 VDD
port 41 nsew
rlabel metal1 s 5249 -59803 5295 -59603 8 VDD
port 41 nsew
rlabel metal1 s 29520 -59592 30919 -59510 8 VDD
port 41 nsew
rlabel metal1 s 30823 -59510 30919 -59481 8 VDD
port 41 nsew
rlabel metal1 s 29520 -59510 29703 -59469 8 VDD
port 41 nsew
rlabel metal1 s 75231 -59443 75327 -59414 8 VDD
port 41 nsew
rlabel metal1 s 84595 -59405 84691 -59376 8 VDD
port 41 nsew
rlabel metal1 s 83292 -59405 83475 -59364 8 VDD
port 41 nsew
rlabel metal1 s 73928 -59443 74111 -59402 8 VDD
port 41 nsew
rlabel metal1 s 66078 -59460 66174 -59431 8 VDD
port 41 nsew
rlabel metal1 s 64775 -59460 64958 -59419 8 VDD
port 41 nsew
rlabel metal1 s 87955 -59162 88001 -59062 8 VDD
port 41 nsew
rlabel metal1 s 87759 -59162 87805 -59062 8 VDD
port 41 nsew
rlabel metal1 s 87563 -59162 87609 -59062 8 VDD
port 41 nsew
rlabel metal1 s 87367 -59162 87413 -59062 8 VDD
port 41 nsew
rlabel metal1 s 87150 -59161 87196 -58861 8 VDD
port 41 nsew
rlabel metal1 s 86954 -59161 87000 -58861 8 VDD
port 41 nsew
rlabel metal1 s 86758 -59161 86804 -58861 8 VDD
port 41 nsew
rlabel metal1 s 86373 -59032 86419 -58832 8 VDD
port 41 nsew
rlabel metal1 s 86177 -59032 86223 -58832 8 VDD
port 41 nsew
rlabel metal1 s 85981 -59032 86027 -58832 8 VDD
port 41 nsew
rlabel metal1 s 85785 -59032 85831 -58832 8 VDD
port 41 nsew
rlabel metal1 s 84287 -59131 84333 -59031 8 VDD
port 41 nsew
rlabel metal1 s 84091 -59131 84137 -59031 8 VDD
port 41 nsew
rlabel metal1 s 83895 -59131 83941 -59031 8 VDD
port 41 nsew
rlabel metal1 s 83699 -59131 83745 -59031 8 VDD
port 41 nsew
rlabel metal1 s 83482 -59130 83528 -58830 8 VDD
port 41 nsew
rlabel metal1 s 83286 -59130 83332 -58830 8 VDD
port 41 nsew
rlabel metal1 s 83090 -59130 83136 -58830 8 VDD
port 41 nsew
rlabel metal1 s 78591 -59200 78637 -59100 8 VDD
port 41 nsew
rlabel metal1 s 78395 -59200 78441 -59100 8 VDD
port 41 nsew
rlabel metal1 s 78199 -59200 78245 -59100 8 VDD
port 41 nsew
rlabel metal1 s 78003 -59200 78049 -59100 8 VDD
port 41 nsew
rlabel metal1 s 82705 -59001 82751 -58801 8 VDD
port 41 nsew
rlabel metal1 s 82509 -59001 82555 -58801 8 VDD
port 41 nsew
rlabel metal1 s 82313 -59001 82359 -58801 8 VDD
port 41 nsew
rlabel metal1 s 82117 -59001 82163 -58801 8 VDD
port 41 nsew
rlabel metal1 s 77786 -59199 77832 -58899 8 VDD
port 41 nsew
rlabel metal1 s 77590 -59199 77636 -58899 8 VDD
port 41 nsew
rlabel metal1 s 77394 -59199 77440 -58899 8 VDD
port 41 nsew
rlabel metal1 s 77009 -59070 77055 -58870 8 VDD
port 41 nsew
rlabel metal1 s 76813 -59070 76859 -58870 8 VDD
port 41 nsew
rlabel metal1 s 76617 -59070 76663 -58870 8 VDD
port 41 nsew
rlabel metal1 s 76421 -59070 76467 -58870 8 VDD
port 41 nsew
rlabel metal1 s 74923 -59169 74969 -59069 8 VDD
port 41 nsew
rlabel metal1 s 74727 -59169 74773 -59069 8 VDD
port 41 nsew
rlabel metal1 s 74531 -59169 74577 -59069 8 VDD
port 41 nsew
rlabel metal1 s 74335 -59169 74381 -59069 8 VDD
port 41 nsew
rlabel metal1 s 74118 -59168 74164 -58868 8 VDD
port 41 nsew
rlabel metal1 s 73922 -59168 73968 -58868 8 VDD
port 41 nsew
rlabel metal1 s 73726 -59168 73772 -58868 8 VDD
port 41 nsew
rlabel metal1 s 69438 -59217 69484 -59117 8 VDD
port 41 nsew
rlabel metal1 s 69242 -59217 69288 -59117 8 VDD
port 41 nsew
rlabel metal1 s 69046 -59217 69092 -59117 8 VDD
port 41 nsew
rlabel metal1 s 68850 -59217 68896 -59117 8 VDD
port 41 nsew
rlabel metal1 s 73341 -59039 73387 -58839 8 VDD
port 41 nsew
rlabel metal1 s 73145 -59039 73191 -58839 8 VDD
port 41 nsew
rlabel metal1 s 72949 -59039 72995 -58839 8 VDD
port 41 nsew
rlabel metal1 s 72753 -59039 72799 -58839 8 VDD
port 41 nsew
rlabel metal1 s 68633 -59216 68679 -58916 8 VDD
port 41 nsew
rlabel metal1 s 68437 -59216 68483 -58916 8 VDD
port 41 nsew
rlabel metal1 s 68241 -59216 68287 -58916 8 VDD
port 41 nsew
rlabel metal1 s 67856 -59087 67902 -58887 8 VDD
port 41 nsew
rlabel metal1 s 67660 -59087 67706 -58887 8 VDD
port 41 nsew
rlabel metal1 s 67464 -59087 67510 -58887 8 VDD
port 41 nsew
rlabel metal1 s 67268 -59087 67314 -58887 8 VDD
port 41 nsew
rlabel metal1 s 65770 -59186 65816 -59086 8 VDD
port 41 nsew
rlabel metal1 s 65574 -59186 65620 -59086 8 VDD
port 41 nsew
rlabel metal1 s 65378 -59186 65424 -59086 8 VDD
port 41 nsew
rlabel metal1 s 65182 -59186 65228 -59086 8 VDD
port 41 nsew
rlabel metal1 s 64965 -59185 65011 -58885 8 VDD
port 41 nsew
rlabel metal1 s 64769 -59185 64815 -58885 8 VDD
port 41 nsew
rlabel metal1 s 64573 -59185 64619 -58885 8 VDD
port 41 nsew
rlabel metal1 s 60684 -59283 60730 -59183 8 VDD
port 41 nsew
rlabel metal1 s 60488 -59283 60534 -59183 8 VDD
port 41 nsew
rlabel metal1 s 60292 -59283 60338 -59183 8 VDD
port 41 nsew
rlabel metal1 s 60096 -59283 60142 -59183 8 VDD
port 41 nsew
rlabel metal1 s 64188 -59056 64234 -58856 8 VDD
port 41 nsew
rlabel metal1 s 63992 -59056 64038 -58856 8 VDD
port 41 nsew
rlabel metal1 s 63796 -59056 63842 -58856 8 VDD
port 41 nsew
rlabel metal1 s 63600 -59056 63646 -58856 8 VDD
port 41 nsew
rlabel metal1 s 59879 -59282 59925 -58982 8 VDD
port 41 nsew
rlabel metal1 s 59683 -59282 59729 -58982 8 VDD
port 41 nsew
rlabel metal1 s 59487 -59282 59533 -58982 8 VDD
port 41 nsew
rlabel metal1 s 59102 -59153 59148 -58953 8 VDD
port 41 nsew
rlabel metal1 s 58906 -59153 58952 -58953 8 VDD
port 41 nsew
rlabel metal1 s 58710 -59153 58756 -58953 8 VDD
port 41 nsew
rlabel metal1 s 58514 -59153 58560 -58953 8 VDD
port 41 nsew
rlabel metal1 s 57016 -59252 57062 -59152 8 VDD
port 41 nsew
rlabel metal1 s 56820 -59252 56866 -59152 8 VDD
port 41 nsew
rlabel metal1 s 56624 -59252 56670 -59152 8 VDD
port 41 nsew
rlabel metal1 s 56428 -59252 56474 -59152 8 VDD
port 41 nsew
rlabel metal1 s 56211 -59251 56257 -58951 8 VDD
port 41 nsew
rlabel metal1 s 56015 -59251 56061 -58951 8 VDD
port 41 nsew
rlabel metal1 s 55819 -59251 55865 -58951 8 VDD
port 41 nsew
rlabel metal1 s 51486 -59317 51532 -59217 8 VDD
port 41 nsew
rlabel metal1 s 51290 -59317 51336 -59217 8 VDD
port 41 nsew
rlabel metal1 s 51094 -59317 51140 -59217 8 VDD
port 41 nsew
rlabel metal1 s 50898 -59317 50944 -59217 8 VDD
port 41 nsew
rlabel metal1 s 55434 -59122 55480 -58922 8 VDD
port 41 nsew
rlabel metal1 s 55238 -59122 55284 -58922 8 VDD
port 41 nsew
rlabel metal1 s 55042 -59122 55088 -58922 8 VDD
port 41 nsew
rlabel metal1 s 54846 -59122 54892 -58922 8 VDD
port 41 nsew
rlabel metal1 s 50681 -59316 50727 -59016 8 VDD
port 41 nsew
rlabel metal1 s 50485 -59316 50531 -59016 8 VDD
port 41 nsew
rlabel metal1 s 50289 -59316 50335 -59016 8 VDD
port 41 nsew
rlabel metal1 s 49904 -59187 49950 -58987 8 VDD
port 41 nsew
rlabel metal1 s 49708 -59187 49754 -58987 8 VDD
port 41 nsew
rlabel metal1 s 49512 -59187 49558 -58987 8 VDD
port 41 nsew
rlabel metal1 s 49316 -59187 49362 -58987 8 VDD
port 41 nsew
rlabel metal1 s 47818 -59286 47864 -59186 8 VDD
port 41 nsew
rlabel metal1 s 47622 -59286 47668 -59186 8 VDD
port 41 nsew
rlabel metal1 s 47426 -59286 47472 -59186 8 VDD
port 41 nsew
rlabel metal1 s 47230 -59286 47276 -59186 8 VDD
port 41 nsew
rlabel metal1 s 47013 -59285 47059 -58985 8 VDD
port 41 nsew
rlabel metal1 s 46817 -59285 46863 -58985 8 VDD
port 41 nsew
rlabel metal1 s 46621 -59285 46667 -58985 8 VDD
port 41 nsew
rlabel metal1 s 42623 -59278 42669 -59178 8 VDD
port 41 nsew
rlabel metal1 s 42427 -59278 42473 -59178 8 VDD
port 41 nsew
rlabel metal1 s 42231 -59278 42277 -59178 8 VDD
port 41 nsew
rlabel metal1 s 42035 -59278 42081 -59178 8 VDD
port 41 nsew
rlabel metal1 s 46236 -59156 46282 -58956 8 VDD
port 41 nsew
rlabel metal1 s 46040 -59156 46086 -58956 8 VDD
port 41 nsew
rlabel metal1 s 45844 -59156 45890 -58956 8 VDD
port 41 nsew
rlabel metal1 s 45648 -59156 45694 -58956 8 VDD
port 41 nsew
rlabel metal1 s 41818 -59277 41864 -58977 8 VDD
port 41 nsew
rlabel metal1 s 41622 -59277 41668 -58977 8 VDD
port 41 nsew
rlabel metal1 s 41426 -59277 41472 -58977 8 VDD
port 41 nsew
rlabel metal1 s 41041 -59148 41087 -58948 8 VDD
port 41 nsew
rlabel metal1 s 40845 -59148 40891 -58948 8 VDD
port 41 nsew
rlabel metal1 s 40649 -59148 40695 -58948 8 VDD
port 41 nsew
rlabel metal1 s 40453 -59148 40499 -58948 8 VDD
port 41 nsew
rlabel metal1 s 38955 -59247 39001 -59147 8 VDD
port 41 nsew
rlabel metal1 s 38759 -59247 38805 -59147 8 VDD
port 41 nsew
rlabel metal1 s 38563 -59247 38609 -59147 8 VDD
port 41 nsew
rlabel metal1 s 38367 -59247 38413 -59147 8 VDD
port 41 nsew
rlabel metal1 s 38150 -59246 38196 -58946 8 VDD
port 41 nsew
rlabel metal1 s 37954 -59246 38000 -58946 8 VDD
port 41 nsew
rlabel metal1 s 37758 -59246 37804 -58946 8 VDD
port 41 nsew
rlabel metal1 s 34183 -59267 34229 -59167 8 VDD
port 41 nsew
rlabel metal1 s 33987 -59267 34033 -59167 8 VDD
port 41 nsew
rlabel metal1 s 33791 -59267 33837 -59167 8 VDD
port 41 nsew
rlabel metal1 s 33595 -59267 33641 -59167 8 VDD
port 41 nsew
rlabel metal1 s 37373 -59117 37419 -58917 8 VDD
port 41 nsew
rlabel metal1 s 37177 -59117 37223 -58917 8 VDD
port 41 nsew
rlabel metal1 s 36981 -59117 37027 -58917 8 VDD
port 41 nsew
rlabel metal1 s 36785 -59117 36831 -58917 8 VDD
port 41 nsew
rlabel metal1 s 33378 -59266 33424 -58966 8 VDD
port 41 nsew
rlabel metal1 s 33182 -59266 33228 -58966 8 VDD
port 41 nsew
rlabel metal1 s 32986 -59266 33032 -58966 8 VDD
port 41 nsew
rlabel metal1 s 32601 -59137 32647 -58937 8 VDD
port 41 nsew
rlabel metal1 s 32405 -59137 32451 -58937 8 VDD
port 41 nsew
rlabel metal1 s 32209 -59137 32255 -58937 8 VDD
port 41 nsew
rlabel metal1 s 32013 -59137 32059 -58937 8 VDD
port 41 nsew
rlabel metal1 s 30515 -59236 30561 -59136 8 VDD
port 41 nsew
rlabel metal1 s 30319 -59236 30365 -59136 8 VDD
port 41 nsew
rlabel metal1 s 30123 -59236 30169 -59136 8 VDD
port 41 nsew
rlabel metal1 s 29927 -59236 29973 -59136 8 VDD
port 41 nsew
rlabel metal1 s 29710 -59235 29756 -58935 8 VDD
port 41 nsew
rlabel metal1 s 29514 -59235 29560 -58935 8 VDD
port 41 nsew
rlabel metal1 s 29318 -59235 29364 -58935 8 VDD
port 41 nsew
rlabel metal1 s 28933 -59106 28979 -58906 8 VDD
port 41 nsew
rlabel metal1 s 28737 -59106 28783 -58906 8 VDD
port 41 nsew
rlabel metal1 s 28541 -59106 28587 -58906 8 VDD
port 41 nsew
rlabel metal1 s 28345 -59106 28391 -58906 8 VDD
port 41 nsew
rlabel metal1 s 25966 -59506 26012 -58806 8 VDD
port 41 nsew
rlabel metal1 s 25770 -59506 25816 -58806 8 VDD
port 41 nsew
rlabel metal1 s 25566 -59506 25612 -58806 8 VDD
port 41 nsew
rlabel metal1 s 25370 -59506 25416 -58806 8 VDD
port 41 nsew
rlabel metal1 s 24966 -59506 25012 -58806 8 VDD
port 41 nsew
rlabel metal1 s 24770 -59506 24816 -58806 8 VDD
port 41 nsew
rlabel metal1 s 24566 -59506 24612 -58806 8 VDD
port 41 nsew
rlabel metal1 s 24370 -59506 24416 -58806 8 VDD
port 41 nsew
rlabel metal1 s 23966 -59506 24012 -58806 8 VDD
port 41 nsew
rlabel metal1 s 23770 -59506 23816 -58806 8 VDD
port 41 nsew
rlabel metal1 s 23566 -59506 23612 -58806 8 VDD
port 41 nsew
rlabel metal1 s 23370 -59506 23416 -58806 8 VDD
port 41 nsew
rlabel metal1 s 22882 -59577 22928 -59377 8 VDD
port 41 nsew
rlabel metal1 s 22686 -59577 22732 -59377 8 VDD
port 41 nsew
rlabel metal1 s 22490 -59577 22536 -59377 8 VDD
port 41 nsew
rlabel metal1 s 21957 -59584 22003 -59384 8 VDD
port 41 nsew
rlabel metal1 s 21761 -59584 21807 -59384 8 VDD
port 41 nsew
rlabel metal1 s 21219 -59584 21265 -59384 8 VDD
port 41 nsew
rlabel metal1 s 21023 -59584 21069 -59384 8 VDD
port 41 nsew
rlabel metal1 s 20827 -59584 20873 -59384 8 VDD
port 41 nsew
rlabel metal1 s 20631 -59584 20677 -59384 8 VDD
port 41 nsew
rlabel metal1 s 19911 -59550 19957 -59150 8 VDD
port 41 nsew
rlabel metal1 s 19715 -59550 19761 -59150 8 VDD
port 41 nsew
rlabel metal1 s 18965 -59550 19011 -59150 8 VDD
port 41 nsew
rlabel metal1 s 18769 -59550 18815 -59150 8 VDD
port 41 nsew
rlabel metal1 s 4822 -59778 4868 -59478 8 VDD
port 41 nsew
rlabel metal1 s 4626 -59778 4672 -59478 8 VDD
port 41 nsew
rlabel metal1 s 4430 -59778 4476 -59478 8 VDD
port 41 nsew
rlabel metal1 s 4213 -59779 4259 -59679 8 VDD
port 41 nsew
rlabel metal1 s 4017 -59779 4063 -59679 8 VDD
port 41 nsew
rlabel metal1 s 3821 -59779 3867 -59679 8 VDD
port 41 nsew
rlabel metal1 s 3625 -59779 3671 -59679 8 VDD
port 41 nsew
rlabel metal1 s 3217 -59780 3263 -59480 8 VDD
port 41 nsew
rlabel metal1 s 3021 -59780 3067 -59480 8 VDD
port 41 nsew
rlabel metal1 s 2825 -59780 2871 -59480 8 VDD
port 41 nsew
rlabel metal1 s 2608 -59781 2654 -59681 8 VDD
port 41 nsew
rlabel metal1 s 2412 -59781 2458 -59681 8 VDD
port 41 nsew
rlabel metal1 s 2216 -59781 2262 -59681 8 VDD
port 41 nsew
rlabel metal1 s 2020 -59781 2066 -59681 8 VDD
port 41 nsew
rlabel metal1 s 1613 -59794 1659 -59594 8 VDD
port 41 nsew
rlabel metal1 s 1417 -59794 1463 -59594 8 VDD
port 41 nsew
rlabel metal1 s 1221 -59794 1267 -59594 8 VDD
port 41 nsew
rlabel metal1 s 1025 -59794 1071 -59594 8 VDD
port 41 nsew
rlabel metal1 s 483 -59794 529 -59594 8 VDD
port 41 nsew
rlabel metal1 s 287 -59794 333 -59594 8 VDD
port 41 nsew
rlabel metal1 s -55 -59811 -9 -59611 2 VDD
port 41 nsew
rlabel metal1 s -251 -59811 -205 -59611 2 VDD
port 41 nsew
rlabel metal1 s -447 -59811 -401 -59611 2 VDD
port 41 nsew
rlabel metal1 s -937 -59811 -891 -59611 2 VDD
port 41 nsew
rlabel metal1 s -1133 -59811 -1087 -59611 2 VDD
port 41 nsew
rlabel metal1 s -1329 -59811 -1283 -59611 2 VDD
port 41 nsew
rlabel metal1 s -2680 -59811 -2634 -59611 2 VDD
port 41 nsew
rlabel metal1 s -2876 -59811 -2830 -59611 2 VDD
port 41 nsew
rlabel metal1 s -3072 -59811 -3026 -59611 2 VDD
port 41 nsew
rlabel metal1 s -3637 -59811 -3591 -59611 2 VDD
port 41 nsew
rlabel metal1 s -3833 -59811 -3787 -59611 2 VDD
port 41 nsew
rlabel metal1 s -4029 -59811 -3983 -59611 2 VDD
port 41 nsew
rlabel metal1 s -5380 -59811 -5334 -59611 2 VDD
port 41 nsew
rlabel metal1 s -5576 -59811 -5530 -59611 2 VDD
port 41 nsew
rlabel metal1 s -5772 -59811 -5726 -59611 2 VDD
port 41 nsew
rlabel metal1 s -15642 -60359 -15596 -59759 2 VDD
port 41 nsew
rlabel metal1 s -16065 -60359 -16019 -59759 2 VDD
port 41 nsew
rlabel metal1 s -16261 -60359 -16215 -59759 2 VDD
port 41 nsew
rlabel metal1 s -16511 -60271 -16465 -60171 2 VDD
port 41 nsew
rlabel metal1 s -16707 -60271 -16661 -60171 2 VDD
port 41 nsew
rlabel metal1 s -16903 -60271 -16857 -60171 2 VDD
port 41 nsew
rlabel metal1 s -17099 -60271 -17053 -60171 2 VDD
port 41 nsew
rlabel metal1 s -17316 -60270 -17270 -59970 2 VDD
port 41 nsew
rlabel metal1 s -17512 -60270 -17466 -59970 2 VDD
port 41 nsew
rlabel metal1 s -17708 -60270 -17662 -59970 2 VDD
port 41 nsew
rlabel metal1 s -7929 -59544 -7883 -59344 2 VDD
port 41 nsew
rlabel metal1 s -8125 -59544 -8079 -59344 2 VDD
port 41 nsew
rlabel metal1 s -8321 -59544 -8275 -59344 2 VDD
port 41 nsew
rlabel metal1 s -8811 -59544 -8765 -59344 2 VDD
port 41 nsew
rlabel metal1 s -9007 -59544 -8961 -59344 2 VDD
port 41 nsew
rlabel metal1 s -9203 -59544 -9157 -59344 2 VDD
port 41 nsew
rlabel metal1 s -10554 -59544 -10508 -59344 2 VDD
port 41 nsew
rlabel metal1 s -10750 -59544 -10704 -59344 2 VDD
port 41 nsew
rlabel metal1 s -10946 -59544 -10900 -59344 2 VDD
port 41 nsew
rlabel metal1 s -11511 -59544 -11465 -59344 2 VDD
port 41 nsew
rlabel metal1 s -11707 -59544 -11661 -59344 2 VDD
port 41 nsew
rlabel metal1 s -11903 -59544 -11857 -59344 2 VDD
port 41 nsew
rlabel metal1 s -13254 -59544 -13208 -59344 2 VDD
port 41 nsew
rlabel metal1 s -13450 -59544 -13404 -59344 2 VDD
port 41 nsew
rlabel metal1 s -13646 -59544 -13600 -59344 2 VDD
port 41 nsew
rlabel metal1 s -18142 -60495 -18016 -58731 2 VDD
port 41 nsew
rlabel metal1 s -18914 -59441 -18868 -59041 2 VDD
port 41 nsew
rlabel metal1 s -19110 -59441 -19064 -59041 2 VDD
port 41 nsew
rlabel metal1 s -19819 -59440 -19773 -59040 2 VDD
port 41 nsew
rlabel metal1 s -20015 -59440 -19969 -59040 2 VDD
port 41 nsew
rlabel metal1 s -21025 -59711 -20979 -59111 2 VDD
port 41 nsew
rlabel metal1 s -21221 -59711 -21175 -59111 2 VDD
port 41 nsew
rlabel metal1 s -27832 -59674 -27432 -59628 2 VDD
port 41 nsew
rlabel metal1 s -27832 -59438 -27432 -59392 2 VDD
port 41 nsew
rlabel metal1 s -27832 -59202 -27432 -59156 2 VDD
port 41 nsew
rlabel metal1 s -27832 -59072 -27432 -59026 2 VDD
port 41 nsew
rlabel metal1 s -27832 -58836 -27432 -58790 2 VDD
port 41 nsew
rlabel metal1 s -1941 -58493 -1895 -58293 2 VDD
port 41 nsew
rlabel metal1 s -2137 -58493 -2091 -58293 2 VDD
port 41 nsew
rlabel metal1 s -2333 -58493 -2287 -58293 2 VDD
port 41 nsew
rlabel metal1 s -2778 -58493 -2732 -58293 2 VDD
port 41 nsew
rlabel metal1 s -2974 -58493 -2928 -58293 2 VDD
port 41 nsew
rlabel metal1 s -3170 -58493 -3124 -58293 2 VDD
port 41 nsew
rlabel metal1 s -4641 -58493 -4595 -58293 2 VDD
port 41 nsew
rlabel metal1 s -4837 -58493 -4791 -58293 2 VDD
port 41 nsew
rlabel metal1 s -5033 -58493 -4987 -58293 2 VDD
port 41 nsew
rlabel metal1 s -5478 -58493 -5432 -58293 2 VDD
port 41 nsew
rlabel metal1 s -5674 -58493 -5628 -58293 2 VDD
port 41 nsew
rlabel metal1 s -5870 -58493 -5824 -58293 2 VDD
port 41 nsew
rlabel metal1 s 22932 -58276 22978 -57876 8 VDD
port 41 nsew
rlabel metal1 s 22736 -58276 22782 -57876 8 VDD
port 41 nsew
rlabel metal1 s 22540 -58276 22586 -57876 8 VDD
port 41 nsew
rlabel metal1 s -6736 -58643 -6690 -58043 2 VDD
port 41 nsew
rlabel metal1 s -6932 -58643 -6886 -58043 2 VDD
port 41 nsew
rlabel metal1 s -7355 -58643 -7309 -58043 2 VDD
port 41 nsew
rlabel metal1 s -18169 -58731 -17990 -58564 2 VDD
port 41 nsew
rlabel metal1 s -27832 -58600 -27432 -58554 2 VDD
port 41 nsew
rlabel metal1 s -27832 -58364 -27432 -58318 2 VDD
port 41 nsew
rlabel metal1 s -9815 -58226 -9769 -58026 2 VDD
port 41 nsew
rlabel metal1 s -10011 -58226 -9965 -58026 2 VDD
port 41 nsew
rlabel metal1 s -10207 -58226 -10161 -58026 2 VDD
port 41 nsew
rlabel metal1 s -10652 -58226 -10606 -58026 2 VDD
port 41 nsew
rlabel metal1 s -10848 -58226 -10802 -58026 2 VDD
port 41 nsew
rlabel metal1 s -11044 -58226 -10998 -58026 2 VDD
port 41 nsew
rlabel metal1 s -12515 -58226 -12469 -58026 2 VDD
port 41 nsew
rlabel metal1 s -12711 -58226 -12665 -58026 2 VDD
port 41 nsew
rlabel metal1 s -12907 -58226 -12861 -58026 2 VDD
port 41 nsew
rlabel metal1 s -13352 -58226 -13306 -58026 2 VDD
port 41 nsew
rlabel metal1 s -13548 -58226 -13502 -58026 2 VDD
port 41 nsew
rlabel metal1 s -13744 -58226 -13698 -58026 2 VDD
port 41 nsew
rlabel metal1 s -27832 -58128 -27432 -58082 2 VDD
port 41 nsew
rlabel metal1 s -27832 -57998 -27432 -57952 2 VDD
port 41 nsew
rlabel metal1 s -27832 -57762 -27432 -57716 2 VDD
port 41 nsew
rlabel metal1 s -27832 -57526 -27432 -57480 2 VDD
port 41 nsew
rlabel metal1 s 25812 -57324 25858 -57124 8 VDD
port 41 nsew
rlabel metal1 s 25616 -57324 25662 -57124 8 VDD
port 41 nsew
rlabel metal1 s 25420 -57324 25466 -57124 8 VDD
port 41 nsew
rlabel metal1 s 24069 -57324 24115 -57124 8 VDD
port 41 nsew
rlabel metal1 s 23873 -57324 23919 -57124 8 VDD
port 41 nsew
rlabel metal1 s 23677 -57324 23723 -57124 8 VDD
port 41 nsew
rlabel metal1 s 23112 -57324 23158 -57124 8 VDD
port 41 nsew
rlabel metal1 s 22916 -57324 22962 -57124 8 VDD
port 41 nsew
rlabel metal1 s 22720 -57324 22766 -57124 8 VDD
port 41 nsew
rlabel metal1 s 21369 -57324 21415 -57124 8 VDD
port 41 nsew
rlabel metal1 s 21173 -57324 21219 -57124 8 VDD
port 41 nsew
rlabel metal1 s 20977 -57324 21023 -57124 8 VDD
port 41 nsew
rlabel metal1 s 20487 -57324 20533 -57124 8 VDD
port 41 nsew
rlabel metal1 s 20291 -57324 20337 -57124 8 VDD
port 41 nsew
rlabel metal1 s 20095 -57324 20141 -57124 8 VDD
port 41 nsew
rlabel metal1 s -27832 -57290 -27432 -57244 2 VDD
port 41 nsew
rlabel metal1 s 86883 -56346 86929 -56046 8 VDD
port 41 nsew
rlabel metal1 s 86687 -56346 86733 -56046 8 VDD
port 41 nsew
rlabel metal1 s 86459 -56546 86505 -56046 8 VDD
port 41 nsew
rlabel metal1 s 86329 -56546 86375 -56046 8 VDD
port 41 nsew
rlabel metal1 s 85734 -56546 85780 -56046 8 VDD
port 41 nsew
rlabel metal1 s 85538 -56546 85584 -56046 8 VDD
port 41 nsew
rlabel metal1 s 84165 -56788 84211 -56188 8 VDD
port 41 nsew
rlabel metal1 s 83742 -56788 83788 -56188 8 VDD
port 41 nsew
rlabel metal1 s 83546 -56788 83592 -56188 8 VDD
port 41 nsew
rlabel metal1 s 83296 -56376 83342 -56276 8 VDD
port 41 nsew
rlabel metal1 s 83100 -56376 83146 -56276 8 VDD
port 41 nsew
rlabel metal1 s 82904 -56376 82950 -56276 8 VDD
port 41 nsew
rlabel metal1 s 82708 -56376 82754 -56276 8 VDD
port 41 nsew
rlabel metal1 s 82491 -56577 82537 -56277 8 VDD
port 41 nsew
rlabel metal1 s 82295 -56577 82341 -56277 8 VDD
port 41 nsew
rlabel metal1 s 82099 -56577 82145 -56277 8 VDD
port 41 nsew
rlabel metal1 s 84605 -56107 84715 -56089 8 VDD
port 41 nsew
rlabel metal1 s 84377 -56095 84451 -56089 8 VDD
port 41 nsew
rlabel metal1 s 84377 -56089 84715 -55993 8 VDD
port 41 nsew
rlabel metal1 s 77519 -56384 77565 -56084 8 VDD
port 41 nsew
rlabel metal1 s 77323 -56384 77369 -56084 8 VDD
port 41 nsew
rlabel metal1 s 77095 -56584 77141 -56084 8 VDD
port 41 nsew
rlabel metal1 s 76965 -56584 77011 -56084 8 VDD
port 41 nsew
rlabel metal1 s 76370 -56584 76416 -56084 8 VDD
port 41 nsew
rlabel metal1 s 76174 -56584 76220 -56084 8 VDD
port 41 nsew
rlabel metal1 s 74801 -56826 74847 -56226 8 VDD
port 41 nsew
rlabel metal1 s 74378 -56826 74424 -56226 8 VDD
port 41 nsew
rlabel metal1 s 74182 -56826 74228 -56226 8 VDD
port 41 nsew
rlabel metal1 s 73932 -56414 73978 -56314 8 VDD
port 41 nsew
rlabel metal1 s 73736 -56414 73782 -56314 8 VDD
port 41 nsew
rlabel metal1 s 73540 -56414 73586 -56314 8 VDD
port 41 nsew
rlabel metal1 s 73344 -56414 73390 -56314 8 VDD
port 41 nsew
rlabel metal1 s 73127 -56615 73173 -56315 8 VDD
port 41 nsew
rlabel metal1 s 72931 -56615 72977 -56315 8 VDD
port 41 nsew
rlabel metal1 s 72735 -56615 72781 -56315 8 VDD
port 41 nsew
rlabel metal1 s 75241 -56145 75351 -56127 8 VDD
port 41 nsew
rlabel metal1 s 75013 -56133 75087 -56127 8 VDD
port 41 nsew
rlabel metal1 s 75013 -56127 75351 -56031 8 VDD
port 41 nsew
rlabel metal1 s 68366 -56401 68412 -56101 8 VDD
port 41 nsew
rlabel metal1 s 68170 -56401 68216 -56101 8 VDD
port 41 nsew
rlabel metal1 s 67942 -56601 67988 -56101 8 VDD
port 41 nsew
rlabel metal1 s 67812 -56601 67858 -56101 8 VDD
port 41 nsew
rlabel metal1 s 67217 -56601 67263 -56101 8 VDD
port 41 nsew
rlabel metal1 s 67021 -56601 67067 -56101 8 VDD
port 41 nsew
rlabel metal1 s 65648 -56843 65694 -56243 8 VDD
port 41 nsew
rlabel metal1 s 65225 -56843 65271 -56243 8 VDD
port 41 nsew
rlabel metal1 s 65029 -56843 65075 -56243 8 VDD
port 41 nsew
rlabel metal1 s 64779 -56431 64825 -56331 8 VDD
port 41 nsew
rlabel metal1 s 64583 -56431 64629 -56331 8 VDD
port 41 nsew
rlabel metal1 s 64387 -56431 64433 -56331 8 VDD
port 41 nsew
rlabel metal1 s 64191 -56431 64237 -56331 8 VDD
port 41 nsew
rlabel metal1 s 63974 -56632 64020 -56332 8 VDD
port 41 nsew
rlabel metal1 s 63778 -56632 63824 -56332 8 VDD
port 41 nsew
rlabel metal1 s 63582 -56632 63628 -56332 8 VDD
port 41 nsew
rlabel metal1 s 59612 -56467 59658 -56167 8 VDD
port 41 nsew
rlabel metal1 s 59416 -56467 59462 -56167 8 VDD
port 41 nsew
rlabel metal1 s 59188 -56667 59234 -56167 8 VDD
port 41 nsew
rlabel metal1 s 59058 -56667 59104 -56167 8 VDD
port 41 nsew
rlabel metal1 s 58463 -56667 58509 -56167 8 VDD
port 41 nsew
rlabel metal1 s 58267 -56667 58313 -56167 8 VDD
port 41 nsew
rlabel metal1 s 56894 -56909 56940 -56309 8 VDD
port 41 nsew
rlabel metal1 s 56471 -56909 56517 -56309 8 VDD
port 41 nsew
rlabel metal1 s 56275 -56909 56321 -56309 8 VDD
port 41 nsew
rlabel metal1 s 56025 -56497 56071 -56397 8 VDD
port 41 nsew
rlabel metal1 s 55829 -56497 55875 -56397 8 VDD
port 41 nsew
rlabel metal1 s 55633 -56497 55679 -56397 8 VDD
port 41 nsew
rlabel metal1 s 55437 -56497 55483 -56397 8 VDD
port 41 nsew
rlabel metal1 s 55220 -56698 55266 -56398 8 VDD
port 41 nsew
rlabel metal1 s 55024 -56698 55070 -56398 8 VDD
port 41 nsew
rlabel metal1 s 54828 -56698 54874 -56398 8 VDD
port 41 nsew
rlabel metal1 s 57334 -56228 57444 -56210 8 VDD
port 41 nsew
rlabel metal1 s 57106 -56216 57180 -56210 8 VDD
port 41 nsew
rlabel metal1 s 66088 -56162 66198 -56144 8 VDD
port 41 nsew
rlabel metal1 s 65860 -56150 65934 -56144 8 VDD
port 41 nsew
rlabel metal1 s 75241 -56031 75351 -55995 8 VDD
port 41 nsew
rlabel metal1 s 75013 -56031 75087 -56015 8 VDD
port 41 nsew
rlabel metal1 s 65860 -56144 66198 -56048 8 VDD
port 41 nsew
rlabel metal1 s 57106 -56210 57444 -56114 8 VDD
port 41 nsew
rlabel metal1 s 50414 -56501 50460 -56201 8 VDD
port 41 nsew
rlabel metal1 s 50218 -56501 50264 -56201 8 VDD
port 41 nsew
rlabel metal1 s 49990 -56701 50036 -56201 8 VDD
port 41 nsew
rlabel metal1 s 49860 -56701 49906 -56201 8 VDD
port 41 nsew
rlabel metal1 s 49265 -56701 49311 -56201 8 VDD
port 41 nsew
rlabel metal1 s 49069 -56701 49115 -56201 8 VDD
port 41 nsew
rlabel metal1 s 47696 -56943 47742 -56343 8 VDD
port 41 nsew
rlabel metal1 s 47273 -56943 47319 -56343 8 VDD
port 41 nsew
rlabel metal1 s 47077 -56943 47123 -56343 8 VDD
port 41 nsew
rlabel metal1 s 46827 -56531 46873 -56431 8 VDD
port 41 nsew
rlabel metal1 s 46631 -56531 46677 -56431 8 VDD
port 41 nsew
rlabel metal1 s 46435 -56531 46481 -56431 8 VDD
port 41 nsew
rlabel metal1 s 46239 -56531 46285 -56431 8 VDD
port 41 nsew
rlabel metal1 s 46022 -56732 46068 -56432 8 VDD
port 41 nsew
rlabel metal1 s 45826 -56732 45872 -56432 8 VDD
port 41 nsew
rlabel metal1 s 45630 -56732 45676 -56432 8 VDD
port 41 nsew
rlabel metal1 s 48136 -56262 48246 -56244 8 VDD
port 41 nsew
rlabel metal1 s 47908 -56250 47982 -56244 8 VDD
port 41 nsew
rlabel metal1 s 57334 -56114 57444 -56078 8 VDD
port 41 nsew
rlabel metal1 s 57106 -56114 57180 -56098 8 VDD
port 41 nsew
rlabel metal1 s 47908 -56244 48246 -56148 8 VDD
port 41 nsew
rlabel metal1 s 41551 -56462 41597 -56162 8 VDD
port 41 nsew
rlabel metal1 s 41355 -56462 41401 -56162 8 VDD
port 41 nsew
rlabel metal1 s 41127 -56662 41173 -56162 8 VDD
port 41 nsew
rlabel metal1 s 40997 -56662 41043 -56162 8 VDD
port 41 nsew
rlabel metal1 s 40402 -56662 40448 -56162 8 VDD
port 41 nsew
rlabel metal1 s 40206 -56662 40252 -56162 8 VDD
port 41 nsew
rlabel metal1 s 38833 -56904 38879 -56304 8 VDD
port 41 nsew
rlabel metal1 s 38410 -56904 38456 -56304 8 VDD
port 41 nsew
rlabel metal1 s 38214 -56904 38260 -56304 8 VDD
port 41 nsew
rlabel metal1 s 37964 -56492 38010 -56392 8 VDD
port 41 nsew
rlabel metal1 s 37768 -56492 37814 -56392 8 VDD
port 41 nsew
rlabel metal1 s 37572 -56492 37618 -56392 8 VDD
port 41 nsew
rlabel metal1 s 37376 -56492 37422 -56392 8 VDD
port 41 nsew
rlabel metal1 s 37159 -56693 37205 -56393 8 VDD
port 41 nsew
rlabel metal1 s 36963 -56693 37009 -56393 8 VDD
port 41 nsew
rlabel metal1 s 36767 -56693 36813 -56393 8 VDD
port 41 nsew
rlabel metal1 s 39273 -56223 39383 -56205 8 VDD
port 41 nsew
rlabel metal1 s 39045 -56211 39119 -56205 8 VDD
port 41 nsew
rlabel metal1 s 48136 -56148 48246 -56112 8 VDD
port 41 nsew
rlabel metal1 s 47908 -56148 47982 -56132 8 VDD
port 41 nsew
rlabel metal1 s 39045 -56205 39383 -56109 8 VDD
port 41 nsew
rlabel metal1 s 33111 -56451 33157 -56151 8 VDD
port 41 nsew
rlabel metal1 s 32915 -56451 32961 -56151 8 VDD
port 41 nsew
rlabel metal1 s 32687 -56651 32733 -56151 8 VDD
port 41 nsew
rlabel metal1 s 32557 -56651 32603 -56151 8 VDD
port 41 nsew
rlabel metal1 s 31962 -56651 32008 -56151 8 VDD
port 41 nsew
rlabel metal1 s 31766 -56651 31812 -56151 8 VDD
port 41 nsew
rlabel metal1 s 30393 -56893 30439 -56293 8 VDD
port 41 nsew
rlabel metal1 s 29970 -56893 30016 -56293 8 VDD
port 41 nsew
rlabel metal1 s 29774 -56893 29820 -56293 8 VDD
port 41 nsew
rlabel metal1 s 29524 -56481 29570 -56381 8 VDD
port 41 nsew
rlabel metal1 s 29328 -56481 29374 -56381 8 VDD
port 41 nsew
rlabel metal1 s 29132 -56481 29178 -56381 8 VDD
port 41 nsew
rlabel metal1 s 28936 -56481 28982 -56381 8 VDD
port 41 nsew
rlabel metal1 s 28719 -56682 28765 -56382 8 VDD
port 41 nsew
rlabel metal1 s 28523 -56682 28569 -56382 8 VDD
port 41 nsew
rlabel metal1 s 28327 -56682 28373 -56382 8 VDD
port 41 nsew
rlabel metal1 s 18970 -57204 19016 -56604 8 VDD
port 41 nsew
rlabel metal1 s 18774 -57204 18820 -56604 8 VDD
port 41 nsew
rlabel metal1 s -1941 -57055 -1895 -56855 2 VDD
port 41 nsew
rlabel metal1 s -2137 -57055 -2091 -56855 2 VDD
port 41 nsew
rlabel metal1 s -2333 -57055 -2287 -56855 2 VDD
port 41 nsew
rlabel metal1 s -2778 -57055 -2732 -56855 2 VDD
port 41 nsew
rlabel metal1 s -2974 -57055 -2928 -56855 2 VDD
port 41 nsew
rlabel metal1 s -3170 -57055 -3124 -56855 2 VDD
port 41 nsew
rlabel metal1 s -4641 -57055 -4595 -56855 2 VDD
port 41 nsew
rlabel metal1 s -4837 -57055 -4791 -56855 2 VDD
port 41 nsew
rlabel metal1 s -5033 -57055 -4987 -56855 2 VDD
port 41 nsew
rlabel metal1 s -5478 -57055 -5432 -56855 2 VDD
port 41 nsew
rlabel metal1 s -5674 -57055 -5628 -56855 2 VDD
port 41 nsew
rlabel metal1 s -5870 -57055 -5824 -56855 2 VDD
port 41 nsew
rlabel metal1 s -10523 -56945 -10477 -56845 2 VDD
port 41 nsew
rlabel metal1 s -10719 -56945 -10673 -56845 2 VDD
port 41 nsew
rlabel metal1 s -10915 -56945 -10869 -56845 2 VDD
port 41 nsew
rlabel metal1 s -11111 -56945 -11065 -56845 2 VDD
port 41 nsew
rlabel metal1 s -11328 -57146 -11282 -56846 2 VDD
port 41 nsew
rlabel metal1 s -11524 -57146 -11478 -56846 2 VDD
port 41 nsew
rlabel metal1 s -11720 -57146 -11674 -56846 2 VDD
port 41 nsew
rlabel metal1 s -12105 -57175 -12059 -56975 2 VDD
port 41 nsew
rlabel metal1 s -12301 -57175 -12255 -56975 2 VDD
port 41 nsew
rlabel metal1 s -12497 -57175 -12451 -56975 2 VDD
port 41 nsew
rlabel metal1 s -12693 -57175 -12647 -56975 2 VDD
port 41 nsew
rlabel metal1 s -27832 -57054 -27432 -57008 2 VDD
port 41 nsew
rlabel metal1 s -27832 -56818 -27432 -56772 2 VDD
port 41 nsew
rlabel metal1 s -27832 -56582 -27432 -56536 2 VDD
port 41 nsew
rlabel metal1 s 30833 -56212 30943 -56194 8 VDD
port 41 nsew
rlabel metal1 s 30605 -56200 30679 -56194 8 VDD
port 41 nsew
rlabel metal1 s 39273 -56109 39383 -56073 8 VDD
port 41 nsew
rlabel metal1 s 39045 -56109 39119 -56093 8 VDD
port 41 nsew
rlabel metal1 s 30605 -56194 30943 -56098 8 VDD
port 41 nsew
rlabel metal1 s 30833 -56098 30943 -56062 8 VDD
port 41 nsew
rlabel metal1 s 30605 -56098 30679 -56082 8 VDD
port 41 nsew
rlabel metal1 s 66088 -56048 66198 -56012 8 VDD
port 41 nsew
rlabel metal1 s 65860 -56048 65934 -56032 8 VDD
port 41 nsew
rlabel metal1 s 84605 -55993 84715 -55957 8 VDD
port 41 nsew
rlabel metal1 s 84377 -55993 84451 -55977 8 VDD
port 41 nsew
rlabel metal1 s 84295 -55678 84341 -55578 8 VDD
port 41 nsew
rlabel metal1 s 84099 -55678 84145 -55578 8 VDD
port 41 nsew
rlabel metal1 s 83903 -55678 83949 -55578 8 VDD
port 41 nsew
rlabel metal1 s 83707 -55678 83753 -55578 8 VDD
port 41 nsew
rlabel metal1 s 83490 -55677 83536 -55377 8 VDD
port 41 nsew
rlabel metal1 s 83294 -55677 83340 -55377 8 VDD
port 41 nsew
rlabel metal1 s 83098 -55677 83144 -55377 8 VDD
port 41 nsew
rlabel metal1 s 74931 -55716 74977 -55616 8 VDD
port 41 nsew
rlabel metal1 s 74735 -55716 74781 -55616 8 VDD
port 41 nsew
rlabel metal1 s 74539 -55716 74585 -55616 8 VDD
port 41 nsew
rlabel metal1 s 74343 -55716 74389 -55616 8 VDD
port 41 nsew
rlabel metal1 s 82713 -55548 82759 -55348 8 VDD
port 41 nsew
rlabel metal1 s 82517 -55548 82563 -55348 8 VDD
port 41 nsew
rlabel metal1 s 82321 -55548 82367 -55348 8 VDD
port 41 nsew
rlabel metal1 s 82125 -55548 82171 -55348 8 VDD
port 41 nsew
rlabel metal1 s 74126 -55715 74172 -55415 8 VDD
port 41 nsew
rlabel metal1 s 73930 -55715 73976 -55415 8 VDD
port 41 nsew
rlabel metal1 s 73734 -55715 73780 -55415 8 VDD
port 41 nsew
rlabel metal1 s 65778 -55733 65824 -55633 8 VDD
port 41 nsew
rlabel metal1 s 65582 -55733 65628 -55633 8 VDD
port 41 nsew
rlabel metal1 s 65386 -55733 65432 -55633 8 VDD
port 41 nsew
rlabel metal1 s 65190 -55733 65236 -55633 8 VDD
port 41 nsew
rlabel metal1 s 73349 -55586 73395 -55386 8 VDD
port 41 nsew
rlabel metal1 s 73153 -55586 73199 -55386 8 VDD
port 41 nsew
rlabel metal1 s 72957 -55586 73003 -55386 8 VDD
port 41 nsew
rlabel metal1 s 72761 -55586 72807 -55386 8 VDD
port 41 nsew
rlabel metal1 s 64973 -55732 65019 -55432 8 VDD
port 41 nsew
rlabel metal1 s 64777 -55732 64823 -55432 8 VDD
port 41 nsew
rlabel metal1 s 64581 -55732 64627 -55432 8 VDD
port 41 nsew
rlabel metal1 s 57024 -55799 57070 -55699 8 VDD
port 41 nsew
rlabel metal1 s 56828 -55799 56874 -55699 8 VDD
port 41 nsew
rlabel metal1 s 56632 -55799 56678 -55699 8 VDD
port 41 nsew
rlabel metal1 s 56436 -55799 56482 -55699 8 VDD
port 41 nsew
rlabel metal1 s 64196 -55603 64242 -55403 8 VDD
port 41 nsew
rlabel metal1 s 64000 -55603 64046 -55403 8 VDD
port 41 nsew
rlabel metal1 s 63804 -55603 63850 -55403 8 VDD
port 41 nsew
rlabel metal1 s 63608 -55603 63654 -55403 8 VDD
port 41 nsew
rlabel metal1 s 56219 -55798 56265 -55498 8 VDD
port 41 nsew
rlabel metal1 s 56023 -55798 56069 -55498 8 VDD
port 41 nsew
rlabel metal1 s 55827 -55798 55873 -55498 8 VDD
port 41 nsew
rlabel metal1 s 47826 -55833 47872 -55733 8 VDD
port 41 nsew
rlabel metal1 s 47630 -55833 47676 -55733 8 VDD
port 41 nsew
rlabel metal1 s 47434 -55833 47480 -55733 8 VDD
port 41 nsew
rlabel metal1 s 47238 -55833 47284 -55733 8 VDD
port 41 nsew
rlabel metal1 s 55442 -55669 55488 -55469 8 VDD
port 41 nsew
rlabel metal1 s 55246 -55669 55292 -55469 8 VDD
port 41 nsew
rlabel metal1 s 55050 -55669 55096 -55469 8 VDD
port 41 nsew
rlabel metal1 s 54854 -55669 54900 -55469 8 VDD
port 41 nsew
rlabel metal1 s 47021 -55832 47067 -55532 8 VDD
port 41 nsew
rlabel metal1 s 46825 -55832 46871 -55532 8 VDD
port 41 nsew
rlabel metal1 s 46629 -55832 46675 -55532 8 VDD
port 41 nsew
rlabel metal1 s 25910 -56006 25956 -55806 8 VDD
port 41 nsew
rlabel metal1 s 25714 -56006 25760 -55806 8 VDD
port 41 nsew
rlabel metal1 s 25518 -56006 25564 -55806 8 VDD
port 41 nsew
rlabel metal1 s 25073 -56006 25119 -55806 8 VDD
port 41 nsew
rlabel metal1 s 24877 -56006 24923 -55806 8 VDD
port 41 nsew
rlabel metal1 s 24681 -56006 24727 -55806 8 VDD
port 41 nsew
rlabel metal1 s 23210 -56006 23256 -55806 8 VDD
port 41 nsew
rlabel metal1 s 23014 -56006 23060 -55806 8 VDD
port 41 nsew
rlabel metal1 s 22818 -56006 22864 -55806 8 VDD
port 41 nsew
rlabel metal1 s 22373 -56006 22419 -55806 8 VDD
port 41 nsew
rlabel metal1 s 22177 -56006 22223 -55806 8 VDD
port 41 nsew
rlabel metal1 s 21981 -56006 22027 -55806 8 VDD
port 41 nsew
rlabel metal1 s 46244 -55703 46290 -55503 8 VDD
port 41 nsew
rlabel metal1 s 46048 -55703 46094 -55503 8 VDD
port 41 nsew
rlabel metal1 s 45852 -55703 45898 -55503 8 VDD
port 41 nsew
rlabel metal1 s 45656 -55703 45702 -55503 8 VDD
port 41 nsew
rlabel metal1 s 38963 -55794 39009 -55694 8 VDD
port 41 nsew
rlabel metal1 s 38767 -55794 38813 -55694 8 VDD
port 41 nsew
rlabel metal1 s 38571 -55794 38617 -55694 8 VDD
port 41 nsew
rlabel metal1 s 38375 -55794 38421 -55694 8 VDD
port 41 nsew
rlabel metal1 s 38158 -55793 38204 -55493 8 VDD
port 41 nsew
rlabel metal1 s 37962 -55793 38008 -55493 8 VDD
port 41 nsew
rlabel metal1 s 37766 -55793 37812 -55493 8 VDD
port 41 nsew
rlabel metal1 s 30523 -55783 30569 -55683 8 VDD
port 41 nsew
rlabel metal1 s 30327 -55783 30373 -55683 8 VDD
port 41 nsew
rlabel metal1 s 30131 -55783 30177 -55683 8 VDD
port 41 nsew
rlabel metal1 s 29935 -55783 29981 -55683 8 VDD
port 41 nsew
rlabel metal1 s 37381 -55664 37427 -55464 8 VDD
port 41 nsew
rlabel metal1 s 37185 -55664 37231 -55464 8 VDD
port 41 nsew
rlabel metal1 s 36989 -55664 37035 -55464 8 VDD
port 41 nsew
rlabel metal1 s 36793 -55664 36839 -55464 8 VDD
port 41 nsew
rlabel metal1 s 29718 -55782 29764 -55482 8 VDD
port 41 nsew
rlabel metal1 s 29522 -55782 29568 -55482 8 VDD
port 41 nsew
rlabel metal1 s 29326 -55782 29372 -55482 8 VDD
port 41 nsew
rlabel metal1 s 28941 -55653 28987 -55453 8 VDD
port 41 nsew
rlabel metal1 s 28745 -55653 28791 -55453 8 VDD
port 41 nsew
rlabel metal1 s 28549 -55653 28595 -55453 8 VDD
port 41 nsew
rlabel metal1 s 28353 -55653 28399 -55453 8 VDD
port 41 nsew
rlabel metal1 s 8747 -55756 8793 -55556 8 VDD
port 41 nsew
rlabel metal1 s 8551 -55756 8597 -55556 8 VDD
port 41 nsew
rlabel metal1 s 8438 -55756 8484 -55556 8 VDD
port 41 nsew
rlabel metal1 s 8242 -55756 8288 -55556 8 VDD
port 41 nsew
rlabel metal1 s 8128 -55756 8174 -55556 8 VDD
port 41 nsew
rlabel metal1 s 7932 -55756 7978 -55556 8 VDD
port 41 nsew
rlabel metal1 s 7736 -55756 7782 -55556 8 VDD
port 41 nsew
rlabel metal1 s 6575 -55745 6621 -55545 8 VDD
port 41 nsew
rlabel metal1 s 6379 -55745 6425 -55545 8 VDD
port 41 nsew
rlabel metal1 s 6183 -55745 6229 -55545 8 VDD
port 41 nsew
rlabel metal1 s 5987 -55745 6033 -55545 8 VDD
port 41 nsew
rlabel metal1 s 5445 -55745 5491 -55545 8 VDD
port 41 nsew
rlabel metal1 s 5249 -55745 5295 -55545 8 VDD
port 41 nsew
rlabel metal1 s 4822 -55870 4868 -55570 8 VDD
port 41 nsew
rlabel metal1 s 4626 -55870 4672 -55570 8 VDD
port 41 nsew
rlabel metal1 s 4430 -55870 4476 -55570 8 VDD
port 41 nsew
rlabel metal1 s 4213 -55669 4259 -55569 8 VDD
port 41 nsew
rlabel metal1 s 4017 -55669 4063 -55569 8 VDD
port 41 nsew
rlabel metal1 s 3821 -55669 3867 -55569 8 VDD
port 41 nsew
rlabel metal1 s 3625 -55669 3671 -55569 8 VDD
port 41 nsew
rlabel metal1 s 3217 -55868 3263 -55568 8 VDD
port 41 nsew
rlabel metal1 s 3021 -55868 3067 -55568 8 VDD
port 41 nsew
rlabel metal1 s 2825 -55868 2871 -55568 8 VDD
port 41 nsew
rlabel metal1 s 2608 -55667 2654 -55567 8 VDD
port 41 nsew
rlabel metal1 s 2412 -55667 2458 -55567 8 VDD
port 41 nsew
rlabel metal1 s 2216 -55667 2262 -55567 8 VDD
port 41 nsew
rlabel metal1 s 2020 -55667 2066 -55567 8 VDD
port 41 nsew
rlabel metal1 s 1613 -55754 1659 -55554 8 VDD
port 41 nsew
rlabel metal1 s 1417 -55754 1463 -55554 8 VDD
port 41 nsew
rlabel metal1 s 1221 -55754 1267 -55554 8 VDD
port 41 nsew
rlabel metal1 s 1025 -55754 1071 -55554 8 VDD
port 41 nsew
rlabel metal1 s 483 -55754 529 -55554 8 VDD
port 41 nsew
rlabel metal1 s 287 -55754 333 -55554 8 VDD
port 41 nsew
rlabel metal1 s -55 -55737 -9 -55537 2 VDD
port 41 nsew
rlabel metal1 s -251 -55737 -205 -55537 2 VDD
port 41 nsew
rlabel metal1 s -447 -55737 -401 -55537 2 VDD
port 41 nsew
rlabel metal1 s -937 -55737 -891 -55537 2 VDD
port 41 nsew
rlabel metal1 s -1133 -55737 -1087 -55537 2 VDD
port 41 nsew
rlabel metal1 s -1329 -55737 -1283 -55537 2 VDD
port 41 nsew
rlabel metal1 s -2680 -55737 -2634 -55537 2 VDD
port 41 nsew
rlabel metal1 s -2876 -55737 -2830 -55537 2 VDD
port 41 nsew
rlabel metal1 s -3072 -55737 -3026 -55537 2 VDD
port 41 nsew
rlabel metal1 s -3637 -55737 -3591 -55537 2 VDD
port 41 nsew
rlabel metal1 s -3833 -55737 -3787 -55537 2 VDD
port 41 nsew
rlabel metal1 s -4029 -55737 -3983 -55537 2 VDD
port 41 nsew
rlabel metal1 s -5380 -55737 -5334 -55537 2 VDD
port 41 nsew
rlabel metal1 s -5576 -55737 -5530 -55537 2 VDD
port 41 nsew
rlabel metal1 s -5772 -55737 -5726 -55537 2 VDD
port 41 nsew
rlabel metal1 s -10653 -56335 -10607 -55735 2 VDD
port 41 nsew
rlabel metal1 s -11076 -56335 -11030 -55735 2 VDD
port 41 nsew
rlabel metal1 s -11272 -56335 -11226 -55735 2 VDD
port 41 nsew
rlabel metal1 s -27832 -56346 -27432 -56300 2 VDD
port 41 nsew
rlabel metal1 s -11522 -56247 -11476 -56147 2 VDD
port 41 nsew
rlabel metal1 s -11718 -56247 -11672 -56147 2 VDD
port 41 nsew
rlabel metal1 s -11914 -56247 -11868 -56147 2 VDD
port 41 nsew
rlabel metal1 s -12110 -56247 -12064 -56147 2 VDD
port 41 nsew
rlabel metal1 s -12327 -56246 -12281 -55946 2 VDD
port 41 nsew
rlabel metal1 s -12523 -56246 -12477 -55946 2 VDD
port 41 nsew
rlabel metal1 s -12719 -56246 -12673 -55946 2 VDD
port 41 nsew
rlabel metal1 s -15512 -55969 -15466 -55869 2 VDD
port 41 nsew
rlabel metal1 s -15708 -55969 -15662 -55869 2 VDD
port 41 nsew
rlabel metal1 s -15904 -55969 -15858 -55869 2 VDD
port 41 nsew
rlabel metal1 s -16100 -55969 -16054 -55869 2 VDD
port 41 nsew
rlabel metal1 s -16317 -56170 -16271 -55870 2 VDD
port 41 nsew
rlabel metal1 s -16513 -56170 -16467 -55870 2 VDD
port 41 nsew
rlabel metal1 s -16709 -56170 -16663 -55870 2 VDD
port 41 nsew
rlabel metal1 s -17094 -56199 -17048 -55999 2 VDD
port 41 nsew
rlabel metal1 s -17290 -56199 -17244 -55999 2 VDD
port 41 nsew
rlabel metal1 s -17486 -56199 -17440 -55999 2 VDD
port 41 nsew
rlabel metal1 s -17682 -56199 -17636 -55999 2 VDD
port 41 nsew
rlabel metal1 s -18187 -56022 -18141 -55822 2 VDD
port 41 nsew
rlabel metal1 s -18383 -56022 -18337 -55822 2 VDD
port 41 nsew
rlabel metal1 s -18925 -56022 -18879 -55822 2 VDD
port 41 nsew
rlabel metal1 s -19121 -56022 -19075 -55822 2 VDD
port 41 nsew
rlabel metal1 s -19317 -56022 -19271 -55822 2 VDD
port 41 nsew
rlabel metal1 s -19513 -56022 -19467 -55822 2 VDD
port 41 nsew
rlabel metal1 s -20089 -56016 -20043 -55916 2 VDD
port 41 nsew
rlabel metal1 s -20285 -56016 -20239 -55916 2 VDD
port 41 nsew
rlabel metal1 s -20481 -56016 -20435 -55916 2 VDD
port 41 nsew
rlabel metal1 s -20677 -56016 -20631 -55916 2 VDD
port 41 nsew
rlabel metal1 s -20894 -56217 -20848 -55917 2 VDD
port 41 nsew
rlabel metal1 s -21090 -56217 -21044 -55917 2 VDD
port 41 nsew
rlabel metal1 s -21286 -56217 -21240 -55917 2 VDD
port 41 nsew
rlabel metal1 s -27832 -56110 -27432 -56064 2 VDD
port 41 nsew
rlabel metal1 s -27832 -55862 -27432 -55816 2 VDD
port 41 nsew
rlabel metal1 s -27832 -55626 -27432 -55580 2 VDD
port 41 nsew
rlabel metal1 s 3540 -55507 3663 -55494 8 VDD
port 41 nsew
rlabel metal1 s 3151 -55508 3274 -55494 8 VDD
port 41 nsew
rlabel metal1 s 7741 -55488 7864 -55469 8 VDD
port 41 nsew
rlabel metal1 s 6525 -55487 6648 -55469 8 VDD
port 41 nsew
rlabel metal1 s 6525 -55469 7864 -55364 8 VDD
port 41 nsew
rlabel metal1 s 7741 -55364 7864 -55352 8 VDD
port 41 nsew
rlabel metal1 s 6525 -55364 6648 -55351 8 VDD
port 41 nsew
rlabel metal1 s 5169 -55482 5292 -55464 8 VDD
port 41 nsew
rlabel metal1 s 4768 -55484 4891 -55464 8 VDD
port 41 nsew
rlabel metal1 s 4768 -55464 5292 -55357 8 VDD
port 41 nsew
rlabel metal1 s 3151 -55494 3663 -55387 8 VDD
port 41 nsew
rlabel metal1 s 3540 -55387 3663 -55371 8 VDD
port 41 nsew
rlabel metal1 s 3151 -55387 3274 -55372 8 VDD
port 41 nsew
rlabel metal1 s 173 -55495 296 -55487 8 VDD
port 41 nsew
rlabel metal1 s -121 -55496 2 -55487 2 VDD
port 41 nsew
rlabel metal1 s -121 -55487 296 -55372 8 VDD
port 41 nsew
rlabel metal1 s 173 -55372 296 -55359 8 VDD
port 41 nsew
rlabel metal1 s -121 -55372 2 -55360 2 VDD
port 41 nsew
rlabel metal1 s 5169 -55357 5292 -55346 8 VDD
port 41 nsew
rlabel metal1 s 4768 -55357 4891 -55348 8 VDD
port 41 nsew
rlabel metal1 s -3947 -54830 -3824 -54694 2 VDD
port 41 nsew
rlabel metal1 s 1103 -54578 1409 -54516 8 VDD
port 41 nsew
rlabel metal1 s -1380 -54686 -1257 -54550 2 VDD
port 41 nsew
rlabel metal1 s 1103 -54516 1226 -54515 8 VDD
port 41 nsew
rlabel metal1 s 1108 -54515 1222 -54098 8 VDD
port 41 nsew
rlabel metal1 s -1375 -54550 -1261 -54098 2 VDD
port 41 nsew
rlabel metal1 s 1104 -54098 1227 -53962 8 VDD
port 41 nsew
rlabel metal1 s -1379 -54098 -1256 -53962 2 VDD
port 41 nsew
rlabel metal1 s -3942 -54694 -3828 -54063 2 VDD
port 41 nsew
rlabel metal1 s -5221 -54834 -5175 -54634 2 VDD
port 41 nsew
rlabel metal1 s -5417 -54834 -5371 -54634 2 VDD
port 41 nsew
rlabel metal1 s -5613 -54834 -5567 -54634 2 VDD
port 41 nsew
rlabel metal1 s -15642 -55359 -15596 -54759 2 VDD
port 41 nsew
rlabel metal1 s -16065 -55359 -16019 -54759 2 VDD
port 41 nsew
rlabel metal1 s -16261 -55359 -16215 -54759 2 VDD
port 41 nsew
rlabel metal1 s -27832 -55390 -27432 -55344 2 VDD
port 41 nsew
rlabel metal1 s -16511 -55271 -16465 -55171 2 VDD
port 41 nsew
rlabel metal1 s -16707 -55271 -16661 -55171 2 VDD
port 41 nsew
rlabel metal1 s -16903 -55271 -16857 -55171 2 VDD
port 41 nsew
rlabel metal1 s -17099 -55271 -17053 -55171 2 VDD
port 41 nsew
rlabel metal1 s -17316 -55270 -17270 -54970 2 VDD
port 41 nsew
rlabel metal1 s -17512 -55270 -17466 -54970 2 VDD
port 41 nsew
rlabel metal1 s -17708 -55270 -17662 -54970 2 VDD
port 41 nsew
rlabel metal1 s -27832 -55154 -27432 -55108 2 VDD
port 41 nsew
rlabel metal1 s -27832 -54918 -27432 -54872 2 VDD
port 41 nsew
rlabel metal1 s -27832 -54682 -27432 -54636 2 VDD
port 41 nsew
rlabel metal1 s -7929 -54617 -7883 -54417 2 VDD
port 41 nsew
rlabel metal1 s -8125 -54617 -8079 -54417 2 VDD
port 41 nsew
rlabel metal1 s -8321 -54617 -8275 -54417 2 VDD
port 41 nsew
rlabel metal1 s -8811 -54617 -8765 -54417 2 VDD
port 41 nsew
rlabel metal1 s -9007 -54617 -8961 -54417 2 VDD
port 41 nsew
rlabel metal1 s -9203 -54617 -9157 -54417 2 VDD
port 41 nsew
rlabel metal1 s -10554 -54617 -10508 -54417 2 VDD
port 41 nsew
rlabel metal1 s -10750 -54617 -10704 -54417 2 VDD
port 41 nsew
rlabel metal1 s -10946 -54617 -10900 -54417 2 VDD
port 41 nsew
rlabel metal1 s -11511 -54617 -11465 -54417 2 VDD
port 41 nsew
rlabel metal1 s -11707 -54617 -11661 -54417 2 VDD
port 41 nsew
rlabel metal1 s -11903 -54617 -11857 -54417 2 VDD
port 41 nsew
rlabel metal1 s -13254 -54617 -13208 -54417 2 VDD
port 41 nsew
rlabel metal1 s -13450 -54617 -13404 -54417 2 VDD
port 41 nsew
rlabel metal1 s -13646 -54617 -13600 -54417 2 VDD
port 41 nsew
rlabel metal1 s -27832 -54446 -27432 -54400 2 VDD
port 41 nsew
rlabel metal1 s -3946 -54063 -3823 -53927 2 VDD
port 41 nsew
rlabel metal1 s -18147 -54107 -18101 -54007 2 VDD
port 41 nsew
rlabel metal1 s -18343 -54107 -18297 -54007 2 VDD
port 41 nsew
rlabel metal1 s -18539 -54107 -18493 -54007 2 VDD
port 41 nsew
rlabel metal1 s -18735 -54107 -18689 -54007 2 VDD
port 41 nsew
rlabel metal1 s -18952 -54308 -18906 -54008 2 VDD
port 41 nsew
rlabel metal1 s -19148 -54308 -19102 -54008 2 VDD
port 41 nsew
rlabel metal1 s -19344 -54308 -19298 -54008 2 VDD
port 41 nsew
rlabel metal1 s -27832 -54210 -27432 -54164 2 VDD
port 41 nsew
rlabel metal1 s -20017 -54086 -19971 -53886 2 VDD
port 41 nsew
rlabel metal1 s -20213 -54086 -20167 -53886 2 VDD
port 41 nsew
rlabel metal1 s -20755 -54086 -20709 -53886 2 VDD
port 41 nsew
rlabel metal1 s -20951 -54086 -20905 -53886 2 VDD
port 41 nsew
rlabel metal1 s -21147 -54086 -21101 -53886 2 VDD
port 41 nsew
rlabel metal1 s -21343 -54086 -21297 -53886 2 VDD
port 41 nsew
rlabel metal1 s -27832 -53974 -27432 -53928 2 VDD
port 41 nsew
rlabel metal1 s 8737 -53505 8783 -53305 8 VDD
port 41 nsew
rlabel metal1 s 8541 -53505 8587 -53305 8 VDD
port 41 nsew
rlabel metal1 s 8428 -53505 8474 -53305 8 VDD
port 41 nsew
rlabel metal1 s 8232 -53505 8278 -53305 8 VDD
port 41 nsew
rlabel metal1 s 8118 -53505 8164 -53305 8 VDD
port 41 nsew
rlabel metal1 s 7922 -53505 7968 -53305 8 VDD
port 41 nsew
rlabel metal1 s 7726 -53505 7772 -53305 8 VDD
port 41 nsew
rlabel metal1 s 5737 -53505 5783 -53305 8 VDD
port 41 nsew
rlabel metal1 s 5541 -53505 5587 -53305 8 VDD
port 41 nsew
rlabel metal1 s 5428 -53505 5474 -53305 8 VDD
port 41 nsew
rlabel metal1 s 5232 -53505 5278 -53305 8 VDD
port 41 nsew
rlabel metal1 s 5118 -53505 5164 -53305 8 VDD
port 41 nsew
rlabel metal1 s 4922 -53505 4968 -53305 8 VDD
port 41 nsew
rlabel metal1 s 4726 -53505 4772 -53305 8 VDD
port 41 nsew
rlabel metal1 s 3237 -53505 3283 -53305 8 VDD
port 41 nsew
rlabel metal1 s 3041 -53505 3087 -53305 8 VDD
port 41 nsew
rlabel metal1 s 2928 -53505 2974 -53305 8 VDD
port 41 nsew
rlabel metal1 s 2732 -53505 2778 -53305 8 VDD
port 41 nsew
rlabel metal1 s 2618 -53505 2664 -53305 8 VDD
port 41 nsew
rlabel metal1 s 2422 -53505 2468 -53305 8 VDD
port 41 nsew
rlabel metal1 s 2226 -53505 2272 -53305 8 VDD
port 41 nsew
rlabel metal1 s 737 -53505 783 -53305 8 VDD
port 41 nsew
rlabel metal1 s 541 -53505 587 -53305 8 VDD
port 41 nsew
rlabel metal1 s 428 -53505 474 -53305 8 VDD
port 41 nsew
rlabel metal1 s 232 -53505 278 -53305 8 VDD
port 41 nsew
rlabel metal1 s 118 -53505 164 -53305 8 VDD
port 41 nsew
rlabel metal1 s -78 -53505 -32 -53305 2 VDD
port 41 nsew
rlabel metal1 s -274 -53505 -228 -53305 2 VDD
port 41 nsew
rlabel metal1 s -1763 -53505 -1717 -53305 2 VDD
port 41 nsew
rlabel metal1 s -1959 -53505 -1913 -53305 2 VDD
port 41 nsew
rlabel metal1 s -2072 -53505 -2026 -53305 2 VDD
port 41 nsew
rlabel metal1 s -2268 -53505 -2222 -53305 2 VDD
port 41 nsew
rlabel metal1 s -2382 -53505 -2336 -53305 2 VDD
port 41 nsew
rlabel metal1 s -2578 -53505 -2532 -53305 2 VDD
port 41 nsew
rlabel metal1 s -2774 -53505 -2728 -53305 2 VDD
port 41 nsew
rlabel metal1 s -4263 -53505 -4217 -53305 2 VDD
port 41 nsew
rlabel metal1 s -4459 -53505 -4413 -53305 2 VDD
port 41 nsew
rlabel metal1 s -4572 -53505 -4526 -53305 2 VDD
port 41 nsew
rlabel metal1 s -4768 -53505 -4722 -53305 2 VDD
port 41 nsew
rlabel metal1 s -4882 -53505 -4836 -53305 2 VDD
port 41 nsew
rlabel metal1 s -5078 -53505 -5032 -53305 2 VDD
port 41 nsew
rlabel metal1 s -5274 -53505 -5228 -53305 2 VDD
port 41 nsew
rlabel metal1 s -6763 -53709 -6717 -53109 2 VDD
port 41 nsew
rlabel metal1 s -6959 -53709 -6913 -53109 2 VDD
port 41 nsew
rlabel metal1 s -7382 -53709 -7336 -53109 2 VDD
port 41 nsew
rlabel metal1 s -27832 -53738 -27432 -53692 2 VDD
port 41 nsew
rlabel metal1 s -27832 -53502 -27432 -53456 2 VDD
port 41 nsew
rlabel metal1 s -9815 -53299 -9769 -53099 2 VDD
port 41 nsew
rlabel metal1 s -10011 -53299 -9965 -53099 2 VDD
port 41 nsew
rlabel metal1 s -10207 -53299 -10161 -53099 2 VDD
port 41 nsew
rlabel metal1 s -10652 -53299 -10606 -53099 2 VDD
port 41 nsew
rlabel metal1 s -10848 -53299 -10802 -53099 2 VDD
port 41 nsew
rlabel metal1 s -11044 -53299 -10998 -53099 2 VDD
port 41 nsew
rlabel metal1 s -12515 -53299 -12469 -53099 2 VDD
port 41 nsew
rlabel metal1 s -12711 -53299 -12665 -53099 2 VDD
port 41 nsew
rlabel metal1 s -12907 -53299 -12861 -53099 2 VDD
port 41 nsew
rlabel metal1 s -13352 -53299 -13306 -53099 2 VDD
port 41 nsew
rlabel metal1 s -13548 -53299 -13502 -53099 2 VDD
port 41 nsew
rlabel metal1 s -13744 -53299 -13698 -53099 2 VDD
port 41 nsew
rlabel metal1 s -27832 -53266 -27432 -53220 2 VDD
port 41 nsew
rlabel metal1 s -27832 -53030 -27432 -52984 2 VDD
port 41 nsew
rlabel metal1 s -27832 -52794 -27432 -52748 2 VDD
port 41 nsew
rlabel metal1 s -27832 -52558 -27432 -52512 2 VDD
port 41 nsew
rlabel metal1 s -27832 -52322 -27432 -52276 2 VDD
port 41 nsew
rlabel metal1 s 17079 -43769 17125 -43569 8 VDD
port 41 nsew
rlabel metal1 s 16883 -43769 16929 -43569 8 VDD
port 41 nsew
rlabel metal1 s 16687 -43769 16733 -43569 8 VDD
port 41 nsew
rlabel metal1 s 16242 -43769 16288 -43569 8 VDD
port 41 nsew
rlabel metal1 s 16046 -43769 16092 -43569 8 VDD
port 41 nsew
rlabel metal1 s 15850 -43769 15896 -43569 8 VDD
port 41 nsew
rlabel metal1 s 14379 -43769 14425 -43569 8 VDD
port 41 nsew
rlabel metal1 s 14183 -43769 14229 -43569 8 VDD
port 41 nsew
rlabel metal1 s 13987 -43769 14033 -43569 8 VDD
port 41 nsew
rlabel metal1 s 13542 -43769 13588 -43569 8 VDD
port 41 nsew
rlabel metal1 s 13346 -43769 13392 -43569 8 VDD
port 41 nsew
rlabel metal1 s 13150 -43769 13196 -43569 8 VDD
port 41 nsew
rlabel metal1 s 8034 -43932 8080 -43732 8 VDD
port 41 nsew
rlabel metal1 s 7838 -43932 7884 -43732 8 VDD
port 41 nsew
rlabel metal1 s 7725 -43932 7771 -43732 8 VDD
port 41 nsew
rlabel metal1 s 7529 -43932 7575 -43732 8 VDD
port 41 nsew
rlabel metal1 s 7415 -43932 7461 -43732 8 VDD
port 41 nsew
rlabel metal1 s 7219 -43932 7265 -43732 8 VDD
port 41 nsew
rlabel metal1 s 7023 -43932 7069 -43732 8 VDD
port 41 nsew
rlabel metal1 s 5034 -43932 5080 -43732 8 VDD
port 41 nsew
rlabel metal1 s 4838 -43932 4884 -43732 8 VDD
port 41 nsew
rlabel metal1 s 4725 -43932 4771 -43732 8 VDD
port 41 nsew
rlabel metal1 s 4529 -43932 4575 -43732 8 VDD
port 41 nsew
rlabel metal1 s 4415 -43932 4461 -43732 8 VDD
port 41 nsew
rlabel metal1 s 4219 -43932 4265 -43732 8 VDD
port 41 nsew
rlabel metal1 s 4023 -43932 4069 -43732 8 VDD
port 41 nsew
rlabel metal1 s 2534 -43932 2580 -43732 8 VDD
port 41 nsew
rlabel metal1 s 2338 -43932 2384 -43732 8 VDD
port 41 nsew
rlabel metal1 s 2225 -43932 2271 -43732 8 VDD
port 41 nsew
rlabel metal1 s 2029 -43932 2075 -43732 8 VDD
port 41 nsew
rlabel metal1 s 1915 -43932 1961 -43732 8 VDD
port 41 nsew
rlabel metal1 s 1719 -43932 1765 -43732 8 VDD
port 41 nsew
rlabel metal1 s 1523 -43932 1569 -43732 8 VDD
port 41 nsew
rlabel metal1 s 34 -43932 80 -43732 8 VDD
port 41 nsew
rlabel metal1 s -162 -43932 -116 -43732 2 VDD
port 41 nsew
rlabel metal1 s -275 -43932 -229 -43732 2 VDD
port 41 nsew
rlabel metal1 s -471 -43932 -425 -43732 2 VDD
port 41 nsew
rlabel metal1 s -585 -43932 -539 -43732 2 VDD
port 41 nsew
rlabel metal1 s -781 -43932 -735 -43732 2 VDD
port 41 nsew
rlabel metal1 s -977 -43932 -931 -43732 2 VDD
port 41 nsew
rlabel metal1 s -2466 -43932 -2420 -43732 2 VDD
port 41 nsew
rlabel metal1 s -2662 -43932 -2616 -43732 2 VDD
port 41 nsew
rlabel metal1 s -2775 -43932 -2729 -43732 2 VDD
port 41 nsew
rlabel metal1 s -2971 -43932 -2925 -43732 2 VDD
port 41 nsew
rlabel metal1 s -3085 -43932 -3039 -43732 2 VDD
port 41 nsew
rlabel metal1 s -3281 -43932 -3235 -43732 2 VDD
port 41 nsew
rlabel metal1 s -3477 -43932 -3431 -43732 2 VDD
port 41 nsew
rlabel metal1 s -4966 -43932 -4920 -43732 2 VDD
port 41 nsew
rlabel metal1 s -5162 -43932 -5116 -43732 2 VDD
port 41 nsew
rlabel metal1 s -5275 -43932 -5229 -43732 2 VDD
port 41 nsew
rlabel metal1 s -5471 -43932 -5425 -43732 2 VDD
port 41 nsew
rlabel metal1 s -5585 -43932 -5539 -43732 2 VDD
port 41 nsew
rlabel metal1 s -5781 -43932 -5735 -43732 2 VDD
port 41 nsew
rlabel metal1 s -5977 -43932 -5931 -43732 2 VDD
port 41 nsew
rlabel metal1 s -19651 -44182 -19475 -43551 2 VDD
port 41 nsew
rlabel metal1 s -20935 -44018 -20889 -43818 2 VDD
port 41 nsew
rlabel metal1 s -21131 -44018 -21085 -43818 2 VDD
port 41 nsew
rlabel metal1 s -21327 -44018 -21281 -43818 2 VDD
port 41 nsew
rlabel metal1 s -21523 -44018 -21477 -43818 2 VDD
port 41 nsew
rlabel metal1 s -22065 -44018 -22019 -43818 2 VDD
port 41 nsew
rlabel metal1 s -22261 -44018 -22215 -43818 2 VDD
port 41 nsew
rlabel metal1 s 401 -43275 524 -43139 8 VDD
port 41 nsew
rlabel metal1 s -2082 -43275 -1959 -43139 2 VDD
port 41 nsew
rlabel metal1 s -4649 -43310 -4526 -43174 2 VDD
port 41 nsew
rlabel metal1 s 405 -43139 519 -42722 8 VDD
port 41 nsew
rlabel metal1 s 400 -42722 523 -42721 8 VDD
port 41 nsew
rlabel metal1 s 400 -42721 706 -42659 8 VDD
port 41 nsew
rlabel metal1 s -2078 -43139 -1964 -42687 2 VDD
port 41 nsew
rlabel metal1 s -2083 -42687 -1960 -42551 2 VDD
port 41 nsew
rlabel metal1 s -4645 -43174 -4531 -42543 2 VDD
port 41 nsew
rlabel metal1 s -16215 -42858 -16169 -42758 2 VDD
port 41 nsew
rlabel metal1 s -16411 -42858 -16365 -42758 2 VDD
port 41 nsew
rlabel metal1 s -16607 -42858 -16561 -42758 2 VDD
port 41 nsew
rlabel metal1 s -16803 -42858 -16757 -42758 2 VDD
port 41 nsew
rlabel metal1 s -17020 -43059 -16974 -42759 2 VDD
port 41 nsew
rlabel metal1 s -17216 -43059 -17170 -42759 2 VDD
port 41 nsew
rlabel metal1 s -17412 -43059 -17366 -42759 2 VDD
port 41 nsew
rlabel metal1 s -17797 -43088 -17751 -42888 2 VDD
port 41 nsew
rlabel metal1 s -17993 -43088 -17947 -42888 2 VDD
port 41 nsew
rlabel metal1 s -18189 -43088 -18143 -42888 2 VDD
port 41 nsew
rlabel metal1 s -18385 -43088 -18339 -42888 2 VDD
port 41 nsew
rlabel metal1 s 87122 -42161 87168 -41561 8 VDD
port 41 nsew
rlabel metal1 s 86699 -42161 86745 -41561 8 VDD
port 41 nsew
rlabel metal1 s 86503 -42161 86549 -41561 8 VDD
port 41 nsew
rlabel metal1 s 86253 -41749 86299 -41649 8 VDD
port 41 nsew
rlabel metal1 s 86057 -41749 86103 -41649 8 VDD
port 41 nsew
rlabel metal1 s 85861 -41749 85907 -41649 8 VDD
port 41 nsew
rlabel metal1 s 85665 -41749 85711 -41649 8 VDD
port 41 nsew
rlabel metal1 s 85448 -41950 85494 -41650 8 VDD
port 41 nsew
rlabel metal1 s 85252 -41950 85298 -41650 8 VDD
port 41 nsew
rlabel metal1 s 85056 -41950 85102 -41650 8 VDD
port 41 nsew
rlabel metal1 s 83454 -42130 83500 -41530 8 VDD
port 41 nsew
rlabel metal1 s 83031 -42130 83077 -41530 8 VDD
port 41 nsew
rlabel metal1 s 82835 -42130 82881 -41530 8 VDD
port 41 nsew
rlabel metal1 s 82585 -41718 82631 -41618 8 VDD
port 41 nsew
rlabel metal1 s 82389 -41718 82435 -41618 8 VDD
port 41 nsew
rlabel metal1 s 82193 -41718 82239 -41618 8 VDD
port 41 nsew
rlabel metal1 s 81997 -41718 82043 -41618 8 VDD
port 41 nsew
rlabel metal1 s 81780 -41919 81826 -41619 8 VDD
port 41 nsew
rlabel metal1 s 81584 -41919 81630 -41619 8 VDD
port 41 nsew
rlabel metal1 s 81388 -41919 81434 -41619 8 VDD
port 41 nsew
rlabel metal1 s 77758 -42199 77804 -41599 8 VDD
port 41 nsew
rlabel metal1 s 77335 -42199 77381 -41599 8 VDD
port 41 nsew
rlabel metal1 s 77139 -42199 77185 -41599 8 VDD
port 41 nsew
rlabel metal1 s 76889 -41787 76935 -41687 8 VDD
port 41 nsew
rlabel metal1 s 76693 -41787 76739 -41687 8 VDD
port 41 nsew
rlabel metal1 s 76497 -41787 76543 -41687 8 VDD
port 41 nsew
rlabel metal1 s 76301 -41787 76347 -41687 8 VDD
port 41 nsew
rlabel metal1 s 76084 -41988 76130 -41688 8 VDD
port 41 nsew
rlabel metal1 s 75888 -41988 75934 -41688 8 VDD
port 41 nsew
rlabel metal1 s 75692 -41988 75738 -41688 8 VDD
port 41 nsew
rlabel metal1 s 74090 -42168 74136 -41568 8 VDD
port 41 nsew
rlabel metal1 s 73667 -42168 73713 -41568 8 VDD
port 41 nsew
rlabel metal1 s 73471 -42168 73517 -41568 8 VDD
port 41 nsew
rlabel metal1 s 73221 -41756 73267 -41656 8 VDD
port 41 nsew
rlabel metal1 s 73025 -41756 73071 -41656 8 VDD
port 41 nsew
rlabel metal1 s 72829 -41756 72875 -41656 8 VDD
port 41 nsew
rlabel metal1 s 72633 -41756 72679 -41656 8 VDD
port 41 nsew
rlabel metal1 s 72416 -41957 72462 -41657 8 VDD
port 41 nsew
rlabel metal1 s 72220 -41957 72266 -41657 8 VDD
port 41 nsew
rlabel metal1 s 72024 -41957 72070 -41657 8 VDD
port 41 nsew
rlabel metal1 s 68605 -42216 68651 -41616 8 VDD
port 41 nsew
rlabel metal1 s 68182 -42216 68228 -41616 8 VDD
port 41 nsew
rlabel metal1 s 67986 -42216 68032 -41616 8 VDD
port 41 nsew
rlabel metal1 s 67736 -41804 67782 -41704 8 VDD
port 41 nsew
rlabel metal1 s 67540 -41804 67586 -41704 8 VDD
port 41 nsew
rlabel metal1 s 67344 -41804 67390 -41704 8 VDD
port 41 nsew
rlabel metal1 s 67148 -41804 67194 -41704 8 VDD
port 41 nsew
rlabel metal1 s 66931 -42005 66977 -41705 8 VDD
port 41 nsew
rlabel metal1 s 66735 -42005 66781 -41705 8 VDD
port 41 nsew
rlabel metal1 s 66539 -42005 66585 -41705 8 VDD
port 41 nsew
rlabel metal1 s 64937 -42185 64983 -41585 8 VDD
port 41 nsew
rlabel metal1 s 64514 -42185 64560 -41585 8 VDD
port 41 nsew
rlabel metal1 s 64318 -42185 64364 -41585 8 VDD
port 41 nsew
rlabel metal1 s 64068 -41773 64114 -41673 8 VDD
port 41 nsew
rlabel metal1 s 63872 -41773 63918 -41673 8 VDD
port 41 nsew
rlabel metal1 s 63676 -41773 63722 -41673 8 VDD
port 41 nsew
rlabel metal1 s 63480 -41773 63526 -41673 8 VDD
port 41 nsew
rlabel metal1 s 63263 -41974 63309 -41674 8 VDD
port 41 nsew
rlabel metal1 s 63067 -41974 63113 -41674 8 VDD
port 41 nsew
rlabel metal1 s 62871 -41974 62917 -41674 8 VDD
port 41 nsew
rlabel metal1 s 59851 -42282 59897 -41682 8 VDD
port 41 nsew
rlabel metal1 s 59428 -42282 59474 -41682 8 VDD
port 41 nsew
rlabel metal1 s 59232 -42282 59278 -41682 8 VDD
port 41 nsew
rlabel metal1 s 58982 -41870 59028 -41770 8 VDD
port 41 nsew
rlabel metal1 s 58786 -41870 58832 -41770 8 VDD
port 41 nsew
rlabel metal1 s 58590 -41870 58636 -41770 8 VDD
port 41 nsew
rlabel metal1 s 58394 -41870 58440 -41770 8 VDD
port 41 nsew
rlabel metal1 s 58177 -42071 58223 -41771 8 VDD
port 41 nsew
rlabel metal1 s 57981 -42071 58027 -41771 8 VDD
port 41 nsew
rlabel metal1 s 57785 -42071 57831 -41771 8 VDD
port 41 nsew
rlabel metal1 s 56183 -42251 56229 -41651 8 VDD
port 41 nsew
rlabel metal1 s 55760 -42251 55806 -41651 8 VDD
port 41 nsew
rlabel metal1 s 55564 -42251 55610 -41651 8 VDD
port 41 nsew
rlabel metal1 s 55314 -41839 55360 -41739 8 VDD
port 41 nsew
rlabel metal1 s 55118 -41839 55164 -41739 8 VDD
port 41 nsew
rlabel metal1 s 54922 -41839 54968 -41739 8 VDD
port 41 nsew
rlabel metal1 s 54726 -41839 54772 -41739 8 VDD
port 41 nsew
rlabel metal1 s 54509 -42040 54555 -41740 8 VDD
port 41 nsew
rlabel metal1 s 54313 -42040 54359 -41740 8 VDD
port 41 nsew
rlabel metal1 s 54117 -42040 54163 -41740 8 VDD
port 41 nsew
rlabel metal1 s 50653 -42316 50699 -41716 8 VDD
port 41 nsew
rlabel metal1 s 50230 -42316 50276 -41716 8 VDD
port 41 nsew
rlabel metal1 s 50034 -42316 50080 -41716 8 VDD
port 41 nsew
rlabel metal1 s 49784 -41904 49830 -41804 8 VDD
port 41 nsew
rlabel metal1 s 49588 -41904 49634 -41804 8 VDD
port 41 nsew
rlabel metal1 s 49392 -41904 49438 -41804 8 VDD
port 41 nsew
rlabel metal1 s 49196 -41904 49242 -41804 8 VDD
port 41 nsew
rlabel metal1 s 48979 -42105 49025 -41805 8 VDD
port 41 nsew
rlabel metal1 s 48783 -42105 48829 -41805 8 VDD
port 41 nsew
rlabel metal1 s 48587 -42105 48633 -41805 8 VDD
port 41 nsew
rlabel metal1 s 46985 -42285 47031 -41685 8 VDD
port 41 nsew
rlabel metal1 s 46562 -42285 46608 -41685 8 VDD
port 41 nsew
rlabel metal1 s 46366 -42285 46412 -41685 8 VDD
port 41 nsew
rlabel metal1 s 46116 -41873 46162 -41773 8 VDD
port 41 nsew
rlabel metal1 s 45920 -41873 45966 -41773 8 VDD
port 41 nsew
rlabel metal1 s 45724 -41873 45770 -41773 8 VDD
port 41 nsew
rlabel metal1 s 45528 -41873 45574 -41773 8 VDD
port 41 nsew
rlabel metal1 s 45311 -42074 45357 -41774 8 VDD
port 41 nsew
rlabel metal1 s 45115 -42074 45161 -41774 8 VDD
port 41 nsew
rlabel metal1 s 44919 -42074 44965 -41774 8 VDD
port 41 nsew
rlabel metal1 s 41790 -42277 41836 -41677 8 VDD
port 41 nsew
rlabel metal1 s 41367 -42277 41413 -41677 8 VDD
port 41 nsew
rlabel metal1 s 41171 -42277 41217 -41677 8 VDD
port 41 nsew
rlabel metal1 s 40921 -41865 40967 -41765 8 VDD
port 41 nsew
rlabel metal1 s 40725 -41865 40771 -41765 8 VDD
port 41 nsew
rlabel metal1 s 40529 -41865 40575 -41765 8 VDD
port 41 nsew
rlabel metal1 s 40333 -41865 40379 -41765 8 VDD
port 41 nsew
rlabel metal1 s 40116 -42066 40162 -41766 8 VDD
port 41 nsew
rlabel metal1 s 39920 -42066 39966 -41766 8 VDD
port 41 nsew
rlabel metal1 s 39724 -42066 39770 -41766 8 VDD
port 41 nsew
rlabel metal1 s 38122 -42246 38168 -41646 8 VDD
port 41 nsew
rlabel metal1 s 37699 -42246 37745 -41646 8 VDD
port 41 nsew
rlabel metal1 s 37503 -42246 37549 -41646 8 VDD
port 41 nsew
rlabel metal1 s 37253 -41834 37299 -41734 8 VDD
port 41 nsew
rlabel metal1 s 37057 -41834 37103 -41734 8 VDD
port 41 nsew
rlabel metal1 s 36861 -41834 36907 -41734 8 VDD
port 41 nsew
rlabel metal1 s 36665 -41834 36711 -41734 8 VDD
port 41 nsew
rlabel metal1 s 36448 -42035 36494 -41735 8 VDD
port 41 nsew
rlabel metal1 s 36252 -42035 36298 -41735 8 VDD
port 41 nsew
rlabel metal1 s 36056 -42035 36102 -41735 8 VDD
port 41 nsew
rlabel metal1 s 33350 -42266 33396 -41666 8 VDD
port 41 nsew
rlabel metal1 s 32927 -42266 32973 -41666 8 VDD
port 41 nsew
rlabel metal1 s 32731 -42266 32777 -41666 8 VDD
port 41 nsew
rlabel metal1 s 16981 -42451 17027 -42251 8 VDD
port 41 nsew
rlabel metal1 s 16785 -42451 16831 -42251 8 VDD
port 41 nsew
rlabel metal1 s 16589 -42451 16635 -42251 8 VDD
port 41 nsew
rlabel metal1 s 15238 -42451 15284 -42251 8 VDD
port 41 nsew
rlabel metal1 s 15042 -42451 15088 -42251 8 VDD
port 41 nsew
rlabel metal1 s 14846 -42451 14892 -42251 8 VDD
port 41 nsew
rlabel metal1 s 14281 -42451 14327 -42251 8 VDD
port 41 nsew
rlabel metal1 s 14085 -42451 14131 -42251 8 VDD
port 41 nsew
rlabel metal1 s 13889 -42451 13935 -42251 8 VDD
port 41 nsew
rlabel metal1 s 12538 -42451 12584 -42251 8 VDD
port 41 nsew
rlabel metal1 s 12342 -42451 12388 -42251 8 VDD
port 41 nsew
rlabel metal1 s 12146 -42451 12192 -42251 8 VDD
port 41 nsew
rlabel metal1 s 11656 -42451 11702 -42251 8 VDD
port 41 nsew
rlabel metal1 s 11460 -42451 11506 -42251 8 VDD
port 41 nsew
rlabel metal1 s 11264 -42451 11310 -42251 8 VDD
port 41 nsew
rlabel metal1 s -4650 -42543 -4527 -42407 2 VDD
port 41 nsew
rlabel metal1 s -18846 -42556 -18654 -42384 2 VDD
port 41 nsew
rlabel metal1 s 32481 -41854 32527 -41754 8 VDD
port 41 nsew
rlabel metal1 s 32285 -41854 32331 -41754 8 VDD
port 41 nsew
rlabel metal1 s 32089 -41854 32135 -41754 8 VDD
port 41 nsew
rlabel metal1 s 31893 -41854 31939 -41754 8 VDD
port 41 nsew
rlabel metal1 s 31676 -42055 31722 -41755 8 VDD
port 41 nsew
rlabel metal1 s 31480 -42055 31526 -41755 8 VDD
port 41 nsew
rlabel metal1 s 31284 -42055 31330 -41755 8 VDD
port 41 nsew
rlabel metal1 s 29682 -42235 29728 -41635 8 VDD
port 41 nsew
rlabel metal1 s 29259 -42235 29305 -41635 8 VDD
port 41 nsew
rlabel metal1 s 29063 -42235 29109 -41635 8 VDD
port 41 nsew
rlabel metal1 s 28813 -41823 28859 -41723 8 VDD
port 41 nsew
rlabel metal1 s 28617 -41823 28663 -41723 8 VDD
port 41 nsew
rlabel metal1 s 28421 -41823 28467 -41723 8 VDD
port 41 nsew
rlabel metal1 s 28225 -41823 28271 -41723 8 VDD
port 41 nsew
rlabel metal1 s 28008 -42024 28054 -41724 8 VDD
port 41 nsew
rlabel metal1 s 27812 -42024 27858 -41724 8 VDD
port 41 nsew
rlabel metal1 s 27616 -42024 27662 -41724 8 VDD
port 41 nsew
rlabel metal1 s 7038 -41885 7161 -41873 8 VDD
port 41 nsew
rlabel metal1 s 5822 -41886 5945 -41873 8 VDD
port 41 nsew
rlabel metal1 s 5822 -41873 7161 -41768 8 VDD
port 41 nsew
rlabel metal1 s 7038 -41768 7161 -41749 8 VDD
port 41 nsew
rlabel metal1 s 5822 -41768 5945 -41750 8 VDD
port 41 nsew
rlabel metal1 s 4466 -41891 4589 -41880 8 VDD
port 41 nsew
rlabel metal1 s 4065 -41889 4188 -41880 8 VDD
port 41 nsew
rlabel metal1 s 4065 -41880 4589 -41773 8 VDD
port 41 nsew
rlabel metal1 s 4466 -41773 4589 -41755 8 VDD
port 41 nsew
rlabel metal1 s 4065 -41773 4188 -41753 8 VDD
port 41 nsew
rlabel metal1 s 2837 -41866 2960 -41850 8 VDD
port 41 nsew
rlabel metal1 s -530 -41878 -407 -41865 2 VDD
port 41 nsew
rlabel metal1 s -824 -41877 -701 -41865 2 VDD
port 41 nsew
rlabel metal1 s 2448 -41865 2571 -41850 8 VDD
port 41 nsew
rlabel metal1 s 2448 -41850 2960 -41743 8 VDD
port 41 nsew
rlabel metal1 s 2837 -41743 2960 -41730 8 VDD
port 41 nsew
rlabel metal1 s 2448 -41743 2571 -41729 8 VDD
port 41 nsew
rlabel metal1 s -824 -41865 -407 -41750 2 VDD
port 41 nsew
rlabel metal1 s -530 -41750 -407 -41742 2 VDD
port 41 nsew
rlabel metal1 s -824 -41750 -701 -41741 2 VDD
port 41 nsew
rlabel metal1 s 51093 -41635 51244 -41610 8 VDD
port 41 nsew
rlabel metal1 s 50843 -41622 50934 -41610 8 VDD
port 41 nsew
rlabel metal1 s 60291 -41601 60442 -41576 8 VDD
port 41 nsew
rlabel metal1 s 60041 -41588 60132 -41576 8 VDD
port 41 nsew
rlabel metal1 s 78198 -41518 78349 -41493 8 VDD
port 41 nsew
rlabel metal1 s 69045 -41535 69196 -41510 8 VDD
port 41 nsew
rlabel metal1 s 68795 -41522 68886 -41510 8 VDD
port 41 nsew
rlabel metal1 s 77948 -41505 78039 -41493 8 VDD
port 41 nsew
rlabel metal1 s 87562 -41480 87713 -41455 8 VDD
port 41 nsew
rlabel metal1 s 87312 -41467 87403 -41455 8 VDD
port 41 nsew
rlabel metal1 s 87312 -41455 87713 -41316 8 VDD
port 41 nsew
rlabel metal1 s 87562 -41316 87713 -41289 8 VDD
port 41 nsew
rlabel metal1 s 87312 -41316 87403 -41304 8 VDD
port 41 nsew
rlabel metal1 s 83892 -41402 83988 -41376 8 VDD
port 41 nsew
rlabel metal1 s 82589 -41383 82772 -41376 8 VDD
port 41 nsew
rlabel metal1 s 82589 -41376 83988 -41294 8 VDD
port 41 nsew
rlabel metal1 s 77948 -41493 78349 -41354 8 VDD
port 41 nsew
rlabel metal1 s 78198 -41354 78349 -41327 8 VDD
port 41 nsew
rlabel metal1 s 77948 -41354 78039 -41342 8 VDD
port 41 nsew
rlabel metal1 s 74528 -41440 74624 -41414 8 VDD
port 41 nsew
rlabel metal1 s 73225 -41421 73408 -41414 8 VDD
port 41 nsew
rlabel metal1 s 73225 -41414 74624 -41332 8 VDD
port 41 nsew
rlabel metal1 s 68795 -41510 69196 -41371 8 VDD
port 41 nsew
rlabel metal1 s 69045 -41371 69196 -41344 8 VDD
port 41 nsew
rlabel metal1 s 68795 -41371 68886 -41359 8 VDD
port 41 nsew
rlabel metal1 s 65375 -41457 65471 -41431 8 VDD
port 41 nsew
rlabel metal1 s 64072 -41438 64255 -41431 8 VDD
port 41 nsew
rlabel metal1 s 64072 -41431 65471 -41349 8 VDD
port 41 nsew
rlabel metal1 s 60041 -41576 60442 -41437 8 VDD
port 41 nsew
rlabel metal1 s 60291 -41437 60442 -41410 8 VDD
port 41 nsew
rlabel metal1 s 60041 -41437 60132 -41425 8 VDD
port 41 nsew
rlabel metal1 s 56621 -41523 56717 -41497 8 VDD
port 41 nsew
rlabel metal1 s 55318 -41504 55501 -41497 8 VDD
port 41 nsew
rlabel metal1 s 55318 -41497 56717 -41415 8 VDD
port 41 nsew
rlabel metal1 s 50843 -41610 51244 -41471 8 VDD
port 41 nsew
rlabel metal1 s 42230 -41596 42381 -41571 8 VDD
port 41 nsew
rlabel metal1 s 41980 -41583 42071 -41571 8 VDD
port 41 nsew
rlabel metal1 s 51093 -41471 51244 -41444 8 VDD
port 41 nsew
rlabel metal1 s 50843 -41471 50934 -41459 8 VDD
port 41 nsew
rlabel metal1 s 47423 -41557 47519 -41531 8 VDD
port 41 nsew
rlabel metal1 s 46120 -41538 46303 -41531 8 VDD
port 41 nsew
rlabel metal1 s 46120 -41531 47519 -41449 8 VDD
port 41 nsew
rlabel metal1 s 47423 -41449 47519 -41420 8 VDD
port 41 nsew
rlabel metal1 s 56621 -41415 56717 -41386 8 VDD
port 41 nsew
rlabel metal1 s 55318 -41415 55501 -41374 8 VDD
port 41 nsew
rlabel metal1 s 46120 -41449 46303 -41408 8 VDD
port 41 nsew
rlabel metal1 s 41980 -41571 42381 -41432 8 VDD
port 41 nsew
rlabel metal1 s 33790 -41585 33941 -41560 8 VDD
port 41 nsew
rlabel metal1 s 33540 -41572 33631 -41560 8 VDD
port 41 nsew
rlabel metal1 s 42230 -41432 42381 -41405 8 VDD
port 41 nsew
rlabel metal1 s 41980 -41432 42071 -41420 8 VDD
port 41 nsew
rlabel metal1 s 38560 -41518 38656 -41492 8 VDD
port 41 nsew
rlabel metal1 s 37257 -41499 37440 -41492 8 VDD
port 41 nsew
rlabel metal1 s 37257 -41492 38656 -41410 8 VDD
port 41 nsew
rlabel metal1 s 38560 -41410 38656 -41381 8 VDD
port 41 nsew
rlabel metal1 s 37257 -41410 37440 -41369 8 VDD
port 41 nsew
rlabel metal1 s 33540 -41560 33941 -41421 8 VDD
port 41 nsew
rlabel metal1 s 33790 -41421 33941 -41394 8 VDD
port 41 nsew
rlabel metal1 s 33540 -41421 33631 -41409 8 VDD
port 41 nsew
rlabel metal1 s 30120 -41507 30216 -41481 8 VDD
port 41 nsew
rlabel metal1 s 28817 -41488 29000 -41481 8 VDD
port 41 nsew
rlabel metal1 s 8044 -41681 8090 -41481 8 VDD
port 41 nsew
rlabel metal1 s 7848 -41681 7894 -41481 8 VDD
port 41 nsew
rlabel metal1 s 7735 -41681 7781 -41481 8 VDD
port 41 nsew
rlabel metal1 s 7539 -41681 7585 -41481 8 VDD
port 41 nsew
rlabel metal1 s 7425 -41681 7471 -41481 8 VDD
port 41 nsew
rlabel metal1 s 7229 -41681 7275 -41481 8 VDD
port 41 nsew
rlabel metal1 s 7033 -41681 7079 -41481 8 VDD
port 41 nsew
rlabel metal1 s 5872 -41692 5918 -41492 8 VDD
port 41 nsew
rlabel metal1 s 5676 -41692 5722 -41492 8 VDD
port 41 nsew
rlabel metal1 s 5480 -41692 5526 -41492 8 VDD
port 41 nsew
rlabel metal1 s 5284 -41692 5330 -41492 8 VDD
port 41 nsew
rlabel metal1 s 4742 -41692 4788 -41492 8 VDD
port 41 nsew
rlabel metal1 s 4546 -41692 4592 -41492 8 VDD
port 41 nsew
rlabel metal1 s 28817 -41481 30216 -41399 8 VDD
port 41 nsew
rlabel metal1 s 30120 -41399 30216 -41370 8 VDD
port 41 nsew
rlabel metal1 s 28817 -41399 29000 -41358 8 VDD
port 41 nsew
rlabel metal1 s 74528 -41332 74624 -41303 8 VDD
port 41 nsew
rlabel metal1 s 83892 -41294 83988 -41265 8 VDD
port 41 nsew
rlabel metal1 s 82589 -41294 82772 -41253 8 VDD
port 41 nsew
rlabel metal1 s 73225 -41332 73408 -41291 8 VDD
port 41 nsew
rlabel metal1 s 65375 -41349 65471 -41320 8 VDD
port 41 nsew
rlabel metal1 s 64072 -41349 64255 -41308 8 VDD
port 41 nsew
rlabel metal1 s 87252 -41051 87298 -40951 8 VDD
port 41 nsew
rlabel metal1 s 87056 -41051 87102 -40951 8 VDD
port 41 nsew
rlabel metal1 s 86860 -41051 86906 -40951 8 VDD
port 41 nsew
rlabel metal1 s 86664 -41051 86710 -40951 8 VDD
port 41 nsew
rlabel metal1 s 86447 -41050 86493 -40750 8 VDD
port 41 nsew
rlabel metal1 s 86251 -41050 86297 -40750 8 VDD
port 41 nsew
rlabel metal1 s 86055 -41050 86101 -40750 8 VDD
port 41 nsew
rlabel metal1 s 85670 -40921 85716 -40721 8 VDD
port 41 nsew
rlabel metal1 s 85474 -40921 85520 -40721 8 VDD
port 41 nsew
rlabel metal1 s 85278 -40921 85324 -40721 8 VDD
port 41 nsew
rlabel metal1 s 85082 -40921 85128 -40721 8 VDD
port 41 nsew
rlabel metal1 s 83584 -41020 83630 -40920 8 VDD
port 41 nsew
rlabel metal1 s 83388 -41020 83434 -40920 8 VDD
port 41 nsew
rlabel metal1 s 83192 -41020 83238 -40920 8 VDD
port 41 nsew
rlabel metal1 s 82996 -41020 83042 -40920 8 VDD
port 41 nsew
rlabel metal1 s 82779 -41019 82825 -40719 8 VDD
port 41 nsew
rlabel metal1 s 82583 -41019 82629 -40719 8 VDD
port 41 nsew
rlabel metal1 s 82387 -41019 82433 -40719 8 VDD
port 41 nsew
rlabel metal1 s 77888 -41089 77934 -40989 8 VDD
port 41 nsew
rlabel metal1 s 77692 -41089 77738 -40989 8 VDD
port 41 nsew
rlabel metal1 s 77496 -41089 77542 -40989 8 VDD
port 41 nsew
rlabel metal1 s 77300 -41089 77346 -40989 8 VDD
port 41 nsew
rlabel metal1 s 82002 -40890 82048 -40690 8 VDD
port 41 nsew
rlabel metal1 s 81806 -40890 81852 -40690 8 VDD
port 41 nsew
rlabel metal1 s 81610 -40890 81656 -40690 8 VDD
port 41 nsew
rlabel metal1 s 81414 -40890 81460 -40690 8 VDD
port 41 nsew
rlabel metal1 s 77083 -41088 77129 -40788 8 VDD
port 41 nsew
rlabel metal1 s 76887 -41088 76933 -40788 8 VDD
port 41 nsew
rlabel metal1 s 76691 -41088 76737 -40788 8 VDD
port 41 nsew
rlabel metal1 s 76306 -40959 76352 -40759 8 VDD
port 41 nsew
rlabel metal1 s 76110 -40959 76156 -40759 8 VDD
port 41 nsew
rlabel metal1 s 75914 -40959 75960 -40759 8 VDD
port 41 nsew
rlabel metal1 s 75718 -40959 75764 -40759 8 VDD
port 41 nsew
rlabel metal1 s 74220 -41058 74266 -40958 8 VDD
port 41 nsew
rlabel metal1 s 74024 -41058 74070 -40958 8 VDD
port 41 nsew
rlabel metal1 s 73828 -41058 73874 -40958 8 VDD
port 41 nsew
rlabel metal1 s 73632 -41058 73678 -40958 8 VDD
port 41 nsew
rlabel metal1 s 73415 -41057 73461 -40757 8 VDD
port 41 nsew
rlabel metal1 s 73219 -41057 73265 -40757 8 VDD
port 41 nsew
rlabel metal1 s 73023 -41057 73069 -40757 8 VDD
port 41 nsew
rlabel metal1 s 68735 -41106 68781 -41006 8 VDD
port 41 nsew
rlabel metal1 s 68539 -41106 68585 -41006 8 VDD
port 41 nsew
rlabel metal1 s 68343 -41106 68389 -41006 8 VDD
port 41 nsew
rlabel metal1 s 68147 -41106 68193 -41006 8 VDD
port 41 nsew
rlabel metal1 s 72638 -40928 72684 -40728 8 VDD
port 41 nsew
rlabel metal1 s 72442 -40928 72488 -40728 8 VDD
port 41 nsew
rlabel metal1 s 72246 -40928 72292 -40728 8 VDD
port 41 nsew
rlabel metal1 s 72050 -40928 72096 -40728 8 VDD
port 41 nsew
rlabel metal1 s 67930 -41105 67976 -40805 8 VDD
port 41 nsew
rlabel metal1 s 67734 -41105 67780 -40805 8 VDD
port 41 nsew
rlabel metal1 s 67538 -41105 67584 -40805 8 VDD
port 41 nsew
rlabel metal1 s 67153 -40976 67199 -40776 8 VDD
port 41 nsew
rlabel metal1 s 66957 -40976 67003 -40776 8 VDD
port 41 nsew
rlabel metal1 s 66761 -40976 66807 -40776 8 VDD
port 41 nsew
rlabel metal1 s 66565 -40976 66611 -40776 8 VDD
port 41 nsew
rlabel metal1 s 65067 -41075 65113 -40975 8 VDD
port 41 nsew
rlabel metal1 s 64871 -41075 64917 -40975 8 VDD
port 41 nsew
rlabel metal1 s 64675 -41075 64721 -40975 8 VDD
port 41 nsew
rlabel metal1 s 64479 -41075 64525 -40975 8 VDD
port 41 nsew
rlabel metal1 s 64262 -41074 64308 -40774 8 VDD
port 41 nsew
rlabel metal1 s 64066 -41074 64112 -40774 8 VDD
port 41 nsew
rlabel metal1 s 63870 -41074 63916 -40774 8 VDD
port 41 nsew
rlabel metal1 s 59981 -41172 60027 -41072 8 VDD
port 41 nsew
rlabel metal1 s 59785 -41172 59831 -41072 8 VDD
port 41 nsew
rlabel metal1 s 59589 -41172 59635 -41072 8 VDD
port 41 nsew
rlabel metal1 s 59393 -41172 59439 -41072 8 VDD
port 41 nsew
rlabel metal1 s 63485 -40945 63531 -40745 8 VDD
port 41 nsew
rlabel metal1 s 63289 -40945 63335 -40745 8 VDD
port 41 nsew
rlabel metal1 s 63093 -40945 63139 -40745 8 VDD
port 41 nsew
rlabel metal1 s 62897 -40945 62943 -40745 8 VDD
port 41 nsew
rlabel metal1 s 59176 -41171 59222 -40871 8 VDD
port 41 nsew
rlabel metal1 s 58980 -41171 59026 -40871 8 VDD
port 41 nsew
rlabel metal1 s 58784 -41171 58830 -40871 8 VDD
port 41 nsew
rlabel metal1 s 58399 -41042 58445 -40842 8 VDD
port 41 nsew
rlabel metal1 s 58203 -41042 58249 -40842 8 VDD
port 41 nsew
rlabel metal1 s 58007 -41042 58053 -40842 8 VDD
port 41 nsew
rlabel metal1 s 57811 -41042 57857 -40842 8 VDD
port 41 nsew
rlabel metal1 s 56313 -41141 56359 -41041 8 VDD
port 41 nsew
rlabel metal1 s 56117 -41141 56163 -41041 8 VDD
port 41 nsew
rlabel metal1 s 55921 -41141 55967 -41041 8 VDD
port 41 nsew
rlabel metal1 s 55725 -41141 55771 -41041 8 VDD
port 41 nsew
rlabel metal1 s 55508 -41140 55554 -40840 8 VDD
port 41 nsew
rlabel metal1 s 55312 -41140 55358 -40840 8 VDD
port 41 nsew
rlabel metal1 s 55116 -41140 55162 -40840 8 VDD
port 41 nsew
rlabel metal1 s 50783 -41206 50829 -41106 8 VDD
port 41 nsew
rlabel metal1 s 50587 -41206 50633 -41106 8 VDD
port 41 nsew
rlabel metal1 s 50391 -41206 50437 -41106 8 VDD
port 41 nsew
rlabel metal1 s 50195 -41206 50241 -41106 8 VDD
port 41 nsew
rlabel metal1 s 54731 -41011 54777 -40811 8 VDD
port 41 nsew
rlabel metal1 s 54535 -41011 54581 -40811 8 VDD
port 41 nsew
rlabel metal1 s 54339 -41011 54385 -40811 8 VDD
port 41 nsew
rlabel metal1 s 54143 -41011 54189 -40811 8 VDD
port 41 nsew
rlabel metal1 s 49978 -41205 50024 -40905 8 VDD
port 41 nsew
rlabel metal1 s 49782 -41205 49828 -40905 8 VDD
port 41 nsew
rlabel metal1 s 49586 -41205 49632 -40905 8 VDD
port 41 nsew
rlabel metal1 s 49201 -41076 49247 -40876 8 VDD
port 41 nsew
rlabel metal1 s 49005 -41076 49051 -40876 8 VDD
port 41 nsew
rlabel metal1 s 48809 -41076 48855 -40876 8 VDD
port 41 nsew
rlabel metal1 s 48613 -41076 48659 -40876 8 VDD
port 41 nsew
rlabel metal1 s 47115 -41175 47161 -41075 8 VDD
port 41 nsew
rlabel metal1 s 46919 -41175 46965 -41075 8 VDD
port 41 nsew
rlabel metal1 s 46723 -41175 46769 -41075 8 VDD
port 41 nsew
rlabel metal1 s 46527 -41175 46573 -41075 8 VDD
port 41 nsew
rlabel metal1 s 46310 -41174 46356 -40874 8 VDD
port 41 nsew
rlabel metal1 s 46114 -41174 46160 -40874 8 VDD
port 41 nsew
rlabel metal1 s 45918 -41174 45964 -40874 8 VDD
port 41 nsew
rlabel metal1 s 41920 -41167 41966 -41067 8 VDD
port 41 nsew
rlabel metal1 s 41724 -41167 41770 -41067 8 VDD
port 41 nsew
rlabel metal1 s 41528 -41167 41574 -41067 8 VDD
port 41 nsew
rlabel metal1 s 41332 -41167 41378 -41067 8 VDD
port 41 nsew
rlabel metal1 s 45533 -41045 45579 -40845 8 VDD
port 41 nsew
rlabel metal1 s 45337 -41045 45383 -40845 8 VDD
port 41 nsew
rlabel metal1 s 45141 -41045 45187 -40845 8 VDD
port 41 nsew
rlabel metal1 s 44945 -41045 44991 -40845 8 VDD
port 41 nsew
rlabel metal1 s 41115 -41166 41161 -40866 8 VDD
port 41 nsew
rlabel metal1 s 40919 -41166 40965 -40866 8 VDD
port 41 nsew
rlabel metal1 s 40723 -41166 40769 -40866 8 VDD
port 41 nsew
rlabel metal1 s 40338 -41037 40384 -40837 8 VDD
port 41 nsew
rlabel metal1 s 40142 -41037 40188 -40837 8 VDD
port 41 nsew
rlabel metal1 s 39946 -41037 39992 -40837 8 VDD
port 41 nsew
rlabel metal1 s 39750 -41037 39796 -40837 8 VDD
port 41 nsew
rlabel metal1 s 38252 -41136 38298 -41036 8 VDD
port 41 nsew
rlabel metal1 s 38056 -41136 38102 -41036 8 VDD
port 41 nsew
rlabel metal1 s 37860 -41136 37906 -41036 8 VDD
port 41 nsew
rlabel metal1 s 37664 -41136 37710 -41036 8 VDD
port 41 nsew
rlabel metal1 s 37447 -41135 37493 -40835 8 VDD
port 41 nsew
rlabel metal1 s 37251 -41135 37297 -40835 8 VDD
port 41 nsew
rlabel metal1 s 37055 -41135 37101 -40835 8 VDD
port 41 nsew
rlabel metal1 s 33480 -41156 33526 -41056 8 VDD
port 41 nsew
rlabel metal1 s 33284 -41156 33330 -41056 8 VDD
port 41 nsew
rlabel metal1 s 33088 -41156 33134 -41056 8 VDD
port 41 nsew
rlabel metal1 s 32892 -41156 32938 -41056 8 VDD
port 41 nsew
rlabel metal1 s 36670 -41006 36716 -40806 8 VDD
port 41 nsew
rlabel metal1 s 36474 -41006 36520 -40806 8 VDD
port 41 nsew
rlabel metal1 s 36278 -41006 36324 -40806 8 VDD
port 41 nsew
rlabel metal1 s 36082 -41006 36128 -40806 8 VDD
port 41 nsew
rlabel metal1 s 32675 -41155 32721 -40855 8 VDD
port 41 nsew
rlabel metal1 s 32479 -41155 32525 -40855 8 VDD
port 41 nsew
rlabel metal1 s 32283 -41155 32329 -40855 8 VDD
port 41 nsew
rlabel metal1 s 31898 -41026 31944 -40826 8 VDD
port 41 nsew
rlabel metal1 s 31702 -41026 31748 -40826 8 VDD
port 41 nsew
rlabel metal1 s 31506 -41026 31552 -40826 8 VDD
port 41 nsew
rlabel metal1 s 31310 -41026 31356 -40826 8 VDD
port 41 nsew
rlabel metal1 s 29812 -41125 29858 -41025 8 VDD
port 41 nsew
rlabel metal1 s 29616 -41125 29662 -41025 8 VDD
port 41 nsew
rlabel metal1 s 29420 -41125 29466 -41025 8 VDD
port 41 nsew
rlabel metal1 s 29224 -41125 29270 -41025 8 VDD
port 41 nsew
rlabel metal1 s 29007 -41124 29053 -40824 8 VDD
port 41 nsew
rlabel metal1 s 28811 -41124 28857 -40824 8 VDD
port 41 nsew
rlabel metal1 s 28615 -41124 28661 -40824 8 VDD
port 41 nsew
rlabel metal1 s 28230 -40995 28276 -40795 8 VDD
port 41 nsew
rlabel metal1 s 28034 -40995 28080 -40795 8 VDD
port 41 nsew
rlabel metal1 s 27838 -40995 27884 -40795 8 VDD
port 41 nsew
rlabel metal1 s 27642 -40995 27688 -40795 8 VDD
port 41 nsew
rlabel metal1 s 25263 -41395 25309 -40695 8 VDD
port 41 nsew
rlabel metal1 s 25067 -41395 25113 -40695 8 VDD
port 41 nsew
rlabel metal1 s 24863 -41395 24909 -40695 8 VDD
port 41 nsew
rlabel metal1 s 24667 -41395 24713 -40695 8 VDD
port 41 nsew
rlabel metal1 s 24263 -41395 24309 -40695 8 VDD
port 41 nsew
rlabel metal1 s 24067 -41395 24113 -40695 8 VDD
port 41 nsew
rlabel metal1 s 23863 -41395 23909 -40695 8 VDD
port 41 nsew
rlabel metal1 s 23667 -41395 23713 -40695 8 VDD
port 41 nsew
rlabel metal1 s 23263 -41395 23309 -40695 8 VDD
port 41 nsew
rlabel metal1 s 23067 -41395 23113 -40695 8 VDD
port 41 nsew
rlabel metal1 s 22863 -41395 22909 -40695 8 VDD
port 41 nsew
rlabel metal1 s 22667 -41395 22713 -40695 8 VDD
port 41 nsew
rlabel metal1 s 22179 -41466 22225 -41266 8 VDD
port 41 nsew
rlabel metal1 s 21983 -41466 22029 -41266 8 VDD
port 41 nsew
rlabel metal1 s 21787 -41466 21833 -41266 8 VDD
port 41 nsew
rlabel metal1 s 21254 -41473 21300 -41273 8 VDD
port 41 nsew
rlabel metal1 s 21058 -41473 21104 -41273 8 VDD
port 41 nsew
rlabel metal1 s 20516 -41473 20562 -41273 8 VDD
port 41 nsew
rlabel metal1 s 20320 -41473 20366 -41273 8 VDD
port 41 nsew
rlabel metal1 s 20124 -41473 20170 -41273 8 VDD
port 41 nsew
rlabel metal1 s 19928 -41473 19974 -41273 8 VDD
port 41 nsew
rlabel metal1 s 19208 -41439 19254 -41039 8 VDD
port 41 nsew
rlabel metal1 s 19012 -41439 19058 -41039 8 VDD
port 41 nsew
rlabel metal1 s 18262 -41439 18308 -41039 8 VDD
port 41 nsew
rlabel metal1 s 18066 -41439 18112 -41039 8 VDD
port 41 nsew
rlabel metal1 s 4119 -41667 4165 -41367 8 VDD
port 41 nsew
rlabel metal1 s 3923 -41667 3969 -41367 8 VDD
port 41 nsew
rlabel metal1 s 3727 -41667 3773 -41367 8 VDD
port 41 nsew
rlabel metal1 s 3510 -41668 3556 -41568 8 VDD
port 41 nsew
rlabel metal1 s 3314 -41668 3360 -41568 8 VDD
port 41 nsew
rlabel metal1 s 3118 -41668 3164 -41568 8 VDD
port 41 nsew
rlabel metal1 s 2922 -41668 2968 -41568 8 VDD
port 41 nsew
rlabel metal1 s 2514 -41669 2560 -41369 8 VDD
port 41 nsew
rlabel metal1 s 2318 -41669 2364 -41369 8 VDD
port 41 nsew
rlabel metal1 s 2122 -41669 2168 -41369 8 VDD
port 41 nsew
rlabel metal1 s 1905 -41670 1951 -41570 8 VDD
port 41 nsew
rlabel metal1 s 1709 -41670 1755 -41570 8 VDD
port 41 nsew
rlabel metal1 s 1513 -41670 1559 -41570 8 VDD
port 41 nsew
rlabel metal1 s 1317 -41670 1363 -41570 8 VDD
port 41 nsew
rlabel metal1 s 910 -41683 956 -41483 8 VDD
port 41 nsew
rlabel metal1 s 714 -41683 760 -41483 8 VDD
port 41 nsew
rlabel metal1 s 518 -41683 564 -41483 8 VDD
port 41 nsew
rlabel metal1 s 322 -41683 368 -41483 8 VDD
port 41 nsew
rlabel metal1 s -220 -41683 -174 -41483 2 VDD
port 41 nsew
rlabel metal1 s -416 -41683 -370 -41483 2 VDD
port 41 nsew
rlabel metal1 s -758 -41700 -712 -41500 2 VDD
port 41 nsew
rlabel metal1 s -954 -41700 -908 -41500 2 VDD
port 41 nsew
rlabel metal1 s -1150 -41700 -1104 -41500 2 VDD
port 41 nsew
rlabel metal1 s -1640 -41700 -1594 -41500 2 VDD
port 41 nsew
rlabel metal1 s -1836 -41700 -1790 -41500 2 VDD
port 41 nsew
rlabel metal1 s -2032 -41700 -1986 -41500 2 VDD
port 41 nsew
rlabel metal1 s -3383 -41700 -3337 -41500 2 VDD
port 41 nsew
rlabel metal1 s -3579 -41700 -3533 -41500 2 VDD
port 41 nsew
rlabel metal1 s -3775 -41700 -3729 -41500 2 VDD
port 41 nsew
rlabel metal1 s -4340 -41700 -4294 -41500 2 VDD
port 41 nsew
rlabel metal1 s -4536 -41700 -4490 -41500 2 VDD
port 41 nsew
rlabel metal1 s -4732 -41700 -4686 -41500 2 VDD
port 41 nsew
rlabel metal1 s -6083 -41700 -6037 -41500 2 VDD
port 41 nsew
rlabel metal1 s -6279 -41700 -6233 -41500 2 VDD
port 41 nsew
rlabel metal1 s -6475 -41700 -6429 -41500 2 VDD
port 41 nsew
rlabel metal1 s -16345 -42248 -16299 -41648 2 VDD
port 41 nsew
rlabel metal1 s -16768 -42248 -16722 -41648 2 VDD
port 41 nsew
rlabel metal1 s -16964 -42248 -16918 -41648 2 VDD
port 41 nsew
rlabel metal1 s -17214 -42160 -17168 -42060 2 VDD
port 41 nsew
rlabel metal1 s -17410 -42160 -17364 -42060 2 VDD
port 41 nsew
rlabel metal1 s -17606 -42160 -17560 -42060 2 VDD
port 41 nsew
rlabel metal1 s -17802 -42160 -17756 -42060 2 VDD
port 41 nsew
rlabel metal1 s -18019 -42159 -17973 -41859 2 VDD
port 41 nsew
rlabel metal1 s -18215 -42159 -18169 -41859 2 VDD
port 41 nsew
rlabel metal1 s -18411 -42159 -18365 -41859 2 VDD
port 41 nsew
rlabel metal1 s -8632 -41433 -8586 -41233 2 VDD
port 41 nsew
rlabel metal1 s -8828 -41433 -8782 -41233 2 VDD
port 41 nsew
rlabel metal1 s -9024 -41433 -8978 -41233 2 VDD
port 41 nsew
rlabel metal1 s -9514 -41433 -9468 -41233 2 VDD
port 41 nsew
rlabel metal1 s -9710 -41433 -9664 -41233 2 VDD
port 41 nsew
rlabel metal1 s -9906 -41433 -9860 -41233 2 VDD
port 41 nsew
rlabel metal1 s -11257 -41433 -11211 -41233 2 VDD
port 41 nsew
rlabel metal1 s -11453 -41433 -11407 -41233 2 VDD
port 41 nsew
rlabel metal1 s -11649 -41433 -11603 -41233 2 VDD
port 41 nsew
rlabel metal1 s -12214 -41433 -12168 -41233 2 VDD
port 41 nsew
rlabel metal1 s -12410 -41433 -12364 -41233 2 VDD
port 41 nsew
rlabel metal1 s -12606 -41433 -12560 -41233 2 VDD
port 41 nsew
rlabel metal1 s -13957 -41433 -13911 -41233 2 VDD
port 41 nsew
rlabel metal1 s -14153 -41433 -14107 -41233 2 VDD
port 41 nsew
rlabel metal1 s -14349 -41433 -14303 -41233 2 VDD
port 41 nsew
rlabel metal1 s -18845 -42384 -18719 -40620 2 VDD
port 41 nsew
rlabel metal1 s -19617 -41330 -19571 -40930 2 VDD
port 41 nsew
rlabel metal1 s -19813 -41330 -19767 -40930 2 VDD
port 41 nsew
rlabel metal1 s -20522 -41329 -20476 -40929 2 VDD
port 41 nsew
rlabel metal1 s -20718 -41329 -20672 -40929 2 VDD
port 41 nsew
rlabel metal1 s -21728 -41600 -21682 -41000 2 VDD
port 41 nsew
rlabel metal1 s -21924 -41600 -21878 -41000 2 VDD
port 41 nsew
rlabel metal1 s -26012 -41529 -25612 -41483 2 VDD
port 41 nsew
rlabel metal1 s -26012 -41293 -25612 -41247 2 VDD
port 41 nsew
rlabel metal1 s -26012 -41057 -25612 -41011 2 VDD
port 41 nsew
rlabel metal1 s -26012 -40927 -25612 -40881 2 VDD
port 41 nsew
rlabel metal1 s -26012 -40691 -25612 -40645 2 VDD
port 41 nsew
rlabel metal1 s -2644 -40382 -2598 -40182 2 VDD
port 41 nsew
rlabel metal1 s -2840 -40382 -2794 -40182 2 VDD
port 41 nsew
rlabel metal1 s -3036 -40382 -2990 -40182 2 VDD
port 41 nsew
rlabel metal1 s -3481 -40382 -3435 -40182 2 VDD
port 41 nsew
rlabel metal1 s -3677 -40382 -3631 -40182 2 VDD
port 41 nsew
rlabel metal1 s -3873 -40382 -3827 -40182 2 VDD
port 41 nsew
rlabel metal1 s -5344 -40382 -5298 -40182 2 VDD
port 41 nsew
rlabel metal1 s -5540 -40382 -5494 -40182 2 VDD
port 41 nsew
rlabel metal1 s -5736 -40382 -5690 -40182 2 VDD
port 41 nsew
rlabel metal1 s -6181 -40382 -6135 -40182 2 VDD
port 41 nsew
rlabel metal1 s -6377 -40382 -6331 -40182 2 VDD
port 41 nsew
rlabel metal1 s -6573 -40382 -6527 -40182 2 VDD
port 41 nsew
rlabel metal1 s 22229 -40165 22275 -39765 8 VDD
port 41 nsew
rlabel metal1 s 22033 -40165 22079 -39765 8 VDD
port 41 nsew
rlabel metal1 s 21837 -40165 21883 -39765 8 VDD
port 41 nsew
rlabel metal1 s -7439 -40532 -7393 -39932 2 VDD
port 41 nsew
rlabel metal1 s -7635 -40532 -7589 -39932 2 VDD
port 41 nsew
rlabel metal1 s -8058 -40532 -8012 -39932 2 VDD
port 41 nsew
rlabel metal1 s -18872 -40620 -18693 -40453 2 VDD
port 41 nsew
rlabel metal1 s -26012 -40455 -25612 -40409 2 VDD
port 41 nsew
rlabel metal1 s -26012 -40219 -25612 -40173 2 VDD
port 41 nsew
rlabel metal1 s -10518 -40115 -10472 -39915 2 VDD
port 41 nsew
rlabel metal1 s -10714 -40115 -10668 -39915 2 VDD
port 41 nsew
rlabel metal1 s -10910 -40115 -10864 -39915 2 VDD
port 41 nsew
rlabel metal1 s -11355 -40115 -11309 -39915 2 VDD
port 41 nsew
rlabel metal1 s -11551 -40115 -11505 -39915 2 VDD
port 41 nsew
rlabel metal1 s -11747 -40115 -11701 -39915 2 VDD
port 41 nsew
rlabel metal1 s -13218 -40115 -13172 -39915 2 VDD
port 41 nsew
rlabel metal1 s -13414 -40115 -13368 -39915 2 VDD
port 41 nsew
rlabel metal1 s -13610 -40115 -13564 -39915 2 VDD
port 41 nsew
rlabel metal1 s -14055 -40115 -14009 -39915 2 VDD
port 41 nsew
rlabel metal1 s -14251 -40115 -14205 -39915 2 VDD
port 41 nsew
rlabel metal1 s -14447 -40115 -14401 -39915 2 VDD
port 41 nsew
rlabel metal1 s -26012 -39983 -25612 -39937 2 VDD
port 41 nsew
rlabel metal1 s -26012 -39853 -25612 -39807 2 VDD
port 41 nsew
rlabel metal1 s -26012 -39617 -25612 -39571 2 VDD
port 41 nsew
rlabel metal1 s -26012 -39381 -25612 -39335 2 VDD
port 41 nsew
rlabel metal1 s 25109 -39213 25155 -39013 8 VDD
port 41 nsew
rlabel metal1 s 24913 -39213 24959 -39013 8 VDD
port 41 nsew
rlabel metal1 s 24717 -39213 24763 -39013 8 VDD
port 41 nsew
rlabel metal1 s 23366 -39213 23412 -39013 8 VDD
port 41 nsew
rlabel metal1 s 23170 -39213 23216 -39013 8 VDD
port 41 nsew
rlabel metal1 s 22974 -39213 23020 -39013 8 VDD
port 41 nsew
rlabel metal1 s 22409 -39213 22455 -39013 8 VDD
port 41 nsew
rlabel metal1 s 22213 -39213 22259 -39013 8 VDD
port 41 nsew
rlabel metal1 s 22017 -39213 22063 -39013 8 VDD
port 41 nsew
rlabel metal1 s 20666 -39213 20712 -39013 8 VDD
port 41 nsew
rlabel metal1 s 20470 -39213 20516 -39013 8 VDD
port 41 nsew
rlabel metal1 s 20274 -39213 20320 -39013 8 VDD
port 41 nsew
rlabel metal1 s 19784 -39213 19830 -39013 8 VDD
port 41 nsew
rlabel metal1 s 19588 -39213 19634 -39013 8 VDD
port 41 nsew
rlabel metal1 s 19392 -39213 19438 -39013 8 VDD
port 41 nsew
rlabel metal1 s -26012 -39145 -25612 -39099 2 VDD
port 41 nsew
rlabel metal1 s 86180 -38235 86226 -37935 8 VDD
port 41 nsew
rlabel metal1 s 85984 -38235 86030 -37935 8 VDD
port 41 nsew
rlabel metal1 s 85756 -38435 85802 -37935 8 VDD
port 41 nsew
rlabel metal1 s 85626 -38435 85672 -37935 8 VDD
port 41 nsew
rlabel metal1 s 85031 -38435 85077 -37935 8 VDD
port 41 nsew
rlabel metal1 s 84835 -38435 84881 -37935 8 VDD
port 41 nsew
rlabel metal1 s 83462 -38677 83508 -38077 8 VDD
port 41 nsew
rlabel metal1 s 83039 -38677 83085 -38077 8 VDD
port 41 nsew
rlabel metal1 s 82843 -38677 82889 -38077 8 VDD
port 41 nsew
rlabel metal1 s 82593 -38265 82639 -38165 8 VDD
port 41 nsew
rlabel metal1 s 82397 -38265 82443 -38165 8 VDD
port 41 nsew
rlabel metal1 s 82201 -38265 82247 -38165 8 VDD
port 41 nsew
rlabel metal1 s 82005 -38265 82051 -38165 8 VDD
port 41 nsew
rlabel metal1 s 81788 -38466 81834 -38166 8 VDD
port 41 nsew
rlabel metal1 s 81592 -38466 81638 -38166 8 VDD
port 41 nsew
rlabel metal1 s 81396 -38466 81442 -38166 8 VDD
port 41 nsew
rlabel metal1 s 83902 -37996 84012 -37978 8 VDD
port 41 nsew
rlabel metal1 s 83674 -37984 83748 -37978 8 VDD
port 41 nsew
rlabel metal1 s 83674 -37978 84012 -37882 8 VDD
port 41 nsew
rlabel metal1 s 76816 -38273 76862 -37973 8 VDD
port 41 nsew
rlabel metal1 s 76620 -38273 76666 -37973 8 VDD
port 41 nsew
rlabel metal1 s 76392 -38473 76438 -37973 8 VDD
port 41 nsew
rlabel metal1 s 76262 -38473 76308 -37973 8 VDD
port 41 nsew
rlabel metal1 s 75667 -38473 75713 -37973 8 VDD
port 41 nsew
rlabel metal1 s 75471 -38473 75517 -37973 8 VDD
port 41 nsew
rlabel metal1 s 74098 -38715 74144 -38115 8 VDD
port 41 nsew
rlabel metal1 s 73675 -38715 73721 -38115 8 VDD
port 41 nsew
rlabel metal1 s 73479 -38715 73525 -38115 8 VDD
port 41 nsew
rlabel metal1 s 73229 -38303 73275 -38203 8 VDD
port 41 nsew
rlabel metal1 s 73033 -38303 73079 -38203 8 VDD
port 41 nsew
rlabel metal1 s 72837 -38303 72883 -38203 8 VDD
port 41 nsew
rlabel metal1 s 72641 -38303 72687 -38203 8 VDD
port 41 nsew
rlabel metal1 s 72424 -38504 72470 -38204 8 VDD
port 41 nsew
rlabel metal1 s 72228 -38504 72274 -38204 8 VDD
port 41 nsew
rlabel metal1 s 72032 -38504 72078 -38204 8 VDD
port 41 nsew
rlabel metal1 s 74538 -38034 74648 -38016 8 VDD
port 41 nsew
rlabel metal1 s 74310 -38022 74384 -38016 8 VDD
port 41 nsew
rlabel metal1 s 74310 -38016 74648 -37920 8 VDD
port 41 nsew
rlabel metal1 s 67663 -38290 67709 -37990 8 VDD
port 41 nsew
rlabel metal1 s 67467 -38290 67513 -37990 8 VDD
port 41 nsew
rlabel metal1 s 67239 -38490 67285 -37990 8 VDD
port 41 nsew
rlabel metal1 s 67109 -38490 67155 -37990 8 VDD
port 41 nsew
rlabel metal1 s 66514 -38490 66560 -37990 8 VDD
port 41 nsew
rlabel metal1 s 66318 -38490 66364 -37990 8 VDD
port 41 nsew
rlabel metal1 s 64945 -38732 64991 -38132 8 VDD
port 41 nsew
rlabel metal1 s 64522 -38732 64568 -38132 8 VDD
port 41 nsew
rlabel metal1 s 64326 -38732 64372 -38132 8 VDD
port 41 nsew
rlabel metal1 s 64076 -38320 64122 -38220 8 VDD
port 41 nsew
rlabel metal1 s 63880 -38320 63926 -38220 8 VDD
port 41 nsew
rlabel metal1 s 63684 -38320 63730 -38220 8 VDD
port 41 nsew
rlabel metal1 s 63488 -38320 63534 -38220 8 VDD
port 41 nsew
rlabel metal1 s 63271 -38521 63317 -38221 8 VDD
port 41 nsew
rlabel metal1 s 63075 -38521 63121 -38221 8 VDD
port 41 nsew
rlabel metal1 s 62879 -38521 62925 -38221 8 VDD
port 41 nsew
rlabel metal1 s 58909 -38356 58955 -38056 8 VDD
port 41 nsew
rlabel metal1 s 58713 -38356 58759 -38056 8 VDD
port 41 nsew
rlabel metal1 s 58485 -38556 58531 -38056 8 VDD
port 41 nsew
rlabel metal1 s 58355 -38556 58401 -38056 8 VDD
port 41 nsew
rlabel metal1 s 57760 -38556 57806 -38056 8 VDD
port 41 nsew
rlabel metal1 s 57564 -38556 57610 -38056 8 VDD
port 41 nsew
rlabel metal1 s 56191 -38798 56237 -38198 8 VDD
port 41 nsew
rlabel metal1 s 55768 -38798 55814 -38198 8 VDD
port 41 nsew
rlabel metal1 s 55572 -38798 55618 -38198 8 VDD
port 41 nsew
rlabel metal1 s 55322 -38386 55368 -38286 8 VDD
port 41 nsew
rlabel metal1 s 55126 -38386 55172 -38286 8 VDD
port 41 nsew
rlabel metal1 s 54930 -38386 54976 -38286 8 VDD
port 41 nsew
rlabel metal1 s 54734 -38386 54780 -38286 8 VDD
port 41 nsew
rlabel metal1 s 54517 -38587 54563 -38287 8 VDD
port 41 nsew
rlabel metal1 s 54321 -38587 54367 -38287 8 VDD
port 41 nsew
rlabel metal1 s 54125 -38587 54171 -38287 8 VDD
port 41 nsew
rlabel metal1 s 56631 -38117 56741 -38099 8 VDD
port 41 nsew
rlabel metal1 s 56403 -38105 56477 -38099 8 VDD
port 41 nsew
rlabel metal1 s 65385 -38051 65495 -38033 8 VDD
port 41 nsew
rlabel metal1 s 65157 -38039 65231 -38033 8 VDD
port 41 nsew
rlabel metal1 s 74538 -37920 74648 -37884 8 VDD
port 41 nsew
rlabel metal1 s 74310 -37920 74384 -37904 8 VDD
port 41 nsew
rlabel metal1 s 65157 -38033 65495 -37937 8 VDD
port 41 nsew
rlabel metal1 s 56403 -38099 56741 -38003 8 VDD
port 41 nsew
rlabel metal1 s 49711 -38390 49757 -38090 8 VDD
port 41 nsew
rlabel metal1 s 49515 -38390 49561 -38090 8 VDD
port 41 nsew
rlabel metal1 s 49287 -38590 49333 -38090 8 VDD
port 41 nsew
rlabel metal1 s 49157 -38590 49203 -38090 8 VDD
port 41 nsew
rlabel metal1 s 48562 -38590 48608 -38090 8 VDD
port 41 nsew
rlabel metal1 s 48366 -38590 48412 -38090 8 VDD
port 41 nsew
rlabel metal1 s 46993 -38832 47039 -38232 8 VDD
port 41 nsew
rlabel metal1 s 46570 -38832 46616 -38232 8 VDD
port 41 nsew
rlabel metal1 s 46374 -38832 46420 -38232 8 VDD
port 41 nsew
rlabel metal1 s 46124 -38420 46170 -38320 8 VDD
port 41 nsew
rlabel metal1 s 45928 -38420 45974 -38320 8 VDD
port 41 nsew
rlabel metal1 s 45732 -38420 45778 -38320 8 VDD
port 41 nsew
rlabel metal1 s 45536 -38420 45582 -38320 8 VDD
port 41 nsew
rlabel metal1 s 45319 -38621 45365 -38321 8 VDD
port 41 nsew
rlabel metal1 s 45123 -38621 45169 -38321 8 VDD
port 41 nsew
rlabel metal1 s 44927 -38621 44973 -38321 8 VDD
port 41 nsew
rlabel metal1 s 47433 -38151 47543 -38133 8 VDD
port 41 nsew
rlabel metal1 s 47205 -38139 47279 -38133 8 VDD
port 41 nsew
rlabel metal1 s 56631 -38003 56741 -37967 8 VDD
port 41 nsew
rlabel metal1 s 56403 -38003 56477 -37987 8 VDD
port 41 nsew
rlabel metal1 s 47205 -38133 47543 -38037 8 VDD
port 41 nsew
rlabel metal1 s 40848 -38351 40894 -38051 8 VDD
port 41 nsew
rlabel metal1 s 40652 -38351 40698 -38051 8 VDD
port 41 nsew
rlabel metal1 s 40424 -38551 40470 -38051 8 VDD
port 41 nsew
rlabel metal1 s 40294 -38551 40340 -38051 8 VDD
port 41 nsew
rlabel metal1 s 39699 -38551 39745 -38051 8 VDD
port 41 nsew
rlabel metal1 s 39503 -38551 39549 -38051 8 VDD
port 41 nsew
rlabel metal1 s 38130 -38793 38176 -38193 8 VDD
port 41 nsew
rlabel metal1 s 37707 -38793 37753 -38193 8 VDD
port 41 nsew
rlabel metal1 s 37511 -38793 37557 -38193 8 VDD
port 41 nsew
rlabel metal1 s 37261 -38381 37307 -38281 8 VDD
port 41 nsew
rlabel metal1 s 37065 -38381 37111 -38281 8 VDD
port 41 nsew
rlabel metal1 s 36869 -38381 36915 -38281 8 VDD
port 41 nsew
rlabel metal1 s 36673 -38381 36719 -38281 8 VDD
port 41 nsew
rlabel metal1 s 36456 -38582 36502 -38282 8 VDD
port 41 nsew
rlabel metal1 s 36260 -38582 36306 -38282 8 VDD
port 41 nsew
rlabel metal1 s 36064 -38582 36110 -38282 8 VDD
port 41 nsew
rlabel metal1 s 38570 -38112 38680 -38094 8 VDD
port 41 nsew
rlabel metal1 s 38342 -38100 38416 -38094 8 VDD
port 41 nsew
rlabel metal1 s 47433 -38037 47543 -38001 8 VDD
port 41 nsew
rlabel metal1 s 47205 -38037 47279 -38021 8 VDD
port 41 nsew
rlabel metal1 s 38342 -38094 38680 -37998 8 VDD
port 41 nsew
rlabel metal1 s 32408 -38340 32454 -38040 8 VDD
port 41 nsew
rlabel metal1 s 32212 -38340 32258 -38040 8 VDD
port 41 nsew
rlabel metal1 s 31984 -38540 32030 -38040 8 VDD
port 41 nsew
rlabel metal1 s 31854 -38540 31900 -38040 8 VDD
port 41 nsew
rlabel metal1 s 31259 -38540 31305 -38040 8 VDD
port 41 nsew
rlabel metal1 s 31063 -38540 31109 -38040 8 VDD
port 41 nsew
rlabel metal1 s 29690 -38782 29736 -38182 8 VDD
port 41 nsew
rlabel metal1 s 29267 -38782 29313 -38182 8 VDD
port 41 nsew
rlabel metal1 s 29071 -38782 29117 -38182 8 VDD
port 41 nsew
rlabel metal1 s 28821 -38370 28867 -38270 8 VDD
port 41 nsew
rlabel metal1 s 28625 -38370 28671 -38270 8 VDD
port 41 nsew
rlabel metal1 s 28429 -38370 28475 -38270 8 VDD
port 41 nsew
rlabel metal1 s 28233 -38370 28279 -38270 8 VDD
port 41 nsew
rlabel metal1 s 28016 -38571 28062 -38271 8 VDD
port 41 nsew
rlabel metal1 s 27820 -38571 27866 -38271 8 VDD
port 41 nsew
rlabel metal1 s 27624 -38571 27670 -38271 8 VDD
port 41 nsew
rlabel metal1 s 18267 -39093 18313 -38493 8 VDD
port 41 nsew
rlabel metal1 s 18071 -39093 18117 -38493 8 VDD
port 41 nsew
rlabel metal1 s -2644 -38944 -2598 -38744 2 VDD
port 41 nsew
rlabel metal1 s -2840 -38944 -2794 -38744 2 VDD
port 41 nsew
rlabel metal1 s -3036 -38944 -2990 -38744 2 VDD
port 41 nsew
rlabel metal1 s -3481 -38944 -3435 -38744 2 VDD
port 41 nsew
rlabel metal1 s -3677 -38944 -3631 -38744 2 VDD
port 41 nsew
rlabel metal1 s -3873 -38944 -3827 -38744 2 VDD
port 41 nsew
rlabel metal1 s -5344 -38944 -5298 -38744 2 VDD
port 41 nsew
rlabel metal1 s -5540 -38944 -5494 -38744 2 VDD
port 41 nsew
rlabel metal1 s -5736 -38944 -5690 -38744 2 VDD
port 41 nsew
rlabel metal1 s -6181 -38944 -6135 -38744 2 VDD
port 41 nsew
rlabel metal1 s -6377 -38944 -6331 -38744 2 VDD
port 41 nsew
rlabel metal1 s -6573 -38944 -6527 -38744 2 VDD
port 41 nsew
rlabel metal1 s -11226 -38834 -11180 -38734 2 VDD
port 41 nsew
rlabel metal1 s -11422 -38834 -11376 -38734 2 VDD
port 41 nsew
rlabel metal1 s -11618 -38834 -11572 -38734 2 VDD
port 41 nsew
rlabel metal1 s -11814 -38834 -11768 -38734 2 VDD
port 41 nsew
rlabel metal1 s -12031 -39035 -11985 -38735 2 VDD
port 41 nsew
rlabel metal1 s -12227 -39035 -12181 -38735 2 VDD
port 41 nsew
rlabel metal1 s -12423 -39035 -12377 -38735 2 VDD
port 41 nsew
rlabel metal1 s -12808 -39064 -12762 -38864 2 VDD
port 41 nsew
rlabel metal1 s -13004 -39064 -12958 -38864 2 VDD
port 41 nsew
rlabel metal1 s -13200 -39064 -13154 -38864 2 VDD
port 41 nsew
rlabel metal1 s -13396 -39064 -13350 -38864 2 VDD
port 41 nsew
rlabel metal1 s -26012 -38909 -25612 -38863 2 VDD
port 41 nsew
rlabel metal1 s -26012 -38673 -25612 -38627 2 VDD
port 41 nsew
rlabel metal1 s -26012 -38437 -25612 -38391 2 VDD
port 41 nsew
rlabel metal1 s 30130 -38101 30240 -38083 8 VDD
port 41 nsew
rlabel metal1 s 29902 -38089 29976 -38083 8 VDD
port 41 nsew
rlabel metal1 s 38570 -37998 38680 -37962 8 VDD
port 41 nsew
rlabel metal1 s 38342 -37998 38416 -37982 8 VDD
port 41 nsew
rlabel metal1 s 29902 -38083 30240 -37987 8 VDD
port 41 nsew
rlabel metal1 s 30130 -37987 30240 -37951 8 VDD
port 41 nsew
rlabel metal1 s 29902 -37987 29976 -37971 8 VDD
port 41 nsew
rlabel metal1 s 65385 -37937 65495 -37901 8 VDD
port 41 nsew
rlabel metal1 s 65157 -37937 65231 -37921 8 VDD
port 41 nsew
rlabel metal1 s 83902 -37882 84012 -37846 8 VDD
port 41 nsew
rlabel metal1 s 83674 -37882 83748 -37866 8 VDD
port 41 nsew
rlabel metal1 s 83592 -37567 83638 -37467 8 VDD
port 41 nsew
rlabel metal1 s 83396 -37567 83442 -37467 8 VDD
port 41 nsew
rlabel metal1 s 83200 -37567 83246 -37467 8 VDD
port 41 nsew
rlabel metal1 s 83004 -37567 83050 -37467 8 VDD
port 41 nsew
rlabel metal1 s 82787 -37566 82833 -37266 8 VDD
port 41 nsew
rlabel metal1 s 82591 -37566 82637 -37266 8 VDD
port 41 nsew
rlabel metal1 s 82395 -37566 82441 -37266 8 VDD
port 41 nsew
rlabel metal1 s 74228 -37605 74274 -37505 8 VDD
port 41 nsew
rlabel metal1 s 74032 -37605 74078 -37505 8 VDD
port 41 nsew
rlabel metal1 s 73836 -37605 73882 -37505 8 VDD
port 41 nsew
rlabel metal1 s 73640 -37605 73686 -37505 8 VDD
port 41 nsew
rlabel metal1 s 82010 -37437 82056 -37237 8 VDD
port 41 nsew
rlabel metal1 s 81814 -37437 81860 -37237 8 VDD
port 41 nsew
rlabel metal1 s 81618 -37437 81664 -37237 8 VDD
port 41 nsew
rlabel metal1 s 81422 -37437 81468 -37237 8 VDD
port 41 nsew
rlabel metal1 s 73423 -37604 73469 -37304 8 VDD
port 41 nsew
rlabel metal1 s 73227 -37604 73273 -37304 8 VDD
port 41 nsew
rlabel metal1 s 73031 -37604 73077 -37304 8 VDD
port 41 nsew
rlabel metal1 s 65075 -37622 65121 -37522 8 VDD
port 41 nsew
rlabel metal1 s 64879 -37622 64925 -37522 8 VDD
port 41 nsew
rlabel metal1 s 64683 -37622 64729 -37522 8 VDD
port 41 nsew
rlabel metal1 s 64487 -37622 64533 -37522 8 VDD
port 41 nsew
rlabel metal1 s 72646 -37475 72692 -37275 8 VDD
port 41 nsew
rlabel metal1 s 72450 -37475 72496 -37275 8 VDD
port 41 nsew
rlabel metal1 s 72254 -37475 72300 -37275 8 VDD
port 41 nsew
rlabel metal1 s 72058 -37475 72104 -37275 8 VDD
port 41 nsew
rlabel metal1 s 64270 -37621 64316 -37321 8 VDD
port 41 nsew
rlabel metal1 s 64074 -37621 64120 -37321 8 VDD
port 41 nsew
rlabel metal1 s 63878 -37621 63924 -37321 8 VDD
port 41 nsew
rlabel metal1 s 56321 -37688 56367 -37588 8 VDD
port 41 nsew
rlabel metal1 s 56125 -37688 56171 -37588 8 VDD
port 41 nsew
rlabel metal1 s 55929 -37688 55975 -37588 8 VDD
port 41 nsew
rlabel metal1 s 55733 -37688 55779 -37588 8 VDD
port 41 nsew
rlabel metal1 s 63493 -37492 63539 -37292 8 VDD
port 41 nsew
rlabel metal1 s 63297 -37492 63343 -37292 8 VDD
port 41 nsew
rlabel metal1 s 63101 -37492 63147 -37292 8 VDD
port 41 nsew
rlabel metal1 s 62905 -37492 62951 -37292 8 VDD
port 41 nsew
rlabel metal1 s 55516 -37687 55562 -37387 8 VDD
port 41 nsew
rlabel metal1 s 55320 -37687 55366 -37387 8 VDD
port 41 nsew
rlabel metal1 s 55124 -37687 55170 -37387 8 VDD
port 41 nsew
rlabel metal1 s 47123 -37722 47169 -37622 8 VDD
port 41 nsew
rlabel metal1 s 46927 -37722 46973 -37622 8 VDD
port 41 nsew
rlabel metal1 s 46731 -37722 46777 -37622 8 VDD
port 41 nsew
rlabel metal1 s 46535 -37722 46581 -37622 8 VDD
port 41 nsew
rlabel metal1 s 54739 -37558 54785 -37358 8 VDD
port 41 nsew
rlabel metal1 s 54543 -37558 54589 -37358 8 VDD
port 41 nsew
rlabel metal1 s 54347 -37558 54393 -37358 8 VDD
port 41 nsew
rlabel metal1 s 54151 -37558 54197 -37358 8 VDD
port 41 nsew
rlabel metal1 s 46318 -37721 46364 -37421 8 VDD
port 41 nsew
rlabel metal1 s 46122 -37721 46168 -37421 8 VDD
port 41 nsew
rlabel metal1 s 45926 -37721 45972 -37421 8 VDD
port 41 nsew
rlabel metal1 s 25207 -37895 25253 -37695 8 VDD
port 41 nsew
rlabel metal1 s 25011 -37895 25057 -37695 8 VDD
port 41 nsew
rlabel metal1 s 24815 -37895 24861 -37695 8 VDD
port 41 nsew
rlabel metal1 s 24370 -37895 24416 -37695 8 VDD
port 41 nsew
rlabel metal1 s 24174 -37895 24220 -37695 8 VDD
port 41 nsew
rlabel metal1 s 23978 -37895 24024 -37695 8 VDD
port 41 nsew
rlabel metal1 s 22507 -37895 22553 -37695 8 VDD
port 41 nsew
rlabel metal1 s 22311 -37895 22357 -37695 8 VDD
port 41 nsew
rlabel metal1 s 22115 -37895 22161 -37695 8 VDD
port 41 nsew
rlabel metal1 s 21670 -37895 21716 -37695 8 VDD
port 41 nsew
rlabel metal1 s 21474 -37895 21520 -37695 8 VDD
port 41 nsew
rlabel metal1 s 21278 -37895 21324 -37695 8 VDD
port 41 nsew
rlabel metal1 s 45541 -37592 45587 -37392 8 VDD
port 41 nsew
rlabel metal1 s 45345 -37592 45391 -37392 8 VDD
port 41 nsew
rlabel metal1 s 45149 -37592 45195 -37392 8 VDD
port 41 nsew
rlabel metal1 s 44953 -37592 44999 -37392 8 VDD
port 41 nsew
rlabel metal1 s 38260 -37683 38306 -37583 8 VDD
port 41 nsew
rlabel metal1 s 38064 -37683 38110 -37583 8 VDD
port 41 nsew
rlabel metal1 s 37868 -37683 37914 -37583 8 VDD
port 41 nsew
rlabel metal1 s 37672 -37683 37718 -37583 8 VDD
port 41 nsew
rlabel metal1 s 37455 -37682 37501 -37382 8 VDD
port 41 nsew
rlabel metal1 s 37259 -37682 37305 -37382 8 VDD
port 41 nsew
rlabel metal1 s 37063 -37682 37109 -37382 8 VDD
port 41 nsew
rlabel metal1 s 29820 -37672 29866 -37572 8 VDD
port 41 nsew
rlabel metal1 s 29624 -37672 29670 -37572 8 VDD
port 41 nsew
rlabel metal1 s 29428 -37672 29474 -37572 8 VDD
port 41 nsew
rlabel metal1 s 29232 -37672 29278 -37572 8 VDD
port 41 nsew
rlabel metal1 s 36678 -37553 36724 -37353 8 VDD
port 41 nsew
rlabel metal1 s 36482 -37553 36528 -37353 8 VDD
port 41 nsew
rlabel metal1 s 36286 -37553 36332 -37353 8 VDD
port 41 nsew
rlabel metal1 s 36090 -37553 36136 -37353 8 VDD
port 41 nsew
rlabel metal1 s 29015 -37671 29061 -37371 8 VDD
port 41 nsew
rlabel metal1 s 28819 -37671 28865 -37371 8 VDD
port 41 nsew
rlabel metal1 s 28623 -37671 28669 -37371 8 VDD
port 41 nsew
rlabel metal1 s 28238 -37542 28284 -37342 8 VDD
port 41 nsew
rlabel metal1 s 28042 -37542 28088 -37342 8 VDD
port 41 nsew
rlabel metal1 s 27846 -37542 27892 -37342 8 VDD
port 41 nsew
rlabel metal1 s 27650 -37542 27696 -37342 8 VDD
port 41 nsew
rlabel metal1 s 8044 -37645 8090 -37445 8 VDD
port 41 nsew
rlabel metal1 s 7848 -37645 7894 -37445 8 VDD
port 41 nsew
rlabel metal1 s 7735 -37645 7781 -37445 8 VDD
port 41 nsew
rlabel metal1 s 7539 -37645 7585 -37445 8 VDD
port 41 nsew
rlabel metal1 s 7425 -37645 7471 -37445 8 VDD
port 41 nsew
rlabel metal1 s 7229 -37645 7275 -37445 8 VDD
port 41 nsew
rlabel metal1 s 7033 -37645 7079 -37445 8 VDD
port 41 nsew
rlabel metal1 s 5872 -37634 5918 -37434 8 VDD
port 41 nsew
rlabel metal1 s 5676 -37634 5722 -37434 8 VDD
port 41 nsew
rlabel metal1 s 5480 -37634 5526 -37434 8 VDD
port 41 nsew
rlabel metal1 s 5284 -37634 5330 -37434 8 VDD
port 41 nsew
rlabel metal1 s 4742 -37634 4788 -37434 8 VDD
port 41 nsew
rlabel metal1 s 4546 -37634 4592 -37434 8 VDD
port 41 nsew
rlabel metal1 s 4119 -37759 4165 -37459 8 VDD
port 41 nsew
rlabel metal1 s 3923 -37759 3969 -37459 8 VDD
port 41 nsew
rlabel metal1 s 3727 -37759 3773 -37459 8 VDD
port 41 nsew
rlabel metal1 s 3510 -37558 3556 -37458 8 VDD
port 41 nsew
rlabel metal1 s 3314 -37558 3360 -37458 8 VDD
port 41 nsew
rlabel metal1 s 3118 -37558 3164 -37458 8 VDD
port 41 nsew
rlabel metal1 s 2922 -37558 2968 -37458 8 VDD
port 41 nsew
rlabel metal1 s 2514 -37757 2560 -37457 8 VDD
port 41 nsew
rlabel metal1 s 2318 -37757 2364 -37457 8 VDD
port 41 nsew
rlabel metal1 s 2122 -37757 2168 -37457 8 VDD
port 41 nsew
rlabel metal1 s 1905 -37556 1951 -37456 8 VDD
port 41 nsew
rlabel metal1 s 1709 -37556 1755 -37456 8 VDD
port 41 nsew
rlabel metal1 s 1513 -37556 1559 -37456 8 VDD
port 41 nsew
rlabel metal1 s 1317 -37556 1363 -37456 8 VDD
port 41 nsew
rlabel metal1 s 910 -37643 956 -37443 8 VDD
port 41 nsew
rlabel metal1 s 714 -37643 760 -37443 8 VDD
port 41 nsew
rlabel metal1 s 518 -37643 564 -37443 8 VDD
port 41 nsew
rlabel metal1 s 322 -37643 368 -37443 8 VDD
port 41 nsew
rlabel metal1 s -220 -37643 -174 -37443 2 VDD
port 41 nsew
rlabel metal1 s -416 -37643 -370 -37443 2 VDD
port 41 nsew
rlabel metal1 s -758 -37626 -712 -37426 2 VDD
port 41 nsew
rlabel metal1 s -954 -37626 -908 -37426 2 VDD
port 41 nsew
rlabel metal1 s -1150 -37626 -1104 -37426 2 VDD
port 41 nsew
rlabel metal1 s -1640 -37626 -1594 -37426 2 VDD
port 41 nsew
rlabel metal1 s -1836 -37626 -1790 -37426 2 VDD
port 41 nsew
rlabel metal1 s -2032 -37626 -1986 -37426 2 VDD
port 41 nsew
rlabel metal1 s -3383 -37626 -3337 -37426 2 VDD
port 41 nsew
rlabel metal1 s -3579 -37626 -3533 -37426 2 VDD
port 41 nsew
rlabel metal1 s -3775 -37626 -3729 -37426 2 VDD
port 41 nsew
rlabel metal1 s -4340 -37626 -4294 -37426 2 VDD
port 41 nsew
rlabel metal1 s -4536 -37626 -4490 -37426 2 VDD
port 41 nsew
rlabel metal1 s -4732 -37626 -4686 -37426 2 VDD
port 41 nsew
rlabel metal1 s -6083 -37626 -6037 -37426 2 VDD
port 41 nsew
rlabel metal1 s -6279 -37626 -6233 -37426 2 VDD
port 41 nsew
rlabel metal1 s -6475 -37626 -6429 -37426 2 VDD
port 41 nsew
rlabel metal1 s -11356 -38224 -11310 -37624 2 VDD
port 41 nsew
rlabel metal1 s -11779 -38224 -11733 -37624 2 VDD
port 41 nsew
rlabel metal1 s -11975 -38224 -11929 -37624 2 VDD
port 41 nsew
rlabel metal1 s -26012 -38201 -25612 -38155 2 VDD
port 41 nsew
rlabel metal1 s -12225 -38136 -12179 -38036 2 VDD
port 41 nsew
rlabel metal1 s -12421 -38136 -12375 -38036 2 VDD
port 41 nsew
rlabel metal1 s -12617 -38136 -12571 -38036 2 VDD
port 41 nsew
rlabel metal1 s -12813 -38136 -12767 -38036 2 VDD
port 41 nsew
rlabel metal1 s -13030 -38135 -12984 -37835 2 VDD
port 41 nsew
rlabel metal1 s -13226 -38135 -13180 -37835 2 VDD
port 41 nsew
rlabel metal1 s -13422 -38135 -13376 -37835 2 VDD
port 41 nsew
rlabel metal1 s -16215 -37858 -16169 -37758 2 VDD
port 41 nsew
rlabel metal1 s -16411 -37858 -16365 -37758 2 VDD
port 41 nsew
rlabel metal1 s -16607 -37858 -16561 -37758 2 VDD
port 41 nsew
rlabel metal1 s -16803 -37858 -16757 -37758 2 VDD
port 41 nsew
rlabel metal1 s -17020 -38059 -16974 -37759 2 VDD
port 41 nsew
rlabel metal1 s -17216 -38059 -17170 -37759 2 VDD
port 41 nsew
rlabel metal1 s -17412 -38059 -17366 -37759 2 VDD
port 41 nsew
rlabel metal1 s -17797 -38088 -17751 -37888 2 VDD
port 41 nsew
rlabel metal1 s -17993 -38088 -17947 -37888 2 VDD
port 41 nsew
rlabel metal1 s -18189 -38088 -18143 -37888 2 VDD
port 41 nsew
rlabel metal1 s -18385 -38088 -18339 -37888 2 VDD
port 41 nsew
rlabel metal1 s -18890 -37911 -18844 -37711 2 VDD
port 41 nsew
rlabel metal1 s -19086 -37911 -19040 -37711 2 VDD
port 41 nsew
rlabel metal1 s -19628 -37911 -19582 -37711 2 VDD
port 41 nsew
rlabel metal1 s -19824 -37911 -19778 -37711 2 VDD
port 41 nsew
rlabel metal1 s -20020 -37911 -19974 -37711 2 VDD
port 41 nsew
rlabel metal1 s -20216 -37911 -20170 -37711 2 VDD
port 41 nsew
rlabel metal1 s -20792 -37905 -20746 -37805 2 VDD
port 41 nsew
rlabel metal1 s -20988 -37905 -20942 -37805 2 VDD
port 41 nsew
rlabel metal1 s -21184 -37905 -21138 -37805 2 VDD
port 41 nsew
rlabel metal1 s -21380 -37905 -21334 -37805 2 VDD
port 41 nsew
rlabel metal1 s -21597 -38106 -21551 -37806 2 VDD
port 41 nsew
rlabel metal1 s -21793 -38106 -21747 -37806 2 VDD
port 41 nsew
rlabel metal1 s -21989 -38106 -21943 -37806 2 VDD
port 41 nsew
rlabel metal1 s -26012 -37965 -25612 -37919 2 VDD
port 41 nsew
rlabel metal1 s -26012 -37717 -25612 -37671 2 VDD
port 41 nsew
rlabel metal1 s -26012 -37481 -25612 -37435 2 VDD
port 41 nsew
rlabel metal1 s 2837 -37396 2960 -37383 8 VDD
port 41 nsew
rlabel metal1 s 2448 -37397 2571 -37383 8 VDD
port 41 nsew
rlabel metal1 s 7038 -37377 7161 -37358 8 VDD
port 41 nsew
rlabel metal1 s 5822 -37376 5945 -37358 8 VDD
port 41 nsew
rlabel metal1 s 5822 -37358 7161 -37253 8 VDD
port 41 nsew
rlabel metal1 s 7038 -37253 7161 -37241 8 VDD
port 41 nsew
rlabel metal1 s 5822 -37253 5945 -37240 8 VDD
port 41 nsew
rlabel metal1 s 4466 -37371 4589 -37353 8 VDD
port 41 nsew
rlabel metal1 s 4065 -37373 4188 -37353 8 VDD
port 41 nsew
rlabel metal1 s 4065 -37353 4589 -37246 8 VDD
port 41 nsew
rlabel metal1 s 2448 -37383 2960 -37276 8 VDD
port 41 nsew
rlabel metal1 s 2837 -37276 2960 -37260 8 VDD
port 41 nsew
rlabel metal1 s 2448 -37276 2571 -37261 8 VDD
port 41 nsew
rlabel metal1 s -530 -37384 -407 -37376 2 VDD
port 41 nsew
rlabel metal1 s -824 -37385 -701 -37376 2 VDD
port 41 nsew
rlabel metal1 s -824 -37376 -407 -37261 2 VDD
port 41 nsew
rlabel metal1 s -530 -37261 -407 -37248 2 VDD
port 41 nsew
rlabel metal1 s -824 -37261 -701 -37249 2 VDD
port 41 nsew
rlabel metal1 s 4466 -37246 4589 -37235 8 VDD
port 41 nsew
rlabel metal1 s 4065 -37246 4188 -37237 8 VDD
port 41 nsew
rlabel metal1 s -4650 -36719 -4527 -36583 2 VDD
port 41 nsew
rlabel metal1 s 400 -36467 706 -36405 8 VDD
port 41 nsew
rlabel metal1 s -2083 -36575 -1960 -36439 2 VDD
port 41 nsew
rlabel metal1 s 400 -36405 523 -36404 8 VDD
port 41 nsew
rlabel metal1 s 405 -36404 519 -35987 8 VDD
port 41 nsew
rlabel metal1 s -2078 -36439 -1964 -35987 2 VDD
port 41 nsew
rlabel metal1 s 401 -35987 524 -35851 8 VDD
port 41 nsew
rlabel metal1 s -2082 -35987 -1959 -35851 2 VDD
port 41 nsew
rlabel metal1 s -4645 -36583 -4531 -35952 2 VDD
port 41 nsew
rlabel metal1 s -5924 -36723 -5878 -36523 2 VDD
port 41 nsew
rlabel metal1 s -6120 -36723 -6074 -36523 2 VDD
port 41 nsew
rlabel metal1 s -6316 -36723 -6270 -36523 2 VDD
port 41 nsew
rlabel metal1 s -16345 -37248 -16299 -36648 2 VDD
port 41 nsew
rlabel metal1 s -16768 -37248 -16722 -36648 2 VDD
port 41 nsew
rlabel metal1 s -16964 -37248 -16918 -36648 2 VDD
port 41 nsew
rlabel metal1 s -26012 -37245 -25612 -37199 2 VDD
port 41 nsew
rlabel metal1 s -17214 -37160 -17168 -37060 2 VDD
port 41 nsew
rlabel metal1 s -17410 -37160 -17364 -37060 2 VDD
port 41 nsew
rlabel metal1 s -17606 -37160 -17560 -37060 2 VDD
port 41 nsew
rlabel metal1 s -17802 -37160 -17756 -37060 2 VDD
port 41 nsew
rlabel metal1 s -18019 -37159 -17973 -36859 2 VDD
port 41 nsew
rlabel metal1 s -18215 -37159 -18169 -36859 2 VDD
port 41 nsew
rlabel metal1 s -18411 -37159 -18365 -36859 2 VDD
port 41 nsew
rlabel metal1 s -26012 -37009 -25612 -36963 2 VDD
port 41 nsew
rlabel metal1 s -26012 -36773 -25612 -36727 2 VDD
port 41 nsew
rlabel metal1 s -8632 -36506 -8586 -36306 2 VDD
port 41 nsew
rlabel metal1 s -8828 -36506 -8782 -36306 2 VDD
port 41 nsew
rlabel metal1 s -9024 -36506 -8978 -36306 2 VDD
port 41 nsew
rlabel metal1 s -9514 -36506 -9468 -36306 2 VDD
port 41 nsew
rlabel metal1 s -9710 -36506 -9664 -36306 2 VDD
port 41 nsew
rlabel metal1 s -9906 -36506 -9860 -36306 2 VDD
port 41 nsew
rlabel metal1 s -11257 -36506 -11211 -36306 2 VDD
port 41 nsew
rlabel metal1 s -11453 -36506 -11407 -36306 2 VDD
port 41 nsew
rlabel metal1 s -11649 -36506 -11603 -36306 2 VDD
port 41 nsew
rlabel metal1 s -12214 -36506 -12168 -36306 2 VDD
port 41 nsew
rlabel metal1 s -12410 -36506 -12364 -36306 2 VDD
port 41 nsew
rlabel metal1 s -12606 -36506 -12560 -36306 2 VDD
port 41 nsew
rlabel metal1 s -13957 -36506 -13911 -36306 2 VDD
port 41 nsew
rlabel metal1 s -14153 -36506 -14107 -36306 2 VDD
port 41 nsew
rlabel metal1 s -14349 -36506 -14303 -36306 2 VDD
port 41 nsew
rlabel metal1 s -26012 -36537 -25612 -36491 2 VDD
port 41 nsew
rlabel metal1 s -26012 -36301 -25612 -36255 2 VDD
port 41 nsew
rlabel metal1 s -4649 -35952 -4526 -35816 2 VDD
port 41 nsew
rlabel metal1 s -18850 -35996 -18804 -35896 2 VDD
port 41 nsew
rlabel metal1 s -19046 -35996 -19000 -35896 2 VDD
port 41 nsew
rlabel metal1 s -19242 -35996 -19196 -35896 2 VDD
port 41 nsew
rlabel metal1 s -19438 -35996 -19392 -35896 2 VDD
port 41 nsew
rlabel metal1 s -19655 -36197 -19609 -35897 2 VDD
port 41 nsew
rlabel metal1 s -19851 -36197 -19805 -35897 2 VDD
port 41 nsew
rlabel metal1 s -20047 -36197 -20001 -35897 2 VDD
port 41 nsew
rlabel metal1 s -26012 -36065 -25612 -36019 2 VDD
port 41 nsew
rlabel metal1 s -20720 -35975 -20674 -35775 2 VDD
port 41 nsew
rlabel metal1 s -20916 -35975 -20870 -35775 2 VDD
port 41 nsew
rlabel metal1 s -21458 -35975 -21412 -35775 2 VDD
port 41 nsew
rlabel metal1 s -21654 -35975 -21608 -35775 2 VDD
port 41 nsew
rlabel metal1 s -21850 -35975 -21804 -35775 2 VDD
port 41 nsew
rlabel metal1 s -22046 -35975 -22000 -35775 2 VDD
port 41 nsew
rlabel metal1 s -26012 -35829 -25612 -35783 2 VDD
port 41 nsew
rlabel metal1 s 8034 -35394 8080 -35194 8 VDD
port 41 nsew
rlabel metal1 s 7838 -35394 7884 -35194 8 VDD
port 41 nsew
rlabel metal1 s 7725 -35394 7771 -35194 8 VDD
port 41 nsew
rlabel metal1 s 7529 -35394 7575 -35194 8 VDD
port 41 nsew
rlabel metal1 s 7415 -35394 7461 -35194 8 VDD
port 41 nsew
rlabel metal1 s 7219 -35394 7265 -35194 8 VDD
port 41 nsew
rlabel metal1 s 7023 -35394 7069 -35194 8 VDD
port 41 nsew
rlabel metal1 s 5034 -35394 5080 -35194 8 VDD
port 41 nsew
rlabel metal1 s 4838 -35394 4884 -35194 8 VDD
port 41 nsew
rlabel metal1 s 4725 -35394 4771 -35194 8 VDD
port 41 nsew
rlabel metal1 s 4529 -35394 4575 -35194 8 VDD
port 41 nsew
rlabel metal1 s 4415 -35394 4461 -35194 8 VDD
port 41 nsew
rlabel metal1 s 4219 -35394 4265 -35194 8 VDD
port 41 nsew
rlabel metal1 s 4023 -35394 4069 -35194 8 VDD
port 41 nsew
rlabel metal1 s 2534 -35394 2580 -35194 8 VDD
port 41 nsew
rlabel metal1 s 2338 -35394 2384 -35194 8 VDD
port 41 nsew
rlabel metal1 s 2225 -35394 2271 -35194 8 VDD
port 41 nsew
rlabel metal1 s 2029 -35394 2075 -35194 8 VDD
port 41 nsew
rlabel metal1 s 1915 -35394 1961 -35194 8 VDD
port 41 nsew
rlabel metal1 s 1719 -35394 1765 -35194 8 VDD
port 41 nsew
rlabel metal1 s 1523 -35394 1569 -35194 8 VDD
port 41 nsew
rlabel metal1 s 34 -35394 80 -35194 8 VDD
port 41 nsew
rlabel metal1 s -162 -35394 -116 -35194 2 VDD
port 41 nsew
rlabel metal1 s -275 -35394 -229 -35194 2 VDD
port 41 nsew
rlabel metal1 s -471 -35394 -425 -35194 2 VDD
port 41 nsew
rlabel metal1 s -585 -35394 -539 -35194 2 VDD
port 41 nsew
rlabel metal1 s -781 -35394 -735 -35194 2 VDD
port 41 nsew
rlabel metal1 s -977 -35394 -931 -35194 2 VDD
port 41 nsew
rlabel metal1 s -2466 -35394 -2420 -35194 2 VDD
port 41 nsew
rlabel metal1 s -2662 -35394 -2616 -35194 2 VDD
port 41 nsew
rlabel metal1 s -2775 -35394 -2729 -35194 2 VDD
port 41 nsew
rlabel metal1 s -2971 -35394 -2925 -35194 2 VDD
port 41 nsew
rlabel metal1 s -3085 -35394 -3039 -35194 2 VDD
port 41 nsew
rlabel metal1 s -3281 -35394 -3235 -35194 2 VDD
port 41 nsew
rlabel metal1 s -3477 -35394 -3431 -35194 2 VDD
port 41 nsew
rlabel metal1 s -4966 -35394 -4920 -35194 2 VDD
port 41 nsew
rlabel metal1 s -5162 -35394 -5116 -35194 2 VDD
port 41 nsew
rlabel metal1 s -5275 -35394 -5229 -35194 2 VDD
port 41 nsew
rlabel metal1 s -5471 -35394 -5425 -35194 2 VDD
port 41 nsew
rlabel metal1 s -5585 -35394 -5539 -35194 2 VDD
port 41 nsew
rlabel metal1 s -5781 -35394 -5735 -35194 2 VDD
port 41 nsew
rlabel metal1 s -5977 -35394 -5931 -35194 2 VDD
port 41 nsew
rlabel metal1 s -7466 -35598 -7420 -34998 2 VDD
port 41 nsew
rlabel metal1 s -7662 -35598 -7616 -34998 2 VDD
port 41 nsew
rlabel metal1 s -8085 -35598 -8039 -34998 2 VDD
port 41 nsew
rlabel metal1 s -26012 -35593 -25612 -35547 2 VDD
port 41 nsew
rlabel metal1 s -26012 -35357 -25612 -35311 2 VDD
port 41 nsew
rlabel metal1 s -10518 -35188 -10472 -34988 2 VDD
port 41 nsew
rlabel metal1 s -10714 -35188 -10668 -34988 2 VDD
port 41 nsew
rlabel metal1 s -10910 -35188 -10864 -34988 2 VDD
port 41 nsew
rlabel metal1 s -11355 -35188 -11309 -34988 2 VDD
port 41 nsew
rlabel metal1 s -11551 -35188 -11505 -34988 2 VDD
port 41 nsew
rlabel metal1 s -11747 -35188 -11701 -34988 2 VDD
port 41 nsew
rlabel metal1 s -13218 -35188 -13172 -34988 2 VDD
port 41 nsew
rlabel metal1 s -13414 -35188 -13368 -34988 2 VDD
port 41 nsew
rlabel metal1 s -13610 -35188 -13564 -34988 2 VDD
port 41 nsew
rlabel metal1 s -14055 -35188 -14009 -34988 2 VDD
port 41 nsew
rlabel metal1 s -14251 -35188 -14205 -34988 2 VDD
port 41 nsew
rlabel metal1 s -14447 -35188 -14401 -34988 2 VDD
port 41 nsew
rlabel metal1 s -26012 -35121 -25612 -35075 2 VDD
port 41 nsew
rlabel metal1 s -26012 -34885 -25612 -34839 2 VDD
port 41 nsew
rlabel metal1 s -26012 -34649 -25612 -34603 2 VDD
port 41 nsew
rlabel metal1 s -26012 -34413 -25612 -34367 2 VDD
port 41 nsew
rlabel metal1 s -26012 -34177 -25612 -34131 2 VDD
port 41 nsew
rlabel metal1 s 16381 -27178 16427 -26978 8 VDD
port 41 nsew
rlabel metal1 s 16185 -27178 16231 -26978 8 VDD
port 41 nsew
rlabel metal1 s 15989 -27178 16035 -26978 8 VDD
port 41 nsew
rlabel metal1 s 15544 -27178 15590 -26978 8 VDD
port 41 nsew
rlabel metal1 s 15348 -27178 15394 -26978 8 VDD
port 41 nsew
rlabel metal1 s 15152 -27178 15198 -26978 8 VDD
port 41 nsew
rlabel metal1 s 13681 -27178 13727 -26978 8 VDD
port 41 nsew
rlabel metal1 s 13485 -27178 13531 -26978 8 VDD
port 41 nsew
rlabel metal1 s 13289 -27178 13335 -26978 8 VDD
port 41 nsew
rlabel metal1 s 12844 -27178 12890 -26978 8 VDD
port 41 nsew
rlabel metal1 s 12648 -27178 12694 -26978 8 VDD
port 41 nsew
rlabel metal1 s 12452 -27178 12498 -26978 8 VDD
port 41 nsew
rlabel metal1 s 7336 -27341 7382 -27141 8 VDD
port 41 nsew
rlabel metal1 s 7140 -27341 7186 -27141 8 VDD
port 41 nsew
rlabel metal1 s 7027 -27341 7073 -27141 8 VDD
port 41 nsew
rlabel metal1 s 6831 -27341 6877 -27141 8 VDD
port 41 nsew
rlabel metal1 s 6717 -27341 6763 -27141 8 VDD
port 41 nsew
rlabel metal1 s 6521 -27341 6567 -27141 8 VDD
port 41 nsew
rlabel metal1 s 6325 -27341 6371 -27141 8 VDD
port 41 nsew
rlabel metal1 s 4336 -27341 4382 -27141 8 VDD
port 41 nsew
rlabel metal1 s 4140 -27341 4186 -27141 8 VDD
port 41 nsew
rlabel metal1 s 4027 -27341 4073 -27141 8 VDD
port 41 nsew
rlabel metal1 s 3831 -27341 3877 -27141 8 VDD
port 41 nsew
rlabel metal1 s 3717 -27341 3763 -27141 8 VDD
port 41 nsew
rlabel metal1 s 3521 -27341 3567 -27141 8 VDD
port 41 nsew
rlabel metal1 s 3325 -27341 3371 -27141 8 VDD
port 41 nsew
rlabel metal1 s 1836 -27341 1882 -27141 8 VDD
port 41 nsew
rlabel metal1 s 1640 -27341 1686 -27141 8 VDD
port 41 nsew
rlabel metal1 s 1527 -27341 1573 -27141 8 VDD
port 41 nsew
rlabel metal1 s 1331 -27341 1377 -27141 8 VDD
port 41 nsew
rlabel metal1 s 1217 -27341 1263 -27141 8 VDD
port 41 nsew
rlabel metal1 s 1021 -27341 1067 -27141 8 VDD
port 41 nsew
rlabel metal1 s 825 -27341 871 -27141 8 VDD
port 41 nsew
rlabel metal1 s -664 -27341 -618 -27141 2 VDD
port 41 nsew
rlabel metal1 s -860 -27341 -814 -27141 2 VDD
port 41 nsew
rlabel metal1 s -973 -27341 -927 -27141 2 VDD
port 41 nsew
rlabel metal1 s -1169 -27341 -1123 -27141 2 VDD
port 41 nsew
rlabel metal1 s -1283 -27341 -1237 -27141 2 VDD
port 41 nsew
rlabel metal1 s -1479 -27341 -1433 -27141 2 VDD
port 41 nsew
rlabel metal1 s -1675 -27341 -1629 -27141 2 VDD
port 41 nsew
rlabel metal1 s -3164 -27341 -3118 -27141 2 VDD
port 41 nsew
rlabel metal1 s -3360 -27341 -3314 -27141 2 VDD
port 41 nsew
rlabel metal1 s -3473 -27341 -3427 -27141 2 VDD
port 41 nsew
rlabel metal1 s -3669 -27341 -3623 -27141 2 VDD
port 41 nsew
rlabel metal1 s -3783 -27341 -3737 -27141 2 VDD
port 41 nsew
rlabel metal1 s -3979 -27341 -3933 -27141 2 VDD
port 41 nsew
rlabel metal1 s -4175 -27341 -4129 -27141 2 VDD
port 41 nsew
rlabel metal1 s -5664 -27341 -5618 -27141 2 VDD
port 41 nsew
rlabel metal1 s -5860 -27341 -5814 -27141 2 VDD
port 41 nsew
rlabel metal1 s -5973 -27341 -5927 -27141 2 VDD
port 41 nsew
rlabel metal1 s -6169 -27341 -6123 -27141 2 VDD
port 41 nsew
rlabel metal1 s -6283 -27341 -6237 -27141 2 VDD
port 41 nsew
rlabel metal1 s -6479 -27341 -6433 -27141 2 VDD
port 41 nsew
rlabel metal1 s -6675 -27341 -6629 -27141 2 VDD
port 41 nsew
rlabel metal1 s -20349 -27591 -20173 -26960 2 VDD
port 41 nsew
rlabel metal1 s -21633 -27427 -21587 -27227 2 VDD
port 41 nsew
rlabel metal1 s -21829 -27427 -21783 -27227 2 VDD
port 41 nsew
rlabel metal1 s -22025 -27427 -21979 -27227 2 VDD
port 41 nsew
rlabel metal1 s -22221 -27427 -22175 -27227 2 VDD
port 41 nsew
rlabel metal1 s -22763 -27427 -22717 -27227 2 VDD
port 41 nsew
rlabel metal1 s -22959 -27427 -22913 -27227 2 VDD
port 41 nsew
rlabel metal1 s -297 -26684 -174 -26548 2 VDD
port 41 nsew
rlabel metal1 s -2780 -26684 -2657 -26548 2 VDD
port 41 nsew
rlabel metal1 s -5347 -26719 -5224 -26583 2 VDD
port 41 nsew
rlabel metal1 s -293 -26548 -179 -26131 2 VDD
port 41 nsew
rlabel metal1 s -298 -26131 -175 -26130 2 VDD
port 41 nsew
rlabel metal1 s -298 -26130 8 -26068 2 VDD
port 41 nsew
rlabel metal1 s -2776 -26548 -2662 -26096 2 VDD
port 41 nsew
rlabel metal1 s -2781 -26096 -2658 -25960 2 VDD
port 41 nsew
rlabel metal1 s -5343 -26583 -5229 -25952 2 VDD
port 41 nsew
rlabel metal1 s -16913 -26267 -16867 -26167 2 VDD
port 41 nsew
rlabel metal1 s -17109 -26267 -17063 -26167 2 VDD
port 41 nsew
rlabel metal1 s -17305 -26267 -17259 -26167 2 VDD
port 41 nsew
rlabel metal1 s -17501 -26267 -17455 -26167 2 VDD
port 41 nsew
rlabel metal1 s -17718 -26468 -17672 -26168 2 VDD
port 41 nsew
rlabel metal1 s -17914 -26468 -17868 -26168 2 VDD
port 41 nsew
rlabel metal1 s -18110 -26468 -18064 -26168 2 VDD
port 41 nsew
rlabel metal1 s -18495 -26497 -18449 -26297 2 VDD
port 41 nsew
rlabel metal1 s -18691 -26497 -18645 -26297 2 VDD
port 41 nsew
rlabel metal1 s -18887 -26497 -18841 -26297 2 VDD
port 41 nsew
rlabel metal1 s -19083 -26497 -19037 -26297 2 VDD
port 41 nsew
rlabel metal1 s 86424 -25570 86470 -24970 8 VDD
port 41 nsew
rlabel metal1 s 86001 -25570 86047 -24970 8 VDD
port 41 nsew
rlabel metal1 s 85805 -25570 85851 -24970 8 VDD
port 41 nsew
rlabel metal1 s 85555 -25158 85601 -25058 8 VDD
port 41 nsew
rlabel metal1 s 85359 -25158 85405 -25058 8 VDD
port 41 nsew
rlabel metal1 s 85163 -25158 85209 -25058 8 VDD
port 41 nsew
rlabel metal1 s 84967 -25158 85013 -25058 8 VDD
port 41 nsew
rlabel metal1 s 84750 -25359 84796 -25059 8 VDD
port 41 nsew
rlabel metal1 s 84554 -25359 84600 -25059 8 VDD
port 41 nsew
rlabel metal1 s 84358 -25359 84404 -25059 8 VDD
port 41 nsew
rlabel metal1 s 82756 -25539 82802 -24939 8 VDD
port 41 nsew
rlabel metal1 s 82333 -25539 82379 -24939 8 VDD
port 41 nsew
rlabel metal1 s 82137 -25539 82183 -24939 8 VDD
port 41 nsew
rlabel metal1 s 81887 -25127 81933 -25027 8 VDD
port 41 nsew
rlabel metal1 s 81691 -25127 81737 -25027 8 VDD
port 41 nsew
rlabel metal1 s 81495 -25127 81541 -25027 8 VDD
port 41 nsew
rlabel metal1 s 81299 -25127 81345 -25027 8 VDD
port 41 nsew
rlabel metal1 s 81082 -25328 81128 -25028 8 VDD
port 41 nsew
rlabel metal1 s 80886 -25328 80932 -25028 8 VDD
port 41 nsew
rlabel metal1 s 80690 -25328 80736 -25028 8 VDD
port 41 nsew
rlabel metal1 s 77060 -25608 77106 -25008 8 VDD
port 41 nsew
rlabel metal1 s 76637 -25608 76683 -25008 8 VDD
port 41 nsew
rlabel metal1 s 76441 -25608 76487 -25008 8 VDD
port 41 nsew
rlabel metal1 s 76191 -25196 76237 -25096 8 VDD
port 41 nsew
rlabel metal1 s 75995 -25196 76041 -25096 8 VDD
port 41 nsew
rlabel metal1 s 75799 -25196 75845 -25096 8 VDD
port 41 nsew
rlabel metal1 s 75603 -25196 75649 -25096 8 VDD
port 41 nsew
rlabel metal1 s 75386 -25397 75432 -25097 8 VDD
port 41 nsew
rlabel metal1 s 75190 -25397 75236 -25097 8 VDD
port 41 nsew
rlabel metal1 s 74994 -25397 75040 -25097 8 VDD
port 41 nsew
rlabel metal1 s 73392 -25577 73438 -24977 8 VDD
port 41 nsew
rlabel metal1 s 72969 -25577 73015 -24977 8 VDD
port 41 nsew
rlabel metal1 s 72773 -25577 72819 -24977 8 VDD
port 41 nsew
rlabel metal1 s 72523 -25165 72569 -25065 8 VDD
port 41 nsew
rlabel metal1 s 72327 -25165 72373 -25065 8 VDD
port 41 nsew
rlabel metal1 s 72131 -25165 72177 -25065 8 VDD
port 41 nsew
rlabel metal1 s 71935 -25165 71981 -25065 8 VDD
port 41 nsew
rlabel metal1 s 71718 -25366 71764 -25066 8 VDD
port 41 nsew
rlabel metal1 s 71522 -25366 71568 -25066 8 VDD
port 41 nsew
rlabel metal1 s 71326 -25366 71372 -25066 8 VDD
port 41 nsew
rlabel metal1 s 67907 -25625 67953 -25025 8 VDD
port 41 nsew
rlabel metal1 s 67484 -25625 67530 -25025 8 VDD
port 41 nsew
rlabel metal1 s 67288 -25625 67334 -25025 8 VDD
port 41 nsew
rlabel metal1 s 67038 -25213 67084 -25113 8 VDD
port 41 nsew
rlabel metal1 s 66842 -25213 66888 -25113 8 VDD
port 41 nsew
rlabel metal1 s 66646 -25213 66692 -25113 8 VDD
port 41 nsew
rlabel metal1 s 66450 -25213 66496 -25113 8 VDD
port 41 nsew
rlabel metal1 s 66233 -25414 66279 -25114 8 VDD
port 41 nsew
rlabel metal1 s 66037 -25414 66083 -25114 8 VDD
port 41 nsew
rlabel metal1 s 65841 -25414 65887 -25114 8 VDD
port 41 nsew
rlabel metal1 s 64239 -25594 64285 -24994 8 VDD
port 41 nsew
rlabel metal1 s 63816 -25594 63862 -24994 8 VDD
port 41 nsew
rlabel metal1 s 63620 -25594 63666 -24994 8 VDD
port 41 nsew
rlabel metal1 s 63370 -25182 63416 -25082 8 VDD
port 41 nsew
rlabel metal1 s 63174 -25182 63220 -25082 8 VDD
port 41 nsew
rlabel metal1 s 62978 -25182 63024 -25082 8 VDD
port 41 nsew
rlabel metal1 s 62782 -25182 62828 -25082 8 VDD
port 41 nsew
rlabel metal1 s 62565 -25383 62611 -25083 8 VDD
port 41 nsew
rlabel metal1 s 62369 -25383 62415 -25083 8 VDD
port 41 nsew
rlabel metal1 s 62173 -25383 62219 -25083 8 VDD
port 41 nsew
rlabel metal1 s 59153 -25691 59199 -25091 8 VDD
port 41 nsew
rlabel metal1 s 58730 -25691 58776 -25091 8 VDD
port 41 nsew
rlabel metal1 s 58534 -25691 58580 -25091 8 VDD
port 41 nsew
rlabel metal1 s 58284 -25279 58330 -25179 8 VDD
port 41 nsew
rlabel metal1 s 58088 -25279 58134 -25179 8 VDD
port 41 nsew
rlabel metal1 s 57892 -25279 57938 -25179 8 VDD
port 41 nsew
rlabel metal1 s 57696 -25279 57742 -25179 8 VDD
port 41 nsew
rlabel metal1 s 57479 -25480 57525 -25180 8 VDD
port 41 nsew
rlabel metal1 s 57283 -25480 57329 -25180 8 VDD
port 41 nsew
rlabel metal1 s 57087 -25480 57133 -25180 8 VDD
port 41 nsew
rlabel metal1 s 55485 -25660 55531 -25060 8 VDD
port 41 nsew
rlabel metal1 s 55062 -25660 55108 -25060 8 VDD
port 41 nsew
rlabel metal1 s 54866 -25660 54912 -25060 8 VDD
port 41 nsew
rlabel metal1 s 54616 -25248 54662 -25148 8 VDD
port 41 nsew
rlabel metal1 s 54420 -25248 54466 -25148 8 VDD
port 41 nsew
rlabel metal1 s 54224 -25248 54270 -25148 8 VDD
port 41 nsew
rlabel metal1 s 54028 -25248 54074 -25148 8 VDD
port 41 nsew
rlabel metal1 s 53811 -25449 53857 -25149 8 VDD
port 41 nsew
rlabel metal1 s 53615 -25449 53661 -25149 8 VDD
port 41 nsew
rlabel metal1 s 53419 -25449 53465 -25149 8 VDD
port 41 nsew
rlabel metal1 s 49955 -25725 50001 -25125 8 VDD
port 41 nsew
rlabel metal1 s 49532 -25725 49578 -25125 8 VDD
port 41 nsew
rlabel metal1 s 49336 -25725 49382 -25125 8 VDD
port 41 nsew
rlabel metal1 s 49086 -25313 49132 -25213 8 VDD
port 41 nsew
rlabel metal1 s 48890 -25313 48936 -25213 8 VDD
port 41 nsew
rlabel metal1 s 48694 -25313 48740 -25213 8 VDD
port 41 nsew
rlabel metal1 s 48498 -25313 48544 -25213 8 VDD
port 41 nsew
rlabel metal1 s 48281 -25514 48327 -25214 8 VDD
port 41 nsew
rlabel metal1 s 48085 -25514 48131 -25214 8 VDD
port 41 nsew
rlabel metal1 s 47889 -25514 47935 -25214 8 VDD
port 41 nsew
rlabel metal1 s 46287 -25694 46333 -25094 8 VDD
port 41 nsew
rlabel metal1 s 45864 -25694 45910 -25094 8 VDD
port 41 nsew
rlabel metal1 s 45668 -25694 45714 -25094 8 VDD
port 41 nsew
rlabel metal1 s 45418 -25282 45464 -25182 8 VDD
port 41 nsew
rlabel metal1 s 45222 -25282 45268 -25182 8 VDD
port 41 nsew
rlabel metal1 s 45026 -25282 45072 -25182 8 VDD
port 41 nsew
rlabel metal1 s 44830 -25282 44876 -25182 8 VDD
port 41 nsew
rlabel metal1 s 44613 -25483 44659 -25183 8 VDD
port 41 nsew
rlabel metal1 s 44417 -25483 44463 -25183 8 VDD
port 41 nsew
rlabel metal1 s 44221 -25483 44267 -25183 8 VDD
port 41 nsew
rlabel metal1 s 41092 -25686 41138 -25086 8 VDD
port 41 nsew
rlabel metal1 s 40669 -25686 40715 -25086 8 VDD
port 41 nsew
rlabel metal1 s 40473 -25686 40519 -25086 8 VDD
port 41 nsew
rlabel metal1 s 40223 -25274 40269 -25174 8 VDD
port 41 nsew
rlabel metal1 s 40027 -25274 40073 -25174 8 VDD
port 41 nsew
rlabel metal1 s 39831 -25274 39877 -25174 8 VDD
port 41 nsew
rlabel metal1 s 39635 -25274 39681 -25174 8 VDD
port 41 nsew
rlabel metal1 s 39418 -25475 39464 -25175 8 VDD
port 41 nsew
rlabel metal1 s 39222 -25475 39268 -25175 8 VDD
port 41 nsew
rlabel metal1 s 39026 -25475 39072 -25175 8 VDD
port 41 nsew
rlabel metal1 s 37424 -25655 37470 -25055 8 VDD
port 41 nsew
rlabel metal1 s 37001 -25655 37047 -25055 8 VDD
port 41 nsew
rlabel metal1 s 36805 -25655 36851 -25055 8 VDD
port 41 nsew
rlabel metal1 s 36555 -25243 36601 -25143 8 VDD
port 41 nsew
rlabel metal1 s 36359 -25243 36405 -25143 8 VDD
port 41 nsew
rlabel metal1 s 36163 -25243 36209 -25143 8 VDD
port 41 nsew
rlabel metal1 s 35967 -25243 36013 -25143 8 VDD
port 41 nsew
rlabel metal1 s 35750 -25444 35796 -25144 8 VDD
port 41 nsew
rlabel metal1 s 35554 -25444 35600 -25144 8 VDD
port 41 nsew
rlabel metal1 s 35358 -25444 35404 -25144 8 VDD
port 41 nsew
rlabel metal1 s 32652 -25675 32698 -25075 8 VDD
port 41 nsew
rlabel metal1 s 32229 -25675 32275 -25075 8 VDD
port 41 nsew
rlabel metal1 s 32033 -25675 32079 -25075 8 VDD
port 41 nsew
rlabel metal1 s 16283 -25860 16329 -25660 8 VDD
port 41 nsew
rlabel metal1 s 16087 -25860 16133 -25660 8 VDD
port 41 nsew
rlabel metal1 s 15891 -25860 15937 -25660 8 VDD
port 41 nsew
rlabel metal1 s 14540 -25860 14586 -25660 8 VDD
port 41 nsew
rlabel metal1 s 14344 -25860 14390 -25660 8 VDD
port 41 nsew
rlabel metal1 s 14148 -25860 14194 -25660 8 VDD
port 41 nsew
rlabel metal1 s 13583 -25860 13629 -25660 8 VDD
port 41 nsew
rlabel metal1 s 13387 -25860 13433 -25660 8 VDD
port 41 nsew
rlabel metal1 s 13191 -25860 13237 -25660 8 VDD
port 41 nsew
rlabel metal1 s 11840 -25860 11886 -25660 8 VDD
port 41 nsew
rlabel metal1 s 11644 -25860 11690 -25660 8 VDD
port 41 nsew
rlabel metal1 s 11448 -25860 11494 -25660 8 VDD
port 41 nsew
rlabel metal1 s 10958 -25860 11004 -25660 8 VDD
port 41 nsew
rlabel metal1 s 10762 -25860 10808 -25660 8 VDD
port 41 nsew
rlabel metal1 s 10566 -25860 10612 -25660 8 VDD
port 41 nsew
rlabel metal1 s -5348 -25952 -5225 -25816 2 VDD
port 41 nsew
rlabel metal1 s -19544 -25965 -19352 -25793 2 VDD
port 41 nsew
rlabel metal1 s 31783 -25263 31829 -25163 8 VDD
port 41 nsew
rlabel metal1 s 31587 -25263 31633 -25163 8 VDD
port 41 nsew
rlabel metal1 s 31391 -25263 31437 -25163 8 VDD
port 41 nsew
rlabel metal1 s 31195 -25263 31241 -25163 8 VDD
port 41 nsew
rlabel metal1 s 30978 -25464 31024 -25164 8 VDD
port 41 nsew
rlabel metal1 s 30782 -25464 30828 -25164 8 VDD
port 41 nsew
rlabel metal1 s 30586 -25464 30632 -25164 8 VDD
port 41 nsew
rlabel metal1 s 28984 -25644 29030 -25044 8 VDD
port 41 nsew
rlabel metal1 s 28561 -25644 28607 -25044 8 VDD
port 41 nsew
rlabel metal1 s 28365 -25644 28411 -25044 8 VDD
port 41 nsew
rlabel metal1 s 28115 -25232 28161 -25132 8 VDD
port 41 nsew
rlabel metal1 s 27919 -25232 27965 -25132 8 VDD
port 41 nsew
rlabel metal1 s 27723 -25232 27769 -25132 8 VDD
port 41 nsew
rlabel metal1 s 27527 -25232 27573 -25132 8 VDD
port 41 nsew
rlabel metal1 s 27310 -25433 27356 -25133 8 VDD
port 41 nsew
rlabel metal1 s 27114 -25433 27160 -25133 8 VDD
port 41 nsew
rlabel metal1 s 26918 -25433 26964 -25133 8 VDD
port 41 nsew
rlabel metal1 s 6340 -25294 6463 -25282 8 VDD
port 41 nsew
rlabel metal1 s 5124 -25295 5247 -25282 8 VDD
port 41 nsew
rlabel metal1 s 5124 -25282 6463 -25177 8 VDD
port 41 nsew
rlabel metal1 s 6340 -25177 6463 -25158 8 VDD
port 41 nsew
rlabel metal1 s 5124 -25177 5247 -25159 8 VDD
port 41 nsew
rlabel metal1 s 3768 -25300 3891 -25289 8 VDD
port 41 nsew
rlabel metal1 s 3367 -25298 3490 -25289 8 VDD
port 41 nsew
rlabel metal1 s 3367 -25289 3891 -25182 8 VDD
port 41 nsew
rlabel metal1 s 3768 -25182 3891 -25164 8 VDD
port 41 nsew
rlabel metal1 s 3367 -25182 3490 -25162 8 VDD
port 41 nsew
rlabel metal1 s 2139 -25275 2262 -25259 8 VDD
port 41 nsew
rlabel metal1 s -1228 -25287 -1105 -25274 2 VDD
port 41 nsew
rlabel metal1 s -1522 -25286 -1399 -25274 2 VDD
port 41 nsew
rlabel metal1 s 1750 -25274 1873 -25259 8 VDD
port 41 nsew
rlabel metal1 s 1750 -25259 2262 -25152 8 VDD
port 41 nsew
rlabel metal1 s 2139 -25152 2262 -25139 8 VDD
port 41 nsew
rlabel metal1 s 1750 -25152 1873 -25138 8 VDD
port 41 nsew
rlabel metal1 s -1522 -25274 -1105 -25159 2 VDD
port 41 nsew
rlabel metal1 s -1228 -25159 -1105 -25151 2 VDD
port 41 nsew
rlabel metal1 s -1522 -25159 -1399 -25150 2 VDD
port 41 nsew
rlabel metal1 s 50395 -25044 50546 -25019 8 VDD
port 41 nsew
rlabel metal1 s 50145 -25031 50236 -25019 8 VDD
port 41 nsew
rlabel metal1 s 59593 -25010 59744 -24985 8 VDD
port 41 nsew
rlabel metal1 s 59343 -24997 59434 -24985 8 VDD
port 41 nsew
rlabel metal1 s 77500 -24927 77651 -24902 8 VDD
port 41 nsew
rlabel metal1 s 68347 -24944 68498 -24919 8 VDD
port 41 nsew
rlabel metal1 s 68097 -24931 68188 -24919 8 VDD
port 41 nsew
rlabel metal1 s 77250 -24914 77341 -24902 8 VDD
port 41 nsew
rlabel metal1 s 86864 -24889 87015 -24864 8 VDD
port 41 nsew
rlabel metal1 s 86614 -24876 86705 -24864 8 VDD
port 41 nsew
rlabel metal1 s 86614 -24864 87015 -24725 8 VDD
port 41 nsew
rlabel metal1 s 86864 -24725 87015 -24698 8 VDD
port 41 nsew
rlabel metal1 s 86614 -24725 86705 -24713 8 VDD
port 41 nsew
rlabel metal1 s 83194 -24811 83290 -24785 8 VDD
port 41 nsew
rlabel metal1 s 81891 -24792 82074 -24785 8 VDD
port 41 nsew
rlabel metal1 s 81891 -24785 83290 -24703 8 VDD
port 41 nsew
rlabel metal1 s 77250 -24902 77651 -24763 8 VDD
port 41 nsew
rlabel metal1 s 77500 -24763 77651 -24736 8 VDD
port 41 nsew
rlabel metal1 s 77250 -24763 77341 -24751 8 VDD
port 41 nsew
rlabel metal1 s 73830 -24849 73926 -24823 8 VDD
port 41 nsew
rlabel metal1 s 72527 -24830 72710 -24823 8 VDD
port 41 nsew
rlabel metal1 s 72527 -24823 73926 -24741 8 VDD
port 41 nsew
rlabel metal1 s 68097 -24919 68498 -24780 8 VDD
port 41 nsew
rlabel metal1 s 68347 -24780 68498 -24753 8 VDD
port 41 nsew
rlabel metal1 s 68097 -24780 68188 -24768 8 VDD
port 41 nsew
rlabel metal1 s 64677 -24866 64773 -24840 8 VDD
port 41 nsew
rlabel metal1 s 63374 -24847 63557 -24840 8 VDD
port 41 nsew
rlabel metal1 s 63374 -24840 64773 -24758 8 VDD
port 41 nsew
rlabel metal1 s 59343 -24985 59744 -24846 8 VDD
port 41 nsew
rlabel metal1 s 59593 -24846 59744 -24819 8 VDD
port 41 nsew
rlabel metal1 s 59343 -24846 59434 -24834 8 VDD
port 41 nsew
rlabel metal1 s 55923 -24932 56019 -24906 8 VDD
port 41 nsew
rlabel metal1 s 54620 -24913 54803 -24906 8 VDD
port 41 nsew
rlabel metal1 s 54620 -24906 56019 -24824 8 VDD
port 41 nsew
rlabel metal1 s 50145 -25019 50546 -24880 8 VDD
port 41 nsew
rlabel metal1 s 41532 -25005 41683 -24980 8 VDD
port 41 nsew
rlabel metal1 s 41282 -24992 41373 -24980 8 VDD
port 41 nsew
rlabel metal1 s 50395 -24880 50546 -24853 8 VDD
port 41 nsew
rlabel metal1 s 50145 -24880 50236 -24868 8 VDD
port 41 nsew
rlabel metal1 s 46725 -24966 46821 -24940 8 VDD
port 41 nsew
rlabel metal1 s 45422 -24947 45605 -24940 8 VDD
port 41 nsew
rlabel metal1 s 45422 -24940 46821 -24858 8 VDD
port 41 nsew
rlabel metal1 s 46725 -24858 46821 -24829 8 VDD
port 41 nsew
rlabel metal1 s 55923 -24824 56019 -24795 8 VDD
port 41 nsew
rlabel metal1 s 54620 -24824 54803 -24783 8 VDD
port 41 nsew
rlabel metal1 s 45422 -24858 45605 -24817 8 VDD
port 41 nsew
rlabel metal1 s 41282 -24980 41683 -24841 8 VDD
port 41 nsew
rlabel metal1 s 33092 -24994 33243 -24969 8 VDD
port 41 nsew
rlabel metal1 s 32842 -24981 32933 -24969 8 VDD
port 41 nsew
rlabel metal1 s 41532 -24841 41683 -24814 8 VDD
port 41 nsew
rlabel metal1 s 41282 -24841 41373 -24829 8 VDD
port 41 nsew
rlabel metal1 s 37862 -24927 37958 -24901 8 VDD
port 41 nsew
rlabel metal1 s 36559 -24908 36742 -24901 8 VDD
port 41 nsew
rlabel metal1 s 36559 -24901 37958 -24819 8 VDD
port 41 nsew
rlabel metal1 s 37862 -24819 37958 -24790 8 VDD
port 41 nsew
rlabel metal1 s 36559 -24819 36742 -24778 8 VDD
port 41 nsew
rlabel metal1 s 32842 -24969 33243 -24830 8 VDD
port 41 nsew
rlabel metal1 s 33092 -24830 33243 -24803 8 VDD
port 41 nsew
rlabel metal1 s 32842 -24830 32933 -24818 8 VDD
port 41 nsew
rlabel metal1 s 29422 -24916 29518 -24890 8 VDD
port 41 nsew
rlabel metal1 s 28119 -24897 28302 -24890 8 VDD
port 41 nsew
rlabel metal1 s 7346 -25090 7392 -24890 8 VDD
port 41 nsew
rlabel metal1 s 7150 -25090 7196 -24890 8 VDD
port 41 nsew
rlabel metal1 s 7037 -25090 7083 -24890 8 VDD
port 41 nsew
rlabel metal1 s 6841 -25090 6887 -24890 8 VDD
port 41 nsew
rlabel metal1 s 6727 -25090 6773 -24890 8 VDD
port 41 nsew
rlabel metal1 s 6531 -25090 6577 -24890 8 VDD
port 41 nsew
rlabel metal1 s 6335 -25090 6381 -24890 8 VDD
port 41 nsew
rlabel metal1 s 5174 -25101 5220 -24901 8 VDD
port 41 nsew
rlabel metal1 s 4978 -25101 5024 -24901 8 VDD
port 41 nsew
rlabel metal1 s 4782 -25101 4828 -24901 8 VDD
port 41 nsew
rlabel metal1 s 4586 -25101 4632 -24901 8 VDD
port 41 nsew
rlabel metal1 s 4044 -25101 4090 -24901 8 VDD
port 41 nsew
rlabel metal1 s 3848 -25101 3894 -24901 8 VDD
port 41 nsew
rlabel metal1 s 28119 -24890 29518 -24808 8 VDD
port 41 nsew
rlabel metal1 s 29422 -24808 29518 -24779 8 VDD
port 41 nsew
rlabel metal1 s 28119 -24808 28302 -24767 8 VDD
port 41 nsew
rlabel metal1 s 73830 -24741 73926 -24712 8 VDD
port 41 nsew
rlabel metal1 s 83194 -24703 83290 -24674 8 VDD
port 41 nsew
rlabel metal1 s 81891 -24703 82074 -24662 8 VDD
port 41 nsew
rlabel metal1 s 72527 -24741 72710 -24700 8 VDD
port 41 nsew
rlabel metal1 s 64677 -24758 64773 -24729 8 VDD
port 41 nsew
rlabel metal1 s 63374 -24758 63557 -24717 8 VDD
port 41 nsew
rlabel metal1 s 86554 -24460 86600 -24360 8 VDD
port 41 nsew
rlabel metal1 s 86358 -24460 86404 -24360 8 VDD
port 41 nsew
rlabel metal1 s 86162 -24460 86208 -24360 8 VDD
port 41 nsew
rlabel metal1 s 85966 -24460 86012 -24360 8 VDD
port 41 nsew
rlabel metal1 s 85749 -24459 85795 -24159 8 VDD
port 41 nsew
rlabel metal1 s 85553 -24459 85599 -24159 8 VDD
port 41 nsew
rlabel metal1 s 85357 -24459 85403 -24159 8 VDD
port 41 nsew
rlabel metal1 s 84972 -24330 85018 -24130 8 VDD
port 41 nsew
rlabel metal1 s 84776 -24330 84822 -24130 8 VDD
port 41 nsew
rlabel metal1 s 84580 -24330 84626 -24130 8 VDD
port 41 nsew
rlabel metal1 s 84384 -24330 84430 -24130 8 VDD
port 41 nsew
rlabel metal1 s 82886 -24429 82932 -24329 8 VDD
port 41 nsew
rlabel metal1 s 82690 -24429 82736 -24329 8 VDD
port 41 nsew
rlabel metal1 s 82494 -24429 82540 -24329 8 VDD
port 41 nsew
rlabel metal1 s 82298 -24429 82344 -24329 8 VDD
port 41 nsew
rlabel metal1 s 82081 -24428 82127 -24128 8 VDD
port 41 nsew
rlabel metal1 s 81885 -24428 81931 -24128 8 VDD
port 41 nsew
rlabel metal1 s 81689 -24428 81735 -24128 8 VDD
port 41 nsew
rlabel metal1 s 77190 -24498 77236 -24398 8 VDD
port 41 nsew
rlabel metal1 s 76994 -24498 77040 -24398 8 VDD
port 41 nsew
rlabel metal1 s 76798 -24498 76844 -24398 8 VDD
port 41 nsew
rlabel metal1 s 76602 -24498 76648 -24398 8 VDD
port 41 nsew
rlabel metal1 s 81304 -24299 81350 -24099 8 VDD
port 41 nsew
rlabel metal1 s 81108 -24299 81154 -24099 8 VDD
port 41 nsew
rlabel metal1 s 80912 -24299 80958 -24099 8 VDD
port 41 nsew
rlabel metal1 s 80716 -24299 80762 -24099 8 VDD
port 41 nsew
rlabel metal1 s 76385 -24497 76431 -24197 8 VDD
port 41 nsew
rlabel metal1 s 76189 -24497 76235 -24197 8 VDD
port 41 nsew
rlabel metal1 s 75993 -24497 76039 -24197 8 VDD
port 41 nsew
rlabel metal1 s 75608 -24368 75654 -24168 8 VDD
port 41 nsew
rlabel metal1 s 75412 -24368 75458 -24168 8 VDD
port 41 nsew
rlabel metal1 s 75216 -24368 75262 -24168 8 VDD
port 41 nsew
rlabel metal1 s 75020 -24368 75066 -24168 8 VDD
port 41 nsew
rlabel metal1 s 73522 -24467 73568 -24367 8 VDD
port 41 nsew
rlabel metal1 s 73326 -24467 73372 -24367 8 VDD
port 41 nsew
rlabel metal1 s 73130 -24467 73176 -24367 8 VDD
port 41 nsew
rlabel metal1 s 72934 -24467 72980 -24367 8 VDD
port 41 nsew
rlabel metal1 s 72717 -24466 72763 -24166 8 VDD
port 41 nsew
rlabel metal1 s 72521 -24466 72567 -24166 8 VDD
port 41 nsew
rlabel metal1 s 72325 -24466 72371 -24166 8 VDD
port 41 nsew
rlabel metal1 s 68037 -24515 68083 -24415 8 VDD
port 41 nsew
rlabel metal1 s 67841 -24515 67887 -24415 8 VDD
port 41 nsew
rlabel metal1 s 67645 -24515 67691 -24415 8 VDD
port 41 nsew
rlabel metal1 s 67449 -24515 67495 -24415 8 VDD
port 41 nsew
rlabel metal1 s 71940 -24337 71986 -24137 8 VDD
port 41 nsew
rlabel metal1 s 71744 -24337 71790 -24137 8 VDD
port 41 nsew
rlabel metal1 s 71548 -24337 71594 -24137 8 VDD
port 41 nsew
rlabel metal1 s 71352 -24337 71398 -24137 8 VDD
port 41 nsew
rlabel metal1 s 67232 -24514 67278 -24214 8 VDD
port 41 nsew
rlabel metal1 s 67036 -24514 67082 -24214 8 VDD
port 41 nsew
rlabel metal1 s 66840 -24514 66886 -24214 8 VDD
port 41 nsew
rlabel metal1 s 66455 -24385 66501 -24185 8 VDD
port 41 nsew
rlabel metal1 s 66259 -24385 66305 -24185 8 VDD
port 41 nsew
rlabel metal1 s 66063 -24385 66109 -24185 8 VDD
port 41 nsew
rlabel metal1 s 65867 -24385 65913 -24185 8 VDD
port 41 nsew
rlabel metal1 s 64369 -24484 64415 -24384 8 VDD
port 41 nsew
rlabel metal1 s 64173 -24484 64219 -24384 8 VDD
port 41 nsew
rlabel metal1 s 63977 -24484 64023 -24384 8 VDD
port 41 nsew
rlabel metal1 s 63781 -24484 63827 -24384 8 VDD
port 41 nsew
rlabel metal1 s 63564 -24483 63610 -24183 8 VDD
port 41 nsew
rlabel metal1 s 63368 -24483 63414 -24183 8 VDD
port 41 nsew
rlabel metal1 s 63172 -24483 63218 -24183 8 VDD
port 41 nsew
rlabel metal1 s 59283 -24581 59329 -24481 8 VDD
port 41 nsew
rlabel metal1 s 59087 -24581 59133 -24481 8 VDD
port 41 nsew
rlabel metal1 s 58891 -24581 58937 -24481 8 VDD
port 41 nsew
rlabel metal1 s 58695 -24581 58741 -24481 8 VDD
port 41 nsew
rlabel metal1 s 62787 -24354 62833 -24154 8 VDD
port 41 nsew
rlabel metal1 s 62591 -24354 62637 -24154 8 VDD
port 41 nsew
rlabel metal1 s 62395 -24354 62441 -24154 8 VDD
port 41 nsew
rlabel metal1 s 62199 -24354 62245 -24154 8 VDD
port 41 nsew
rlabel metal1 s 58478 -24580 58524 -24280 8 VDD
port 41 nsew
rlabel metal1 s 58282 -24580 58328 -24280 8 VDD
port 41 nsew
rlabel metal1 s 58086 -24580 58132 -24280 8 VDD
port 41 nsew
rlabel metal1 s 57701 -24451 57747 -24251 8 VDD
port 41 nsew
rlabel metal1 s 57505 -24451 57551 -24251 8 VDD
port 41 nsew
rlabel metal1 s 57309 -24451 57355 -24251 8 VDD
port 41 nsew
rlabel metal1 s 57113 -24451 57159 -24251 8 VDD
port 41 nsew
rlabel metal1 s 55615 -24550 55661 -24450 8 VDD
port 41 nsew
rlabel metal1 s 55419 -24550 55465 -24450 8 VDD
port 41 nsew
rlabel metal1 s 55223 -24550 55269 -24450 8 VDD
port 41 nsew
rlabel metal1 s 55027 -24550 55073 -24450 8 VDD
port 41 nsew
rlabel metal1 s 54810 -24549 54856 -24249 8 VDD
port 41 nsew
rlabel metal1 s 54614 -24549 54660 -24249 8 VDD
port 41 nsew
rlabel metal1 s 54418 -24549 54464 -24249 8 VDD
port 41 nsew
rlabel metal1 s 50085 -24615 50131 -24515 8 VDD
port 41 nsew
rlabel metal1 s 49889 -24615 49935 -24515 8 VDD
port 41 nsew
rlabel metal1 s 49693 -24615 49739 -24515 8 VDD
port 41 nsew
rlabel metal1 s 49497 -24615 49543 -24515 8 VDD
port 41 nsew
rlabel metal1 s 54033 -24420 54079 -24220 8 VDD
port 41 nsew
rlabel metal1 s 53837 -24420 53883 -24220 8 VDD
port 41 nsew
rlabel metal1 s 53641 -24420 53687 -24220 8 VDD
port 41 nsew
rlabel metal1 s 53445 -24420 53491 -24220 8 VDD
port 41 nsew
rlabel metal1 s 49280 -24614 49326 -24314 8 VDD
port 41 nsew
rlabel metal1 s 49084 -24614 49130 -24314 8 VDD
port 41 nsew
rlabel metal1 s 48888 -24614 48934 -24314 8 VDD
port 41 nsew
rlabel metal1 s 48503 -24485 48549 -24285 8 VDD
port 41 nsew
rlabel metal1 s 48307 -24485 48353 -24285 8 VDD
port 41 nsew
rlabel metal1 s 48111 -24485 48157 -24285 8 VDD
port 41 nsew
rlabel metal1 s 47915 -24485 47961 -24285 8 VDD
port 41 nsew
rlabel metal1 s 46417 -24584 46463 -24484 8 VDD
port 41 nsew
rlabel metal1 s 46221 -24584 46267 -24484 8 VDD
port 41 nsew
rlabel metal1 s 46025 -24584 46071 -24484 8 VDD
port 41 nsew
rlabel metal1 s 45829 -24584 45875 -24484 8 VDD
port 41 nsew
rlabel metal1 s 45612 -24583 45658 -24283 8 VDD
port 41 nsew
rlabel metal1 s 45416 -24583 45462 -24283 8 VDD
port 41 nsew
rlabel metal1 s 45220 -24583 45266 -24283 8 VDD
port 41 nsew
rlabel metal1 s 41222 -24576 41268 -24476 8 VDD
port 41 nsew
rlabel metal1 s 41026 -24576 41072 -24476 8 VDD
port 41 nsew
rlabel metal1 s 40830 -24576 40876 -24476 8 VDD
port 41 nsew
rlabel metal1 s 40634 -24576 40680 -24476 8 VDD
port 41 nsew
rlabel metal1 s 44835 -24454 44881 -24254 8 VDD
port 41 nsew
rlabel metal1 s 44639 -24454 44685 -24254 8 VDD
port 41 nsew
rlabel metal1 s 44443 -24454 44489 -24254 8 VDD
port 41 nsew
rlabel metal1 s 44247 -24454 44293 -24254 8 VDD
port 41 nsew
rlabel metal1 s 40417 -24575 40463 -24275 8 VDD
port 41 nsew
rlabel metal1 s 40221 -24575 40267 -24275 8 VDD
port 41 nsew
rlabel metal1 s 40025 -24575 40071 -24275 8 VDD
port 41 nsew
rlabel metal1 s 39640 -24446 39686 -24246 8 VDD
port 41 nsew
rlabel metal1 s 39444 -24446 39490 -24246 8 VDD
port 41 nsew
rlabel metal1 s 39248 -24446 39294 -24246 8 VDD
port 41 nsew
rlabel metal1 s 39052 -24446 39098 -24246 8 VDD
port 41 nsew
rlabel metal1 s 37554 -24545 37600 -24445 8 VDD
port 41 nsew
rlabel metal1 s 37358 -24545 37404 -24445 8 VDD
port 41 nsew
rlabel metal1 s 37162 -24545 37208 -24445 8 VDD
port 41 nsew
rlabel metal1 s 36966 -24545 37012 -24445 8 VDD
port 41 nsew
rlabel metal1 s 36749 -24544 36795 -24244 8 VDD
port 41 nsew
rlabel metal1 s 36553 -24544 36599 -24244 8 VDD
port 41 nsew
rlabel metal1 s 36357 -24544 36403 -24244 8 VDD
port 41 nsew
rlabel metal1 s 32782 -24565 32828 -24465 8 VDD
port 41 nsew
rlabel metal1 s 32586 -24565 32632 -24465 8 VDD
port 41 nsew
rlabel metal1 s 32390 -24565 32436 -24465 8 VDD
port 41 nsew
rlabel metal1 s 32194 -24565 32240 -24465 8 VDD
port 41 nsew
rlabel metal1 s 35972 -24415 36018 -24215 8 VDD
port 41 nsew
rlabel metal1 s 35776 -24415 35822 -24215 8 VDD
port 41 nsew
rlabel metal1 s 35580 -24415 35626 -24215 8 VDD
port 41 nsew
rlabel metal1 s 35384 -24415 35430 -24215 8 VDD
port 41 nsew
rlabel metal1 s 31977 -24564 32023 -24264 8 VDD
port 41 nsew
rlabel metal1 s 31781 -24564 31827 -24264 8 VDD
port 41 nsew
rlabel metal1 s 31585 -24564 31631 -24264 8 VDD
port 41 nsew
rlabel metal1 s 31200 -24435 31246 -24235 8 VDD
port 41 nsew
rlabel metal1 s 31004 -24435 31050 -24235 8 VDD
port 41 nsew
rlabel metal1 s 30808 -24435 30854 -24235 8 VDD
port 41 nsew
rlabel metal1 s 30612 -24435 30658 -24235 8 VDD
port 41 nsew
rlabel metal1 s 29114 -24534 29160 -24434 8 VDD
port 41 nsew
rlabel metal1 s 28918 -24534 28964 -24434 8 VDD
port 41 nsew
rlabel metal1 s 28722 -24534 28768 -24434 8 VDD
port 41 nsew
rlabel metal1 s 28526 -24534 28572 -24434 8 VDD
port 41 nsew
rlabel metal1 s 28309 -24533 28355 -24233 8 VDD
port 41 nsew
rlabel metal1 s 28113 -24533 28159 -24233 8 VDD
port 41 nsew
rlabel metal1 s 27917 -24533 27963 -24233 8 VDD
port 41 nsew
rlabel metal1 s 27532 -24404 27578 -24204 8 VDD
port 41 nsew
rlabel metal1 s 27336 -24404 27382 -24204 8 VDD
port 41 nsew
rlabel metal1 s 27140 -24404 27186 -24204 8 VDD
port 41 nsew
rlabel metal1 s 26944 -24404 26990 -24204 8 VDD
port 41 nsew
rlabel metal1 s 24565 -24804 24611 -24104 8 VDD
port 41 nsew
rlabel metal1 s 24369 -24804 24415 -24104 8 VDD
port 41 nsew
rlabel metal1 s 24165 -24804 24211 -24104 8 VDD
port 41 nsew
rlabel metal1 s 23969 -24804 24015 -24104 8 VDD
port 41 nsew
rlabel metal1 s 23565 -24804 23611 -24104 8 VDD
port 41 nsew
rlabel metal1 s 23369 -24804 23415 -24104 8 VDD
port 41 nsew
rlabel metal1 s 23165 -24804 23211 -24104 8 VDD
port 41 nsew
rlabel metal1 s 22969 -24804 23015 -24104 8 VDD
port 41 nsew
rlabel metal1 s 22565 -24804 22611 -24104 8 VDD
port 41 nsew
rlabel metal1 s 22369 -24804 22415 -24104 8 VDD
port 41 nsew
rlabel metal1 s 22165 -24804 22211 -24104 8 VDD
port 41 nsew
rlabel metal1 s 21969 -24804 22015 -24104 8 VDD
port 41 nsew
rlabel metal1 s 21481 -24875 21527 -24675 8 VDD
port 41 nsew
rlabel metal1 s 21285 -24875 21331 -24675 8 VDD
port 41 nsew
rlabel metal1 s 21089 -24875 21135 -24675 8 VDD
port 41 nsew
rlabel metal1 s 20556 -24882 20602 -24682 8 VDD
port 41 nsew
rlabel metal1 s 20360 -24882 20406 -24682 8 VDD
port 41 nsew
rlabel metal1 s 19818 -24882 19864 -24682 8 VDD
port 41 nsew
rlabel metal1 s 19622 -24882 19668 -24682 8 VDD
port 41 nsew
rlabel metal1 s 19426 -24882 19472 -24682 8 VDD
port 41 nsew
rlabel metal1 s 19230 -24882 19276 -24682 8 VDD
port 41 nsew
rlabel metal1 s 18510 -24848 18556 -24448 8 VDD
port 41 nsew
rlabel metal1 s 18314 -24848 18360 -24448 8 VDD
port 41 nsew
rlabel metal1 s 17564 -24848 17610 -24448 8 VDD
port 41 nsew
rlabel metal1 s 17368 -24848 17414 -24448 8 VDD
port 41 nsew
rlabel metal1 s 3421 -25076 3467 -24776 8 VDD
port 41 nsew
rlabel metal1 s 3225 -25076 3271 -24776 8 VDD
port 41 nsew
rlabel metal1 s 3029 -25076 3075 -24776 8 VDD
port 41 nsew
rlabel metal1 s 2812 -25077 2858 -24977 8 VDD
port 41 nsew
rlabel metal1 s 2616 -25077 2662 -24977 8 VDD
port 41 nsew
rlabel metal1 s 2420 -25077 2466 -24977 8 VDD
port 41 nsew
rlabel metal1 s 2224 -25077 2270 -24977 8 VDD
port 41 nsew
rlabel metal1 s 1816 -25078 1862 -24778 8 VDD
port 41 nsew
rlabel metal1 s 1620 -25078 1666 -24778 8 VDD
port 41 nsew
rlabel metal1 s 1424 -25078 1470 -24778 8 VDD
port 41 nsew
rlabel metal1 s 1207 -25079 1253 -24979 8 VDD
port 41 nsew
rlabel metal1 s 1011 -25079 1057 -24979 8 VDD
port 41 nsew
rlabel metal1 s 815 -25079 861 -24979 8 VDD
port 41 nsew
rlabel metal1 s 619 -25079 665 -24979 8 VDD
port 41 nsew
rlabel metal1 s 212 -25092 258 -24892 8 VDD
port 41 nsew
rlabel metal1 s 16 -25092 62 -24892 8 VDD
port 41 nsew
rlabel metal1 s -180 -25092 -134 -24892 2 VDD
port 41 nsew
rlabel metal1 s -376 -25092 -330 -24892 2 VDD
port 41 nsew
rlabel metal1 s -918 -25092 -872 -24892 2 VDD
port 41 nsew
rlabel metal1 s -1114 -25092 -1068 -24892 2 VDD
port 41 nsew
rlabel metal1 s -1456 -25109 -1410 -24909 2 VDD
port 41 nsew
rlabel metal1 s -1652 -25109 -1606 -24909 2 VDD
port 41 nsew
rlabel metal1 s -1848 -25109 -1802 -24909 2 VDD
port 41 nsew
rlabel metal1 s -2338 -25109 -2292 -24909 2 VDD
port 41 nsew
rlabel metal1 s -2534 -25109 -2488 -24909 2 VDD
port 41 nsew
rlabel metal1 s -2730 -25109 -2684 -24909 2 VDD
port 41 nsew
rlabel metal1 s -4081 -25109 -4035 -24909 2 VDD
port 41 nsew
rlabel metal1 s -4277 -25109 -4231 -24909 2 VDD
port 41 nsew
rlabel metal1 s -4473 -25109 -4427 -24909 2 VDD
port 41 nsew
rlabel metal1 s -5038 -25109 -4992 -24909 2 VDD
port 41 nsew
rlabel metal1 s -5234 -25109 -5188 -24909 2 VDD
port 41 nsew
rlabel metal1 s -5430 -25109 -5384 -24909 2 VDD
port 41 nsew
rlabel metal1 s -6781 -25109 -6735 -24909 2 VDD
port 41 nsew
rlabel metal1 s -6977 -25109 -6931 -24909 2 VDD
port 41 nsew
rlabel metal1 s -7173 -25109 -7127 -24909 2 VDD
port 41 nsew
rlabel metal1 s -17043 -25657 -16997 -25057 2 VDD
port 41 nsew
rlabel metal1 s -17466 -25657 -17420 -25057 2 VDD
port 41 nsew
rlabel metal1 s -17662 -25657 -17616 -25057 2 VDD
port 41 nsew
rlabel metal1 s -17912 -25569 -17866 -25469 2 VDD
port 41 nsew
rlabel metal1 s -18108 -25569 -18062 -25469 2 VDD
port 41 nsew
rlabel metal1 s -18304 -25569 -18258 -25469 2 VDD
port 41 nsew
rlabel metal1 s -18500 -25569 -18454 -25469 2 VDD
port 41 nsew
rlabel metal1 s -18717 -25568 -18671 -25268 2 VDD
port 41 nsew
rlabel metal1 s -18913 -25568 -18867 -25268 2 VDD
port 41 nsew
rlabel metal1 s -19109 -25568 -19063 -25268 2 VDD
port 41 nsew
rlabel metal1 s -9330 -24842 -9284 -24642 2 VDD
port 41 nsew
rlabel metal1 s -9526 -24842 -9480 -24642 2 VDD
port 41 nsew
rlabel metal1 s -9722 -24842 -9676 -24642 2 VDD
port 41 nsew
rlabel metal1 s -10212 -24842 -10166 -24642 2 VDD
port 41 nsew
rlabel metal1 s -10408 -24842 -10362 -24642 2 VDD
port 41 nsew
rlabel metal1 s -10604 -24842 -10558 -24642 2 VDD
port 41 nsew
rlabel metal1 s -11955 -24842 -11909 -24642 2 VDD
port 41 nsew
rlabel metal1 s -12151 -24842 -12105 -24642 2 VDD
port 41 nsew
rlabel metal1 s -12347 -24842 -12301 -24642 2 VDD
port 41 nsew
rlabel metal1 s -12912 -24842 -12866 -24642 2 VDD
port 41 nsew
rlabel metal1 s -13108 -24842 -13062 -24642 2 VDD
port 41 nsew
rlabel metal1 s -13304 -24842 -13258 -24642 2 VDD
port 41 nsew
rlabel metal1 s -14655 -24842 -14609 -24642 2 VDD
port 41 nsew
rlabel metal1 s -14851 -24842 -14805 -24642 2 VDD
port 41 nsew
rlabel metal1 s -15047 -24842 -15001 -24642 2 VDD
port 41 nsew
rlabel metal1 s -19543 -25793 -19417 -24029 2 VDD
port 41 nsew
rlabel metal1 s -20315 -24739 -20269 -24339 2 VDD
port 41 nsew
rlabel metal1 s -20511 -24739 -20465 -24339 2 VDD
port 41 nsew
rlabel metal1 s -21220 -24738 -21174 -24338 2 VDD
port 41 nsew
rlabel metal1 s -21416 -24738 -21370 -24338 2 VDD
port 41 nsew
rlabel metal1 s -22426 -25009 -22380 -24409 2 VDD
port 41 nsew
rlabel metal1 s -22622 -25009 -22576 -24409 2 VDD
port 41 nsew
rlabel metal1 s -3342 -23791 -3296 -23591 2 VDD
port 41 nsew
rlabel metal1 s -3538 -23791 -3492 -23591 2 VDD
port 41 nsew
rlabel metal1 s -3734 -23791 -3688 -23591 2 VDD
port 41 nsew
rlabel metal1 s -4179 -23791 -4133 -23591 2 VDD
port 41 nsew
rlabel metal1 s -4375 -23791 -4329 -23591 2 VDD
port 41 nsew
rlabel metal1 s -4571 -23791 -4525 -23591 2 VDD
port 41 nsew
rlabel metal1 s -6042 -23791 -5996 -23591 2 VDD
port 41 nsew
rlabel metal1 s -6238 -23791 -6192 -23591 2 VDD
port 41 nsew
rlabel metal1 s -6434 -23791 -6388 -23591 2 VDD
port 41 nsew
rlabel metal1 s -6879 -23791 -6833 -23591 2 VDD
port 41 nsew
rlabel metal1 s -7075 -23791 -7029 -23591 2 VDD
port 41 nsew
rlabel metal1 s -7271 -23791 -7225 -23591 2 VDD
port 41 nsew
rlabel metal1 s 21531 -23574 21577 -23174 8 VDD
port 41 nsew
rlabel metal1 s 21335 -23574 21381 -23174 8 VDD
port 41 nsew
rlabel metal1 s 21139 -23574 21185 -23174 8 VDD
port 41 nsew
rlabel metal1 s -8137 -23941 -8091 -23341 2 VDD
port 41 nsew
rlabel metal1 s -8333 -23941 -8287 -23341 2 VDD
port 41 nsew
rlabel metal1 s -8756 -23941 -8710 -23341 2 VDD
port 41 nsew
rlabel metal1 s -19570 -24029 -19391 -23862 2 VDD
port 41 nsew
rlabel metal1 s -11216 -23524 -11170 -23324 2 VDD
port 41 nsew
rlabel metal1 s -11412 -23524 -11366 -23324 2 VDD
port 41 nsew
rlabel metal1 s -11608 -23524 -11562 -23324 2 VDD
port 41 nsew
rlabel metal1 s -12053 -23524 -12007 -23324 2 VDD
port 41 nsew
rlabel metal1 s -12249 -23524 -12203 -23324 2 VDD
port 41 nsew
rlabel metal1 s -12445 -23524 -12399 -23324 2 VDD
port 41 nsew
rlabel metal1 s -13916 -23524 -13870 -23324 2 VDD
port 41 nsew
rlabel metal1 s -14112 -23524 -14066 -23324 2 VDD
port 41 nsew
rlabel metal1 s -14308 -23524 -14262 -23324 2 VDD
port 41 nsew
rlabel metal1 s -14753 -23524 -14707 -23324 2 VDD
port 41 nsew
rlabel metal1 s -14949 -23524 -14903 -23324 2 VDD
port 41 nsew
rlabel metal1 s -15145 -23524 -15099 -23324 2 VDD
port 41 nsew
rlabel metal1 s 24411 -22622 24457 -22422 8 VDD
port 41 nsew
rlabel metal1 s 24215 -22622 24261 -22422 8 VDD
port 41 nsew
rlabel metal1 s 24019 -22622 24065 -22422 8 VDD
port 41 nsew
rlabel metal1 s 22668 -22622 22714 -22422 8 VDD
port 41 nsew
rlabel metal1 s 22472 -22622 22518 -22422 8 VDD
port 41 nsew
rlabel metal1 s 22276 -22622 22322 -22422 8 VDD
port 41 nsew
rlabel metal1 s 21711 -22622 21757 -22422 8 VDD
port 41 nsew
rlabel metal1 s 21515 -22622 21561 -22422 8 VDD
port 41 nsew
rlabel metal1 s 21319 -22622 21365 -22422 8 VDD
port 41 nsew
rlabel metal1 s 19968 -22622 20014 -22422 8 VDD
port 41 nsew
rlabel metal1 s 19772 -22622 19818 -22422 8 VDD
port 41 nsew
rlabel metal1 s 19576 -22622 19622 -22422 8 VDD
port 41 nsew
rlabel metal1 s 19086 -22622 19132 -22422 8 VDD
port 41 nsew
rlabel metal1 s 18890 -22622 18936 -22422 8 VDD
port 41 nsew
rlabel metal1 s 18694 -22622 18740 -22422 8 VDD
port 41 nsew
rlabel metal1 s 85482 -21644 85528 -21344 8 VDD
port 41 nsew
rlabel metal1 s 85286 -21644 85332 -21344 8 VDD
port 41 nsew
rlabel metal1 s 85058 -21844 85104 -21344 8 VDD
port 41 nsew
rlabel metal1 s 84928 -21844 84974 -21344 8 VDD
port 41 nsew
rlabel metal1 s 84333 -21844 84379 -21344 8 VDD
port 41 nsew
rlabel metal1 s 84137 -21844 84183 -21344 8 VDD
port 41 nsew
rlabel metal1 s 82764 -22086 82810 -21486 8 VDD
port 41 nsew
rlabel metal1 s 82341 -22086 82387 -21486 8 VDD
port 41 nsew
rlabel metal1 s 82145 -22086 82191 -21486 8 VDD
port 41 nsew
rlabel metal1 s 81895 -21674 81941 -21574 8 VDD
port 41 nsew
rlabel metal1 s 81699 -21674 81745 -21574 8 VDD
port 41 nsew
rlabel metal1 s 81503 -21674 81549 -21574 8 VDD
port 41 nsew
rlabel metal1 s 81307 -21674 81353 -21574 8 VDD
port 41 nsew
rlabel metal1 s 81090 -21875 81136 -21575 8 VDD
port 41 nsew
rlabel metal1 s 80894 -21875 80940 -21575 8 VDD
port 41 nsew
rlabel metal1 s 80698 -21875 80744 -21575 8 VDD
port 41 nsew
rlabel metal1 s 83204 -21405 83314 -21387 8 VDD
port 41 nsew
rlabel metal1 s 82976 -21393 83050 -21387 8 VDD
port 41 nsew
rlabel metal1 s 82976 -21387 83314 -21291 8 VDD
port 41 nsew
rlabel metal1 s 76118 -21682 76164 -21382 8 VDD
port 41 nsew
rlabel metal1 s 75922 -21682 75968 -21382 8 VDD
port 41 nsew
rlabel metal1 s 75694 -21882 75740 -21382 8 VDD
port 41 nsew
rlabel metal1 s 75564 -21882 75610 -21382 8 VDD
port 41 nsew
rlabel metal1 s 74969 -21882 75015 -21382 8 VDD
port 41 nsew
rlabel metal1 s 74773 -21882 74819 -21382 8 VDD
port 41 nsew
rlabel metal1 s 73400 -22124 73446 -21524 8 VDD
port 41 nsew
rlabel metal1 s 72977 -22124 73023 -21524 8 VDD
port 41 nsew
rlabel metal1 s 72781 -22124 72827 -21524 8 VDD
port 41 nsew
rlabel metal1 s 72531 -21712 72577 -21612 8 VDD
port 41 nsew
rlabel metal1 s 72335 -21712 72381 -21612 8 VDD
port 41 nsew
rlabel metal1 s 72139 -21712 72185 -21612 8 VDD
port 41 nsew
rlabel metal1 s 71943 -21712 71989 -21612 8 VDD
port 41 nsew
rlabel metal1 s 71726 -21913 71772 -21613 8 VDD
port 41 nsew
rlabel metal1 s 71530 -21913 71576 -21613 8 VDD
port 41 nsew
rlabel metal1 s 71334 -21913 71380 -21613 8 VDD
port 41 nsew
rlabel metal1 s 73840 -21443 73950 -21425 8 VDD
port 41 nsew
rlabel metal1 s 73612 -21431 73686 -21425 8 VDD
port 41 nsew
rlabel metal1 s 73612 -21425 73950 -21329 8 VDD
port 41 nsew
rlabel metal1 s 66965 -21699 67011 -21399 8 VDD
port 41 nsew
rlabel metal1 s 66769 -21699 66815 -21399 8 VDD
port 41 nsew
rlabel metal1 s 66541 -21899 66587 -21399 8 VDD
port 41 nsew
rlabel metal1 s 66411 -21899 66457 -21399 8 VDD
port 41 nsew
rlabel metal1 s 65816 -21899 65862 -21399 8 VDD
port 41 nsew
rlabel metal1 s 65620 -21899 65666 -21399 8 VDD
port 41 nsew
rlabel metal1 s 64247 -22141 64293 -21541 8 VDD
port 41 nsew
rlabel metal1 s 63824 -22141 63870 -21541 8 VDD
port 41 nsew
rlabel metal1 s 63628 -22141 63674 -21541 8 VDD
port 41 nsew
rlabel metal1 s 63378 -21729 63424 -21629 8 VDD
port 41 nsew
rlabel metal1 s 63182 -21729 63228 -21629 8 VDD
port 41 nsew
rlabel metal1 s 62986 -21729 63032 -21629 8 VDD
port 41 nsew
rlabel metal1 s 62790 -21729 62836 -21629 8 VDD
port 41 nsew
rlabel metal1 s 62573 -21930 62619 -21630 8 VDD
port 41 nsew
rlabel metal1 s 62377 -21930 62423 -21630 8 VDD
port 41 nsew
rlabel metal1 s 62181 -21930 62227 -21630 8 VDD
port 41 nsew
rlabel metal1 s 58211 -21765 58257 -21465 8 VDD
port 41 nsew
rlabel metal1 s 58015 -21765 58061 -21465 8 VDD
port 41 nsew
rlabel metal1 s 57787 -21965 57833 -21465 8 VDD
port 41 nsew
rlabel metal1 s 57657 -21965 57703 -21465 8 VDD
port 41 nsew
rlabel metal1 s 57062 -21965 57108 -21465 8 VDD
port 41 nsew
rlabel metal1 s 56866 -21965 56912 -21465 8 VDD
port 41 nsew
rlabel metal1 s 55493 -22207 55539 -21607 8 VDD
port 41 nsew
rlabel metal1 s 55070 -22207 55116 -21607 8 VDD
port 41 nsew
rlabel metal1 s 54874 -22207 54920 -21607 8 VDD
port 41 nsew
rlabel metal1 s 54624 -21795 54670 -21695 8 VDD
port 41 nsew
rlabel metal1 s 54428 -21795 54474 -21695 8 VDD
port 41 nsew
rlabel metal1 s 54232 -21795 54278 -21695 8 VDD
port 41 nsew
rlabel metal1 s 54036 -21795 54082 -21695 8 VDD
port 41 nsew
rlabel metal1 s 53819 -21996 53865 -21696 8 VDD
port 41 nsew
rlabel metal1 s 53623 -21996 53669 -21696 8 VDD
port 41 nsew
rlabel metal1 s 53427 -21996 53473 -21696 8 VDD
port 41 nsew
rlabel metal1 s 55933 -21526 56043 -21508 8 VDD
port 41 nsew
rlabel metal1 s 55705 -21514 55779 -21508 8 VDD
port 41 nsew
rlabel metal1 s 64687 -21460 64797 -21442 8 VDD
port 41 nsew
rlabel metal1 s 64459 -21448 64533 -21442 8 VDD
port 41 nsew
rlabel metal1 s 73840 -21329 73950 -21293 8 VDD
port 41 nsew
rlabel metal1 s 73612 -21329 73686 -21313 8 VDD
port 41 nsew
rlabel metal1 s 64459 -21442 64797 -21346 8 VDD
port 41 nsew
rlabel metal1 s 55705 -21508 56043 -21412 8 VDD
port 41 nsew
rlabel metal1 s 49013 -21799 49059 -21499 8 VDD
port 41 nsew
rlabel metal1 s 48817 -21799 48863 -21499 8 VDD
port 41 nsew
rlabel metal1 s 48589 -21999 48635 -21499 8 VDD
port 41 nsew
rlabel metal1 s 48459 -21999 48505 -21499 8 VDD
port 41 nsew
rlabel metal1 s 47864 -21999 47910 -21499 8 VDD
port 41 nsew
rlabel metal1 s 47668 -21999 47714 -21499 8 VDD
port 41 nsew
rlabel metal1 s 46295 -22241 46341 -21641 8 VDD
port 41 nsew
rlabel metal1 s 45872 -22241 45918 -21641 8 VDD
port 41 nsew
rlabel metal1 s 45676 -22241 45722 -21641 8 VDD
port 41 nsew
rlabel metal1 s 45426 -21829 45472 -21729 8 VDD
port 41 nsew
rlabel metal1 s 45230 -21829 45276 -21729 8 VDD
port 41 nsew
rlabel metal1 s 45034 -21829 45080 -21729 8 VDD
port 41 nsew
rlabel metal1 s 44838 -21829 44884 -21729 8 VDD
port 41 nsew
rlabel metal1 s 44621 -22030 44667 -21730 8 VDD
port 41 nsew
rlabel metal1 s 44425 -22030 44471 -21730 8 VDD
port 41 nsew
rlabel metal1 s 44229 -22030 44275 -21730 8 VDD
port 41 nsew
rlabel metal1 s 46735 -21560 46845 -21542 8 VDD
port 41 nsew
rlabel metal1 s 46507 -21548 46581 -21542 8 VDD
port 41 nsew
rlabel metal1 s 55933 -21412 56043 -21376 8 VDD
port 41 nsew
rlabel metal1 s 55705 -21412 55779 -21396 8 VDD
port 41 nsew
rlabel metal1 s 46507 -21542 46845 -21446 8 VDD
port 41 nsew
rlabel metal1 s 40150 -21760 40196 -21460 8 VDD
port 41 nsew
rlabel metal1 s 39954 -21760 40000 -21460 8 VDD
port 41 nsew
rlabel metal1 s 39726 -21960 39772 -21460 8 VDD
port 41 nsew
rlabel metal1 s 39596 -21960 39642 -21460 8 VDD
port 41 nsew
rlabel metal1 s 39001 -21960 39047 -21460 8 VDD
port 41 nsew
rlabel metal1 s 38805 -21960 38851 -21460 8 VDD
port 41 nsew
rlabel metal1 s 37432 -22202 37478 -21602 8 VDD
port 41 nsew
rlabel metal1 s 37009 -22202 37055 -21602 8 VDD
port 41 nsew
rlabel metal1 s 36813 -22202 36859 -21602 8 VDD
port 41 nsew
rlabel metal1 s 36563 -21790 36609 -21690 8 VDD
port 41 nsew
rlabel metal1 s 36367 -21790 36413 -21690 8 VDD
port 41 nsew
rlabel metal1 s 36171 -21790 36217 -21690 8 VDD
port 41 nsew
rlabel metal1 s 35975 -21790 36021 -21690 8 VDD
port 41 nsew
rlabel metal1 s 35758 -21991 35804 -21691 8 VDD
port 41 nsew
rlabel metal1 s 35562 -21991 35608 -21691 8 VDD
port 41 nsew
rlabel metal1 s 35366 -21991 35412 -21691 8 VDD
port 41 nsew
rlabel metal1 s 37872 -21521 37982 -21503 8 VDD
port 41 nsew
rlabel metal1 s 37644 -21509 37718 -21503 8 VDD
port 41 nsew
rlabel metal1 s 46735 -21446 46845 -21410 8 VDD
port 41 nsew
rlabel metal1 s 46507 -21446 46581 -21430 8 VDD
port 41 nsew
rlabel metal1 s 37644 -21503 37982 -21407 8 VDD
port 41 nsew
rlabel metal1 s 31710 -21749 31756 -21449 8 VDD
port 41 nsew
rlabel metal1 s 31514 -21749 31560 -21449 8 VDD
port 41 nsew
rlabel metal1 s 31286 -21949 31332 -21449 8 VDD
port 41 nsew
rlabel metal1 s 31156 -21949 31202 -21449 8 VDD
port 41 nsew
rlabel metal1 s 30561 -21949 30607 -21449 8 VDD
port 41 nsew
rlabel metal1 s 30365 -21949 30411 -21449 8 VDD
port 41 nsew
rlabel metal1 s 28992 -22191 29038 -21591 8 VDD
port 41 nsew
rlabel metal1 s 28569 -22191 28615 -21591 8 VDD
port 41 nsew
rlabel metal1 s 28373 -22191 28419 -21591 8 VDD
port 41 nsew
rlabel metal1 s 28123 -21779 28169 -21679 8 VDD
port 41 nsew
rlabel metal1 s 27927 -21779 27973 -21679 8 VDD
port 41 nsew
rlabel metal1 s 27731 -21779 27777 -21679 8 VDD
port 41 nsew
rlabel metal1 s 27535 -21779 27581 -21679 8 VDD
port 41 nsew
rlabel metal1 s 27318 -21980 27364 -21680 8 VDD
port 41 nsew
rlabel metal1 s 27122 -21980 27168 -21680 8 VDD
port 41 nsew
rlabel metal1 s 26926 -21980 26972 -21680 8 VDD
port 41 nsew
rlabel metal1 s 17569 -22502 17615 -21902 8 VDD
port 41 nsew
rlabel metal1 s 17373 -22502 17419 -21902 8 VDD
port 41 nsew
rlabel metal1 s -3342 -22353 -3296 -22153 2 VDD
port 41 nsew
rlabel metal1 s -3538 -22353 -3492 -22153 2 VDD
port 41 nsew
rlabel metal1 s -3734 -22353 -3688 -22153 2 VDD
port 41 nsew
rlabel metal1 s -4179 -22353 -4133 -22153 2 VDD
port 41 nsew
rlabel metal1 s -4375 -22353 -4329 -22153 2 VDD
port 41 nsew
rlabel metal1 s -4571 -22353 -4525 -22153 2 VDD
port 41 nsew
rlabel metal1 s -6042 -22353 -5996 -22153 2 VDD
port 41 nsew
rlabel metal1 s -6238 -22353 -6192 -22153 2 VDD
port 41 nsew
rlabel metal1 s -6434 -22353 -6388 -22153 2 VDD
port 41 nsew
rlabel metal1 s -6879 -22353 -6833 -22153 2 VDD
port 41 nsew
rlabel metal1 s -7075 -22353 -7029 -22153 2 VDD
port 41 nsew
rlabel metal1 s -7271 -22353 -7225 -22153 2 VDD
port 41 nsew
rlabel metal1 s -11924 -22243 -11878 -22143 2 VDD
port 41 nsew
rlabel metal1 s -12120 -22243 -12074 -22143 2 VDD
port 41 nsew
rlabel metal1 s -12316 -22243 -12270 -22143 2 VDD
port 41 nsew
rlabel metal1 s -12512 -22243 -12466 -22143 2 VDD
port 41 nsew
rlabel metal1 s -12729 -22444 -12683 -22144 2 VDD
port 41 nsew
rlabel metal1 s -12925 -22444 -12879 -22144 2 VDD
port 41 nsew
rlabel metal1 s -13121 -22444 -13075 -22144 2 VDD
port 41 nsew
rlabel metal1 s -13506 -22473 -13460 -22273 2 VDD
port 41 nsew
rlabel metal1 s -13702 -22473 -13656 -22273 2 VDD
port 41 nsew
rlabel metal1 s -13898 -22473 -13852 -22273 2 VDD
port 41 nsew
rlabel metal1 s -14094 -22473 -14048 -22273 2 VDD
port 41 nsew
rlabel metal1 s 29432 -21510 29542 -21492 8 VDD
port 41 nsew
rlabel metal1 s 29204 -21498 29278 -21492 8 VDD
port 41 nsew
rlabel metal1 s 37872 -21407 37982 -21371 8 VDD
port 41 nsew
rlabel metal1 s 37644 -21407 37718 -21391 8 VDD
port 41 nsew
rlabel metal1 s 29204 -21492 29542 -21396 8 VDD
port 41 nsew
rlabel metal1 s 29432 -21396 29542 -21360 8 VDD
port 41 nsew
rlabel metal1 s 29204 -21396 29278 -21380 8 VDD
port 41 nsew
rlabel metal1 s 64687 -21346 64797 -21310 8 VDD
port 41 nsew
rlabel metal1 s 64459 -21346 64533 -21330 8 VDD
port 41 nsew
rlabel metal1 s 83204 -21291 83314 -21255 8 VDD
port 41 nsew
rlabel metal1 s 82976 -21291 83050 -21275 8 VDD
port 41 nsew
rlabel metal1 s 82894 -20976 82940 -20876 8 VDD
port 41 nsew
rlabel metal1 s 82698 -20976 82744 -20876 8 VDD
port 41 nsew
rlabel metal1 s 82502 -20976 82548 -20876 8 VDD
port 41 nsew
rlabel metal1 s 82306 -20976 82352 -20876 8 VDD
port 41 nsew
rlabel metal1 s 82089 -20975 82135 -20675 8 VDD
port 41 nsew
rlabel metal1 s 81893 -20975 81939 -20675 8 VDD
port 41 nsew
rlabel metal1 s 81697 -20975 81743 -20675 8 VDD
port 41 nsew
rlabel metal1 s 73530 -21014 73576 -20914 8 VDD
port 41 nsew
rlabel metal1 s 73334 -21014 73380 -20914 8 VDD
port 41 nsew
rlabel metal1 s 73138 -21014 73184 -20914 8 VDD
port 41 nsew
rlabel metal1 s 72942 -21014 72988 -20914 8 VDD
port 41 nsew
rlabel metal1 s 81312 -20846 81358 -20646 8 VDD
port 41 nsew
rlabel metal1 s 81116 -20846 81162 -20646 8 VDD
port 41 nsew
rlabel metal1 s 80920 -20846 80966 -20646 8 VDD
port 41 nsew
rlabel metal1 s 80724 -20846 80770 -20646 8 VDD
port 41 nsew
rlabel metal1 s 72725 -21013 72771 -20713 8 VDD
port 41 nsew
rlabel metal1 s 72529 -21013 72575 -20713 8 VDD
port 41 nsew
rlabel metal1 s 72333 -21013 72379 -20713 8 VDD
port 41 nsew
rlabel metal1 s 64377 -21031 64423 -20931 8 VDD
port 41 nsew
rlabel metal1 s 64181 -21031 64227 -20931 8 VDD
port 41 nsew
rlabel metal1 s 63985 -21031 64031 -20931 8 VDD
port 41 nsew
rlabel metal1 s 63789 -21031 63835 -20931 8 VDD
port 41 nsew
rlabel metal1 s 71948 -20884 71994 -20684 8 VDD
port 41 nsew
rlabel metal1 s 71752 -20884 71798 -20684 8 VDD
port 41 nsew
rlabel metal1 s 71556 -20884 71602 -20684 8 VDD
port 41 nsew
rlabel metal1 s 71360 -20884 71406 -20684 8 VDD
port 41 nsew
rlabel metal1 s 63572 -21030 63618 -20730 8 VDD
port 41 nsew
rlabel metal1 s 63376 -21030 63422 -20730 8 VDD
port 41 nsew
rlabel metal1 s 63180 -21030 63226 -20730 8 VDD
port 41 nsew
rlabel metal1 s 55623 -21097 55669 -20997 8 VDD
port 41 nsew
rlabel metal1 s 55427 -21097 55473 -20997 8 VDD
port 41 nsew
rlabel metal1 s 55231 -21097 55277 -20997 8 VDD
port 41 nsew
rlabel metal1 s 55035 -21097 55081 -20997 8 VDD
port 41 nsew
rlabel metal1 s 62795 -20901 62841 -20701 8 VDD
port 41 nsew
rlabel metal1 s 62599 -20901 62645 -20701 8 VDD
port 41 nsew
rlabel metal1 s 62403 -20901 62449 -20701 8 VDD
port 41 nsew
rlabel metal1 s 62207 -20901 62253 -20701 8 VDD
port 41 nsew
rlabel metal1 s 54818 -21096 54864 -20796 8 VDD
port 41 nsew
rlabel metal1 s 54622 -21096 54668 -20796 8 VDD
port 41 nsew
rlabel metal1 s 54426 -21096 54472 -20796 8 VDD
port 41 nsew
rlabel metal1 s 46425 -21131 46471 -21031 8 VDD
port 41 nsew
rlabel metal1 s 46229 -21131 46275 -21031 8 VDD
port 41 nsew
rlabel metal1 s 46033 -21131 46079 -21031 8 VDD
port 41 nsew
rlabel metal1 s 45837 -21131 45883 -21031 8 VDD
port 41 nsew
rlabel metal1 s 54041 -20967 54087 -20767 8 VDD
port 41 nsew
rlabel metal1 s 53845 -20967 53891 -20767 8 VDD
port 41 nsew
rlabel metal1 s 53649 -20967 53695 -20767 8 VDD
port 41 nsew
rlabel metal1 s 53453 -20967 53499 -20767 8 VDD
port 41 nsew
rlabel metal1 s 45620 -21130 45666 -20830 8 VDD
port 41 nsew
rlabel metal1 s 45424 -21130 45470 -20830 8 VDD
port 41 nsew
rlabel metal1 s 45228 -21130 45274 -20830 8 VDD
port 41 nsew
rlabel metal1 s 24509 -21304 24555 -21104 8 VDD
port 41 nsew
rlabel metal1 s 24313 -21304 24359 -21104 8 VDD
port 41 nsew
rlabel metal1 s 24117 -21304 24163 -21104 8 VDD
port 41 nsew
rlabel metal1 s 23672 -21304 23718 -21104 8 VDD
port 41 nsew
rlabel metal1 s 23476 -21304 23522 -21104 8 VDD
port 41 nsew
rlabel metal1 s 23280 -21304 23326 -21104 8 VDD
port 41 nsew
rlabel metal1 s 21809 -21304 21855 -21104 8 VDD
port 41 nsew
rlabel metal1 s 21613 -21304 21659 -21104 8 VDD
port 41 nsew
rlabel metal1 s 21417 -21304 21463 -21104 8 VDD
port 41 nsew
rlabel metal1 s 20972 -21304 21018 -21104 8 VDD
port 41 nsew
rlabel metal1 s 20776 -21304 20822 -21104 8 VDD
port 41 nsew
rlabel metal1 s 20580 -21304 20626 -21104 8 VDD
port 41 nsew
rlabel metal1 s 44843 -21001 44889 -20801 8 VDD
port 41 nsew
rlabel metal1 s 44647 -21001 44693 -20801 8 VDD
port 41 nsew
rlabel metal1 s 44451 -21001 44497 -20801 8 VDD
port 41 nsew
rlabel metal1 s 44255 -21001 44301 -20801 8 VDD
port 41 nsew
rlabel metal1 s 37562 -21092 37608 -20992 8 VDD
port 41 nsew
rlabel metal1 s 37366 -21092 37412 -20992 8 VDD
port 41 nsew
rlabel metal1 s 37170 -21092 37216 -20992 8 VDD
port 41 nsew
rlabel metal1 s 36974 -21092 37020 -20992 8 VDD
port 41 nsew
rlabel metal1 s 36757 -21091 36803 -20791 8 VDD
port 41 nsew
rlabel metal1 s 36561 -21091 36607 -20791 8 VDD
port 41 nsew
rlabel metal1 s 36365 -21091 36411 -20791 8 VDD
port 41 nsew
rlabel metal1 s 29122 -21081 29168 -20981 8 VDD
port 41 nsew
rlabel metal1 s 28926 -21081 28972 -20981 8 VDD
port 41 nsew
rlabel metal1 s 28730 -21081 28776 -20981 8 VDD
port 41 nsew
rlabel metal1 s 28534 -21081 28580 -20981 8 VDD
port 41 nsew
rlabel metal1 s 35980 -20962 36026 -20762 8 VDD
port 41 nsew
rlabel metal1 s 35784 -20962 35830 -20762 8 VDD
port 41 nsew
rlabel metal1 s 35588 -20962 35634 -20762 8 VDD
port 41 nsew
rlabel metal1 s 35392 -20962 35438 -20762 8 VDD
port 41 nsew
rlabel metal1 s 28317 -21080 28363 -20780 8 VDD
port 41 nsew
rlabel metal1 s 28121 -21080 28167 -20780 8 VDD
port 41 nsew
rlabel metal1 s 27925 -21080 27971 -20780 8 VDD
port 41 nsew
rlabel metal1 s 27540 -20951 27586 -20751 8 VDD
port 41 nsew
rlabel metal1 s 27344 -20951 27390 -20751 8 VDD
port 41 nsew
rlabel metal1 s 27148 -20951 27194 -20751 8 VDD
port 41 nsew
rlabel metal1 s 26952 -20951 26998 -20751 8 VDD
port 41 nsew
rlabel metal1 s 7346 -21054 7392 -20854 8 VDD
port 41 nsew
rlabel metal1 s 7150 -21054 7196 -20854 8 VDD
port 41 nsew
rlabel metal1 s 7037 -21054 7083 -20854 8 VDD
port 41 nsew
rlabel metal1 s 6841 -21054 6887 -20854 8 VDD
port 41 nsew
rlabel metal1 s 6727 -21054 6773 -20854 8 VDD
port 41 nsew
rlabel metal1 s 6531 -21054 6577 -20854 8 VDD
port 41 nsew
rlabel metal1 s 6335 -21054 6381 -20854 8 VDD
port 41 nsew
rlabel metal1 s 5174 -21043 5220 -20843 8 VDD
port 41 nsew
rlabel metal1 s 4978 -21043 5024 -20843 8 VDD
port 41 nsew
rlabel metal1 s 4782 -21043 4828 -20843 8 VDD
port 41 nsew
rlabel metal1 s 4586 -21043 4632 -20843 8 VDD
port 41 nsew
rlabel metal1 s 4044 -21043 4090 -20843 8 VDD
port 41 nsew
rlabel metal1 s 3848 -21043 3894 -20843 8 VDD
port 41 nsew
rlabel metal1 s 3421 -21168 3467 -20868 8 VDD
port 41 nsew
rlabel metal1 s 3225 -21168 3271 -20868 8 VDD
port 41 nsew
rlabel metal1 s 3029 -21168 3075 -20868 8 VDD
port 41 nsew
rlabel metal1 s 2812 -20967 2858 -20867 8 VDD
port 41 nsew
rlabel metal1 s 2616 -20967 2662 -20867 8 VDD
port 41 nsew
rlabel metal1 s 2420 -20967 2466 -20867 8 VDD
port 41 nsew
rlabel metal1 s 2224 -20967 2270 -20867 8 VDD
port 41 nsew
rlabel metal1 s 1816 -21166 1862 -20866 8 VDD
port 41 nsew
rlabel metal1 s 1620 -21166 1666 -20866 8 VDD
port 41 nsew
rlabel metal1 s 1424 -21166 1470 -20866 8 VDD
port 41 nsew
rlabel metal1 s 1207 -20965 1253 -20865 8 VDD
port 41 nsew
rlabel metal1 s 1011 -20965 1057 -20865 8 VDD
port 41 nsew
rlabel metal1 s 815 -20965 861 -20865 8 VDD
port 41 nsew
rlabel metal1 s 619 -20965 665 -20865 8 VDD
port 41 nsew
rlabel metal1 s 212 -21052 258 -20852 8 VDD
port 41 nsew
rlabel metal1 s 16 -21052 62 -20852 8 VDD
port 41 nsew
rlabel metal1 s -180 -21052 -134 -20852 2 VDD
port 41 nsew
rlabel metal1 s -376 -21052 -330 -20852 2 VDD
port 41 nsew
rlabel metal1 s -918 -21052 -872 -20852 2 VDD
port 41 nsew
rlabel metal1 s -1114 -21052 -1068 -20852 2 VDD
port 41 nsew
rlabel metal1 s -1456 -21035 -1410 -20835 2 VDD
port 41 nsew
rlabel metal1 s -1652 -21035 -1606 -20835 2 VDD
port 41 nsew
rlabel metal1 s -1848 -21035 -1802 -20835 2 VDD
port 41 nsew
rlabel metal1 s -2338 -21035 -2292 -20835 2 VDD
port 41 nsew
rlabel metal1 s -2534 -21035 -2488 -20835 2 VDD
port 41 nsew
rlabel metal1 s -2730 -21035 -2684 -20835 2 VDD
port 41 nsew
rlabel metal1 s -4081 -21035 -4035 -20835 2 VDD
port 41 nsew
rlabel metal1 s -4277 -21035 -4231 -20835 2 VDD
port 41 nsew
rlabel metal1 s -4473 -21035 -4427 -20835 2 VDD
port 41 nsew
rlabel metal1 s -5038 -21035 -4992 -20835 2 VDD
port 41 nsew
rlabel metal1 s -5234 -21035 -5188 -20835 2 VDD
port 41 nsew
rlabel metal1 s -5430 -21035 -5384 -20835 2 VDD
port 41 nsew
rlabel metal1 s -6781 -21035 -6735 -20835 2 VDD
port 41 nsew
rlabel metal1 s -6977 -21035 -6931 -20835 2 VDD
port 41 nsew
rlabel metal1 s -7173 -21035 -7127 -20835 2 VDD
port 41 nsew
rlabel metal1 s -12054 -21633 -12008 -21033 2 VDD
port 41 nsew
rlabel metal1 s -12477 -21633 -12431 -21033 2 VDD
port 41 nsew
rlabel metal1 s -12673 -21633 -12627 -21033 2 VDD
port 41 nsew
rlabel metal1 s -12923 -21545 -12877 -21445 2 VDD
port 41 nsew
rlabel metal1 s -13119 -21545 -13073 -21445 2 VDD
port 41 nsew
rlabel metal1 s -13315 -21545 -13269 -21445 2 VDD
port 41 nsew
rlabel metal1 s -13511 -21545 -13465 -21445 2 VDD
port 41 nsew
rlabel metal1 s -13728 -21544 -13682 -21244 2 VDD
port 41 nsew
rlabel metal1 s -13924 -21544 -13878 -21244 2 VDD
port 41 nsew
rlabel metal1 s -14120 -21544 -14074 -21244 2 VDD
port 41 nsew
rlabel metal1 s -16913 -21267 -16867 -21167 2 VDD
port 41 nsew
rlabel metal1 s -17109 -21267 -17063 -21167 2 VDD
port 41 nsew
rlabel metal1 s -17305 -21267 -17259 -21167 2 VDD
port 41 nsew
rlabel metal1 s -17501 -21267 -17455 -21167 2 VDD
port 41 nsew
rlabel metal1 s -17718 -21468 -17672 -21168 2 VDD
port 41 nsew
rlabel metal1 s -17914 -21468 -17868 -21168 2 VDD
port 41 nsew
rlabel metal1 s -18110 -21468 -18064 -21168 2 VDD
port 41 nsew
rlabel metal1 s -18495 -21497 -18449 -21297 2 VDD
port 41 nsew
rlabel metal1 s -18691 -21497 -18645 -21297 2 VDD
port 41 nsew
rlabel metal1 s -18887 -21497 -18841 -21297 2 VDD
port 41 nsew
rlabel metal1 s -19083 -21497 -19037 -21297 2 VDD
port 41 nsew
rlabel metal1 s -19588 -21320 -19542 -21120 2 VDD
port 41 nsew
rlabel metal1 s -19784 -21320 -19738 -21120 2 VDD
port 41 nsew
rlabel metal1 s -20326 -21320 -20280 -21120 2 VDD
port 41 nsew
rlabel metal1 s -20522 -21320 -20476 -21120 2 VDD
port 41 nsew
rlabel metal1 s -20718 -21320 -20672 -21120 2 VDD
port 41 nsew
rlabel metal1 s -20914 -21320 -20868 -21120 2 VDD
port 41 nsew
rlabel metal1 s -21490 -21314 -21444 -21214 2 VDD
port 41 nsew
rlabel metal1 s -21686 -21314 -21640 -21214 2 VDD
port 41 nsew
rlabel metal1 s -21882 -21314 -21836 -21214 2 VDD
port 41 nsew
rlabel metal1 s -22078 -21314 -22032 -21214 2 VDD
port 41 nsew
rlabel metal1 s -22295 -21515 -22249 -21215 2 VDD
port 41 nsew
rlabel metal1 s -22491 -21515 -22445 -21215 2 VDD
port 41 nsew
rlabel metal1 s -22687 -21515 -22641 -21215 2 VDD
port 41 nsew
rlabel metal1 s 2139 -20805 2262 -20792 8 VDD
port 41 nsew
rlabel metal1 s 1750 -20806 1873 -20792 8 VDD
port 41 nsew
rlabel metal1 s 6340 -20786 6463 -20767 8 VDD
port 41 nsew
rlabel metal1 s 5124 -20785 5247 -20767 8 VDD
port 41 nsew
rlabel metal1 s 5124 -20767 6463 -20662 8 VDD
port 41 nsew
rlabel metal1 s 6340 -20662 6463 -20650 8 VDD
port 41 nsew
rlabel metal1 s 5124 -20662 5247 -20649 8 VDD
port 41 nsew
rlabel metal1 s 3768 -20780 3891 -20762 8 VDD
port 41 nsew
rlabel metal1 s 3367 -20782 3490 -20762 8 VDD
port 41 nsew
rlabel metal1 s 3367 -20762 3891 -20655 8 VDD
port 41 nsew
rlabel metal1 s 1750 -20792 2262 -20685 8 VDD
port 41 nsew
rlabel metal1 s 2139 -20685 2262 -20669 8 VDD
port 41 nsew
rlabel metal1 s 1750 -20685 1873 -20670 8 VDD
port 41 nsew
rlabel metal1 s -1228 -20793 -1105 -20785 2 VDD
port 41 nsew
rlabel metal1 s -1522 -20794 -1399 -20785 2 VDD
port 41 nsew
rlabel metal1 s -1522 -20785 -1105 -20670 2 VDD
port 41 nsew
rlabel metal1 s -1228 -20670 -1105 -20657 2 VDD
port 41 nsew
rlabel metal1 s -1522 -20670 -1399 -20658 2 VDD
port 41 nsew
rlabel metal1 s 3768 -20655 3891 -20644 8 VDD
port 41 nsew
rlabel metal1 s 3367 -20655 3490 -20646 8 VDD
port 41 nsew
rlabel metal1 s -5348 -20128 -5225 -19992 2 VDD
port 41 nsew
rlabel metal1 s -298 -19876 8 -19814 2 VDD
port 41 nsew
rlabel metal1 s -2781 -19984 -2658 -19848 2 VDD
port 41 nsew
rlabel metal1 s -298 -19814 -175 -19813 2 VDD
port 41 nsew
rlabel metal1 s -293 -19813 -179 -19396 2 VDD
port 41 nsew
rlabel metal1 s -2776 -19848 -2662 -19396 2 VDD
port 41 nsew
rlabel metal1 s -297 -19396 -174 -19260 2 VDD
port 41 nsew
rlabel metal1 s -2780 -19396 -2657 -19260 2 VDD
port 41 nsew
rlabel metal1 s -5343 -19992 -5229 -19361 2 VDD
port 41 nsew
rlabel metal1 s -6622 -20132 -6576 -19932 2 VDD
port 41 nsew
rlabel metal1 s -6818 -20132 -6772 -19932 2 VDD
port 41 nsew
rlabel metal1 s -7014 -20132 -6968 -19932 2 VDD
port 41 nsew
rlabel metal1 s -17043 -20657 -16997 -20057 2 VDD
port 41 nsew
rlabel metal1 s -17466 -20657 -17420 -20057 2 VDD
port 41 nsew
rlabel metal1 s -17662 -20657 -17616 -20057 2 VDD
port 41 nsew
rlabel metal1 s -17912 -20569 -17866 -20469 2 VDD
port 41 nsew
rlabel metal1 s -18108 -20569 -18062 -20469 2 VDD
port 41 nsew
rlabel metal1 s -18304 -20569 -18258 -20469 2 VDD
port 41 nsew
rlabel metal1 s -18500 -20569 -18454 -20469 2 VDD
port 41 nsew
rlabel metal1 s -18717 -20568 -18671 -20268 2 VDD
port 41 nsew
rlabel metal1 s -18913 -20568 -18867 -20268 2 VDD
port 41 nsew
rlabel metal1 s -19109 -20568 -19063 -20268 2 VDD
port 41 nsew
rlabel metal1 s -9330 -19915 -9284 -19715 2 VDD
port 41 nsew
rlabel metal1 s -9526 -19915 -9480 -19715 2 VDD
port 41 nsew
rlabel metal1 s -9722 -19915 -9676 -19715 2 VDD
port 41 nsew
rlabel metal1 s -10212 -19915 -10166 -19715 2 VDD
port 41 nsew
rlabel metal1 s -10408 -19915 -10362 -19715 2 VDD
port 41 nsew
rlabel metal1 s -10604 -19915 -10558 -19715 2 VDD
port 41 nsew
rlabel metal1 s -11955 -19915 -11909 -19715 2 VDD
port 41 nsew
rlabel metal1 s -12151 -19915 -12105 -19715 2 VDD
port 41 nsew
rlabel metal1 s -12347 -19915 -12301 -19715 2 VDD
port 41 nsew
rlabel metal1 s -12912 -19915 -12866 -19715 2 VDD
port 41 nsew
rlabel metal1 s -13108 -19915 -13062 -19715 2 VDD
port 41 nsew
rlabel metal1 s -13304 -19915 -13258 -19715 2 VDD
port 41 nsew
rlabel metal1 s -14655 -19915 -14609 -19715 2 VDD
port 41 nsew
rlabel metal1 s -14851 -19915 -14805 -19715 2 VDD
port 41 nsew
rlabel metal1 s -15047 -19915 -15001 -19715 2 VDD
port 41 nsew
rlabel metal1 s -5347 -19361 -5224 -19225 2 VDD
port 41 nsew
rlabel metal1 s -19548 -19405 -19502 -19305 2 VDD
port 41 nsew
rlabel metal1 s -19744 -19405 -19698 -19305 2 VDD
port 41 nsew
rlabel metal1 s -19940 -19405 -19894 -19305 2 VDD
port 41 nsew
rlabel metal1 s -20136 -19405 -20090 -19305 2 VDD
port 41 nsew
rlabel metal1 s -20353 -19606 -20307 -19306 2 VDD
port 41 nsew
rlabel metal1 s -20549 -19606 -20503 -19306 2 VDD
port 41 nsew
rlabel metal1 s -20745 -19606 -20699 -19306 2 VDD
port 41 nsew
rlabel metal1 s -21418 -19384 -21372 -19184 2 VDD
port 41 nsew
rlabel metal1 s -21614 -19384 -21568 -19184 2 VDD
port 41 nsew
rlabel metal1 s -22156 -19384 -22110 -19184 2 VDD
port 41 nsew
rlabel metal1 s -22352 -19384 -22306 -19184 2 VDD
port 41 nsew
rlabel metal1 s -22548 -19384 -22502 -19184 2 VDD
port 41 nsew
rlabel metal1 s -22744 -19384 -22698 -19184 2 VDD
port 41 nsew
rlabel metal1 s 7336 -18803 7382 -18603 8 VDD
port 41 nsew
rlabel metal1 s 7140 -18803 7186 -18603 8 VDD
port 41 nsew
rlabel metal1 s 7027 -18803 7073 -18603 8 VDD
port 41 nsew
rlabel metal1 s 6831 -18803 6877 -18603 8 VDD
port 41 nsew
rlabel metal1 s 6717 -18803 6763 -18603 8 VDD
port 41 nsew
rlabel metal1 s 6521 -18803 6567 -18603 8 VDD
port 41 nsew
rlabel metal1 s 6325 -18803 6371 -18603 8 VDD
port 41 nsew
rlabel metal1 s 4336 -18803 4382 -18603 8 VDD
port 41 nsew
rlabel metal1 s 4140 -18803 4186 -18603 8 VDD
port 41 nsew
rlabel metal1 s 4027 -18803 4073 -18603 8 VDD
port 41 nsew
rlabel metal1 s 3831 -18803 3877 -18603 8 VDD
port 41 nsew
rlabel metal1 s 3717 -18803 3763 -18603 8 VDD
port 41 nsew
rlabel metal1 s 3521 -18803 3567 -18603 8 VDD
port 41 nsew
rlabel metal1 s 3325 -18803 3371 -18603 8 VDD
port 41 nsew
rlabel metal1 s 1836 -18803 1882 -18603 8 VDD
port 41 nsew
rlabel metal1 s 1640 -18803 1686 -18603 8 VDD
port 41 nsew
rlabel metal1 s 1527 -18803 1573 -18603 8 VDD
port 41 nsew
rlabel metal1 s 1331 -18803 1377 -18603 8 VDD
port 41 nsew
rlabel metal1 s 1217 -18803 1263 -18603 8 VDD
port 41 nsew
rlabel metal1 s 1021 -18803 1067 -18603 8 VDD
port 41 nsew
rlabel metal1 s 825 -18803 871 -18603 8 VDD
port 41 nsew
rlabel metal1 s -664 -18803 -618 -18603 2 VDD
port 41 nsew
rlabel metal1 s -860 -18803 -814 -18603 2 VDD
port 41 nsew
rlabel metal1 s -973 -18803 -927 -18603 2 VDD
port 41 nsew
rlabel metal1 s -1169 -18803 -1123 -18603 2 VDD
port 41 nsew
rlabel metal1 s -1283 -18803 -1237 -18603 2 VDD
port 41 nsew
rlabel metal1 s -1479 -18803 -1433 -18603 2 VDD
port 41 nsew
rlabel metal1 s -1675 -18803 -1629 -18603 2 VDD
port 41 nsew
rlabel metal1 s -3164 -18803 -3118 -18603 2 VDD
port 41 nsew
rlabel metal1 s -3360 -18803 -3314 -18603 2 VDD
port 41 nsew
rlabel metal1 s -3473 -18803 -3427 -18603 2 VDD
port 41 nsew
rlabel metal1 s -3669 -18803 -3623 -18603 2 VDD
port 41 nsew
rlabel metal1 s -3783 -18803 -3737 -18603 2 VDD
port 41 nsew
rlabel metal1 s -3979 -18803 -3933 -18603 2 VDD
port 41 nsew
rlabel metal1 s -4175 -18803 -4129 -18603 2 VDD
port 41 nsew
rlabel metal1 s -5664 -18803 -5618 -18603 2 VDD
port 41 nsew
rlabel metal1 s -5860 -18803 -5814 -18603 2 VDD
port 41 nsew
rlabel metal1 s -5973 -18803 -5927 -18603 2 VDD
port 41 nsew
rlabel metal1 s -6169 -18803 -6123 -18603 2 VDD
port 41 nsew
rlabel metal1 s -6283 -18803 -6237 -18603 2 VDD
port 41 nsew
rlabel metal1 s -6479 -18803 -6433 -18603 2 VDD
port 41 nsew
rlabel metal1 s -6675 -18803 -6629 -18603 2 VDD
port 41 nsew
rlabel metal1 s -8164 -19007 -8118 -18407 2 VDD
port 41 nsew
rlabel metal1 s -8360 -19007 -8314 -18407 2 VDD
port 41 nsew
rlabel metal1 s -8783 -19007 -8737 -18407 2 VDD
port 41 nsew
rlabel metal1 s -11216 -18597 -11170 -18397 2 VDD
port 41 nsew
rlabel metal1 s -11412 -18597 -11366 -18397 2 VDD
port 41 nsew
rlabel metal1 s -11608 -18597 -11562 -18397 2 VDD
port 41 nsew
rlabel metal1 s -12053 -18597 -12007 -18397 2 VDD
port 41 nsew
rlabel metal1 s -12249 -18597 -12203 -18397 2 VDD
port 41 nsew
rlabel metal1 s -12445 -18597 -12399 -18397 2 VDD
port 41 nsew
rlabel metal1 s -13916 -18597 -13870 -18397 2 VDD
port 41 nsew
rlabel metal1 s -14112 -18597 -14066 -18397 2 VDD
port 41 nsew
rlabel metal1 s -14308 -18597 -14262 -18397 2 VDD
port 41 nsew
rlabel metal1 s -14753 -18597 -14707 -18397 2 VDD
port 41 nsew
rlabel metal1 s -14949 -18597 -14903 -18397 2 VDD
port 41 nsew
rlabel metal1 s -15145 -18597 -15099 -18397 2 VDD
port 41 nsew
rlabel metal1 s -7585 -16536 -7539 -16136 2 VDD
port 41 nsew
rlabel metal1 s -7821 -16536 -7775 -16136 2 VDD
port 41 nsew
rlabel metal1 s -8057 -16536 -8011 -16136 2 VDD
port 41 nsew
rlabel metal1 s -8187 -16536 -8141 -16136 2 VDD
port 41 nsew
rlabel metal1 s -8423 -16536 -8377 -16136 2 VDD
port 41 nsew
rlabel metal1 s -8659 -16536 -8613 -16136 2 VDD
port 41 nsew
rlabel metal1 s -8895 -16536 -8849 -16136 2 VDD
port 41 nsew
rlabel metal1 s -9131 -16536 -9085 -16136 2 VDD
port 41 nsew
rlabel metal1 s -9261 -16536 -9215 -16136 2 VDD
port 41 nsew
rlabel metal1 s -9497 -16536 -9451 -16136 2 VDD
port 41 nsew
rlabel metal1 s -9733 -16536 -9687 -16136 2 VDD
port 41 nsew
rlabel metal1 s -9969 -16536 -9923 -16136 2 VDD
port 41 nsew
rlabel metal1 s -10205 -16536 -10159 -16136 2 VDD
port 41 nsew
rlabel metal1 s -10441 -16536 -10395 -16136 2 VDD
port 41 nsew
rlabel metal1 s -10677 -16536 -10631 -16136 2 VDD
port 41 nsew
rlabel metal1 s -10913 -16536 -10867 -16136 2 VDD
port 41 nsew
rlabel metal1 s -11149 -16536 -11103 -16136 2 VDD
port 41 nsew
rlabel metal1 s -11397 -16536 -11351 -16136 2 VDD
port 41 nsew
rlabel metal1 s -11633 -16536 -11587 -16136 2 VDD
port 41 nsew
rlabel metal1 s -11869 -16536 -11823 -16136 2 VDD
port 41 nsew
rlabel metal1 s -12105 -16536 -12059 -16136 2 VDD
port 41 nsew
rlabel metal1 s -12341 -16536 -12295 -16136 2 VDD
port 41 nsew
rlabel metal1 s -12577 -16536 -12531 -16136 2 VDD
port 41 nsew
rlabel metal1 s -12813 -16536 -12767 -16136 2 VDD
port 41 nsew
rlabel metal1 s -13049 -16536 -13003 -16136 2 VDD
port 41 nsew
rlabel metal1 s -13285 -16536 -13239 -16136 2 VDD
port 41 nsew
rlabel metal1 s -13521 -16536 -13475 -16136 2 VDD
port 41 nsew
rlabel metal1 s -13757 -16536 -13711 -16136 2 VDD
port 41 nsew
rlabel metal1 s -13993 -16536 -13947 -16136 2 VDD
port 41 nsew
rlabel metal1 s -14229 -16536 -14183 -16136 2 VDD
port 41 nsew
rlabel metal1 s -14465 -16536 -14419 -16136 2 VDD
port 41 nsew
rlabel metal1 s -14701 -16536 -14655 -16136 2 VDD
port 41 nsew
rlabel metal1 s -14937 -16536 -14891 -16136 2 VDD
port 41 nsew
rlabel metal1 s 63629 -4113 63675 -3913 8 VDD
port 41 nsew
rlabel metal1 s 63433 -4113 63479 -3913 8 VDD
port 41 nsew
rlabel metal1 s 63237 -4113 63283 -3913 8 VDD
port 41 nsew
rlabel metal1 s 63629 -3038 63675 -2838 8 VDD
port 41 nsew
rlabel metal1 s 63433 -3038 63479 -2838 8 VDD
port 41 nsew
rlabel metal1 s 63237 -3038 63283 -2838 8 VDD
port 41 nsew
rlabel metal1 s 62779 -3038 62825 -2838 8 VDD
port 41 nsew
rlabel metal1 s 62583 -3038 62629 -2838 8 VDD
port 41 nsew
rlabel metal1 s 62387 -3038 62433 -2838 8 VDD
port 41 nsew
rlabel metal1 s 58039 -3324 58085 -2924 8 VDD
port 41 nsew
rlabel metal1 s 57803 -3324 57849 -2924 8 VDD
port 41 nsew
rlabel metal1 s 57567 -3324 57613 -2924 8 VDD
port 41 nsew
rlabel metal1 s 57331 -3324 57377 -2924 8 VDD
port 41 nsew
rlabel metal1 s 57095 -3324 57141 -2924 8 VDD
port 41 nsew
rlabel metal1 s 56859 -3324 56905 -2924 8 VDD
port 41 nsew
rlabel metal1 s 56623 -3324 56669 -2924 8 VDD
port 41 nsew
rlabel metal1 s 56387 -3324 56433 -2924 8 VDD
port 41 nsew
rlabel metal1 s 56151 -3324 56197 -2924 8 VDD
port 41 nsew
rlabel metal1 s 55915 -3324 55961 -2924 8 VDD
port 41 nsew
rlabel metal1 s 55679 -3324 55725 -2924 8 VDD
port 41 nsew
rlabel metal1 s 55443 -3324 55489 -2924 8 VDD
port 41 nsew
rlabel metal1 s 55207 -3324 55253 -2924 8 VDD
port 41 nsew
rlabel metal1 s 54971 -3324 55017 -2924 8 VDD
port 41 nsew
rlabel metal1 s 54735 -3324 54781 -2924 8 VDD
port 41 nsew
rlabel metal1 s 54499 -3324 54545 -2924 8 VDD
port 41 nsew
rlabel metal1 s 54251 -3324 54297 -2924 8 VDD
port 41 nsew
rlabel metal1 s 54015 -3324 54061 -2924 8 VDD
port 41 nsew
rlabel metal1 s 53779 -3324 53825 -2924 8 VDD
port 41 nsew
rlabel metal1 s 53543 -3324 53589 -2924 8 VDD
port 41 nsew
rlabel metal1 s 53307 -3324 53353 -2924 8 VDD
port 41 nsew
rlabel metal1 s 53071 -3324 53117 -2924 8 VDD
port 41 nsew
rlabel metal1 s 52835 -3324 52881 -2924 8 VDD
port 41 nsew
rlabel metal1 s 52599 -3324 52645 -2924 8 VDD
port 41 nsew
rlabel metal1 s 52363 -3324 52409 -2924 8 VDD
port 41 nsew
rlabel metal1 s 52233 -3324 52279 -2924 8 VDD
port 41 nsew
rlabel metal1 s 51997 -3324 52043 -2924 8 VDD
port 41 nsew
rlabel metal1 s 51761 -3324 51807 -2924 8 VDD
port 41 nsew
rlabel metal1 s 51525 -3324 51571 -2924 8 VDD
port 41 nsew
rlabel metal1 s 51289 -3324 51335 -2924 8 VDD
port 41 nsew
rlabel metal1 s 51159 -3324 51205 -2924 8 VDD
port 41 nsew
rlabel metal1 s 50923 -3324 50969 -2924 8 VDD
port 41 nsew
rlabel metal1 s 50687 -3324 50733 -2924 8 VDD
port 41 nsew
rlabel metal1 s 5766 -1752 5812 -1552 8 VDD
port 41 nsew
rlabel metal1 s 5570 -1752 5616 -1552 8 VDD
port 41 nsew
rlabel metal1 s 5374 -1752 5420 -1552 8 VDD
port 41 nsew
rlabel metal1 s -3816 -1610 -3770 -1410 2 VDD
port 41 nsew
rlabel metal1 s -4012 -1610 -3966 -1410 2 VDD
port 41 nsew
rlabel metal1 s -4208 -1610 -4162 -1410 2 VDD
port 41 nsew
rlabel metal1 s 21202 -1247 21248 -1047 8 VDD
port 41 nsew
rlabel metal1 s 21006 -1247 21052 -1047 8 VDD
port 41 nsew
rlabel metal1 s 20810 -1247 20856 -1047 8 VDD
port 41 nsew
rlabel metal1 s 14923 -899 14969 -499 8 VDD
port 41 nsew
rlabel metal1 s 14687 -899 14733 -499 8 VDD
port 41 nsew
rlabel metal1 s 14451 -899 14497 -499 8 VDD
port 41 nsew
rlabel metal1 s 14215 -899 14261 -499 8 VDD
port 41 nsew
rlabel metal1 s 13979 -899 14025 -499 8 VDD
port 41 nsew
rlabel metal1 s 13743 -899 13789 -499 8 VDD
port 41 nsew
rlabel metal1 s 13507 -899 13553 -499 8 VDD
port 41 nsew
rlabel metal1 s 13271 -899 13317 -499 8 VDD
port 41 nsew
rlabel metal1 s 13035 -899 13081 -499 8 VDD
port 41 nsew
rlabel metal1 s 12799 -899 12845 -499 8 VDD
port 41 nsew
rlabel metal1 s 12563 -899 12609 -499 8 VDD
port 41 nsew
rlabel metal1 s 12327 -899 12373 -499 8 VDD
port 41 nsew
rlabel metal1 s 12091 -899 12137 -499 8 VDD
port 41 nsew
rlabel metal1 s 11855 -899 11901 -499 8 VDD
port 41 nsew
rlabel metal1 s 11619 -899 11665 -499 8 VDD
port 41 nsew
rlabel metal1 s 11383 -899 11429 -499 8 VDD
port 41 nsew
rlabel metal1 s 11135 -899 11181 -499 8 VDD
port 41 nsew
rlabel metal1 s 10899 -899 10945 -499 8 VDD
port 41 nsew
rlabel metal1 s 10663 -899 10709 -499 8 VDD
port 41 nsew
rlabel metal1 s 10427 -899 10473 -499 8 VDD
port 41 nsew
rlabel metal1 s 10191 -899 10237 -499 8 VDD
port 41 nsew
rlabel metal1 s 9955 -899 10001 -499 8 VDD
port 41 nsew
rlabel metal1 s 9719 -899 9765 -499 8 VDD
port 41 nsew
rlabel metal1 s 9483 -899 9529 -499 8 VDD
port 41 nsew
rlabel metal1 s 9247 -899 9293 -499 8 VDD
port 41 nsew
rlabel metal1 s 9117 -899 9163 -499 8 VDD
port 41 nsew
rlabel metal1 s 8881 -899 8927 -499 8 VDD
port 41 nsew
rlabel metal1 s 8645 -899 8691 -499 8 VDD
port 41 nsew
rlabel metal1 s 8409 -899 8455 -499 8 VDD
port 41 nsew
rlabel metal1 s 8173 -899 8219 -499 8 VDD
port 41 nsew
rlabel metal1 s 8043 -899 8089 -499 8 VDD
port 41 nsew
rlabel metal1 s 7807 -899 7853 -499 8 VDD
port 41 nsew
rlabel metal1 s 7571 -899 7617 -499 8 VDD
port 41 nsew
rlabel metal1 s 5766 -677 5812 -477 8 VDD
port 41 nsew
rlabel metal1 s 5570 -677 5616 -477 8 VDD
port 41 nsew
rlabel metal1 s 5374 -677 5420 -477 8 VDD
port 41 nsew
rlabel metal1 s 4916 -677 4962 -477 8 VDD
port 41 nsew
rlabel metal1 s 4720 -677 4766 -477 8 VDD
port 41 nsew
rlabel metal1 s 4524 -677 4570 -477 8 VDD
port 41 nsew
rlabel metal1 s 27390 -386 31946 -306 8 VDD
port 41 nsew
rlabel metal1 s -3816 -535 -3770 -335 2 VDD
port 41 nsew
rlabel metal1 s -4012 -535 -3966 -335 2 VDD
port 41 nsew
rlabel metal1 s -4208 -535 -4162 -335 2 VDD
port 41 nsew
rlabel metal1 s -4666 -535 -4620 -335 2 VDD
port 41 nsew
rlabel metal1 s -4862 -535 -4816 -335 2 VDD
port 41 nsew
rlabel metal1 s -5058 -535 -5012 -335 2 VDD
port 41 nsew
rlabel metal1 s 58039 -277 58085 123 8 VDD
port 41 nsew
rlabel metal1 s 57803 -277 57849 123 8 VDD
port 41 nsew
rlabel metal1 s 57567 -277 57613 123 8 VDD
port 41 nsew
rlabel metal1 s 57331 -277 57377 123 8 VDD
port 41 nsew
rlabel metal1 s 57095 -277 57141 123 8 VDD
port 41 nsew
rlabel metal1 s 56859 -277 56905 123 8 VDD
port 41 nsew
rlabel metal1 s 56623 -277 56669 123 8 VDD
port 41 nsew
rlabel metal1 s 56387 -277 56433 123 8 VDD
port 41 nsew
rlabel metal1 s 56151 -277 56197 123 8 VDD
port 41 nsew
rlabel metal1 s 55915 -277 55961 123 8 VDD
port 41 nsew
rlabel metal1 s 55679 -277 55725 123 8 VDD
port 41 nsew
rlabel metal1 s 55443 -277 55489 123 8 VDD
port 41 nsew
rlabel metal1 s 55207 -277 55253 123 8 VDD
port 41 nsew
rlabel metal1 s 54971 -277 55017 123 8 VDD
port 41 nsew
rlabel metal1 s 54735 -277 54781 123 8 VDD
port 41 nsew
rlabel metal1 s 54499 -277 54545 123 8 VDD
port 41 nsew
rlabel metal1 s 54251 -277 54297 123 8 VDD
port 41 nsew
rlabel metal1 s 54015 -277 54061 123 8 VDD
port 41 nsew
rlabel metal1 s 53779 -277 53825 123 8 VDD
port 41 nsew
rlabel metal1 s 53543 -277 53589 123 8 VDD
port 41 nsew
rlabel metal1 s 53307 -277 53353 123 8 VDD
port 41 nsew
rlabel metal1 s 53071 -277 53117 123 8 VDD
port 41 nsew
rlabel metal1 s 52835 -277 52881 123 8 VDD
port 41 nsew
rlabel metal1 s 52599 -277 52645 123 8 VDD
port 41 nsew
rlabel metal1 s 52363 -277 52409 123 8 VDD
port 41 nsew
rlabel metal1 s 52233 -277 52279 123 8 VDD
port 41 nsew
rlabel metal1 s 51997 -277 52043 123 8 VDD
port 41 nsew
rlabel metal1 s 51761 -277 51807 123 8 VDD
port 41 nsew
rlabel metal1 s 51525 -277 51571 123 8 VDD
port 41 nsew
rlabel metal1 s 51289 -277 51335 123 8 VDD
port 41 nsew
rlabel metal1 s 51159 -277 51205 123 8 VDD
port 41 nsew
rlabel metal1 s 50923 -277 50969 123 8 VDD
port 41 nsew
rlabel metal1 s 50687 -277 50733 123 8 VDD
port 41 nsew
rlabel metal1 s 31866 -306 31946 -152 8 VDD
port 41 nsew
rlabel metal1 s 31866 -152 32623 -72 8 VDD
port 41 nsew
rlabel metal1 s 27390 -306 27470 -149 8 VDD
port 41 nsew
rlabel metal1 s 26988 -166 27304 -149 8 VDD
port 41 nsew
rlabel metal1 s 26988 -149 27767 -69 8 VDD
port 41 nsew
rlabel metal1 s 26988 -69 27304 -38 8 VDD
port 41 nsew
rlabel metal1 s 38044 506 38090 906 6 VDD
port 41 nsew
rlabel metal1 s 37728 506 37774 906 6 VDD
port 41 nsew
rlabel metal1 s 37412 506 37458 906 6 VDD
port 41 nsew
rlabel metal1 s 37096 506 37142 906 6 VDD
port 41 nsew
rlabel metal1 s 36780 506 36826 906 6 VDD
port 41 nsew
rlabel metal1 s 36323 463 36369 863 6 VDD
port 41 nsew
rlabel metal1 s 36007 463 36053 863 6 VDD
port 41 nsew
rlabel metal1 s 35691 463 35737 863 6 VDD
port 41 nsew
rlabel metal1 s 35375 463 35421 863 6 VDD
port 41 nsew
rlabel metal1 s 35059 463 35105 924 6 VDD
port 41 nsew
rlabel metal1 s 31588 440 31634 840 6 VDD
port 41 nsew
rlabel metal1 s 31272 440 31318 840 6 VDD
port 41 nsew
rlabel metal1 s 30956 440 31002 840 6 VDD
port 41 nsew
rlabel metal1 s 30640 440 30686 840 6 VDD
port 41 nsew
rlabel metal1 s 30324 440 30370 840 6 VDD
port 41 nsew
rlabel metal1 s 27052 -38 27180 518 6 VDD
port 41 nsew
rlabel metal1 s 21202 -172 21248 28 8 VDD
port 41 nsew
rlabel metal1 s 21006 -172 21052 28 8 VDD
port 41 nsew
rlabel metal1 s 20810 -172 20856 28 8 VDD
port 41 nsew
rlabel metal1 s 20352 -172 20398 28 8 VDD
port 41 nsew
rlabel metal1 s 20156 -172 20202 28 8 VDD
port 41 nsew
rlabel metal1 s 19960 -172 20006 28 8 VDD
port 41 nsew
rlabel metal1 s 26762 518 27180 646 6 VDD
port 41 nsew
rlabel metal1 s 34550 924 35105 970 6 VDD
port 41 nsew
rlabel metal1 s 45965 1507 46011 1707 6 VDD
port 41 nsew
rlabel metal1 s 45769 1507 45815 1707 6 VDD
port 41 nsew
rlabel metal1 s 45573 1507 45619 1707 6 VDD
port 41 nsew
rlabel metal1 s 44995 1417 45041 1617 6 VDD
port 41 nsew
rlabel metal1 s 44799 1417 44845 1617 6 VDD
port 41 nsew
rlabel metal1 s 44603 1417 44649 1617 6 VDD
port 41 nsew
rlabel metal1 s 44158 1417 44204 1617 6 VDD
port 41 nsew
rlabel metal1 s 43962 1417 44008 1617 6 VDD
port 41 nsew
rlabel metal1 s 43766 1417 43812 1617 6 VDD
port 41 nsew
rlabel metal1 s 42295 1417 42341 1617 6 VDD
port 41 nsew
rlabel metal1 s 42099 1417 42145 1617 6 VDD
port 41 nsew
rlabel metal1 s 41903 1417 41949 1617 6 VDD
port 41 nsew
rlabel metal1 s 41458 1417 41504 1617 6 VDD
port 41 nsew
rlabel metal1 s 41262 1417 41308 1617 6 VDD
port 41 nsew
rlabel metal1 s 41066 1417 41112 1617 6 VDD
port 41 nsew
rlabel metal1 s 38044 1419 38090 1819 6 VDD
port 41 nsew
rlabel metal1 s 37728 1419 37774 1819 6 VDD
port 41 nsew
rlabel metal1 s 37412 1419 37458 1819 6 VDD
port 41 nsew
rlabel metal1 s 37096 1419 37142 1819 6 VDD
port 41 nsew
rlabel metal1 s 36780 1419 36826 1819 6 VDD
port 41 nsew
rlabel metal1 s 36323 1462 36369 1862 6 VDD
port 41 nsew
rlabel metal1 s 36007 1462 36053 1862 6 VDD
port 41 nsew
rlabel metal1 s 35691 1462 35737 1862 6 VDD
port 41 nsew
rlabel metal1 s 35375 1462 35421 1862 6 VDD
port 41 nsew
rlabel metal1 s 35059 1462 35105 1862 6 VDD
port 41 nsew
rlabel metal1 s 34550 970 34596 1747 6 VDD
port 41 nsew
rlabel metal1 s 31588 1371 32616 1417 6 VDD
port 41 nsew
rlabel metal1 s 34324 1460 34370 1747 6 VDD
port 41 nsew
rlabel metal1 s 34166 1460 34212 1747 6 VDD
port 41 nsew
rlabel metal1 s 34141 1747 34596 1793 6 VDD
port 41 nsew
rlabel metal1 s 34550 1793 34596 1841 6 VDD
port 41 nsew
rlabel metal1 s 34320 1793 34366 2055 6 VDD
port 41 nsew
rlabel metal1 s 34162 1793 34208 2055 6 VDD
port 41 nsew
rlabel metal1 s 33878 1461 33924 2055 6 VDD
port 41 nsew
rlabel metal1 s 33432 1461 33478 2050 6 VDD
port 41 nsew
rlabel metal1 s 33116 1461 33162 2050 6 VDD
port 41 nsew
rlabel metal1 s 32728 1461 32774 1661 6 VDD
port 41 nsew
rlabel metal1 s 32570 1417 32616 1661 6 VDD
port 41 nsew
rlabel metal1 s 32728 1784 32774 1984 6 VDD
port 41 nsew
rlabel metal1 s 32570 1784 32616 1984 6 VDD
port 41 nsew
rlabel metal1 s 31588 1417 31634 1840 6 VDD
port 41 nsew
rlabel metal1 s 30083 1365 30370 1411 6 VDD
port 41 nsew
rlabel metal1 s 31272 1440 31318 1840 6 VDD
port 41 nsew
rlabel metal1 s 30956 1440 31002 1840 6 VDD
port 41 nsew
rlabel metal1 s 30640 1440 30686 1840 6 VDD
port 41 nsew
rlabel metal1 s 30324 1411 30370 1840 6 VDD
port 41 nsew
rlabel metal1 s 30083 1411 30129 1717 6 VDD
port 41 nsew
rlabel metal1 s 29469 1467 29515 1717 6 VDD
port 41 nsew
rlabel metal1 s 29469 1717 30129 1754 6 VDD
port 41 nsew
rlabel metal1 s 29311 1467 29357 1754 6 VDD
port 41 nsew
rlabel metal1 s 29286 1754 30129 1763 6 VDD
port 41 nsew
rlabel metal1 s 29286 1763 29546 1800 6 VDD
port 41 nsew
rlabel metal1 s 29465 1800 29511 2062 6 VDD
port 41 nsew
rlabel metal1 s 29307 1800 29353 2062 6 VDD
port 41 nsew
rlabel metal1 s 29023 1468 29069 2062 6 VDD
port 41 nsew
rlabel metal1 s 28577 1468 28623 2057 6 VDD
port 41 nsew
rlabel metal1 s 28261 1468 28307 2057 6 VDD
port 41 nsew
rlabel metal1 s 27873 1468 27919 1668 6 VDD
port 41 nsew
rlabel metal1 s 27715 1468 27761 1668 6 VDD
port 41 nsew
rlabel metal1 s 27873 1791 27919 1991 6 VDD
port 41 nsew
rlabel metal1 s 27715 1791 27761 1991 6 VDD
port 41 nsew
rlabel metal1 s 58242 2634 58288 3034 6 VDD
port 41 nsew
rlabel metal1 s 58006 2634 58052 3034 6 VDD
port 41 nsew
rlabel metal1 s 57770 2634 57816 3034 6 VDD
port 41 nsew
rlabel metal1 s 57534 2634 57580 3034 6 VDD
port 41 nsew
rlabel metal1 s 57298 2634 57344 3034 6 VDD
port 41 nsew
rlabel metal1 s 57062 2634 57108 3034 6 VDD
port 41 nsew
rlabel metal1 s 56826 2634 56872 3034 6 VDD
port 41 nsew
rlabel metal1 s 56590 2634 56636 3034 6 VDD
port 41 nsew
rlabel metal1 s 56354 2634 56400 3034 6 VDD
port 41 nsew
rlabel metal1 s 56118 2634 56164 3034 6 VDD
port 41 nsew
rlabel metal1 s 55882 2634 55928 3034 6 VDD
port 41 nsew
rlabel metal1 s 55646 2634 55692 3034 6 VDD
port 41 nsew
rlabel metal1 s 55410 2634 55456 3034 6 VDD
port 41 nsew
rlabel metal1 s 55174 2634 55220 3034 6 VDD
port 41 nsew
rlabel metal1 s 54938 2634 54984 3034 6 VDD
port 41 nsew
rlabel metal1 s 54702 2634 54748 3034 6 VDD
port 41 nsew
rlabel metal1 s 54454 2634 54500 3034 6 VDD
port 41 nsew
rlabel metal1 s 54218 2634 54264 3034 6 VDD
port 41 nsew
rlabel metal1 s 53982 2634 54028 3034 6 VDD
port 41 nsew
rlabel metal1 s 53746 2634 53792 3034 6 VDD
port 41 nsew
rlabel metal1 s 53510 2634 53556 3034 6 VDD
port 41 nsew
rlabel metal1 s 53274 2634 53320 3034 6 VDD
port 41 nsew
rlabel metal1 s 53038 2634 53084 3034 6 VDD
port 41 nsew
rlabel metal1 s 52802 2634 52848 3034 6 VDD
port 41 nsew
rlabel metal1 s 52566 2634 52612 3034 6 VDD
port 41 nsew
rlabel metal1 s 52436 2634 52482 3034 6 VDD
port 41 nsew
rlabel metal1 s 52200 2634 52246 3034 6 VDD
port 41 nsew
rlabel metal1 s 51964 2634 52010 3034 6 VDD
port 41 nsew
rlabel metal1 s 51728 2634 51774 3034 6 VDD
port 41 nsew
rlabel metal1 s 51492 2634 51538 3034 6 VDD
port 41 nsew
rlabel metal1 s 51362 2634 51408 3034 6 VDD
port 41 nsew
rlabel metal1 s 51126 2634 51172 3034 6 VDD
port 41 nsew
rlabel metal1 s 50890 2634 50936 3034 6 VDD
port 41 nsew
rlabel metal1 s 26762 646 26890 2653 6 VDD
port 41 nsew
rlabel metal1 s 21030 2103 21076 2303 6 VDD
port 41 nsew
rlabel metal1 s 20834 2103 20880 2303 6 VDD
port 41 nsew
rlabel metal1 s 20638 2103 20684 2303 6 VDD
port 41 nsew
rlabel metal1 s 44897 2735 44943 2935 6 VDD
port 41 nsew
rlabel metal1 s 44701 2735 44747 2935 6 VDD
port 41 nsew
rlabel metal1 s 44505 2735 44551 2935 6 VDD
port 41 nsew
rlabel metal1 s 43154 2735 43200 2935 6 VDD
port 41 nsew
rlabel metal1 s 42958 2735 43004 2935 6 VDD
port 41 nsew
rlabel metal1 s 42762 2735 42808 2935 6 VDD
port 41 nsew
rlabel metal1 s 42197 2735 42243 2935 6 VDD
port 41 nsew
rlabel metal1 s 42001 2735 42047 2935 6 VDD
port 41 nsew
rlabel metal1 s 41805 2735 41851 2935 6 VDD
port 41 nsew
rlabel metal1 s 40454 2735 40500 2935 6 VDD
port 41 nsew
rlabel metal1 s 40258 2735 40304 2935 6 VDD
port 41 nsew
rlabel metal1 s 40062 2735 40108 2935 6 VDD
port 41 nsew
rlabel metal1 s 39572 2735 39618 2935 6 VDD
port 41 nsew
rlabel metal1 s 39376 2735 39422 2935 6 VDD
port 41 nsew
rlabel metal1 s 39180 2735 39226 2935 6 VDD
port 41 nsew
rlabel metal1 s 26688 2653 26963 2876 6 VDD
port 41 nsew
rlabel metal1 s 41827 3129 44196 3233 6 VDD
port 41 nsew
rlabel metal1 s 43752 3233 44082 4185 6 VDD
port 41 nsew
rlabel metal1 s 43243 3233 43573 4185 6 VDD
port 41 nsew
rlabel metal1 s 42554 3233 42884 4185 6 VDD
port 41 nsew
rlabel metal1 s 41865 3233 42195 4185 6 VDD
port 41 nsew
rlabel metal1 s 21030 3178 21076 3378 6 VDD
port 41 nsew
rlabel metal1 s 20834 3178 20880 3378 6 VDD
port 41 nsew
rlabel metal1 s 20638 3178 20684 3378 6 VDD
port 41 nsew
rlabel metal1 s 20180 3178 20226 3378 6 VDD
port 41 nsew
rlabel metal1 s 19984 3178 20030 3378 6 VDD
port 41 nsew
rlabel metal1 s 19788 3178 19834 3378 6 VDD
port 41 nsew
rlabel metal1 s 15814 -255 16329 3722 6 VDD
port 41 nsew
rlabel metal1 s 5891 -122 6236 223 6 VDD
port 41 nsew
rlabel metal1 s 5943 223 6135 686 6 VDD
port 41 nsew
rlabel metal1 s 5730 686 6208 775 6 VDD
port 41 nsew
rlabel metal1 s 5751 938 5797 1138 6 VDD
port 41 nsew
rlabel metal1 s 5555 938 5601 1138 6 VDD
port 41 nsew
rlabel metal1 s 5359 938 5405 1138 6 VDD
port 41 nsew
rlabel metal1 s -2348 762 -2302 962 4 VDD
port 41 nsew
rlabel metal1 s -2544 762 -2498 962 4 VDD
port 41 nsew
rlabel metal1 s -2740 762 -2694 962 4 VDD
port 41 nsew
rlabel metal1 s 2803 1041 2849 1209 6 VDD
port 41 nsew
rlabel metal1 s 2494 1041 2540 1209 6 VDD
port 41 nsew
rlabel metal1 s 1830 1043 1876 1223 6 VDD
port 41 nsew
rlabel metal1 s 1684 1043 1730 1223 6 VDD
port 41 nsew
rlabel metal1 s 1395 1043 1441 1163 6 VDD
port 41 nsew
rlabel metal1 s 1219 1043 1265 1163 6 VDD
port 41 nsew
rlabel metal1 s 1043 1043 1089 1163 6 VDD
port 41 nsew
rlabel metal1 s 707 1041 753 1209 6 VDD
port 41 nsew
rlabel metal1 s 14964 1857 15010 2257 6 VDD
port 41 nsew
rlabel metal1 s 14728 1857 14774 2257 6 VDD
port 41 nsew
rlabel metal1 s 14492 1857 14538 2257 6 VDD
port 41 nsew
rlabel metal1 s 14256 1857 14302 2257 6 VDD
port 41 nsew
rlabel metal1 s 14020 1857 14066 2257 6 VDD
port 41 nsew
rlabel metal1 s 13784 1857 13830 2257 6 VDD
port 41 nsew
rlabel metal1 s 13548 1857 13594 2257 6 VDD
port 41 nsew
rlabel metal1 s 13312 1857 13358 2257 6 VDD
port 41 nsew
rlabel metal1 s 13076 1857 13122 2257 6 VDD
port 41 nsew
rlabel metal1 s 12840 1857 12886 2257 6 VDD
port 41 nsew
rlabel metal1 s 12604 1857 12650 2257 6 VDD
port 41 nsew
rlabel metal1 s 12368 1857 12414 2257 6 VDD
port 41 nsew
rlabel metal1 s 12132 1857 12178 2257 6 VDD
port 41 nsew
rlabel metal1 s 11896 1857 11942 2257 6 VDD
port 41 nsew
rlabel metal1 s 11660 1857 11706 2257 6 VDD
port 41 nsew
rlabel metal1 s 11424 1857 11470 2257 6 VDD
port 41 nsew
rlabel metal1 s 11176 1857 11222 2257 6 VDD
port 41 nsew
rlabel metal1 s 10940 1857 10986 2257 6 VDD
port 41 nsew
rlabel metal1 s 10704 1857 10750 2257 6 VDD
port 41 nsew
rlabel metal1 s 10468 1857 10514 2257 6 VDD
port 41 nsew
rlabel metal1 s 10232 1857 10278 2257 6 VDD
port 41 nsew
rlabel metal1 s 9996 1857 10042 2257 6 VDD
port 41 nsew
rlabel metal1 s 9760 1857 9806 2257 6 VDD
port 41 nsew
rlabel metal1 s 9524 1857 9570 2257 6 VDD
port 41 nsew
rlabel metal1 s 9288 1857 9334 2257 6 VDD
port 41 nsew
rlabel metal1 s 9158 1857 9204 2257 6 VDD
port 41 nsew
rlabel metal1 s 8922 1857 8968 2257 6 VDD
port 41 nsew
rlabel metal1 s 8686 1857 8732 2257 6 VDD
port 41 nsew
rlabel metal1 s 8450 1857 8496 2257 6 VDD
port 41 nsew
rlabel metal1 s 8214 1857 8260 2257 6 VDD
port 41 nsew
rlabel metal1 s 8084 1857 8130 2257 6 VDD
port 41 nsew
rlabel metal1 s 7848 1857 7894 2257 6 VDD
port 41 nsew
rlabel metal1 s 7612 1857 7658 2257 6 VDD
port 41 nsew
rlabel metal1 s 5751 2013 5797 2213 6 VDD
port 41 nsew
rlabel metal1 s 5555 2013 5601 2213 6 VDD
port 41 nsew
rlabel metal1 s 5359 2013 5405 2213 6 VDD
port 41 nsew
rlabel metal1 s 4901 2013 4947 2213 6 VDD
port 41 nsew
rlabel metal1 s 4705 2013 4751 2213 6 VDD
port 41 nsew
rlabel metal1 s 4509 2013 4555 2213 6 VDD
port 41 nsew
rlabel metal1 s 15814 3722 16331 4171 6 VDD
port 41 nsew
rlabel metal1 s 41672 4185 44640 4844 6 VDD
port 41 nsew
rlabel metal1 s 12616 6696 12662 7496 6 VDD
port 41 nsew
rlabel metal1 s 11700 6696 11746 7496 6 VDD
port 41 nsew
rlabel metal1 s 11570 6696 11616 7496 6 VDD
port 41 nsew
rlabel metal1 s 9854 6696 9900 7496 6 VDD
port 41 nsew
rlabel metal1 s 8138 6696 8184 7496 6 VDD
port 41 nsew
rlabel metal1 s 3500 1279 3875 7565 6 VDD
port 41 nsew
rlabel metal1 s 2803 1653 2849 1821 6 VDD
port 41 nsew
rlabel metal1 s 2494 1653 2540 1821 6 VDD
port 41 nsew
rlabel metal1 s 1830 1639 1876 1819 6 VDD
port 41 nsew
rlabel metal1 s 1684 1639 1730 1819 6 VDD
port 41 nsew
rlabel metal1 s 1395 1699 1441 1819 6 VDD
port 41 nsew
rlabel metal1 s 1219 1699 1265 1819 6 VDD
port 41 nsew
rlabel metal1 s 1043 1699 1089 1819 6 VDD
port 41 nsew
rlabel metal1 s 707 1653 753 1821 6 VDD
port 41 nsew
rlabel metal1 s -2348 1837 -2302 2037 4 VDD
port 41 nsew
rlabel metal1 s -2544 1837 -2498 2037 4 VDD
port 41 nsew
rlabel metal1 s -2740 1837 -2694 2037 4 VDD
port 41 nsew
rlabel metal1 s -3198 1837 -3152 2037 4 VDD
port 41 nsew
rlabel metal1 s -3394 1837 -3348 2037 4 VDD
port 41 nsew
rlabel metal1 s -3590 1837 -3544 2037 4 VDD
port 41 nsew
rlabel metal1 s -5945 1575 -5899 1975 4 VDD
port 41 nsew
rlabel metal1 s -6181 1575 -6135 1975 4 VDD
port 41 nsew
rlabel metal1 s -6417 1575 -6371 1975 4 VDD
port 41 nsew
rlabel metal1 s -6547 1575 -6501 1975 4 VDD
port 41 nsew
rlabel metal1 s -6783 1575 -6737 1975 4 VDD
port 41 nsew
rlabel metal1 s -7019 1575 -6973 1975 4 VDD
port 41 nsew
rlabel metal1 s -7255 1575 -7209 1975 4 VDD
port 41 nsew
rlabel metal1 s -7491 1575 -7445 1975 4 VDD
port 41 nsew
rlabel metal1 s -7621 1575 -7575 1975 4 VDD
port 41 nsew
rlabel metal1 s -7857 1575 -7811 1975 4 VDD
port 41 nsew
rlabel metal1 s -8093 1575 -8047 1975 4 VDD
port 41 nsew
rlabel metal1 s -8329 1575 -8283 1975 4 VDD
port 41 nsew
rlabel metal1 s -8565 1575 -8519 1975 4 VDD
port 41 nsew
rlabel metal1 s -8801 1575 -8755 1975 4 VDD
port 41 nsew
rlabel metal1 s -9037 1575 -8991 1975 4 VDD
port 41 nsew
rlabel metal1 s -9273 1575 -9227 1975 4 VDD
port 41 nsew
rlabel metal1 s -9509 1575 -9463 1975 4 VDD
port 41 nsew
rlabel metal1 s -9757 1575 -9711 1975 4 VDD
port 41 nsew
rlabel metal1 s -9993 1575 -9947 1975 4 VDD
port 41 nsew
rlabel metal1 s -10229 1575 -10183 1975 4 VDD
port 41 nsew
rlabel metal1 s -10465 1575 -10419 1975 4 VDD
port 41 nsew
rlabel metal1 s -10701 1575 -10655 1975 4 VDD
port 41 nsew
rlabel metal1 s -10937 1575 -10891 1975 4 VDD
port 41 nsew
rlabel metal1 s -11173 1575 -11127 1975 4 VDD
port 41 nsew
rlabel metal1 s -11409 1575 -11363 1975 4 VDD
port 41 nsew
rlabel metal1 s -11645 1575 -11599 1975 4 VDD
port 41 nsew
rlabel metal1 s -11881 1575 -11835 1975 4 VDD
port 41 nsew
rlabel metal1 s -12117 1575 -12071 1975 4 VDD
port 41 nsew
rlabel metal1 s -12353 1575 -12307 1975 4 VDD
port 41 nsew
rlabel metal1 s -12589 1575 -12543 1975 4 VDD
port 41 nsew
rlabel metal1 s -12825 1575 -12779 1975 4 VDD
port 41 nsew
rlabel metal1 s -13061 1575 -13015 1975 4 VDD
port 41 nsew
rlabel metal1 s -13297 1575 -13251 1975 4 VDD
port 41 nsew
rlabel metal1 s -13395 2124 -9226 2361 4 VDD
port 41 nsew
rlabel metal1 s -9633 2361 -9285 3329 4 VDD
port 41 nsew
rlabel metal1 s -10239 2361 -9891 3329 4 VDD
port 41 nsew
rlabel metal1 s -11015 2361 -10667 3329 4 VDD
port 41 nsew
rlabel metal1 s -11909 2361 -11561 3329 4 VDD
port 41 nsew
rlabel metal1 s -13011 2361 -12663 3329 4 VDD
port 41 nsew
rlabel metal1 s -13122 3329 -8953 3566 4 VDD
port 41 nsew
rlabel metal1 s 3375 7565 4103 8200 6 VDD
port 41 nsew
rlabel metal1 s 15726 8966 15886 9012 6 VDD
port 41 nsew
rlabel metal1 s 15588 9095 15788 9141 6 VDD
port 41 nsew
rlabel metal1 s 14785 9353 14985 9399 6 VDD
port 41 nsew
rlabel metal1 s 15588 9611 15788 9657 6 VDD
port 41 nsew
rlabel metal1 s 14785 9869 14985 9915 6 VDD
port 41 nsew
rlabel metal1 s 15588 10127 15788 10173 6 VDD
port 41 nsew
rlabel metal1 s -3582 5554 -2367 39356 4 VDD
port 41 nsew
rlabel metal1 s -12975 3566 -11404 6943 4 VDD
port 41 nsew
rlabel metal1 s -13896 10354 -13696 10400 4 VDD
port 41 nsew
rlabel metal1 s -5853 10569 -5653 10615 4 VDD
port 41 nsew
rlabel metal1 s -13896 10550 -13696 10596 4 VDD
port 41 nsew
rlabel metal1 s -7984 10626 -7684 10672 4 VDD
port 41 nsew
rlabel metal1 s -11478 10691 -10878 10737 4 VDD
port 41 nsew
rlabel metal1 s -5853 10765 -5653 10811 4 VDD
port 41 nsew
rlabel metal1 s -7984 10822 -7684 10868 4 VDD
port 41 nsew
rlabel metal1 s -11478 10887 -10878 10933 4 VDD
port 41 nsew
rlabel metal1 s -5853 10961 -5653 11007 4 VDD
port 41 nsew
rlabel metal1 s -7984 11018 -7684 11064 4 VDD
port 41 nsew
rlabel metal1 s -13896 11092 -13696 11138 4 VDD
port 41 nsew
rlabel metal1 s -5853 11157 -5653 11203 4 VDD
port 41 nsew
rlabel metal1 s -7783 11235 -7683 11281 4 VDD
port 41 nsew
rlabel metal1 s -13896 11288 -13696 11334 4 VDD
port 41 nsew
rlabel metal1 s -7783 11431 -7683 11477 4 VDD
port 41 nsew
rlabel metal1 s -13896 11484 -13696 11530 4 VDD
port 41 nsew
rlabel metal1 s -7783 11627 -7683 11673 4 VDD
port 41 nsew
rlabel metal1 s -5853 11699 -5653 11745 4 VDD
port 41 nsew
rlabel metal1 s -13896 11680 -13696 11726 4 VDD
port 41 nsew
rlabel metal1 s -7783 11823 -7683 11869 4 VDD
port 41 nsew
rlabel metal1 s -5853 11895 -5653 11941 4 VDD
port 41 nsew
rlabel metal1 s -11207 11897 -10807 11943 4 VDD
port 41 nsew
rlabel metal1 s -11207 12093 -10807 12139 4 VDD
port 41 nsew
rlabel metal1 s -7789 12399 -7589 12445 4 VDD
port 41 nsew
rlabel metal1 s -6075 12568 -5775 12614 4 VDD
port 41 nsew
rlabel metal1 s -7789 12595 -7589 12641 4 VDD
port 41 nsew
rlabel metal1 s -6075 12764 -5775 12810 4 VDD
port 41 nsew
rlabel metal1 s -7789 12791 -7589 12837 4 VDD
port 41 nsew
rlabel metal1 s -11208 12802 -10808 12848 4 VDD
port 41 nsew
rlabel metal1 s -6075 12960 -5775 13006 4 VDD
port 41 nsew
rlabel metal1 s -7789 12987 -7589 13033 4 VDD
port 41 nsew
rlabel metal1 s -11208 12998 -10808 13044 4 VDD
port 41 nsew
rlabel metal1 s -14060 12964 -13429 13140 4 VDD
port 41 nsew
rlabel metal1 s -5874 13177 -5774 13223 4 VDD
port 41 nsew
rlabel metal1 s -5874 13373 -5774 13419 4 VDD
port 41 nsew
rlabel metal1 s -5874 13569 -5774 13615 4 VDD
port 41 nsew
rlabel metal1 s -7789 13529 -7589 13575 4 VDD
port 41 nsew
rlabel metal1 s -5874 13765 -5774 13811 4 VDD
port 41 nsew
rlabel metal1 s -7789 13725 -7589 13771 4 VDD
port 41 nsew
rlabel metal1 s -10498 13743 -10331 13770 4 VDD
port 41 nsew
rlabel metal1 s -12434 13769 -12262 13770 4 VDD
port 41 nsew
rlabel metal1 s -12434 13770 -10331 13896 4 VDD
port 41 nsew
rlabel metal1 s -10498 13896 -10331 13922 4 VDD
port 41 nsew
rlabel metal1 s -12434 13896 -12262 13961 4 VDD
port 41 nsew
rlabel metal1 s -7037 14204 -6737 14250 4 VDD
port 41 nsew
rlabel metal1 s -7966 14230 -7766 14276 4 VDD
port 41 nsew
rlabel metal1 s -12037 14204 -11737 14250 4 VDD
port 41 nsew
rlabel metal1 s -12966 14230 -12766 14276 4 VDD
port 41 nsew
rlabel metal1 s -7037 14400 -6737 14446 4 VDD
port 41 nsew
rlabel metal1 s -7966 14426 -7766 14472 4 VDD
port 41 nsew
rlabel metal1 s -12037 14400 -11737 14446 4 VDD
port 41 nsew
rlabel metal1 s -12966 14426 -12766 14472 4 VDD
port 41 nsew
rlabel metal1 s -7037 14596 -6737 14642 4 VDD
port 41 nsew
rlabel metal1 s -7966 14622 -7766 14668 4 VDD
port 41 nsew
rlabel metal1 s -12037 14596 -11737 14642 4 VDD
port 41 nsew
rlabel metal1 s -12966 14622 -12766 14668 4 VDD
port 41 nsew
rlabel metal1 s -7038 14813 -6938 14859 4 VDD
port 41 nsew
rlabel metal1 s -7966 14818 -7766 14864 4 VDD
port 41 nsew
rlabel metal1 s -12038 14813 -11938 14859 4 VDD
port 41 nsew
rlabel metal1 s -12966 14818 -12766 14864 4 VDD
port 41 nsew
rlabel metal1 s -7038 15009 -6938 15055 4 VDD
port 41 nsew
rlabel metal1 s -12038 15009 -11938 15055 4 VDD
port 41 nsew
rlabel metal1 s -7038 15205 -6938 15251 4 VDD
port 41 nsew
rlabel metal1 s -7937 15203 -7637 15249 4 VDD
port 41 nsew
rlabel metal1 s -12038 15205 -11938 15251 4 VDD
port 41 nsew
rlabel metal1 s -12937 15203 -12637 15249 4 VDD
port 41 nsew
rlabel metal1 s -7038 15401 -6938 15447 4 VDD
port 41 nsew
rlabel metal1 s -7937 15399 -7637 15445 4 VDD
port 41 nsew
rlabel metal1 s -12038 15401 -11938 15447 4 VDD
port 41 nsew
rlabel metal1 s -12937 15399 -12637 15445 4 VDD
port 41 nsew
rlabel metal1 s -7937 15595 -7637 15641 4 VDD
port 41 nsew
rlabel metal1 s -12937 15595 -12637 15641 4 VDD
port 41 nsew
rlabel metal1 s -7126 15651 -6526 15697 4 VDD
port 41 nsew
rlabel metal1 s -12126 15651 -11526 15697 4 VDD
port 41 nsew
rlabel metal1 s -7126 15847 -6526 15893 4 VDD
port 41 nsew
rlabel metal1 s -7736 15812 -7636 15858 4 VDD
port 41 nsew
rlabel metal1 s -12126 15847 -11526 15893 4 VDD
port 41 nsew
rlabel metal1 s -12736 15812 -12636 15858 4 VDD
port 41 nsew
rlabel metal1 s -7736 16008 -7636 16054 4 VDD
port 41 nsew
rlabel metal1 s -12736 16008 -12636 16054 4 VDD
port 41 nsew
rlabel metal1 s -7736 16204 -7636 16250 4 VDD
port 41 nsew
rlabel metal1 s -12736 16204 -12636 16250 4 VDD
port 41 nsew
rlabel metal1 s -7126 16270 -6526 16316 4 VDD
port 41 nsew
rlabel metal1 s -12126 16270 -11526 16316 4 VDD
port 41 nsew
rlabel metal1 s -7736 16400 -7636 16446 4 VDD
port 41 nsew
rlabel metal1 s -12736 16400 -12636 16446 4 VDD
port 41 nsew
rlabel metal1 s -5066 18168 -4866 18214 4 VDD
port 41 nsew
rlabel metal1 s -9993 18168 -9793 18214 4 VDD
port 41 nsew
rlabel metal1 s -6384 18266 -6184 18312 4 VDD
port 41 nsew
rlabel metal1 s -11311 18266 -11111 18312 4 VDD
port 41 nsew
rlabel metal1 s -5066 18364 -4866 18410 4 VDD
port 41 nsew
rlabel metal1 s -9993 18364 -9793 18410 4 VDD
port 41 nsew
rlabel metal1 s -6384 18462 -6184 18508 4 VDD
port 41 nsew
rlabel metal1 s -11311 18462 -11111 18508 4 VDD
port 41 nsew
rlabel metal1 s -5066 18560 -4866 18606 4 VDD
port 41 nsew
rlabel metal1 s -9993 18560 -9793 18606 4 VDD
port 41 nsew
rlabel metal1 s -6384 18658 -6184 18704 4 VDD
port 41 nsew
rlabel metal1 s -11311 18658 -11111 18704 4 VDD
port 41 nsew
rlabel metal1 s -5066 19005 -4866 19051 4 VDD
port 41 nsew
rlabel metal1 s -9993 19005 -9793 19051 4 VDD
port 41 nsew
rlabel metal1 s -5066 19201 -4866 19247 4 VDD
port 41 nsew
rlabel metal1 s -8013 19193 -7713 19239 4 VDD
port 41 nsew
rlabel metal1 s -8942 19219 -8742 19265 4 VDD
port 41 nsew
rlabel metal1 s -9993 19201 -9793 19247 4 VDD
port 41 nsew
rlabel metal1 s -5066 19397 -4866 19443 4 VDD
port 41 nsew
rlabel metal1 s -8013 19389 -7713 19435 4 VDD
port 41 nsew
rlabel metal1 s -8942 19415 -8742 19461 4 VDD
port 41 nsew
rlabel metal1 s -9993 19397 -9793 19443 4 VDD
port 41 nsew
rlabel metal1 s -8013 19585 -7713 19631 4 VDD
port 41 nsew
rlabel metal1 s -8942 19611 -8742 19657 4 VDD
port 41 nsew
rlabel metal1 s -8014 19802 -7914 19848 4 VDD
port 41 nsew
rlabel metal1 s -8942 19807 -8742 19853 4 VDD
port 41 nsew
rlabel metal1 s -6384 20009 -6184 20055 4 VDD
port 41 nsew
rlabel metal1 s -8014 19998 -7914 20044 4 VDD
port 41 nsew
rlabel metal1 s -11311 20009 -11111 20055 4 VDD
port 41 nsew
rlabel metal1 s -6384 20205 -6184 20251 4 VDD
port 41 nsew
rlabel metal1 s -8014 20194 -7914 20240 4 VDD
port 41 nsew
rlabel metal1 s -8913 20192 -8613 20238 4 VDD
port 41 nsew
rlabel metal1 s -11311 20205 -11111 20251 4 VDD
port 41 nsew
rlabel metal1 s -6384 20401 -6184 20447 4 VDD
port 41 nsew
rlabel metal1 s -8014 20390 -7914 20436 4 VDD
port 41 nsew
rlabel metal1 s -8913 20388 -8613 20434 4 VDD
port 41 nsew
rlabel metal1 s -11311 20401 -11111 20447 4 VDD
port 41 nsew
rlabel metal1 s -8913 20584 -8613 20630 4 VDD
port 41 nsew
rlabel metal1 s -8102 20640 -7502 20686 4 VDD
port 41 nsew
rlabel metal1 s -5066 20868 -4866 20914 4 VDD
port 41 nsew
rlabel metal1 s -8102 20836 -7502 20882 4 VDD
port 41 nsew
rlabel metal1 s -8712 20801 -8612 20847 4 VDD
port 41 nsew
rlabel metal1 s -9993 20868 -9793 20914 4 VDD
port 41 nsew
rlabel metal1 s -6384 20966 -6184 21012 4 VDD
port 41 nsew
rlabel metal1 s -8712 20997 -8612 21043 4 VDD
port 41 nsew
rlabel metal1 s -11311 20966 -11111 21012 4 VDD
port 41 nsew
rlabel metal1 s -5066 21064 -4866 21110 4 VDD
port 41 nsew
rlabel metal1 s -9993 21064 -9793 21110 4 VDD
port 41 nsew
rlabel metal1 s -6384 21162 -6184 21208 4 VDD
port 41 nsew
rlabel metal1 s -8712 21193 -8612 21239 4 VDD
port 41 nsew
rlabel metal1 s -11311 21162 -11111 21208 4 VDD
port 41 nsew
rlabel metal1 s -5066 21260 -4866 21306 4 VDD
port 41 nsew
rlabel metal1 s -8102 21259 -7502 21305 4 VDD
port 41 nsew
rlabel metal1 s -9993 21260 -9793 21306 4 VDD
port 41 nsew
rlabel metal1 s -6384 21358 -6184 21404 4 VDD
port 41 nsew
rlabel metal1 s -8712 21389 -8612 21435 4 VDD
port 41 nsew
rlabel metal1 s -11311 21358 -11111 21404 4 VDD
port 41 nsew
rlabel metal1 s -5066 21705 -4866 21751 4 VDD
port 41 nsew
rlabel metal1 s -9993 21705 -9793 21751 4 VDD
port 41 nsew
rlabel metal1 s -5066 21901 -4866 21947 4 VDD
port 41 nsew
rlabel metal1 s -9993 21901 -9793 21947 4 VDD
port 41 nsew
rlabel metal1 s -5066 22097 -4866 22143 4 VDD
port 41 nsew
rlabel metal1 s -9993 22097 -9793 22143 4 VDD
port 41 nsew
rlabel metal1 s -6384 22709 -6184 22755 4 VDD
port 41 nsew
rlabel metal1 s -11311 22709 -11111 22755 4 VDD
port 41 nsew
rlabel metal1 s -6384 22905 -6184 22951 4 VDD
port 41 nsew
rlabel metal1 s -11311 22905 -11111 22951 4 VDD
port 41 nsew
rlabel metal1 s -6384 23101 -6184 23147 4 VDD
port 41 nsew
rlabel metal1 s -11311 23101 -11111 23147 4 VDD
port 41 nsew
rlabel metal1 s -6384 23591 -6184 23637 4 VDD
port 41 nsew
rlabel metal1 s -11311 23591 -11111 23637 4 VDD
port 41 nsew
rlabel metal1 s -6384 23787 -6184 23833 4 VDD
port 41 nsew
rlabel metal1 s -11311 23787 -11111 23833 4 VDD
port 41 nsew
rlabel metal1 s -6384 23983 -6184 24029 4 VDD
port 41 nsew
rlabel metal1 s -11311 23983 -11111 24029 4 VDD
port 41 nsew
rlabel metal1 s -5476 24530 -4876 24576 4 VDD
port 41 nsew
rlabel metal1 s -10410 24557 -9810 24603 4 VDD
port 41 nsew
rlabel metal1 s -5476 24953 -4876 24999 4 VDD
port 41 nsew
rlabel metal1 s -10410 24980 -9810 25026 4 VDD
port 41 nsew
rlabel metal1 s -5476 25149 -4876 25195 4 VDD
port 41 nsew
rlabel metal1 s -10410 25176 -9810 25222 4 VDD
port 41 nsew
rlabel metal1 s -8822 26042 -8622 26088 4 VDD
port 41 nsew
rlabel metal1 s -10260 26042 -10060 26088 4 VDD
port 41 nsew
rlabel metal1 s -7504 26140 -7304 26186 4 VDD
port 41 nsew
rlabel metal1 s -11578 26140 -11378 26186 4 VDD
port 41 nsew
rlabel metal1 s -8822 26238 -8622 26284 4 VDD
port 41 nsew
rlabel metal1 s -10260 26238 -10060 26284 4 VDD
port 41 nsew
rlabel metal1 s -6601 26299 -6401 26345 4 VDD
port 41 nsew
rlabel metal1 s -7504 26336 -7304 26382 4 VDD
port 41 nsew
rlabel metal1 s -11578 26336 -11378 26382 4 VDD
port 41 nsew
rlabel metal1 s -8822 26434 -8622 26480 4 VDD
port 41 nsew
rlabel metal1 s -10260 26434 -10060 26480 4 VDD
port 41 nsew
rlabel metal1 s -6601 26495 -6401 26541 4 VDD
port 41 nsew
rlabel metal1 s -7504 26532 -7304 26578 4 VDD
port 41 nsew
rlabel metal1 s -11578 26532 -11378 26578 4 VDD
port 41 nsew
rlabel metal1 s -5272 26638 -5072 26684 4 VDD
port 41 nsew
rlabel metal1 s -13810 26638 -13610 26684 4 VDD
port 41 nsew
rlabel metal1 s -6601 26691 -6401 26737 4 VDD
port 41 nsew
rlabel metal1 s -5272 26834 -5072 26880 4 VDD
port 41 nsew
rlabel metal1 s -8822 26879 -8622 26925 4 VDD
port 41 nsew
rlabel metal1 s -10260 26879 -10060 26925 4 VDD
port 41 nsew
rlabel metal1 s -13810 26834 -13610 26880 4 VDD
port 41 nsew
rlabel metal1 s -5272 27030 -5072 27076 4 VDD
port 41 nsew
rlabel metal1 s -8822 27075 -8622 27121 4 VDD
port 41 nsew
rlabel metal1 s -10260 27075 -10060 27121 4 VDD
port 41 nsew
rlabel metal1 s -13810 27030 -13610 27076 4 VDD
port 41 nsew
rlabel metal1 s -5272 27144 -5072 27190 4 VDD
port 41 nsew
rlabel metal1 s -13810 27144 -13610 27190 4 VDD
port 41 nsew
rlabel metal1 s -8822 27271 -8622 27317 4 VDD
port 41 nsew
rlabel metal1 s -10260 27271 -10060 27317 4 VDD
port 41 nsew
rlabel metal1 s -5272 27340 -5072 27386 4 VDD
port 41 nsew
rlabel metal1 s -13810 27340 -13610 27386 4 VDD
port 41 nsew
rlabel metal1 s -5272 27453 -5072 27499 4 VDD
port 41 nsew
rlabel metal1 s -13810 27453 -13610 27499 4 VDD
port 41 nsew
rlabel metal1 s -5272 27649 -5072 27695 4 VDD
port 41 nsew
rlabel metal1 s -13810 27649 -13610 27695 4 VDD
port 41 nsew
rlabel metal1 s -7504 27883 -7304 27929 4 VDD
port 41 nsew
rlabel metal1 s -11578 27883 -11378 27929 4 VDD
port 41 nsew
rlabel metal1 s -5830 27966 -5694 27970 4 VDD
port 41 nsew
rlabel metal1 s -6597 27965 -6461 27970 4 VDD
port 41 nsew
rlabel metal1 s -6597 27970 -5694 28084 4 VDD
port 41 nsew
rlabel metal1 s -12421 27965 -12285 27970 4 VDD
port 41 nsew
rlabel metal1 s -13188 27966 -13052 27970 4 VDD
port 41 nsew
rlabel metal1 s -5830 28084 -5694 28089 4 VDD
port 41 nsew
rlabel metal1 s -6597 28084 -6461 28088 4 VDD
port 41 nsew
rlabel metal1 s -7504 28079 -7304 28125 4 VDD
port 41 nsew
rlabel metal1 s -11578 28079 -11378 28125 4 VDD
port 41 nsew
rlabel metal1 s -13188 27970 -12285 28084 4 VDD
port 41 nsew
rlabel metal1 s -12421 28084 -12285 28088 4 VDD
port 41 nsew
rlabel metal1 s -13188 28084 -13052 28089 4 VDD
port 41 nsew
rlabel metal1 s -7504 28275 -7304 28321 4 VDD
port 41 nsew
rlabel metal1 s -11578 28275 -11378 28321 4 VDD
port 41 nsew
rlabel metal1 s -8822 28742 -8622 28788 4 VDD
port 41 nsew
rlabel metal1 s -10260 28742 -10060 28788 4 VDD
port 41 nsew
rlabel metal1 s -7504 28840 -7304 28886 4 VDD
port 41 nsew
rlabel metal1 s -11578 28840 -11378 28886 4 VDD
port 41 nsew
rlabel metal1 s -8822 28938 -8622 28984 4 VDD
port 41 nsew
rlabel metal1 s -10260 28938 -10060 28984 4 VDD
port 41 nsew
rlabel metal1 s -7504 29036 -7304 29082 4 VDD
port 41 nsew
rlabel metal1 s -11578 29036 -11378 29082 4 VDD
port 41 nsew
rlabel metal1 s -5272 29138 -5072 29184 4 VDD
port 41 nsew
rlabel metal1 s -8822 29134 -8622 29180 4 VDD
port 41 nsew
rlabel metal1 s -10260 29134 -10060 29180 4 VDD
port 41 nsew
rlabel metal1 s -13810 29138 -13610 29184 4 VDD
port 41 nsew
rlabel metal1 s -7504 29232 -7304 29278 4 VDD
port 41 nsew
rlabel metal1 s -11578 29232 -11378 29278 4 VDD
port 41 nsew
rlabel metal1 s -5272 29334 -5072 29380 4 VDD
port 41 nsew
rlabel metal1 s -13810 29334 -13610 29380 4 VDD
port 41 nsew
rlabel metal1 s -5272 29530 -5072 29576 4 VDD
port 41 nsew
rlabel metal1 s -13810 29530 -13610 29576 4 VDD
port 41 nsew
rlabel metal1 s -8822 29579 -8622 29625 4 VDD
port 41 nsew
rlabel metal1 s -10260 29579 -10060 29625 4 VDD
port 41 nsew
rlabel metal1 s -5272 29644 -5072 29690 4 VDD
port 41 nsew
rlabel metal1 s -13810 29644 -13610 29690 4 VDD
port 41 nsew
rlabel metal1 s -8822 29775 -8622 29821 4 VDD
port 41 nsew
rlabel metal1 s -10260 29775 -10060 29821 4 VDD
port 41 nsew
rlabel metal1 s -5272 29840 -5072 29886 4 VDD
port 41 nsew
rlabel metal1 s -13810 29840 -13610 29886 4 VDD
port 41 nsew
rlabel metal1 s -5272 29953 -5072 29999 4 VDD
port 41 nsew
rlabel metal1 s -8822 29971 -8622 30017 4 VDD
port 41 nsew
rlabel metal1 s -10260 29971 -10060 30017 4 VDD
port 41 nsew
rlabel metal1 s -13810 29953 -13610 29999 4 VDD
port 41 nsew
rlabel metal1 s -5272 30149 -5072 30195 4 VDD
port 41 nsew
rlabel metal1 s -13810 30149 -13610 30195 4 VDD
port 41 nsew
rlabel metal1 s -5865 30533 -5729 30537 4 VDD
port 41 nsew
rlabel metal1 s -6453 30532 -6317 30537 4 VDD
port 41 nsew
rlabel metal1 s -6453 30537 -5729 30651 4 VDD
port 41 nsew
rlabel metal1 s -12565 30532 -12429 30537 4 VDD
port 41 nsew
rlabel metal1 s -13153 30533 -13017 30537 4 VDD
port 41 nsew
rlabel metal1 s -7504 30583 -7304 30629 4 VDD
port 41 nsew
rlabel metal1 s -11578 30583 -11378 30629 4 VDD
port 41 nsew
rlabel metal1 s -5865 30651 -5729 30656 4 VDD
port 41 nsew
rlabel metal1 s -6453 30651 -6317 30655 4 VDD
port 41 nsew
rlabel metal1 s -13153 30537 -12429 30651 4 VDD
port 41 nsew
rlabel metal1 s -12565 30651 -12429 30655 4 VDD
port 41 nsew
rlabel metal1 s -13153 30651 -13017 30656 4 VDD
port 41 nsew
rlabel metal1 s -7504 30779 -7304 30825 4 VDD
port 41 nsew
rlabel metal1 s -11578 30779 -11378 30825 4 VDD
port 41 nsew
rlabel metal1 s -7504 30975 -7304 31021 4 VDD
port 41 nsew
rlabel metal1 s -11578 30975 -11378 31021 4 VDD
port 41 nsew
rlabel metal1 s -7504 31465 -7304 31511 4 VDD
port 41 nsew
rlabel metal1 s -11578 31465 -11378 31511 4 VDD
port 41 nsew
rlabel metal1 s -5272 31638 -5072 31684 4 VDD
port 41 nsew
rlabel metal1 s -7504 31661 -7304 31707 4 VDD
port 41 nsew
rlabel metal1 s -11578 31661 -11378 31707 4 VDD
port 41 nsew
rlabel metal1 s -13810 31638 -13610 31684 4 VDD
port 41 nsew
rlabel metal1 s -5272 31834 -5072 31880 4 VDD
port 41 nsew
rlabel metal1 s -7263 31791 -7127 31914 4 VDD
port 41 nsew
rlabel metal1 s -7504 31857 -7304 31903 4 VDD
port 41 nsew
rlabel metal1 s -11578 31857 -11378 31903 4 VDD
port 41 nsew
rlabel metal1 s -11755 31791 -11619 31914 4 VDD
port 41 nsew
rlabel metal1 s -13810 31834 -13610 31880 4 VDD
port 41 nsew
rlabel metal1 s -5272 32030 -5072 32076 4 VDD
port 41 nsew
rlabel metal1 s -7254 31914 -7139 32085 4 VDD
port 41 nsew
rlabel metal1 s -11743 31914 -11628 32085 4 VDD
port 41 nsew
rlabel metal1 s -13810 32030 -13610 32076 4 VDD
port 41 nsew
rlabel metal1 s -5272 32144 -5072 32190 4 VDD
port 41 nsew
rlabel metal1 s -7262 32085 -7126 32208 4 VDD
port 41 nsew
rlabel metal1 s -7521 32199 -7321 32245 4 VDD
port 41 nsew
rlabel metal1 s -11561 32199 -11361 32245 4 VDD
port 41 nsew
rlabel metal1 s -11756 32085 -11620 32208 4 VDD
port 41 nsew
rlabel metal1 s -13810 32144 -13610 32190 4 VDD
port 41 nsew
rlabel metal1 s -5272 32340 -5072 32386 4 VDD
port 41 nsew
rlabel metal1 s -13810 32340 -13610 32386 4 VDD
port 41 nsew
rlabel metal1 s -7521 32395 -7321 32441 4 VDD
port 41 nsew
rlabel metal1 s -11561 32395 -11361 32441 4 VDD
port 41 nsew
rlabel metal1 s -5272 32453 -5072 32499 4 VDD
port 41 nsew
rlabel metal1 s -13810 32453 -13610 32499 4 VDD
port 41 nsew
rlabel metal1 s -5272 32649 -5072 32695 4 VDD
port 41 nsew
rlabel metal1 s -13810 32649 -13610 32695 4 VDD
port 41 nsew
rlabel metal1 s -7521 32937 -7321 32983 4 VDD
port 41 nsew
rlabel metal1 s -11561 32937 -11361 32983 4 VDD
port 41 nsew
rlabel metal1 s -5865 33016 -5729 33020 4 VDD
port 41 nsew
rlabel metal1 s -6345 33015 -6282 33020 4 VDD
port 41 nsew
rlabel metal1 s -6345 33020 -5729 33134 4 VDD
port 41 nsew
rlabel metal1 s -12600 33015 -12537 33020 4 VDD
port 41 nsew
rlabel metal1 s -13153 33016 -13017 33020 4 VDD
port 41 nsew
rlabel metal1 s -5865 33134 -5729 33139 4 VDD
port 41 nsew
rlabel metal1 s -6345 33134 -6282 33138 4 VDD
port 41 nsew
rlabel metal1 s -6345 33138 -6283 33321 4 VDD
port 41 nsew
rlabel metal1 s -7521 33133 -7321 33179 4 VDD
port 41 nsew
rlabel metal1 s -11561 33133 -11361 33179 4 VDD
port 41 nsew
rlabel metal1 s -13153 33020 -12537 33134 4 VDD
port 41 nsew
rlabel metal1 s -12600 33134 -12537 33138 4 VDD
port 41 nsew
rlabel metal1 s -12599 33138 -12537 33321 4 VDD
port 41 nsew
rlabel metal1 s -13153 33134 -13017 33139 4 VDD
port 41 nsew
rlabel metal1 s -7521 33329 -7321 33375 4 VDD
port 41 nsew
rlabel metal1 s -11561 33329 -11361 33375 4 VDD
port 41 nsew
rlabel metal1 s -7521 33525 -7321 33571 4 VDD
port 41 nsew
rlabel metal1 s -11561 33525 -11361 33571 4 VDD
port 41 nsew
rlabel metal1 s -7434 33932 -7334 33978 4 VDD
port 41 nsew
rlabel metal1 s -11548 33932 -11448 33978 4 VDD
port 41 nsew
rlabel metal1 s -5272 34138 -5072 34184 4 VDD
port 41 nsew
rlabel metal1 s -7434 34128 -7334 34174 4 VDD
port 41 nsew
rlabel metal1 s -11548 34128 -11448 34174 4 VDD
port 41 nsew
rlabel metal1 s -13810 34138 -13610 34184 4 VDD
port 41 nsew
rlabel metal1 s -5272 34334 -5072 34380 4 VDD
port 41 nsew
rlabel metal1 s -7434 34324 -7334 34370 4 VDD
port 41 nsew
rlabel metal1 s -11548 34324 -11448 34370 4 VDD
port 41 nsew
rlabel metal1 s -13810 34334 -13610 34380 4 VDD
port 41 nsew
rlabel metal1 s -5272 34530 -5072 34576 4 VDD
port 41 nsew
rlabel metal1 s -7434 34520 -7334 34566 4 VDD
port 41 nsew
rlabel metal1 s -11548 34520 -11448 34566 4 VDD
port 41 nsew
rlabel metal1 s -13810 34530 -13610 34576 4 VDD
port 41 nsew
rlabel metal1 s -5272 34644 -5072 34690 4 VDD
port 41 nsew
rlabel metal1 s -13810 34644 -13610 34690 4 VDD
port 41 nsew
rlabel metal1 s -7635 34737 -7335 34783 4 VDD
port 41 nsew
rlabel metal1 s -11547 34737 -11247 34783 4 VDD
port 41 nsew
rlabel metal1 s -5272 34840 -5072 34886 4 VDD
port 41 nsew
rlabel metal1 s -13810 34840 -13610 34886 4 VDD
port 41 nsew
rlabel metal1 s -5272 34953 -5072 34999 4 VDD
port 41 nsew
rlabel metal1 s -7635 34933 -7335 34979 4 VDD
port 41 nsew
rlabel metal1 s -11547 34933 -11247 34979 4 VDD
port 41 nsew
rlabel metal1 s -13810 34953 -13610 34999 4 VDD
port 41 nsew
rlabel metal1 s -5272 35149 -5072 35195 4 VDD
port 41 nsew
rlabel metal1 s -7275 35063 -7139 35186 4 VDD
port 41 nsew
rlabel metal1 s -7635 35129 -7335 35175 4 VDD
port 41 nsew
rlabel metal1 s -11547 35129 -11247 35175 4 VDD
port 41 nsew
rlabel metal1 s -11743 35063 -11607 35186 4 VDD
port 41 nsew
rlabel metal1 s -7261 35186 -7154 35452 4 VDD
port 41 nsew
rlabel metal1 s -11728 35186 -11621 35452 4 VDD
port 41 nsew
rlabel metal1 s -13810 35149 -13610 35195 4 VDD
port 41 nsew
rlabel metal1 s -7274 35452 -7138 35575 4 VDD
port 41 nsew
rlabel metal1 s -7436 35537 -7336 35583 4 VDD
port 41 nsew
rlabel metal1 s -11546 35537 -11446 35583 4 VDD
port 41 nsew
rlabel metal1 s -11744 35452 -11608 35575 4 VDD
port 41 nsew
rlabel metal1 s -7436 35733 -7336 35779 4 VDD
port 41 nsew
rlabel metal1 s -11546 35733 -11446 35779 4 VDD
port 41 nsew
rlabel metal1 s -7436 35929 -7336 35975 4 VDD
port 41 nsew
rlabel metal1 s -11546 35929 -11446 35975 4 VDD
port 41 nsew
rlabel metal1 s -7436 36125 -7336 36171 4 VDD
port 41 nsew
rlabel metal1 s -11546 36125 -11446 36171 4 VDD
port 41 nsew
rlabel metal1 s -7637 36342 -7337 36388 4 VDD
port 41 nsew
rlabel metal1 s -11545 36342 -11245 36388 4 VDD
port 41 nsew
rlabel metal1 s -7637 36538 -7337 36584 4 VDD
port 41 nsew
rlabel metal1 s -11545 36538 -11245 36584 4 VDD
port 41 nsew
rlabel metal1 s -5272 36638 -5072 36684 4 VDD
port 41 nsew
rlabel metal1 s -7251 36680 -7115 36803 4 VDD
port 41 nsew
rlabel metal1 s -7637 36734 -7337 36780 4 VDD
port 41 nsew
rlabel metal1 s -11545 36734 -11245 36780 4 VDD
port 41 nsew
rlabel metal1 s -11767 36680 -11631 36803 4 VDD
port 41 nsew
rlabel metal1 s -13810 36638 -13610 36684 4 VDD
port 41 nsew
rlabel metal1 s -5272 36834 -5072 36880 4 VDD
port 41 nsew
rlabel metal1 s -5272 37030 -5072 37076 4 VDD
port 41 nsew
rlabel metal1 s -7231 36803 -7124 37081 4 VDD
port 41 nsew
rlabel metal1 s -11758 36803 -11651 37081 4 VDD
port 41 nsew
rlabel metal1 s -13810 36834 -13610 36880 4 VDD
port 41 nsew
rlabel metal1 s -13810 37030 -13610 37076 4 VDD
port 41 nsew
rlabel metal1 s -5272 37144 -5072 37190 4 VDD
port 41 nsew
rlabel metal1 s -7249 37081 -7113 37204 4 VDD
port 41 nsew
rlabel metal1 s -7512 37161 -7312 37207 4 VDD
port 41 nsew
rlabel metal1 s -11570 37161 -11370 37207 4 VDD
port 41 nsew
rlabel metal1 s -11769 37081 -11633 37204 4 VDD
port 41 nsew
rlabel metal1 s -13810 37144 -13610 37190 4 VDD
port 41 nsew
rlabel metal1 s -5272 37340 -5072 37386 4 VDD
port 41 nsew
rlabel metal1 s -7512 37357 -7312 37403 4 VDD
port 41 nsew
rlabel metal1 s -11570 37357 -11370 37403 4 VDD
port 41 nsew
rlabel metal1 s -13810 37340 -13610 37386 4 VDD
port 41 nsew
rlabel metal1 s -5272 37453 -5072 37499 4 VDD
port 41 nsew
rlabel metal1 s -13810 37453 -13610 37499 4 VDD
port 41 nsew
rlabel metal1 s -5272 37649 -5072 37695 4 VDD
port 41 nsew
rlabel metal1 s -13810 37649 -13610 37695 4 VDD
port 41 nsew
rlabel metal1 s -7512 37899 -7312 37945 4 VDD
port 41 nsew
rlabel metal1 s -11570 37899 -11370 37945 4 VDD
port 41 nsew
rlabel metal1 s -7512 38095 -7312 38141 4 VDD
port 41 nsew
rlabel metal1 s -11570 38095 -11370 38141 4 VDD
port 41 nsew
rlabel metal1 s -7512 38291 -7312 38337 4 VDD
port 41 nsew
rlabel metal1 s -11570 38291 -11370 38337 4 VDD
port 41 nsew
rlabel metal1 s -7254 38437 -7118 38560 4 VDD
port 41 nsew
rlabel metal1 s -7512 38487 -7312 38533 4 VDD
port 41 nsew
rlabel metal1 s -11570 38487 -11370 38533 4 VDD
port 41 nsew
rlabel metal1 s -11764 38437 -11628 38560 4 VDD
port 41 nsew
rlabel metal1 s -3742 39356 -2367 40236 4 VDD
port 41 nsew
rlabel metal1 s -5272 39638 -5072 39684 4 VDD
port 41 nsew
rlabel metal1 s -7236 38560 -7131 39653 4 VDD
port 41 nsew
rlabel metal1 s -7255 39653 -7119 39776 4 VDD
port 41 nsew
rlabel metal1 s -7523 39648 -7323 39694 4 VDD
port 41 nsew
rlabel metal1 s -11559 39648 -11359 39694 4 VDD
port 41 nsew
rlabel metal1 s -11751 38560 -11646 39653 4 VDD
port 41 nsew
rlabel metal1 s -11763 39653 -11627 39776 4 VDD
port 41 nsew
rlabel metal1 s -13810 39638 -13610 39684 4 VDD
port 41 nsew
rlabel metal1 s -5272 39834 -5072 39880 4 VDD
port 41 nsew
rlabel metal1 s -7523 39844 -7323 39890 4 VDD
port 41 nsew
rlabel metal1 s -11559 39844 -11359 39890 4 VDD
port 41 nsew
rlabel metal1 s -13810 39834 -13610 39880 4 VDD
port 41 nsew
rlabel metal1 s -5272 40030 -5072 40076 4 VDD
port 41 nsew
rlabel metal1 s -7523 40040 -7323 40086 4 VDD
port 41 nsew
rlabel metal1 s -11559 40040 -11359 40086 4 VDD
port 41 nsew
rlabel metal1 s -13810 40030 -13610 40076 4 VDD
port 41 nsew
rlabel metal1 s -5272 40144 -5072 40190 4 VDD
port 41 nsew
rlabel metal1 s -7523 40154 -7323 40200 4 VDD
port 41 nsew
rlabel metal1 s -11559 40154 -11359 40200 4 VDD
port 41 nsew
rlabel metal1 s -13810 40144 -13610 40190 4 VDD
port 41 nsew
rlabel metal1 s -3742 40236 -2527 40571 4 VDD
port 41 nsew
rlabel metal1 s -5272 40340 -5072 40386 4 VDD
port 41 nsew
rlabel metal1 s -7523 40350 -7323 40396 4 VDD
port 41 nsew
rlabel metal1 s -11559 40350 -11359 40396 4 VDD
port 41 nsew
rlabel metal1 s -13810 40340 -13610 40386 4 VDD
port 41 nsew
rlabel metal1 s -5272 40453 -5072 40499 4 VDD
port 41 nsew
rlabel metal1 s -7523 40463 -7323 40509 4 VDD
port 41 nsew
rlabel metal1 s -11559 40463 -11359 40509 4 VDD
port 41 nsew
rlabel metal1 s -13810 40453 -13610 40499 4 VDD
port 41 nsew
rlabel metal1 s -5272 40649 -5072 40695 4 VDD
port 41 nsew
rlabel metal1 s -7523 40659 -7323 40705 4 VDD
port 41 nsew
rlabel metal1 s -11559 40659 -11359 40705 4 VDD
port 41 nsew
rlabel metal1 s -13810 40649 -13610 40695 4 VDD
port 41 nsew
rlabel metal1 s -12329 43879 -12129 43925 4 VDD
port 41 nsew
rlabel metal1 s -12329 44075 -12129 44121 4 VDD
port 41 nsew
rlabel metal1 s -12329 44271 -12129 44317 4 VDD
port 41 nsew
rlabel metal1 s -12329 44761 -12129 44807 4 VDD
port 41 nsew
rlabel metal1 s -12329 44957 -12129 45003 4 VDD
port 41 nsew
rlabel metal1 s -12329 45153 -12129 45199 4 VDD
port 41 nsew
rlabel metal1 s -13647 45765 -13447 45811 4 VDD
port 41 nsew
rlabel metal1 s -13647 45961 -13447 46007 4 VDD
port 41 nsew
rlabel metal1 s -13647 46157 -13447 46203 4 VDD
port 41 nsew
rlabel metal1 s -12329 46504 -12129 46550 4 VDD
port 41 nsew
rlabel metal1 s -13647 46602 -13447 46648 4 VDD
port 41 nsew
rlabel metal1 s -12329 46700 -12129 46746 4 VDD
port 41 nsew
rlabel metal1 s -13647 46798 -13447 46844 4 VDD
port 41 nsew
rlabel metal1 s -12329 46896 -12129 46942 4 VDD
port 41 nsew
rlabel metal1 s -13647 46994 -13447 47040 4 VDD
port 41 nsew
rlabel metal1 s -12329 47461 -12129 47507 4 VDD
port 41 nsew
rlabel metal1 s -12329 47657 -12129 47703 4 VDD
port 41 nsew
rlabel metal1 s -12329 47853 -12129 47899 4 VDD
port 41 nsew
rlabel metal1 s -13647 48465 -13447 48511 4 VDD
port 41 nsew
rlabel metal1 s -13647 48661 -13447 48707 4 VDD
port 41 nsew
rlabel metal1 s -13647 48857 -13447 48903 4 VDD
port 41 nsew
rlabel metal1 s -12329 49204 -12129 49250 4 VDD
port 41 nsew
rlabel metal1 s -13647 49302 -13447 49348 4 VDD
port 41 nsew
rlabel metal1 s -12329 49400 -12129 49446 4 VDD
port 41 nsew
rlabel metal1 s -13647 49498 -13447 49544 4 VDD
port 41 nsew
rlabel metal1 s -12329 49596 -12129 49642 4 VDD
port 41 nsew
rlabel metal1 s -13647 49694 -13447 49740 4 VDD
port 41 nsew
rlabel metal1 s -8971 50686 -8371 50732 4 VDD
port 41 nsew
rlabel metal1 s -11317 50681 -10917 50727 4 VDD
port 41 nsew
rlabel metal1 s -8971 50882 -8371 50928 4 VDD
port 41 nsew
rlabel metal1 s -11317 50877 -10917 50923 4 VDD
port 41 nsew
rlabel metal1 s -11317 51627 -10917 51673 4 VDD
port 41 nsew
rlabel metal1 s -11317 51823 -10917 51869 4 VDD
port 41 nsew
rlabel metal1 s -9091 52007 -8891 52053 4 VDD
port 41 nsew
rlabel metal1 s -9091 52203 -8891 52249 4 VDD
port 41 nsew
rlabel metal1 s -9091 52399 -8891 52445 4 VDD
port 41 nsew
rlabel metal1 s -11351 52543 -11151 52589 4 VDD
port 41 nsew
rlabel metal1 s -11351 52739 -11151 52785 4 VDD
port 41 nsew
rlabel metal1 s -9091 52889 -8891 52935 4 VDD
port 41 nsew
rlabel metal1 s -11351 52935 -11151 52981 4 VDD
port 41 nsew
rlabel metal1 s -9091 53085 -8891 53131 4 VDD
port 41 nsew
rlabel metal1 s -11351 53131 -11151 53177 4 VDD
port 41 nsew
rlabel metal1 s -9091 53281 -8891 53327 4 VDD
port 41 nsew
rlabel metal1 s -11351 53673 -11151 53719 4 VDD
port 41 nsew
rlabel metal1 s -7773 53893 -7573 53939 4 VDD
port 41 nsew
rlabel metal1 s -11351 53869 -11151 53915 4 VDD
port 41 nsew
rlabel metal1 s -7773 54089 -7573 54135 4 VDD
port 41 nsew
rlabel metal1 s -7773 54285 -7573 54331 4 VDD
port 41 nsew
rlabel metal1 s -11344 54402 -11144 54448 4 VDD
port 41 nsew
rlabel metal1 s -10043 54452 -9643 54498 4 VDD
port 41 nsew
rlabel metal1 s -9091 54632 -8891 54678 4 VDD
port 41 nsew
rlabel metal1 s -11344 54598 -11144 54644 4 VDD
port 41 nsew
rlabel metal1 s -10043 54648 -9643 54694 4 VDD
port 41 nsew
rlabel metal1 s -7773 54730 -7573 54776 4 VDD
port 41 nsew
rlabel metal1 s -9091 54828 -8891 54874 4 VDD
port 41 nsew
rlabel metal1 s -11344 54794 -11144 54840 4 VDD
port 41 nsew
rlabel metal1 s -10043 54844 -9643 54890 4 VDD
port 41 nsew
rlabel metal1 s -7773 54926 -7573 54972 4 VDD
port 41 nsew
rlabel metal1 s -9091 55024 -8891 55070 4 VDD
port 41 nsew
rlabel metal1 s -7773 55122 -7573 55168 4 VDD
port 41 nsew
rlabel metal1 s -11273 55282 -10573 55328 4 VDD
port 41 nsew
rlabel metal1 s -11273 55478 -10573 55524 4 VDD
port 41 nsew
rlabel metal1 s -9091 55589 -8891 55635 4 VDD
port 41 nsew
rlabel metal1 s -11273 55682 -10573 55728 4 VDD
port 41 nsew
rlabel metal1 s -9091 55785 -8891 55831 4 VDD
port 41 nsew
rlabel metal1 s -11273 55878 -10573 55924 4 VDD
port 41 nsew
rlabel metal1 s -9091 55981 -8891 56027 4 VDD
port 41 nsew
rlabel metal1 s -11273 56282 -10573 56328 4 VDD
port 41 nsew
rlabel metal1 s -11273 56478 -10573 56524 4 VDD
port 41 nsew
rlabel metal1 s -7773 56593 -7573 56639 4 VDD
port 41 nsew
rlabel metal1 s -11273 56682 -10573 56728 4 VDD
port 41 nsew
rlabel metal1 s -7773 56789 -7573 56835 4 VDD
port 41 nsew
rlabel metal1 s -11273 56878 -10573 56924 4 VDD
port 41 nsew
rlabel metal1 s -7773 56985 -7573 57031 4 VDD
port 41 nsew
rlabel metal1 s -11273 57282 -10573 57328 4 VDD
port 41 nsew
rlabel metal1 s -9091 57332 -8891 57378 4 VDD
port 41 nsew
rlabel metal1 s -7773 57430 -7573 57476 4 VDD
port 41 nsew
rlabel metal1 s -11273 57478 -10573 57524 4 VDD
port 41 nsew
rlabel metal1 s -9091 57528 -8891 57574 4 VDD
port 41 nsew
rlabel metal1 s -7773 57626 -7573 57672 4 VDD
port 41 nsew
rlabel metal1 s -9091 57724 -8891 57770 4 VDD
port 41 nsew
rlabel metal1 s -11273 57682 -10573 57728 4 VDD
port 41 nsew
rlabel metal1 s -7773 57822 -7573 57868 4 VDD
port 41 nsew
rlabel metal1 s -11273 57878 -10573 57924 4 VDD
port 41 nsew
rlabel metal1 s -7420 60265 -7220 60311 4 VDD
port 41 nsew
rlabel metal1 s -8449 60239 -8149 60285 4 VDD
port 41 nsew
rlabel metal1 s -10873 60257 -10673 60303 4 VDD
port 41 nsew
rlabel metal1 s -11902 60231 -11602 60277 4 VDD
port 41 nsew
rlabel metal1 s -7420 60461 -7220 60507 4 VDD
port 41 nsew
rlabel metal1 s -8449 60435 -8149 60481 4 VDD
port 41 nsew
rlabel metal1 s -10873 60453 -10673 60499 4 VDD
port 41 nsew
rlabel metal1 s -11902 60427 -11602 60473 4 VDD
port 41 nsew
rlabel metal1 s -7420 60657 -7220 60703 4 VDD
port 41 nsew
rlabel metal1 s -8449 60631 -8149 60677 4 VDD
port 41 nsew
rlabel metal1 s -10873 60649 -10673 60695 4 VDD
port 41 nsew
rlabel metal1 s -11902 60623 -11602 60669 4 VDD
port 41 nsew
rlabel metal1 s -7420 60853 -7220 60899 4 VDD
port 41 nsew
rlabel metal1 s -8248 60848 -8148 60894 4 VDD
port 41 nsew
rlabel metal1 s -10873 60845 -10673 60891 4 VDD
port 41 nsew
rlabel metal1 s -11701 60840 -11601 60886 4 VDD
port 41 nsew
rlabel metal1 s -8248 61044 -8148 61090 4 VDD
port 41 nsew
rlabel metal1 s -11701 61036 -11601 61082 4 VDD
port 41 nsew
rlabel metal1 s -7549 61238 -7249 61284 4 VDD
port 41 nsew
rlabel metal1 s -8248 61240 -8148 61286 4 VDD
port 41 nsew
rlabel metal1 s -11002 61230 -10702 61276 4 VDD
port 41 nsew
rlabel metal1 s -11701 61232 -11601 61278 4 VDD
port 41 nsew
rlabel metal1 s -7549 61434 -7249 61480 4 VDD
port 41 nsew
rlabel metal1 s -8248 61436 -8148 61482 4 VDD
port 41 nsew
rlabel metal1 s -11002 61426 -10702 61472 4 VDD
port 41 nsew
rlabel metal1 s -11366 61432 -11236 61615 4 VDD
port 41 nsew
rlabel metal1 s -11701 61428 -11601 61474 4 VDD
port 41 nsew
rlabel metal1 s -7549 61630 -7249 61676 4 VDD
port 41 nsew
rlabel metal1 s -11002 61622 -10702 61668 4 VDD
port 41 nsew
rlabel metal1 s -8660 61686 -8060 61732 4 VDD
port 41 nsew
rlabel metal1 s -7550 61847 -7450 61893 4 VDD
port 41 nsew
rlabel metal1 s -8660 61882 -8060 61928 4 VDD
port 41 nsew
rlabel metal1 s -11003 61839 -10903 61885 4 VDD
port 41 nsew
rlabel metal1 s -7550 62043 -7450 62089 4 VDD
port 41 nsew
rlabel metal1 s -11003 62035 -10903 62081 4 VDD
port 41 nsew
rlabel metal1 s -7550 62239 -7450 62285 4 VDD
port 41 nsew
rlabel metal1 s -11003 62231 -10903 62277 4 VDD
port 41 nsew
rlabel metal1 s -8660 62305 -8060 62351 4 VDD
port 41 nsew
rlabel metal1 s -7550 62435 -7450 62481 4 VDD
port 41 nsew
rlabel metal1 s -11003 62427 -10903 62473 4 VDD
port 41 nsew
rlabel metal1 s -7967 62517 -7849 62591 4 VDD
port 41 nsew
rlabel metal1 s -7961 62591 -7865 62745 4 VDD
port 41 nsew
rlabel metal1 s -11359 61615 -11277 62735 4 VDD
port 41 nsew
rlabel metal1 s -12113 61678 -11513 61724 4 VDD
port 41 nsew
rlabel metal1 s -12113 61874 -11513 61920 4 VDD
port 41 nsew
rlabel metal1 s -12113 62297 -11513 62343 4 VDD
port 41 nsew
rlabel metal1 s -7979 62745 -7829 62855 4 VDD
port 41 nsew
rlabel metal1 s -11385 62735 -11248 62831 4 VDD
port 41 nsew
rlabel metal1 s -8418 63678 -7918 63724 4 VDD
port 41 nsew
rlabel metal1 s -8418 63874 -7918 63920 4 VDD
port 41 nsew
rlabel metal1 s -10904 63925 -10704 63971 4 VDD
port 41 nsew
rlabel metal1 s -11933 63899 -11633 63945 4 VDD
port 41 nsew
rlabel metal1 s -10904 64121 -10704 64167 4 VDD
port 41 nsew
rlabel metal1 s -11933 64095 -11633 64141 4 VDD
port 41 nsew
rlabel metal1 s -10904 64317 -10704 64363 4 VDD
port 41 nsew
rlabel metal1 s -11933 64291 -11633 64337 4 VDD
port 41 nsew
rlabel metal1 s -8418 64469 -7918 64515 4 VDD
port 41 nsew
rlabel metal1 s -10904 64513 -10704 64559 4 VDD
port 41 nsew
rlabel metal1 s -11732 64508 -11632 64554 4 VDD
port 41 nsew
rlabel metal1 s -8418 64599 -7918 64645 4 VDD
port 41 nsew
rlabel metal1 s -11732 64704 -11632 64750 4 VDD
port 41 nsew
rlabel metal1 s -8218 64827 -7918 64873 4 VDD
port 41 nsew
rlabel metal1 s -11033 64898 -10733 64944 4 VDD
port 41 nsew
rlabel metal1 s -11732 64900 -11632 64946 4 VDD
port 41 nsew
rlabel metal1 s -8218 65023 -7918 65069 4 VDD
port 41 nsew
rlabel metal1 s -11033 65094 -10733 65140 4 VDD
port 41 nsew
rlabel metal1 s -11732 65096 -11632 65142 4 VDD
port 41 nsew
rlabel metal1 s -11033 65290 -10733 65336 4 VDD
port 41 nsew
rlabel metal1 s -12144 65346 -11544 65392 4 VDD
port 41 nsew
rlabel metal1 s -11034 65507 -10934 65553 4 VDD
port 41 nsew
rlabel metal1 s -12144 65542 -11544 65588 4 VDD
port 41 nsew
rlabel metal1 s -11034 65703 -10934 65749 4 VDD
port 41 nsew
rlabel metal1 s -11034 65899 -10934 65945 4 VDD
port 41 nsew
rlabel metal1 s -12144 65965 -11544 66011 4 VDD
port 41 nsew
rlabel metal1 s -11034 66095 -10934 66141 4 VDD
port 41 nsew
rlabel metal1 s -11450 66155 -11287 66246 4 VDD
port 41 nsew
rlabel metal1 s -11438 66246 -11299 66405 4 VDD
port 41 nsew
rlabel metal1 s -11463 66405 -11272 66556 4 VDD
port 41 nsew
rlabel metal1 s -7431 68705 -7231 68751 4 VDD
port 41 nsew
rlabel metal1 s -8460 68679 -8160 68725 4 VDD
port 41 nsew
rlabel metal1 s -10884 68697 -10684 68743 4 VDD
port 41 nsew
rlabel metal1 s -11913 68671 -11613 68717 4 VDD
port 41 nsew
rlabel metal1 s -7431 68901 -7231 68947 4 VDD
port 41 nsew
rlabel metal1 s -8460 68875 -8160 68921 4 VDD
port 41 nsew
rlabel metal1 s -10884 68893 -10684 68939 4 VDD
port 41 nsew
rlabel metal1 s -11913 68867 -11613 68913 4 VDD
port 41 nsew
rlabel metal1 s -7431 69097 -7231 69143 4 VDD
port 41 nsew
rlabel metal1 s -8460 69071 -8160 69117 4 VDD
port 41 nsew
rlabel metal1 s -10884 69089 -10684 69135 4 VDD
port 41 nsew
rlabel metal1 s -11913 69063 -11613 69109 4 VDD
port 41 nsew
rlabel metal1 s -7431 69293 -7231 69339 4 VDD
port 41 nsew
rlabel metal1 s -8259 69288 -8159 69334 4 VDD
port 41 nsew
rlabel metal1 s -10884 69285 -10684 69331 4 VDD
port 41 nsew
rlabel metal1 s -11712 69280 -11612 69326 4 VDD
port 41 nsew
rlabel metal1 s -8259 69484 -8159 69530 4 VDD
port 41 nsew
rlabel metal1 s -11712 69476 -11612 69522 4 VDD
port 41 nsew
rlabel metal1 s -7560 69678 -7260 69724 4 VDD
port 41 nsew
rlabel metal1 s -8259 69680 -8159 69726 4 VDD
port 41 nsew
rlabel metal1 s -11013 69670 -10713 69716 4 VDD
port 41 nsew
rlabel metal1 s -11712 69672 -11612 69718 4 VDD
port 41 nsew
rlabel metal1 s -7560 69874 -7260 69920 4 VDD
port 41 nsew
rlabel metal1 s -8259 69876 -8159 69922 4 VDD
port 41 nsew
rlabel metal1 s -11013 69866 -10713 69912 4 VDD
port 41 nsew
rlabel metal1 s -11377 69872 -11247 70055 4 VDD
port 41 nsew
rlabel metal1 s -11712 69868 -11612 69914 4 VDD
port 41 nsew
rlabel metal1 s -7560 70070 -7260 70116 4 VDD
port 41 nsew
rlabel metal1 s -11013 70062 -10713 70108 4 VDD
port 41 nsew
rlabel metal1 s -8671 70126 -8071 70172 4 VDD
port 41 nsew
rlabel metal1 s -7561 70287 -7461 70333 4 VDD
port 41 nsew
rlabel metal1 s -8671 70322 -8071 70368 4 VDD
port 41 nsew
rlabel metal1 s -11014 70279 -10914 70325 4 VDD
port 41 nsew
rlabel metal1 s -7561 70483 -7461 70529 4 VDD
port 41 nsew
rlabel metal1 s -11014 70475 -10914 70521 4 VDD
port 41 nsew
rlabel metal1 s -7561 70679 -7461 70725 4 VDD
port 41 nsew
rlabel metal1 s -11014 70671 -10914 70717 4 VDD
port 41 nsew
rlabel metal1 s -8671 70745 -8071 70791 4 VDD
port 41 nsew
rlabel metal1 s -7561 70875 -7461 70921 4 VDD
port 41 nsew
rlabel metal1 s -11014 70867 -10914 70913 4 VDD
port 41 nsew
rlabel metal1 s -7978 70957 -7860 71031 4 VDD
port 41 nsew
rlabel metal1 s -7972 71031 -7876 71185 4 VDD
port 41 nsew
rlabel metal1 s -11370 70055 -11288 71175 4 VDD
port 41 nsew
rlabel metal1 s -12124 70118 -11524 70164 4 VDD
port 41 nsew
rlabel metal1 s -12124 70314 -11524 70360 4 VDD
port 41 nsew
rlabel metal1 s -12124 70737 -11524 70783 4 VDD
port 41 nsew
rlabel metal1 s -7990 71185 -7840 71295 4 VDD
port 41 nsew
rlabel metal1 s -11396 71175 -11259 71271 4 VDD
port 41 nsew
rlabel metal1 s -8429 72118 -7929 72164 4 VDD
port 41 nsew
rlabel metal1 s -8429 72314 -7929 72360 4 VDD
port 41 nsew
rlabel metal1 s -10915 72365 -10715 72411 4 VDD
port 41 nsew
rlabel metal1 s -11944 72339 -11644 72385 4 VDD
port 41 nsew
rlabel metal1 s -10915 72561 -10715 72607 4 VDD
port 41 nsew
rlabel metal1 s -11944 72535 -11644 72581 4 VDD
port 41 nsew
rlabel metal1 s -10915 72757 -10715 72803 4 VDD
port 41 nsew
rlabel metal1 s -11944 72731 -11644 72777 4 VDD
port 41 nsew
rlabel metal1 s -8429 72909 -7929 72955 4 VDD
port 41 nsew
rlabel metal1 s -10915 72953 -10715 72999 4 VDD
port 41 nsew
rlabel metal1 s -11743 72948 -11643 72994 4 VDD
port 41 nsew
rlabel metal1 s -8429 73039 -7929 73085 4 VDD
port 41 nsew
rlabel metal1 s -11743 73144 -11643 73190 4 VDD
port 41 nsew
rlabel metal1 s -8229 73267 -7929 73313 4 VDD
port 41 nsew
rlabel metal1 s -11044 73338 -10744 73384 4 VDD
port 41 nsew
rlabel metal1 s -11743 73340 -11643 73386 4 VDD
port 41 nsew
rlabel metal1 s -8229 73463 -7929 73509 4 VDD
port 41 nsew
rlabel metal1 s -11044 73534 -10744 73580 4 VDD
port 41 nsew
rlabel metal1 s -11743 73536 -11643 73582 4 VDD
port 41 nsew
rlabel metal1 s -11044 73730 -10744 73776 4 VDD
port 41 nsew
rlabel metal1 s -12155 73786 -11555 73832 4 VDD
port 41 nsew
rlabel metal1 s -11045 73947 -10945 73993 4 VDD
port 41 nsew
rlabel metal1 s -12155 73982 -11555 74028 4 VDD
port 41 nsew
rlabel metal1 s -11045 74143 -10945 74189 4 VDD
port 41 nsew
rlabel metal1 s -11045 74339 -10945 74385 4 VDD
port 41 nsew
rlabel metal1 s -12155 74405 -11555 74451 4 VDD
port 41 nsew
rlabel metal1 s -11045 74535 -10945 74581 4 VDD
port 41 nsew
rlabel metal1 s -11461 74595 -11298 74686 4 VDD
port 41 nsew
rlabel metal1 s -11449 74686 -11310 74845 4 VDD
port 41 nsew
rlabel metal1 s -11474 74845 -11283 74996 4 VDD
port 41 nsew
rlabel metal1 s -7470 77568 -7270 77614 4 VDD
port 41 nsew
rlabel metal1 s -8499 77542 -8199 77588 4 VDD
port 41 nsew
rlabel metal1 s -10923 77560 -10723 77606 4 VDD
port 41 nsew
rlabel metal1 s -11952 77534 -11652 77580 4 VDD
port 41 nsew
rlabel metal1 s -7470 77764 -7270 77810 4 VDD
port 41 nsew
rlabel metal1 s -8499 77738 -8199 77784 4 VDD
port 41 nsew
rlabel metal1 s -10923 77756 -10723 77802 4 VDD
port 41 nsew
rlabel metal1 s -11952 77730 -11652 77776 4 VDD
port 41 nsew
rlabel metal1 s -7470 77960 -7270 78006 4 VDD
port 41 nsew
rlabel metal1 s -8499 77934 -8199 77980 4 VDD
port 41 nsew
rlabel metal1 s -10923 77952 -10723 77998 4 VDD
port 41 nsew
rlabel metal1 s -11952 77926 -11652 77972 4 VDD
port 41 nsew
rlabel metal1 s -7470 78156 -7270 78202 4 VDD
port 41 nsew
rlabel metal1 s -8298 78151 -8198 78197 4 VDD
port 41 nsew
rlabel metal1 s -10923 78148 -10723 78194 4 VDD
port 41 nsew
rlabel metal1 s -11751 78143 -11651 78189 4 VDD
port 41 nsew
rlabel metal1 s -8298 78347 -8198 78393 4 VDD
port 41 nsew
rlabel metal1 s -11751 78339 -11651 78385 4 VDD
port 41 nsew
rlabel metal1 s -7599 78541 -7299 78587 4 VDD
port 41 nsew
rlabel metal1 s -8298 78543 -8198 78589 4 VDD
port 41 nsew
rlabel metal1 s -11052 78533 -10752 78579 4 VDD
port 41 nsew
rlabel metal1 s -11751 78535 -11651 78581 4 VDD
port 41 nsew
rlabel metal1 s -7599 78737 -7299 78783 4 VDD
port 41 nsew
rlabel metal1 s -8298 78739 -8198 78785 4 VDD
port 41 nsew
rlabel metal1 s -11052 78729 -10752 78775 4 VDD
port 41 nsew
rlabel metal1 s -11416 78735 -11286 78918 4 VDD
port 41 nsew
rlabel metal1 s -11751 78731 -11651 78777 4 VDD
port 41 nsew
rlabel metal1 s -7599 78933 -7299 78979 4 VDD
port 41 nsew
rlabel metal1 s -11052 78925 -10752 78971 4 VDD
port 41 nsew
rlabel metal1 s -8710 78989 -8110 79035 4 VDD
port 41 nsew
rlabel metal1 s -7600 79150 -7500 79196 4 VDD
port 41 nsew
rlabel metal1 s -8710 79185 -8110 79231 4 VDD
port 41 nsew
rlabel metal1 s -11053 79142 -10953 79188 4 VDD
port 41 nsew
rlabel metal1 s -7600 79346 -7500 79392 4 VDD
port 41 nsew
rlabel metal1 s -11053 79338 -10953 79384 4 VDD
port 41 nsew
rlabel metal1 s -7600 79542 -7500 79588 4 VDD
port 41 nsew
rlabel metal1 s -11053 79534 -10953 79580 4 VDD
port 41 nsew
rlabel metal1 s -8710 79608 -8110 79654 4 VDD
port 41 nsew
rlabel metal1 s -7600 79738 -7500 79784 4 VDD
port 41 nsew
rlabel metal1 s -11053 79730 -10953 79776 4 VDD
port 41 nsew
rlabel metal1 s -8017 79820 -7899 79894 4 VDD
port 41 nsew
rlabel metal1 s -8011 79894 -7915 80048 4 VDD
port 41 nsew
rlabel metal1 s -11409 78918 -11327 80038 4 VDD
port 41 nsew
rlabel metal1 s -12163 78981 -11563 79027 4 VDD
port 41 nsew
rlabel metal1 s -12163 79177 -11563 79223 4 VDD
port 41 nsew
rlabel metal1 s -12163 79600 -11563 79646 4 VDD
port 41 nsew
rlabel metal1 s -8029 80048 -7879 80158 4 VDD
port 41 nsew
rlabel metal1 s -11435 80038 -11298 80134 4 VDD
port 41 nsew
rlabel metal1 s -8468 80981 -7968 81027 4 VDD
port 41 nsew
rlabel metal1 s -8468 81177 -7968 81223 4 VDD
port 41 nsew
rlabel metal1 s -10954 81228 -10754 81274 4 VDD
port 41 nsew
rlabel metal1 s -11983 81202 -11683 81248 4 VDD
port 41 nsew
rlabel metal1 s -10954 81424 -10754 81470 4 VDD
port 41 nsew
rlabel metal1 s -11983 81398 -11683 81444 4 VDD
port 41 nsew
rlabel metal1 s -10954 81620 -10754 81666 4 VDD
port 41 nsew
rlabel metal1 s -11983 81594 -11683 81640 4 VDD
port 41 nsew
rlabel metal1 s -8468 81772 -7968 81818 4 VDD
port 41 nsew
rlabel metal1 s -10954 81816 -10754 81862 4 VDD
port 41 nsew
rlabel metal1 s -11782 81811 -11682 81857 4 VDD
port 41 nsew
rlabel metal1 s -8468 81902 -7968 81948 4 VDD
port 41 nsew
rlabel metal1 s -11782 82007 -11682 82053 4 VDD
port 41 nsew
rlabel metal1 s -8268 82130 -7968 82176 4 VDD
port 41 nsew
rlabel metal1 s -11083 82201 -10783 82247 4 VDD
port 41 nsew
rlabel metal1 s -11782 82203 -11682 82249 4 VDD
port 41 nsew
rlabel metal1 s -8268 82326 -7968 82372 4 VDD
port 41 nsew
rlabel metal1 s -11083 82397 -10783 82443 4 VDD
port 41 nsew
rlabel metal1 s -11782 82399 -11682 82445 4 VDD
port 41 nsew
rlabel metal1 s -11083 82593 -10783 82639 4 VDD
port 41 nsew
rlabel metal1 s -12194 82649 -11594 82695 4 VDD
port 41 nsew
rlabel metal1 s -11084 82810 -10984 82856 4 VDD
port 41 nsew
rlabel metal1 s -12194 82845 -11594 82891 4 VDD
port 41 nsew
rlabel metal1 s -11084 83006 -10984 83052 4 VDD
port 41 nsew
rlabel metal1 s -11084 83202 -10984 83248 4 VDD
port 41 nsew
rlabel metal1 s -12194 83268 -11594 83314 4 VDD
port 41 nsew
rlabel metal1 s -11084 83398 -10984 83444 4 VDD
port 41 nsew
rlabel metal1 s -11500 83458 -11337 83549 4 VDD
port 41 nsew
rlabel metal1 s -11488 83549 -11349 83708 4 VDD
port 41 nsew
rlabel metal1 s -11513 83708 -11322 83859 4 VDD
port 41 nsew
rlabel metal1 s -7436 86766 -7236 86812 4 VDD
port 41 nsew
rlabel metal1 s -8465 86740 -8165 86786 4 VDD
port 41 nsew
rlabel metal1 s -10889 86758 -10689 86804 4 VDD
port 41 nsew
rlabel metal1 s -11918 86732 -11618 86778 4 VDD
port 41 nsew
rlabel metal1 s -7436 86962 -7236 87008 4 VDD
port 41 nsew
rlabel metal1 s -8465 86936 -8165 86982 4 VDD
port 41 nsew
rlabel metal1 s -10889 86954 -10689 87000 4 VDD
port 41 nsew
rlabel metal1 s -11918 86928 -11618 86974 4 VDD
port 41 nsew
rlabel metal1 s -7436 87158 -7236 87204 4 VDD
port 41 nsew
rlabel metal1 s -8465 87132 -8165 87178 4 VDD
port 41 nsew
rlabel metal1 s -10889 87150 -10689 87196 4 VDD
port 41 nsew
rlabel metal1 s -11918 87124 -11618 87170 4 VDD
port 41 nsew
rlabel metal1 s -7436 87354 -7236 87400 4 VDD
port 41 nsew
rlabel metal1 s -8264 87349 -8164 87395 4 VDD
port 41 nsew
rlabel metal1 s -10889 87346 -10689 87392 4 VDD
port 41 nsew
rlabel metal1 s -11717 87341 -11617 87387 4 VDD
port 41 nsew
rlabel metal1 s -8264 87545 -8164 87591 4 VDD
port 41 nsew
rlabel metal1 s -11717 87537 -11617 87583 4 VDD
port 41 nsew
rlabel metal1 s -7565 87739 -7265 87785 4 VDD
port 41 nsew
rlabel metal1 s -8264 87741 -8164 87787 4 VDD
port 41 nsew
rlabel metal1 s -11018 87731 -10718 87777 4 VDD
port 41 nsew
rlabel metal1 s -11717 87733 -11617 87779 4 VDD
port 41 nsew
rlabel metal1 s -7565 87935 -7265 87981 4 VDD
port 41 nsew
rlabel metal1 s -8264 87937 -8164 87983 4 VDD
port 41 nsew
rlabel metal1 s -11018 87927 -10718 87973 4 VDD
port 41 nsew
rlabel metal1 s -11382 87933 -11252 88116 4 VDD
port 41 nsew
rlabel metal1 s -11717 87929 -11617 87975 4 VDD
port 41 nsew
rlabel metal1 s -7565 88131 -7265 88177 4 VDD
port 41 nsew
rlabel metal1 s -11018 88123 -10718 88169 4 VDD
port 41 nsew
rlabel metal1 s -8676 88187 -8076 88233 4 VDD
port 41 nsew
rlabel metal1 s -7566 88348 -7466 88394 4 VDD
port 41 nsew
rlabel metal1 s -8676 88383 -8076 88429 4 VDD
port 41 nsew
rlabel metal1 s -11019 88340 -10919 88386 4 VDD
port 41 nsew
rlabel metal1 s -7566 88544 -7466 88590 4 VDD
port 41 nsew
rlabel metal1 s -11019 88536 -10919 88582 4 VDD
port 41 nsew
rlabel metal1 s -7566 88740 -7466 88786 4 VDD
port 41 nsew
rlabel metal1 s -11019 88732 -10919 88778 4 VDD
port 41 nsew
rlabel metal1 s -8676 88806 -8076 88852 4 VDD
port 41 nsew
rlabel metal1 s -7566 88936 -7466 88982 4 VDD
port 41 nsew
rlabel metal1 s -11019 88928 -10919 88974 4 VDD
port 41 nsew
rlabel metal1 s -7983 89018 -7865 89092 4 VDD
port 41 nsew
rlabel metal1 s -7977 89092 -7881 89246 4 VDD
port 41 nsew
rlabel metal1 s -11375 88116 -11293 89236 4 VDD
port 41 nsew
rlabel metal1 s -12129 88179 -11529 88225 4 VDD
port 41 nsew
rlabel metal1 s -12129 88375 -11529 88421 4 VDD
port 41 nsew
rlabel metal1 s -12129 88798 -11529 88844 4 VDD
port 41 nsew
rlabel metal1 s -7995 89246 -7845 89356 4 VDD
port 41 nsew
rlabel metal1 s -11401 89236 -11264 89332 4 VDD
port 41 nsew
rlabel metal1 s -8434 90179 -7934 90225 4 VDD
port 41 nsew
rlabel metal1 s -8434 90375 -7934 90421 4 VDD
port 41 nsew
rlabel metal1 s -10920 90426 -10720 90472 4 VDD
port 41 nsew
rlabel metal1 s -11949 90400 -11649 90446 4 VDD
port 41 nsew
rlabel metal1 s -10920 90622 -10720 90668 4 VDD
port 41 nsew
rlabel metal1 s -11949 90596 -11649 90642 4 VDD
port 41 nsew
rlabel metal1 s -10920 90818 -10720 90864 4 VDD
port 41 nsew
rlabel metal1 s -11949 90792 -11649 90838 4 VDD
port 41 nsew
rlabel metal1 s -8434 90970 -7934 91016 4 VDD
port 41 nsew
rlabel metal1 s -10920 91014 -10720 91060 4 VDD
port 41 nsew
rlabel metal1 s -11748 91009 -11648 91055 4 VDD
port 41 nsew
rlabel metal1 s -8434 91100 -7934 91146 4 VDD
port 41 nsew
rlabel metal1 s -11748 91205 -11648 91251 4 VDD
port 41 nsew
rlabel metal1 s -8234 91328 -7934 91374 4 VDD
port 41 nsew
rlabel metal1 s -11049 91399 -10749 91445 4 VDD
port 41 nsew
rlabel metal1 s -11748 91401 -11648 91447 4 VDD
port 41 nsew
rlabel metal1 s -8234 91524 -7934 91570 4 VDD
port 41 nsew
rlabel metal1 s -11049 91595 -10749 91641 4 VDD
port 41 nsew
rlabel metal1 s -11748 91597 -11648 91643 4 VDD
port 41 nsew
rlabel metal1 s -11049 91791 -10749 91837 4 VDD
port 41 nsew
rlabel metal1 s -12160 91847 -11560 91893 4 VDD
port 41 nsew
rlabel metal1 s -11050 92008 -10950 92054 4 VDD
port 41 nsew
rlabel metal1 s -12160 92043 -11560 92089 4 VDD
port 41 nsew
rlabel metal1 s -11050 92204 -10950 92250 4 VDD
port 41 nsew
rlabel metal1 s -11050 92400 -10950 92446 4 VDD
port 41 nsew
rlabel metal1 s -12160 92466 -11560 92512 4 VDD
port 41 nsew
rlabel metal1 s -11050 92596 -10950 92642 4 VDD
port 41 nsew
rlabel metal1 s -11466 92656 -11303 92747 4 VDD
port 41 nsew
rlabel metal1 s -11454 92747 -11315 92906 4 VDD
port 41 nsew
rlabel metal1 s -11479 92906 -11288 93057 4 VDD
port 41 nsew
rlabel metal1 s -7370 95520 -7170 95566 4 VDD
port 41 nsew
rlabel metal1 s -8399 95494 -8099 95540 4 VDD
port 41 nsew
rlabel metal1 s -10823 95512 -10623 95558 4 VDD
port 41 nsew
rlabel metal1 s -11852 95486 -11552 95532 4 VDD
port 41 nsew
rlabel metal1 s -7370 95716 -7170 95762 4 VDD
port 41 nsew
rlabel metal1 s -8399 95690 -8099 95736 4 VDD
port 41 nsew
rlabel metal1 s -10823 95708 -10623 95754 4 VDD
port 41 nsew
rlabel metal1 s -11852 95682 -11552 95728 4 VDD
port 41 nsew
rlabel metal1 s -7370 95912 -7170 95958 4 VDD
port 41 nsew
rlabel metal1 s -8399 95886 -8099 95932 4 VDD
port 41 nsew
rlabel metal1 s -10823 95904 -10623 95950 4 VDD
port 41 nsew
rlabel metal1 s -11852 95878 -11552 95924 4 VDD
port 41 nsew
rlabel metal1 s -7370 96108 -7170 96154 4 VDD
port 41 nsew
rlabel metal1 s -8198 96103 -8098 96149 4 VDD
port 41 nsew
rlabel metal1 s -10823 96100 -10623 96146 4 VDD
port 41 nsew
rlabel metal1 s -11651 96095 -11551 96141 4 VDD
port 41 nsew
rlabel metal1 s -8198 96299 -8098 96345 4 VDD
port 41 nsew
rlabel metal1 s -11651 96291 -11551 96337 4 VDD
port 41 nsew
rlabel metal1 s -7499 96493 -7199 96539 4 VDD
port 41 nsew
rlabel metal1 s -8198 96495 -8098 96541 4 VDD
port 41 nsew
rlabel metal1 s -10952 96485 -10652 96531 4 VDD
port 41 nsew
rlabel metal1 s -11651 96487 -11551 96533 4 VDD
port 41 nsew
rlabel metal1 s -7499 96689 -7199 96735 4 VDD
port 41 nsew
rlabel metal1 s -8198 96691 -8098 96737 4 VDD
port 41 nsew
rlabel metal1 s -10952 96681 -10652 96727 4 VDD
port 41 nsew
rlabel metal1 s -11316 96687 -11186 96870 4 VDD
port 41 nsew
rlabel metal1 s -11651 96683 -11551 96729 4 VDD
port 41 nsew
rlabel metal1 s -7499 96885 -7199 96931 4 VDD
port 41 nsew
rlabel metal1 s -10952 96877 -10652 96923 4 VDD
port 41 nsew
rlabel metal1 s -8610 96941 -8010 96987 4 VDD
port 41 nsew
rlabel metal1 s -7500 97102 -7400 97148 4 VDD
port 41 nsew
rlabel metal1 s -8610 97137 -8010 97183 4 VDD
port 41 nsew
rlabel metal1 s -10953 97094 -10853 97140 4 VDD
port 41 nsew
rlabel metal1 s -7500 97298 -7400 97344 4 VDD
port 41 nsew
rlabel metal1 s -10953 97290 -10853 97336 4 VDD
port 41 nsew
rlabel metal1 s -7500 97494 -7400 97540 4 VDD
port 41 nsew
rlabel metal1 s -10953 97486 -10853 97532 4 VDD
port 41 nsew
rlabel metal1 s -8610 97560 -8010 97606 4 VDD
port 41 nsew
rlabel metal1 s -7500 97690 -7400 97736 4 VDD
port 41 nsew
rlabel metal1 s -10953 97682 -10853 97728 4 VDD
port 41 nsew
rlabel metal1 s -7917 97772 -7799 97846 4 VDD
port 41 nsew
rlabel metal1 s -7911 97846 -7815 98000 4 VDD
port 41 nsew
rlabel metal1 s -11309 96870 -11227 97990 4 VDD
port 41 nsew
rlabel metal1 s -12063 96933 -11463 96979 4 VDD
port 41 nsew
rlabel metal1 s -12063 97129 -11463 97175 4 VDD
port 41 nsew
rlabel metal1 s -12063 97552 -11463 97598 4 VDD
port 41 nsew
rlabel metal1 s -7929 98000 -7779 98110 4 VDD
port 41 nsew
rlabel metal1 s -11335 97990 -11198 98086 4 VDD
port 41 nsew
rlabel metal1 s -8368 98933 -7868 98979 4 VDD
port 41 nsew
rlabel metal1 s -8368 99129 -7868 99175 4 VDD
port 41 nsew
rlabel metal1 s -10854 99180 -10654 99226 4 VDD
port 41 nsew
rlabel metal1 s -11883 99154 -11583 99200 4 VDD
port 41 nsew
rlabel metal1 s -10854 99376 -10654 99422 4 VDD
port 41 nsew
rlabel metal1 s -11883 99350 -11583 99396 4 VDD
port 41 nsew
rlabel metal1 s -10854 99572 -10654 99618 4 VDD
port 41 nsew
rlabel metal1 s -11883 99546 -11583 99592 4 VDD
port 41 nsew
rlabel metal1 s -8368 99724 -7868 99770 4 VDD
port 41 nsew
rlabel metal1 s -10854 99768 -10654 99814 4 VDD
port 41 nsew
rlabel metal1 s -11682 99763 -11582 99809 4 VDD
port 41 nsew
rlabel metal1 s -8368 99854 -7868 99900 4 VDD
port 41 nsew
rlabel metal1 s -11682 99959 -11582 100005 4 VDD
port 41 nsew
rlabel metal1 s -8168 100082 -7868 100128 4 VDD
port 41 nsew
rlabel metal1 s -10983 100153 -10683 100199 4 VDD
port 41 nsew
rlabel metal1 s -11682 100155 -11582 100201 4 VDD
port 41 nsew
rlabel metal1 s -8168 100278 -7868 100324 4 VDD
port 41 nsew
rlabel metal1 s -10983 100349 -10683 100395 4 VDD
port 41 nsew
rlabel metal1 s -11682 100351 -11582 100397 4 VDD
port 41 nsew
rlabel metal1 s -10983 100545 -10683 100591 4 VDD
port 41 nsew
rlabel metal1 s -12094 100601 -11494 100647 4 VDD
port 41 nsew
rlabel metal1 s -10984 100762 -10884 100808 4 VDD
port 41 nsew
rlabel metal1 s -12094 100797 -11494 100843 4 VDD
port 41 nsew
rlabel metal1 s -10984 100958 -10884 101004 4 VDD
port 41 nsew
rlabel metal1 s -10984 101154 -10884 101200 4 VDD
port 41 nsew
rlabel metal1 s -12094 101220 -11494 101266 4 VDD
port 41 nsew
rlabel metal1 s -10984 101350 -10884 101396 4 VDD
port 41 nsew
rlabel metal1 s -11400 101410 -11237 101501 4 VDD
port 41 nsew
rlabel metal1 s -11388 101501 -11249 101660 4 VDD
port 41 nsew
rlabel metal1 s -11413 101660 -11222 101811 4 VDD
port 41 nsew
rlabel metal1 s -7353 104673 -7153 104719 4 VDD
port 41 nsew
rlabel metal1 s -8382 104647 -8082 104693 4 VDD
port 41 nsew
rlabel metal1 s -10806 104665 -10606 104711 4 VDD
port 41 nsew
rlabel metal1 s -11835 104639 -11535 104685 4 VDD
port 41 nsew
rlabel metal1 s -7353 104869 -7153 104915 4 VDD
port 41 nsew
rlabel metal1 s -8382 104843 -8082 104889 4 VDD
port 41 nsew
rlabel metal1 s -10806 104861 -10606 104907 4 VDD
port 41 nsew
rlabel metal1 s -11835 104835 -11535 104881 4 VDD
port 41 nsew
rlabel metal1 s -7353 105065 -7153 105111 4 VDD
port 41 nsew
rlabel metal1 s -8382 105039 -8082 105085 4 VDD
port 41 nsew
rlabel metal1 s -10806 105057 -10606 105103 4 VDD
port 41 nsew
rlabel metal1 s -11835 105031 -11535 105077 4 VDD
port 41 nsew
rlabel metal1 s -7353 105261 -7153 105307 4 VDD
port 41 nsew
rlabel metal1 s -8181 105256 -8081 105302 4 VDD
port 41 nsew
rlabel metal1 s -10806 105253 -10606 105299 4 VDD
port 41 nsew
rlabel metal1 s -11634 105248 -11534 105294 4 VDD
port 41 nsew
rlabel metal1 s -8181 105452 -8081 105498 4 VDD
port 41 nsew
rlabel metal1 s -11634 105444 -11534 105490 4 VDD
port 41 nsew
rlabel metal1 s -7482 105646 -7182 105692 4 VDD
port 41 nsew
rlabel metal1 s -8181 105648 -8081 105694 4 VDD
port 41 nsew
rlabel metal1 s -10935 105638 -10635 105684 4 VDD
port 41 nsew
rlabel metal1 s -11634 105640 -11534 105686 4 VDD
port 41 nsew
rlabel metal1 s -7482 105842 -7182 105888 4 VDD
port 41 nsew
rlabel metal1 s -8181 105844 -8081 105890 4 VDD
port 41 nsew
rlabel metal1 s -10935 105834 -10635 105880 4 VDD
port 41 nsew
rlabel metal1 s -11299 105840 -11169 106023 4 VDD
port 41 nsew
rlabel metal1 s -11634 105836 -11534 105882 4 VDD
port 41 nsew
rlabel metal1 s -7482 106038 -7182 106084 4 VDD
port 41 nsew
rlabel metal1 s -10935 106030 -10635 106076 4 VDD
port 41 nsew
rlabel metal1 s -8593 106094 -7993 106140 4 VDD
port 41 nsew
rlabel metal1 s -7483 106255 -7383 106301 4 VDD
port 41 nsew
rlabel metal1 s -8593 106290 -7993 106336 4 VDD
port 41 nsew
rlabel metal1 s -10936 106247 -10836 106293 4 VDD
port 41 nsew
rlabel metal1 s -7483 106451 -7383 106497 4 VDD
port 41 nsew
rlabel metal1 s -10936 106443 -10836 106489 4 VDD
port 41 nsew
rlabel metal1 s -7483 106647 -7383 106693 4 VDD
port 41 nsew
rlabel metal1 s -10936 106639 -10836 106685 4 VDD
port 41 nsew
rlabel metal1 s -8593 106713 -7993 106759 4 VDD
port 41 nsew
rlabel metal1 s -7483 106843 -7383 106889 4 VDD
port 41 nsew
rlabel metal1 s -10936 106835 -10836 106881 4 VDD
port 41 nsew
rlabel metal1 s -7900 106925 -7782 106999 4 VDD
port 41 nsew
rlabel metal1 s -7894 106999 -7798 107153 4 VDD
port 41 nsew
rlabel metal1 s -11292 106023 -11210 107143 4 VDD
port 41 nsew
rlabel metal1 s -12046 106086 -11446 106132 4 VDD
port 41 nsew
rlabel metal1 s -12046 106282 -11446 106328 4 VDD
port 41 nsew
rlabel metal1 s -12046 106705 -11446 106751 4 VDD
port 41 nsew
rlabel metal1 s -7912 107153 -7762 107263 4 VDD
port 41 nsew
rlabel metal1 s -11318 107143 -11181 107239 4 VDD
port 41 nsew
rlabel metal1 s -8351 108086 -7851 108132 4 VDD
port 41 nsew
rlabel metal1 s -8351 108282 -7851 108328 4 VDD
port 41 nsew
rlabel metal1 s -10837 108333 -10637 108379 4 VDD
port 41 nsew
rlabel metal1 s -11866 108307 -11566 108353 4 VDD
port 41 nsew
rlabel metal1 s -10837 108529 -10637 108575 4 VDD
port 41 nsew
rlabel metal1 s -11866 108503 -11566 108549 4 VDD
port 41 nsew
rlabel metal1 s -10837 108725 -10637 108771 4 VDD
port 41 nsew
rlabel metal1 s -11866 108699 -11566 108745 4 VDD
port 41 nsew
rlabel metal1 s -8351 108877 -7851 108923 4 VDD
port 41 nsew
rlabel metal1 s -10837 108921 -10637 108967 4 VDD
port 41 nsew
rlabel metal1 s -11665 108916 -11565 108962 4 VDD
port 41 nsew
rlabel metal1 s -8351 109007 -7851 109053 4 VDD
port 41 nsew
rlabel metal1 s -11665 109112 -11565 109158 4 VDD
port 41 nsew
rlabel metal1 s -8151 109235 -7851 109281 4 VDD
port 41 nsew
rlabel metal1 s -10966 109306 -10666 109352 4 VDD
port 41 nsew
rlabel metal1 s -11665 109308 -11565 109354 4 VDD
port 41 nsew
rlabel metal1 s -8151 109431 -7851 109477 4 VDD
port 41 nsew
rlabel metal1 s -10966 109502 -10666 109548 4 VDD
port 41 nsew
rlabel metal1 s -11665 109504 -11565 109550 4 VDD
port 41 nsew
rlabel metal1 s -10966 109698 -10666 109744 4 VDD
port 41 nsew
rlabel metal1 s -12077 109754 -11477 109800 4 VDD
port 41 nsew
rlabel metal1 s -10967 109915 -10867 109961 4 VDD
port 41 nsew
rlabel metal1 s -12077 109950 -11477 109996 4 VDD
port 41 nsew
rlabel metal1 s -10967 110111 -10867 110157 4 VDD
port 41 nsew
rlabel metal1 s -10967 110307 -10867 110353 4 VDD
port 41 nsew
rlabel metal1 s -12077 110373 -11477 110419 4 VDD
port 41 nsew
rlabel metal1 s -10967 110503 -10867 110549 4 VDD
port 41 nsew
rlabel metal1 s -11383 110563 -11220 110654 4 VDD
port 41 nsew
rlabel metal1 s -11371 110654 -11232 110813 4 VDD
port 41 nsew
rlabel metal1 s -11396 110813 -11205 110964 4 VDD
port 41 nsew
rlabel metal1 s -7315 114037 -7115 114083 4 VDD
port 41 nsew
rlabel metal1 s -8344 114011 -8044 114057 4 VDD
port 41 nsew
rlabel metal1 s -10768 114029 -10568 114075 4 VDD
port 41 nsew
rlabel metal1 s -11797 114003 -11497 114049 4 VDD
port 41 nsew
rlabel metal1 s -7315 114233 -7115 114279 4 VDD
port 41 nsew
rlabel metal1 s -8344 114207 -8044 114253 4 VDD
port 41 nsew
rlabel metal1 s -10768 114225 -10568 114271 4 VDD
port 41 nsew
rlabel metal1 s -11797 114199 -11497 114245 4 VDD
port 41 nsew
rlabel metal1 s -7315 114429 -7115 114475 4 VDD
port 41 nsew
rlabel metal1 s -8344 114403 -8044 114449 4 VDD
port 41 nsew
rlabel metal1 s -10768 114421 -10568 114467 4 VDD
port 41 nsew
rlabel metal1 s -11797 114395 -11497 114441 4 VDD
port 41 nsew
rlabel metal1 s -7315 114625 -7115 114671 4 VDD
port 41 nsew
rlabel metal1 s -8143 114620 -8043 114666 4 VDD
port 41 nsew
rlabel metal1 s -10768 114617 -10568 114663 4 VDD
port 41 nsew
rlabel metal1 s -11596 114612 -11496 114658 4 VDD
port 41 nsew
rlabel metal1 s -8143 114816 -8043 114862 4 VDD
port 41 nsew
rlabel metal1 s -11596 114808 -11496 114854 4 VDD
port 41 nsew
rlabel metal1 s -7444 115010 -7144 115056 4 VDD
port 41 nsew
rlabel metal1 s -8143 115012 -8043 115058 4 VDD
port 41 nsew
rlabel metal1 s -10897 115002 -10597 115048 4 VDD
port 41 nsew
rlabel metal1 s -11596 115004 -11496 115050 4 VDD
port 41 nsew
rlabel metal1 s -7444 115206 -7144 115252 4 VDD
port 41 nsew
rlabel metal1 s -8143 115208 -8043 115254 4 VDD
port 41 nsew
rlabel metal1 s -10897 115198 -10597 115244 4 VDD
port 41 nsew
rlabel metal1 s -11261 115204 -11131 115387 4 VDD
port 41 nsew
rlabel metal1 s -11596 115200 -11496 115246 4 VDD
port 41 nsew
rlabel metal1 s -7444 115402 -7144 115448 4 VDD
port 41 nsew
rlabel metal1 s -10897 115394 -10597 115440 4 VDD
port 41 nsew
rlabel metal1 s -8555 115458 -7955 115504 4 VDD
port 41 nsew
rlabel metal1 s -7445 115619 -7345 115665 4 VDD
port 41 nsew
rlabel metal1 s -8555 115654 -7955 115700 4 VDD
port 41 nsew
rlabel metal1 s -10898 115611 -10798 115657 4 VDD
port 41 nsew
rlabel metal1 s -7445 115815 -7345 115861 4 VDD
port 41 nsew
rlabel metal1 s -10898 115807 -10798 115853 4 VDD
port 41 nsew
rlabel metal1 s -7445 116011 -7345 116057 4 VDD
port 41 nsew
rlabel metal1 s -10898 116003 -10798 116049 4 VDD
port 41 nsew
rlabel metal1 s -8555 116077 -7955 116123 4 VDD
port 41 nsew
rlabel metal1 s -7445 116207 -7345 116253 4 VDD
port 41 nsew
rlabel metal1 s -10898 116199 -10798 116245 4 VDD
port 41 nsew
rlabel metal1 s -7862 116289 -7744 116363 4 VDD
port 41 nsew
rlabel metal1 s -7856 116363 -7760 116517 4 VDD
port 41 nsew
rlabel metal1 s -11254 115387 -11172 116507 4 VDD
port 41 nsew
rlabel metal1 s -12008 115450 -11408 115496 4 VDD
port 41 nsew
rlabel metal1 s -12008 115646 -11408 115692 4 VDD
port 41 nsew
rlabel metal1 s -12008 116069 -11408 116115 4 VDD
port 41 nsew
rlabel metal1 s -7874 116517 -7724 116627 4 VDD
port 41 nsew
rlabel metal1 s -11280 116507 -11143 116603 4 VDD
port 41 nsew
rlabel metal1 s -8313 117450 -7813 117496 4 VDD
port 41 nsew
rlabel metal1 s -8313 117646 -7813 117692 4 VDD
port 41 nsew
rlabel metal1 s -10799 117697 -10599 117743 4 VDD
port 41 nsew
rlabel metal1 s -11828 117671 -11528 117717 4 VDD
port 41 nsew
rlabel metal1 s -10799 117893 -10599 117939 4 VDD
port 41 nsew
rlabel metal1 s -11828 117867 -11528 117913 4 VDD
port 41 nsew
rlabel metal1 s -10799 118089 -10599 118135 4 VDD
port 41 nsew
rlabel metal1 s -11828 118063 -11528 118109 4 VDD
port 41 nsew
rlabel metal1 s -8313 118241 -7813 118287 4 VDD
port 41 nsew
rlabel metal1 s -10799 118285 -10599 118331 4 VDD
port 41 nsew
rlabel metal1 s -11627 118280 -11527 118326 4 VDD
port 41 nsew
rlabel metal1 s -8313 118371 -7813 118417 4 VDD
port 41 nsew
rlabel metal1 s -11627 118476 -11527 118522 4 VDD
port 41 nsew
rlabel metal1 s -8113 118599 -7813 118645 4 VDD
port 41 nsew
rlabel metal1 s -10928 118670 -10628 118716 4 VDD
port 41 nsew
rlabel metal1 s -11627 118672 -11527 118718 4 VDD
port 41 nsew
rlabel metal1 s -8113 118795 -7813 118841 4 VDD
port 41 nsew
rlabel metal1 s -10928 118866 -10628 118912 4 VDD
port 41 nsew
rlabel metal1 s -11627 118868 -11527 118914 4 VDD
port 41 nsew
rlabel metal1 s -10928 119062 -10628 119108 4 VDD
port 41 nsew
rlabel metal1 s -12039 119118 -11439 119164 4 VDD
port 41 nsew
rlabel metal1 s -10929 119279 -10829 119325 4 VDD
port 41 nsew
rlabel metal1 s -12039 119314 -11439 119360 4 VDD
port 41 nsew
rlabel metal1 s -10929 119475 -10829 119521 4 VDD
port 41 nsew
rlabel metal1 s -10929 119671 -10829 119717 4 VDD
port 41 nsew
rlabel metal1 s -12039 119737 -11439 119783 4 VDD
port 41 nsew
rlabel metal1 s -10929 119867 -10829 119913 4 VDD
port 41 nsew
rlabel metal1 s -11345 119927 -11182 120018 4 VDD
port 41 nsew
rlabel metal1 s -11333 120018 -11194 120177 4 VDD
port 41 nsew
rlabel metal1 s -11358 120177 -11167 120328 4 VDD
port 41 nsew
rlabel locali s -6133 -62451 8829 -62258 8 VDD
port 41 nsew
rlabel locali s -21374 -62293 -18772 -62284 2 VDD
port 41 nsew
rlabel locali s 7732 -62258 8784 -62151 8 VDD
port 41 nsew
rlabel locali s 5009 -62258 5602 -62220 8 VDD
port 41 nsew
rlabel locali s 2596 -62258 3189 -62220 8 VDD
port 41 nsew
rlabel locali s 12846 -62035 18071 -61972 8 VDD
port 41 nsew
rlabel locali s 8738 -62151 8784 -62029 8 VDD
port 41 nsew
rlabel locali s 16498 -61972 18071 -61967 8 VDD
port 41 nsew
rlabel locali s 13798 -61972 15600 -61967 8 VDD
port 41 nsew
rlabel locali s 87831 -60276 87865 -59684 8 VDD
port 41 nsew
rlabel locali s 88271 -59579 88410 -59551 8 VDD
port 41 nsew
rlabel locali s 88271 -59551 88483 -59412 8 VDD
port 41 nsew
rlabel locali s 88021 -59566 88100 -59541 8 VDD
port 41 nsew
rlabel locali s 87824 -59684 87869 -59560 8 VDD
port 41 nsew
rlabel locali s 87408 -60276 87442 -59683 8 VDD
port 41 nsew
rlabel locali s 87212 -60276 87246 -59686 8 VDD
port 41 nsew
rlabel locali s 86962 -59864 86996 -59698 8 VDD
port 41 nsew
rlabel locali s 86766 -59864 86800 -59698 8 VDD
port 41 nsew
rlabel locali s 86570 -59864 86604 -59698 8 VDD
port 41 nsew
rlabel locali s 86374 -59864 86408 -59698 8 VDD
port 41 nsew
rlabel locali s 86157 -60065 86191 -59698 8 VDD
port 41 nsew
rlabel locali s 87402 -59683 87447 -59560 8 VDD
port 41 nsew
rlabel locali s 87207 -59686 87252 -59560 8 VDD
port 41 nsew
rlabel locali s 86157 -59698 87044 -59648 8 VDD
port 41 nsew
rlabel locali s 85961 -60065 85995 -59648 8 VDD
port 41 nsew
rlabel locali s 85765 -60065 85799 -59648 8 VDD
port 41 nsew
rlabel locali s 84163 -60245 84197 -59653 8 VDD
port 41 nsew
rlabel locali s 85755 -59648 87044 -59599 8 VDD
port 41 nsew
rlabel locali s 85755 -59599 86197 -59584 8 VDD
port 41 nsew
rlabel locali s 87201 -59560 87970 -59541 8 VDD
port 41 nsew
rlabel locali s 87201 -59541 88100 -59536 8 VDD
port 41 nsew
rlabel locali s 86194 -59550 86383 -59543 8 VDD
port 41 nsew
rlabel locali s 86157 -59543 86383 -59536 8 VDD
port 41 nsew
rlabel locali s 85755 -59536 88100 -59494 8 VDD
port 41 nsew
rlabel locali s 84156 -59653 84201 -59529 8 VDD
port 41 nsew
rlabel locali s 83740 -60245 83774 -59652 8 VDD
port 41 nsew
rlabel locali s 83544 -60245 83578 -59655 8 VDD
port 41 nsew
rlabel locali s 83294 -59833 83328 -59667 8 VDD
port 41 nsew
rlabel locali s 83098 -59833 83132 -59667 8 VDD
port 41 nsew
rlabel locali s 82902 -59833 82936 -59667 8 VDD
port 41 nsew
rlabel locali s 82706 -59833 82740 -59667 8 VDD
port 41 nsew
rlabel locali s 82489 -60034 82523 -59667 8 VDD
port 41 nsew
rlabel locali s 83734 -59652 83779 -59529 8 VDD
port 41 nsew
rlabel locali s 83539 -59655 83584 -59529 8 VDD
port 41 nsew
rlabel locali s 82489 -59667 83376 -59617 8 VDD
port 41 nsew
rlabel locali s 82293 -60034 82327 -59617 8 VDD
port 41 nsew
rlabel locali s 82097 -60034 82131 -59617 8 VDD
port 41 nsew
rlabel locali s 78467 -60314 78501 -59722 8 VDD
port 41 nsew
rlabel locali s 82087 -59617 83376 -59568 8 VDD
port 41 nsew
rlabel locali s 78907 -59617 79046 -59589 8 VDD
port 41 nsew
rlabel locali s 82087 -59568 82529 -59553 8 VDD
port 41 nsew
rlabel locali s 83533 -59529 84302 -59505 8 VDD
port 41 nsew
rlabel locali s 82526 -59519 82715 -59512 8 VDD
port 41 nsew
rlabel locali s 82489 -59512 82715 -59505 8 VDD
port 41 nsew
rlabel locali s 87921 -59494 88100 -59458 8 VDD
port 41 nsew
rlabel locali s 85755 -59494 87866 -59483 8 VDD
port 41 nsew
rlabel locali s 88021 -59458 88100 -59427 8 VDD
port 41 nsew
rlabel locali s 84954 -59483 87866 -59417 8 VDD
port 41 nsew
rlabel locali s 88361 -59412 88483 -58416 8 VDD
port 41 nsew
rlabel locali s 85755 -59417 87866 -59383 8 VDD
port 41 nsew
rlabel locali s 86753 -59383 87371 -59366 8 VDD
port 41 nsew
rlabel locali s 86753 -59366 87196 -59337 8 VDD
port 41 nsew
rlabel locali s 86754 -59337 87196 -59323 8 VDD
port 41 nsew
rlabel locali s 86754 -59323 88043 -59274 8 VDD
port 41 nsew
rlabel locali s 87156 -59274 88043 -59224 8 VDD
port 41 nsew
rlabel locali s 87961 -59224 87995 -59058 8 VDD
port 41 nsew
rlabel locali s 87765 -59224 87799 -59058 8 VDD
port 41 nsew
rlabel locali s 87569 -59224 87603 -59058 8 VDD
port 41 nsew
rlabel locali s 87373 -59224 87407 -59058 8 VDD
port 41 nsew
rlabel locali s 87156 -59224 87190 -58857 8 VDD
port 41 nsew
rlabel locali s 86960 -59274 86994 -58857 8 VDD
port 41 nsew
rlabel locali s 86764 -59274 86798 -58857 8 VDD
port 41 nsew
rlabel locali s 85925 -59383 86097 -59193 8 VDD
port 41 nsew
rlabel locali s 85743 -59193 86461 -59094 8 VDD
port 41 nsew
rlabel locali s 86379 -59094 86413 -58828 8 VDD
port 41 nsew
rlabel locali s 86183 -59094 86217 -58828 8 VDD
port 41 nsew
rlabel locali s 85987 -59094 86021 -58828 8 VDD
port 41 nsew
rlabel locali s 85791 -59094 85825 -58828 8 VDD
port 41 nsew
rlabel locali s 87851 -58416 88483 -58294 8 VDD
port 41 nsew
rlabel locali s 87851 -58294 87973 -55897 8 VDD
port 41 nsew
rlabel locali s 84954 -59417 85020 -58087 8 VDD
port 41 nsew
rlabel locali s 84601 -59501 84685 -59388 8 VDD
port 41 nsew
rlabel locali s 82087 -59505 84302 -59463 8 VDD
port 41 nsew
rlabel locali s 84618 -59388 84684 -58087 8 VDD
port 41 nsew
rlabel locali s 82087 -59463 84198 -59352 8 VDD
port 41 nsew
rlabel locali s 78907 -59589 79119 -59450 8 VDD
port 41 nsew
rlabel locali s 78657 -59604 78736 -59579 8 VDD
port 41 nsew
rlabel locali s 78460 -59722 78505 -59598 8 VDD
port 41 nsew
rlabel locali s 78044 -60314 78078 -59721 8 VDD
port 41 nsew
rlabel locali s 77848 -60314 77882 -59724 8 VDD
port 41 nsew
rlabel locali s 77598 -59902 77632 -59736 8 VDD
port 41 nsew
rlabel locali s 77402 -59902 77436 -59736 8 VDD
port 41 nsew
rlabel locali s 77206 -59902 77240 -59736 8 VDD
port 41 nsew
rlabel locali s 77010 -59902 77044 -59736 8 VDD
port 41 nsew
rlabel locali s 76793 -60103 76827 -59736 8 VDD
port 41 nsew
rlabel locali s 78038 -59721 78083 -59598 8 VDD
port 41 nsew
rlabel locali s 77843 -59724 77888 -59598 8 VDD
port 41 nsew
rlabel locali s 76793 -59736 77680 -59686 8 VDD
port 41 nsew
rlabel locali s 76597 -60103 76631 -59686 8 VDD
port 41 nsew
rlabel locali s 76401 -60103 76435 -59686 8 VDD
port 41 nsew
rlabel locali s 74799 -60283 74833 -59691 8 VDD
port 41 nsew
rlabel locali s 76391 -59686 77680 -59637 8 VDD
port 41 nsew
rlabel locali s 76391 -59637 76833 -59622 8 VDD
port 41 nsew
rlabel locali s 77837 -59598 78606 -59579 8 VDD
port 41 nsew
rlabel locali s 77837 -59579 78736 -59574 8 VDD
port 41 nsew
rlabel locali s 76830 -59588 77019 -59581 8 VDD
port 41 nsew
rlabel locali s 76793 -59581 77019 -59574 8 VDD
port 41 nsew
rlabel locali s 76391 -59574 78736 -59532 8 VDD
port 41 nsew
rlabel locali s 74792 -59691 74837 -59567 8 VDD
port 41 nsew
rlabel locali s 74376 -60283 74410 -59690 8 VDD
port 41 nsew
rlabel locali s 74180 -60283 74214 -59693 8 VDD
port 41 nsew
rlabel locali s 73930 -59871 73964 -59705 8 VDD
port 41 nsew
rlabel locali s 73734 -59871 73768 -59705 8 VDD
port 41 nsew
rlabel locali s 73538 -59871 73572 -59705 8 VDD
port 41 nsew
rlabel locali s 73342 -59871 73376 -59705 8 VDD
port 41 nsew
rlabel locali s 73125 -60072 73159 -59705 8 VDD
port 41 nsew
rlabel locali s 74370 -59690 74415 -59567 8 VDD
port 41 nsew
rlabel locali s 74175 -59693 74220 -59567 8 VDD
port 41 nsew
rlabel locali s 73125 -59705 74012 -59655 8 VDD
port 41 nsew
rlabel locali s 72929 -60072 72963 -59655 8 VDD
port 41 nsew
rlabel locali s 72733 -60072 72767 -59655 8 VDD
port 41 nsew
rlabel locali s 69314 -60331 69348 -59739 8 VDD
port 41 nsew
rlabel locali s 72723 -59655 74012 -59606 8 VDD
port 41 nsew
rlabel locali s 69754 -59634 69893 -59606 8 VDD
port 41 nsew
rlabel locali s 72723 -59606 73165 -59591 8 VDD
port 41 nsew
rlabel locali s 74169 -59567 74938 -59543 8 VDD
port 41 nsew
rlabel locali s 73162 -59557 73351 -59550 8 VDD
port 41 nsew
rlabel locali s 73125 -59550 73351 -59543 8 VDD
port 41 nsew
rlabel locali s 78557 -59532 78736 -59496 8 VDD
port 41 nsew
rlabel locali s 76391 -59532 78502 -59521 8 VDD
port 41 nsew
rlabel locali s 78657 -59496 78736 -59465 8 VDD
port 41 nsew
rlabel locali s 75590 -59521 78502 -59455 8 VDD
port 41 nsew
rlabel locali s 83085 -59352 83703 -59335 8 VDD
port 41 nsew
rlabel locali s 83085 -59335 83528 -59306 8 VDD
port 41 nsew
rlabel locali s 83086 -59306 83528 -59292 8 VDD
port 41 nsew
rlabel locali s 83086 -59292 84375 -59243 8 VDD
port 41 nsew
rlabel locali s 83488 -59243 84375 -59193 8 VDD
port 41 nsew
rlabel locali s 84293 -59193 84327 -59027 8 VDD
port 41 nsew
rlabel locali s 84097 -59193 84131 -59027 8 VDD
port 41 nsew
rlabel locali s 83901 -59193 83935 -59027 8 VDD
port 41 nsew
rlabel locali s 83705 -59193 83739 -59027 8 VDD
port 41 nsew
rlabel locali s 83488 -59193 83522 -58826 8 VDD
port 41 nsew
rlabel locali s 83292 -59243 83326 -58826 8 VDD
port 41 nsew
rlabel locali s 83096 -59243 83130 -58826 8 VDD
port 41 nsew
rlabel locali s 82257 -59352 82429 -59162 8 VDD
port 41 nsew
rlabel locali s 82075 -59162 82793 -59063 8 VDD
port 41 nsew
rlabel locali s 82711 -59063 82745 -58797 8 VDD
port 41 nsew
rlabel locali s 82515 -59063 82549 -58797 8 VDD
port 41 nsew
rlabel locali s 82319 -59063 82353 -58797 8 VDD
port 41 nsew
rlabel locali s 82123 -59063 82157 -58797 8 VDD
port 41 nsew
rlabel locali s 78997 -59450 79119 -58454 8 VDD
port 41 nsew
rlabel locali s 76391 -59455 78502 -59421 8 VDD
port 41 nsew
rlabel locali s 77389 -59421 78007 -59404 8 VDD
port 41 nsew
rlabel locali s 77389 -59404 77832 -59375 8 VDD
port 41 nsew
rlabel locali s 77390 -59375 77832 -59361 8 VDD
port 41 nsew
rlabel locali s 77390 -59361 78679 -59312 8 VDD
port 41 nsew
rlabel locali s 77792 -59312 78679 -59262 8 VDD
port 41 nsew
rlabel locali s 78597 -59262 78631 -59096 8 VDD
port 41 nsew
rlabel locali s 78401 -59262 78435 -59096 8 VDD
port 41 nsew
rlabel locali s 78205 -59262 78239 -59096 8 VDD
port 41 nsew
rlabel locali s 78009 -59262 78043 -59096 8 VDD
port 41 nsew
rlabel locali s 77792 -59262 77826 -58895 8 VDD
port 41 nsew
rlabel locali s 77596 -59312 77630 -58895 8 VDD
port 41 nsew
rlabel locali s 77400 -59312 77434 -58895 8 VDD
port 41 nsew
rlabel locali s 76561 -59421 76733 -59231 8 VDD
port 41 nsew
rlabel locali s 76379 -59231 77097 -59132 8 VDD
port 41 nsew
rlabel locali s 77015 -59132 77049 -58866 8 VDD
port 41 nsew
rlabel locali s 76819 -59132 76853 -58866 8 VDD
port 41 nsew
rlabel locali s 76623 -59132 76657 -58866 8 VDD
port 41 nsew
rlabel locali s 76427 -59132 76461 -58866 8 VDD
port 41 nsew
rlabel locali s 78487 -58454 79119 -58332 8 VDD
port 41 nsew
rlabel locali s 84618 -58087 85020 -58021 8 VDD
port 41 nsew
rlabel locali s 86889 -56350 86923 -56058 8 VDD
port 41 nsew
rlabel locali s 86693 -56350 86727 -56060 8 VDD
port 41 nsew
rlabel locali s 86465 -56550 86499 -56075 8 VDD
port 41 nsew
rlabel locali s 86335 -56550 86369 -56078 8 VDD
port 41 nsew
rlabel locali s 86884 -56058 86927 -55898 8 VDD
port 41 nsew
rlabel locali s 86687 -56060 86730 -55898 8 VDD
port 41 nsew
rlabel locali s 86456 -56075 86506 -55898 8 VDD
port 41 nsew
rlabel locali s 86330 -56078 86380 -55898 8 VDD
port 41 nsew
rlabel locali s 85740 -56550 85774 -56055 8 VDD
port 41 nsew
rlabel locali s 85544 -56550 85578 -56057 8 VDD
port 41 nsew
rlabel locali s 84171 -56792 84205 -56200 8 VDD
port 41 nsew
rlabel locali s 84611 -56095 84709 -56089 8 VDD
port 41 nsew
rlabel locali s 85738 -56055 85776 -55898 8 VDD
port 41 nsew
rlabel locali s 85541 -56057 85579 -55962 8 VDD
port 41 nsew
rlabel locali s 84611 -56089 85291 -55972 8 VDD
port 41 nsew
rlabel locali s 84383 -56083 84445 -56069 8 VDD
port 41 nsew
rlabel locali s 84164 -56200 84209 -56076 8 VDD
port 41 nsew
rlabel locali s 83748 -56792 83782 -56199 8 VDD
port 41 nsew
rlabel locali s 83552 -56792 83586 -56202 8 VDD
port 41 nsew
rlabel locali s 83302 -56380 83336 -56214 8 VDD
port 41 nsew
rlabel locali s 83106 -56380 83140 -56214 8 VDD
port 41 nsew
rlabel locali s 82910 -56380 82944 -56214 8 VDD
port 41 nsew
rlabel locali s 82714 -56380 82748 -56214 8 VDD
port 41 nsew
rlabel locali s 82497 -56581 82531 -56214 8 VDD
port 41 nsew
rlabel locali s 83742 -56199 83787 -56076 8 VDD
port 41 nsew
rlabel locali s 83547 -56202 83592 -56076 8 VDD
port 41 nsew
rlabel locali s 82497 -56214 83384 -56164 8 VDD
port 41 nsew
rlabel locali s 82301 -56581 82335 -56164 8 VDD
port 41 nsew
rlabel locali s 82105 -56581 82139 -56164 8 VDD
port 41 nsew
rlabel locali s 82095 -56164 83384 -56115 8 VDD
port 41 nsew
rlabel locali s 82095 -56115 82537 -56100 8 VDD
port 41 nsew
rlabel locali s 83541 -56076 84310 -56069 8 VDD
port 41 nsew
rlabel locali s 83541 -56069 84445 -56052 8 VDD
port 41 nsew
rlabel locali s 82534 -56066 82723 -56059 8 VDD
port 41 nsew
rlabel locali s 82497 -56059 82723 -56052 8 VDD
port 41 nsew
rlabel locali s 82095 -56052 84445 -56017 8 VDD
port 41 nsew
rlabel locali s 84383 -56017 84445 -55989 8 VDD
port 41 nsew
rlabel locali s 82095 -56017 84310 -56010 8 VDD
port 41 nsew
rlabel locali s 82095 -56010 84206 -55996 8 VDD
port 41 nsew
rlabel locali s 78487 -58332 78609 -55996 8 VDD
port 41 nsew
rlabel locali s 75590 -59455 75656 -58125 8 VDD
port 41 nsew
rlabel locali s 75237 -59539 75321 -59426 8 VDD
port 41 nsew
rlabel locali s 72723 -59543 74938 -59501 8 VDD
port 41 nsew
rlabel locali s 75254 -59426 75320 -58125 8 VDD
port 41 nsew
rlabel locali s 72723 -59501 74834 -59390 8 VDD
port 41 nsew
rlabel locali s 69754 -59606 69966 -59467 8 VDD
port 41 nsew
rlabel locali s 69504 -59621 69583 -59596 8 VDD
port 41 nsew
rlabel locali s 69307 -59739 69352 -59615 8 VDD
port 41 nsew
rlabel locali s 68891 -60331 68925 -59738 8 VDD
port 41 nsew
rlabel locali s 68695 -60331 68729 -59741 8 VDD
port 41 nsew
rlabel locali s 68445 -59919 68479 -59753 8 VDD
port 41 nsew
rlabel locali s 68249 -59919 68283 -59753 8 VDD
port 41 nsew
rlabel locali s 68053 -59919 68087 -59753 8 VDD
port 41 nsew
rlabel locali s 67857 -59919 67891 -59753 8 VDD
port 41 nsew
rlabel locali s 67640 -60120 67674 -59753 8 VDD
port 41 nsew
rlabel locali s 68885 -59738 68930 -59615 8 VDD
port 41 nsew
rlabel locali s 68690 -59741 68735 -59615 8 VDD
port 41 nsew
rlabel locali s 67640 -59753 68527 -59703 8 VDD
port 41 nsew
rlabel locali s 67444 -60120 67478 -59703 8 VDD
port 41 nsew
rlabel locali s 67248 -60120 67282 -59703 8 VDD
port 41 nsew
rlabel locali s 65646 -60300 65680 -59708 8 VDD
port 41 nsew
rlabel locali s 67238 -59703 68527 -59654 8 VDD
port 41 nsew
rlabel locali s 67238 -59654 67680 -59639 8 VDD
port 41 nsew
rlabel locali s 68684 -59615 69453 -59596 8 VDD
port 41 nsew
rlabel locali s 68684 -59596 69583 -59591 8 VDD
port 41 nsew
rlabel locali s 67677 -59605 67866 -59598 8 VDD
port 41 nsew
rlabel locali s 67640 -59598 67866 -59591 8 VDD
port 41 nsew
rlabel locali s 67238 -59591 69583 -59549 8 VDD
port 41 nsew
rlabel locali s 65639 -59708 65684 -59584 8 VDD
port 41 nsew
rlabel locali s 65223 -60300 65257 -59707 8 VDD
port 41 nsew
rlabel locali s 65027 -60300 65061 -59710 8 VDD
port 41 nsew
rlabel locali s 64777 -59888 64811 -59722 8 VDD
port 41 nsew
rlabel locali s 64581 -59888 64615 -59722 8 VDD
port 41 nsew
rlabel locali s 64385 -59888 64419 -59722 8 VDD
port 41 nsew
rlabel locali s 64189 -59888 64223 -59722 8 VDD
port 41 nsew
rlabel locali s 63972 -60089 64006 -59722 8 VDD
port 41 nsew
rlabel locali s 65217 -59707 65262 -59584 8 VDD
port 41 nsew
rlabel locali s 65022 -59710 65067 -59584 8 VDD
port 41 nsew
rlabel locali s 63972 -59722 64859 -59672 8 VDD
port 41 nsew
rlabel locali s 63776 -60089 63810 -59672 8 VDD
port 41 nsew
rlabel locali s 63580 -60089 63614 -59672 8 VDD
port 41 nsew
rlabel locali s 60560 -60397 60594 -59805 8 VDD
port 41 nsew
rlabel locali s 61000 -59700 61139 -59672 8 VDD
port 41 nsew
rlabel locali s 63570 -59672 64859 -59623 8 VDD
port 41 nsew
rlabel locali s 63570 -59623 64012 -59608 8 VDD
port 41 nsew
rlabel locali s 65016 -59584 65785 -59560 8 VDD
port 41 nsew
rlabel locali s 64009 -59574 64198 -59567 8 VDD
port 41 nsew
rlabel locali s 63972 -59567 64198 -59560 8 VDD
port 41 nsew
rlabel locali s 69404 -59549 69583 -59513 8 VDD
port 41 nsew
rlabel locali s 67238 -59549 69349 -59538 8 VDD
port 41 nsew
rlabel locali s 69504 -59513 69583 -59482 8 VDD
port 41 nsew
rlabel locali s 66437 -59538 69349 -59472 8 VDD
port 41 nsew
rlabel locali s 73721 -59390 74339 -59373 8 VDD
port 41 nsew
rlabel locali s 73721 -59373 74164 -59344 8 VDD
port 41 nsew
rlabel locali s 73722 -59344 74164 -59330 8 VDD
port 41 nsew
rlabel locali s 73722 -59330 75011 -59281 8 VDD
port 41 nsew
rlabel locali s 74124 -59281 75011 -59231 8 VDD
port 41 nsew
rlabel locali s 74929 -59231 74963 -59065 8 VDD
port 41 nsew
rlabel locali s 74733 -59231 74767 -59065 8 VDD
port 41 nsew
rlabel locali s 74537 -59231 74571 -59065 8 VDD
port 41 nsew
rlabel locali s 74341 -59231 74375 -59065 8 VDD
port 41 nsew
rlabel locali s 74124 -59231 74158 -58864 8 VDD
port 41 nsew
rlabel locali s 73928 -59281 73962 -58864 8 VDD
port 41 nsew
rlabel locali s 73732 -59281 73766 -58864 8 VDD
port 41 nsew
rlabel locali s 72893 -59390 73065 -59200 8 VDD
port 41 nsew
rlabel locali s 72711 -59200 73429 -59101 8 VDD
port 41 nsew
rlabel locali s 73347 -59101 73381 -58835 8 VDD
port 41 nsew
rlabel locali s 73151 -59101 73185 -58835 8 VDD
port 41 nsew
rlabel locali s 72955 -59101 72989 -58835 8 VDD
port 41 nsew
rlabel locali s 72759 -59101 72793 -58835 8 VDD
port 41 nsew
rlabel locali s 69844 -59467 69966 -58471 8 VDD
port 41 nsew
rlabel locali s 67238 -59472 69349 -59438 8 VDD
port 41 nsew
rlabel locali s 68236 -59438 68854 -59421 8 VDD
port 41 nsew
rlabel locali s 68236 -59421 68679 -59392 8 VDD
port 41 nsew
rlabel locali s 68237 -59392 68679 -59378 8 VDD
port 41 nsew
rlabel locali s 68237 -59378 69526 -59329 8 VDD
port 41 nsew
rlabel locali s 68639 -59329 69526 -59279 8 VDD
port 41 nsew
rlabel locali s 69444 -59279 69478 -59113 8 VDD
port 41 nsew
rlabel locali s 69248 -59279 69282 -59113 8 VDD
port 41 nsew
rlabel locali s 69052 -59279 69086 -59113 8 VDD
port 41 nsew
rlabel locali s 68856 -59279 68890 -59113 8 VDD
port 41 nsew
rlabel locali s 68639 -59279 68673 -58912 8 VDD
port 41 nsew
rlabel locali s 68443 -59329 68477 -58912 8 VDD
port 41 nsew
rlabel locali s 68247 -59329 68281 -58912 8 VDD
port 41 nsew
rlabel locali s 67408 -59438 67580 -59248 8 VDD
port 41 nsew
rlabel locali s 67226 -59248 67944 -59149 8 VDD
port 41 nsew
rlabel locali s 67862 -59149 67896 -58883 8 VDD
port 41 nsew
rlabel locali s 67666 -59149 67700 -58883 8 VDD
port 41 nsew
rlabel locali s 67470 -59149 67504 -58883 8 VDD
port 41 nsew
rlabel locali s 67274 -59149 67308 -58883 8 VDD
port 41 nsew
rlabel locali s 69334 -58471 69966 -58349 8 VDD
port 41 nsew
rlabel locali s 75254 -58125 75656 -58059 8 VDD
port 41 nsew
rlabel locali s 77525 -56388 77559 -56096 8 VDD
port 41 nsew
rlabel locali s 77329 -56388 77363 -56098 8 VDD
port 41 nsew
rlabel locali s 77101 -56588 77135 -56113 8 VDD
port 41 nsew
rlabel locali s 76971 -56588 77005 -56116 8 VDD
port 41 nsew
rlabel locali s 77520 -56096 77563 -55996 8 VDD
port 41 nsew
rlabel locali s 85174 -55972 85291 -55962 8 VDD
port 41 nsew
rlabel locali s 84611 -55972 84709 -55969 8 VDD
port 41 nsew
rlabel locali s 85174 -55962 85579 -55898 8 VDD
port 41 nsew
rlabel locali s 77520 -55996 84206 -55936 8 VDD
port 41 nsew
rlabel locali s 77323 -56098 77366 -55936 8 VDD
port 41 nsew
rlabel locali s 77092 -56113 77142 -55936 8 VDD
port 41 nsew
rlabel locali s 76966 -56116 77016 -55936 8 VDD
port 41 nsew
rlabel locali s 76376 -56588 76410 -56093 8 VDD
port 41 nsew
rlabel locali s 76180 -56588 76214 -56095 8 VDD
port 41 nsew
rlabel locali s 74807 -56830 74841 -56238 8 VDD
port 41 nsew
rlabel locali s 75247 -56133 75345 -56127 8 VDD
port 41 nsew
rlabel locali s 76374 -56093 76412 -55936 8 VDD
port 41 nsew
rlabel locali s 76177 -56095 76215 -56000 8 VDD
port 41 nsew
rlabel locali s 75247 -56127 75927 -56010 8 VDD
port 41 nsew
rlabel locali s 75019 -56121 75081 -56107 8 VDD
port 41 nsew
rlabel locali s 74800 -56238 74845 -56114 8 VDD
port 41 nsew
rlabel locali s 74384 -56830 74418 -56237 8 VDD
port 41 nsew
rlabel locali s 74188 -56830 74222 -56240 8 VDD
port 41 nsew
rlabel locali s 73938 -56418 73972 -56252 8 VDD
port 41 nsew
rlabel locali s 73742 -56418 73776 -56252 8 VDD
port 41 nsew
rlabel locali s 73546 -56418 73580 -56252 8 VDD
port 41 nsew
rlabel locali s 73350 -56418 73384 -56252 8 VDD
port 41 nsew
rlabel locali s 73133 -56619 73167 -56252 8 VDD
port 41 nsew
rlabel locali s 74378 -56237 74423 -56114 8 VDD
port 41 nsew
rlabel locali s 74183 -56240 74228 -56114 8 VDD
port 41 nsew
rlabel locali s 73133 -56252 74020 -56202 8 VDD
port 41 nsew
rlabel locali s 72937 -56619 72971 -56202 8 VDD
port 41 nsew
rlabel locali s 72741 -56619 72775 -56202 8 VDD
port 41 nsew
rlabel locali s 72731 -56202 74020 -56153 8 VDD
port 41 nsew
rlabel locali s 72731 -56153 73173 -56138 8 VDD
port 41 nsew
rlabel locali s 74177 -56114 74946 -56107 8 VDD
port 41 nsew
rlabel locali s 74177 -56107 75081 -56090 8 VDD
port 41 nsew
rlabel locali s 73170 -56104 73359 -56097 8 VDD
port 41 nsew
rlabel locali s 73133 -56097 73359 -56090 8 VDD
port 41 nsew
rlabel locali s 72731 -56090 75081 -56055 8 VDD
port 41 nsew
rlabel locali s 75019 -56055 75081 -56027 8 VDD
port 41 nsew
rlabel locali s 72731 -56055 74946 -56048 8 VDD
port 41 nsew
rlabel locali s 75810 -56010 75927 -56000 8 VDD
port 41 nsew
rlabel locali s 75247 -56010 75345 -56007 8 VDD
port 41 nsew
rlabel locali s 75810 -56000 76215 -55936 8 VDD
port 41 nsew
rlabel locali s 72731 -56048 74842 -55987 8 VDD
port 41 nsew
rlabel locali s 69334 -58349 69456 -55987 8 VDD
port 41 nsew
rlabel locali s 66437 -59472 66503 -58142 8 VDD
port 41 nsew
rlabel locali s 66084 -59556 66168 -59443 8 VDD
port 41 nsew
rlabel locali s 63570 -59560 65785 -59518 8 VDD
port 41 nsew
rlabel locali s 66101 -59443 66167 -58142 8 VDD
port 41 nsew
rlabel locali s 63570 -59518 65681 -59407 8 VDD
port 41 nsew
rlabel locali s 61000 -59672 61212 -59533 8 VDD
port 41 nsew
rlabel locali s 60750 -59687 60829 -59662 8 VDD
port 41 nsew
rlabel locali s 60553 -59805 60598 -59681 8 VDD
port 41 nsew
rlabel locali s 60137 -60397 60171 -59804 8 VDD
port 41 nsew
rlabel locali s 59941 -60397 59975 -59807 8 VDD
port 41 nsew
rlabel locali s 59691 -59985 59725 -59819 8 VDD
port 41 nsew
rlabel locali s 59495 -59985 59529 -59819 8 VDD
port 41 nsew
rlabel locali s 59299 -59985 59333 -59819 8 VDD
port 41 nsew
rlabel locali s 59103 -59985 59137 -59819 8 VDD
port 41 nsew
rlabel locali s 58886 -60186 58920 -59819 8 VDD
port 41 nsew
rlabel locali s 60131 -59804 60176 -59681 8 VDD
port 41 nsew
rlabel locali s 59936 -59807 59981 -59681 8 VDD
port 41 nsew
rlabel locali s 58886 -59819 59773 -59769 8 VDD
port 41 nsew
rlabel locali s 58690 -60186 58724 -59769 8 VDD
port 41 nsew
rlabel locali s 58494 -60186 58528 -59769 8 VDD
port 41 nsew
rlabel locali s 56892 -60366 56926 -59774 8 VDD
port 41 nsew
rlabel locali s 58484 -59769 59773 -59720 8 VDD
port 41 nsew
rlabel locali s 58484 -59720 58926 -59705 8 VDD
port 41 nsew
rlabel locali s 59930 -59681 60699 -59662 8 VDD
port 41 nsew
rlabel locali s 59930 -59662 60829 -59657 8 VDD
port 41 nsew
rlabel locali s 58923 -59671 59112 -59664 8 VDD
port 41 nsew
rlabel locali s 58886 -59664 59112 -59657 8 VDD
port 41 nsew
rlabel locali s 58484 -59657 60829 -59615 8 VDD
port 41 nsew
rlabel locali s 56885 -59774 56930 -59650 8 VDD
port 41 nsew
rlabel locali s 56469 -60366 56503 -59773 8 VDD
port 41 nsew
rlabel locali s 56273 -60366 56307 -59776 8 VDD
port 41 nsew
rlabel locali s 56023 -59954 56057 -59788 8 VDD
port 41 nsew
rlabel locali s 55827 -59954 55861 -59788 8 VDD
port 41 nsew
rlabel locali s 55631 -59954 55665 -59788 8 VDD
port 41 nsew
rlabel locali s 55435 -59954 55469 -59788 8 VDD
port 41 nsew
rlabel locali s 55218 -60155 55252 -59788 8 VDD
port 41 nsew
rlabel locali s 56463 -59773 56508 -59650 8 VDD
port 41 nsew
rlabel locali s 56268 -59776 56313 -59650 8 VDD
port 41 nsew
rlabel locali s 55218 -59788 56105 -59738 8 VDD
port 41 nsew
rlabel locali s 55022 -60155 55056 -59738 8 VDD
port 41 nsew
rlabel locali s 54826 -60155 54860 -59738 8 VDD
port 41 nsew
rlabel locali s 51362 -60431 51396 -59839 8 VDD
port 41 nsew
rlabel locali s 54816 -59738 56105 -59689 8 VDD
port 41 nsew
rlabel locali s 51802 -59734 51941 -59706 8 VDD
port 41 nsew
rlabel locali s 54816 -59689 55258 -59674 8 VDD
port 41 nsew
rlabel locali s 56262 -59650 57031 -59626 8 VDD
port 41 nsew
rlabel locali s 55255 -59640 55444 -59633 8 VDD
port 41 nsew
rlabel locali s 55218 -59633 55444 -59626 8 VDD
port 41 nsew
rlabel locali s 60650 -59615 60829 -59579 8 VDD
port 41 nsew
rlabel locali s 58484 -59615 60595 -59604 8 VDD
port 41 nsew
rlabel locali s 60750 -59579 60829 -59548 8 VDD
port 41 nsew
rlabel locali s 57683 -59604 60595 -59538 8 VDD
port 41 nsew
rlabel locali s 64568 -59407 65186 -59390 8 VDD
port 41 nsew
rlabel locali s 64568 -59390 65011 -59361 8 VDD
port 41 nsew
rlabel locali s 64569 -59361 65011 -59347 8 VDD
port 41 nsew
rlabel locali s 64569 -59347 65858 -59298 8 VDD
port 41 nsew
rlabel locali s 64971 -59298 65858 -59248 8 VDD
port 41 nsew
rlabel locali s 65776 -59248 65810 -59082 8 VDD
port 41 nsew
rlabel locali s 65580 -59248 65614 -59082 8 VDD
port 41 nsew
rlabel locali s 65384 -59248 65418 -59082 8 VDD
port 41 nsew
rlabel locali s 65188 -59248 65222 -59082 8 VDD
port 41 nsew
rlabel locali s 64971 -59248 65005 -58881 8 VDD
port 41 nsew
rlabel locali s 64775 -59298 64809 -58881 8 VDD
port 41 nsew
rlabel locali s 64579 -59298 64613 -58881 8 VDD
port 41 nsew
rlabel locali s 63740 -59407 63912 -59217 8 VDD
port 41 nsew
rlabel locali s 63558 -59217 64276 -59118 8 VDD
port 41 nsew
rlabel locali s 64194 -59118 64228 -58852 8 VDD
port 41 nsew
rlabel locali s 63998 -59118 64032 -58852 8 VDD
port 41 nsew
rlabel locali s 63802 -59118 63836 -58852 8 VDD
port 41 nsew
rlabel locali s 63606 -59118 63640 -58852 8 VDD
port 41 nsew
rlabel locali s 61090 -59533 61212 -58537 8 VDD
port 41 nsew
rlabel locali s 58484 -59538 60595 -59504 8 VDD
port 41 nsew
rlabel locali s 59482 -59504 60100 -59487 8 VDD
port 41 nsew
rlabel locali s 59482 -59487 59925 -59458 8 VDD
port 41 nsew
rlabel locali s 59483 -59458 59925 -59444 8 VDD
port 41 nsew
rlabel locali s 59483 -59444 60772 -59395 8 VDD
port 41 nsew
rlabel locali s 59885 -59395 60772 -59345 8 VDD
port 41 nsew
rlabel locali s 60690 -59345 60724 -59179 8 VDD
port 41 nsew
rlabel locali s 60494 -59345 60528 -59179 8 VDD
port 41 nsew
rlabel locali s 60298 -59345 60332 -59179 8 VDD
port 41 nsew
rlabel locali s 60102 -59345 60136 -59179 8 VDD
port 41 nsew
rlabel locali s 59885 -59345 59919 -58978 8 VDD
port 41 nsew
rlabel locali s 59689 -59395 59723 -58978 8 VDD
port 41 nsew
rlabel locali s 59493 -59395 59527 -58978 8 VDD
port 41 nsew
rlabel locali s 58654 -59504 58826 -59314 8 VDD
port 41 nsew
rlabel locali s 58472 -59314 59190 -59215 8 VDD
port 41 nsew
rlabel locali s 59108 -59215 59142 -58949 8 VDD
port 41 nsew
rlabel locali s 58912 -59215 58946 -58949 8 VDD
port 41 nsew
rlabel locali s 58716 -59215 58750 -58949 8 VDD
port 41 nsew
rlabel locali s 58520 -59215 58554 -58949 8 VDD
port 41 nsew
rlabel locali s 60580 -58537 61212 -58415 8 VDD
port 41 nsew
rlabel locali s 66101 -58142 66503 -58076 8 VDD
port 41 nsew
rlabel locali s 68372 -56405 68406 -56113 8 VDD
port 41 nsew
rlabel locali s 68176 -56405 68210 -56115 8 VDD
port 41 nsew
rlabel locali s 67948 -56605 67982 -56130 8 VDD
port 41 nsew
rlabel locali s 67818 -56605 67852 -56133 8 VDD
port 41 nsew
rlabel locali s 68367 -56113 68410 -55987 8 VDD
port 41 nsew
rlabel locali s 68362 -55987 74842 -55953 8 VDD
port 41 nsew
rlabel locali s 68170 -56115 68213 -55953 8 VDD
port 41 nsew
rlabel locali s 67939 -56130 67989 -55953 8 VDD
port 41 nsew
rlabel locali s 67813 -56133 67863 -55953 8 VDD
port 41 nsew
rlabel locali s 67223 -56605 67257 -56110 8 VDD
port 41 nsew
rlabel locali s 67027 -56605 67061 -56112 8 VDD
port 41 nsew
rlabel locali s 65654 -56847 65688 -56255 8 VDD
port 41 nsew
rlabel locali s 66094 -56150 66192 -56144 8 VDD
port 41 nsew
rlabel locali s 67221 -56110 67259 -55953 8 VDD
port 41 nsew
rlabel locali s 67024 -56112 67062 -56017 8 VDD
port 41 nsew
rlabel locali s 66094 -56144 66774 -56027 8 VDD
port 41 nsew
rlabel locali s 65866 -56138 65928 -56124 8 VDD
port 41 nsew
rlabel locali s 65647 -56255 65692 -56131 8 VDD
port 41 nsew
rlabel locali s 65231 -56847 65265 -56254 8 VDD
port 41 nsew
rlabel locali s 65035 -56847 65069 -56257 8 VDD
port 41 nsew
rlabel locali s 64785 -56435 64819 -56269 8 VDD
port 41 nsew
rlabel locali s 64589 -56435 64623 -56269 8 VDD
port 41 nsew
rlabel locali s 64393 -56435 64427 -56269 8 VDD
port 41 nsew
rlabel locali s 64197 -56435 64231 -56269 8 VDD
port 41 nsew
rlabel locali s 63980 -56636 64014 -56269 8 VDD
port 41 nsew
rlabel locali s 65225 -56254 65270 -56131 8 VDD
port 41 nsew
rlabel locali s 65030 -56257 65075 -56131 8 VDD
port 41 nsew
rlabel locali s 63980 -56269 64867 -56219 8 VDD
port 41 nsew
rlabel locali s 63784 -56636 63818 -56219 8 VDD
port 41 nsew
rlabel locali s 63588 -56636 63622 -56219 8 VDD
port 41 nsew
rlabel locali s 63578 -56219 64867 -56170 8 VDD
port 41 nsew
rlabel locali s 63578 -56170 64020 -56155 8 VDD
port 41 nsew
rlabel locali s 65024 -56131 65793 -56124 8 VDD
port 41 nsew
rlabel locali s 65024 -56124 65928 -56107 8 VDD
port 41 nsew
rlabel locali s 64017 -56121 64206 -56114 8 VDD
port 41 nsew
rlabel locali s 63980 -56114 64206 -56107 8 VDD
port 41 nsew
rlabel locali s 63578 -56107 65928 -56081 8 VDD
port 41 nsew
rlabel locali s 60580 -58415 60702 -56081 8 VDD
port 41 nsew
rlabel locali s 57683 -59538 57749 -58208 8 VDD
port 41 nsew
rlabel locali s 57330 -59622 57414 -59509 8 VDD
port 41 nsew
rlabel locali s 54816 -59626 57031 -59584 8 VDD
port 41 nsew
rlabel locali s 57347 -59509 57413 -58208 8 VDD
port 41 nsew
rlabel locali s 54816 -59584 56927 -59473 8 VDD
port 41 nsew
rlabel locali s 51802 -59706 52014 -59567 8 VDD
port 41 nsew
rlabel locali s 51552 -59721 51631 -59696 8 VDD
port 41 nsew
rlabel locali s 51355 -59839 51400 -59715 8 VDD
port 41 nsew
rlabel locali s 50939 -60431 50973 -59838 8 VDD
port 41 nsew
rlabel locali s 50743 -60431 50777 -59841 8 VDD
port 41 nsew
rlabel locali s 50493 -60019 50527 -59853 8 VDD
port 41 nsew
rlabel locali s 50297 -60019 50331 -59853 8 VDD
port 41 nsew
rlabel locali s 50101 -60019 50135 -59853 8 VDD
port 41 nsew
rlabel locali s 49905 -60019 49939 -59853 8 VDD
port 41 nsew
rlabel locali s 49688 -60220 49722 -59853 8 VDD
port 41 nsew
rlabel locali s 50933 -59838 50978 -59715 8 VDD
port 41 nsew
rlabel locali s 50738 -59841 50783 -59715 8 VDD
port 41 nsew
rlabel locali s 49688 -59853 50575 -59803 8 VDD
port 41 nsew
rlabel locali s 49492 -60220 49526 -59803 8 VDD
port 41 nsew
rlabel locali s 49296 -60220 49330 -59803 8 VDD
port 41 nsew
rlabel locali s 47694 -60400 47728 -59808 8 VDD
port 41 nsew
rlabel locali s 49286 -59803 50575 -59754 8 VDD
port 41 nsew
rlabel locali s 49286 -59754 49728 -59739 8 VDD
port 41 nsew
rlabel locali s 50732 -59715 51501 -59696 8 VDD
port 41 nsew
rlabel locali s 50732 -59696 51631 -59691 8 VDD
port 41 nsew
rlabel locali s 49725 -59705 49914 -59698 8 VDD
port 41 nsew
rlabel locali s 49688 -59698 49914 -59691 8 VDD
port 41 nsew
rlabel locali s 49286 -59691 51631 -59649 8 VDD
port 41 nsew
rlabel locali s 47687 -59808 47732 -59684 8 VDD
port 41 nsew
rlabel locali s 47271 -60400 47305 -59807 8 VDD
port 41 nsew
rlabel locali s 47075 -60400 47109 -59810 8 VDD
port 41 nsew
rlabel locali s 46825 -59988 46859 -59822 8 VDD
port 41 nsew
rlabel locali s 46629 -59988 46663 -59822 8 VDD
port 41 nsew
rlabel locali s 46433 -59988 46467 -59822 8 VDD
port 41 nsew
rlabel locali s 46237 -59988 46271 -59822 8 VDD
port 41 nsew
rlabel locali s 46020 -60189 46054 -59822 8 VDD
port 41 nsew
rlabel locali s 47265 -59807 47310 -59684 8 VDD
port 41 nsew
rlabel locali s 47070 -59810 47115 -59684 8 VDD
port 41 nsew
rlabel locali s 46020 -59822 46907 -59772 8 VDD
port 41 nsew
rlabel locali s 45824 -60189 45858 -59772 8 VDD
port 41 nsew
rlabel locali s 45628 -60189 45662 -59772 8 VDD
port 41 nsew
rlabel locali s 42499 -60392 42533 -59800 8 VDD
port 41 nsew
rlabel locali s 45618 -59772 46907 -59723 8 VDD
port 41 nsew
rlabel locali s 45618 -59723 46060 -59708 8 VDD
port 41 nsew
rlabel locali s 47064 -59684 47833 -59660 8 VDD
port 41 nsew
rlabel locali s 46057 -59674 46246 -59667 8 VDD
port 41 nsew
rlabel locali s 42939 -59695 43078 -59667 8 VDD
port 41 nsew
rlabel locali s 46020 -59667 46246 -59660 8 VDD
port 41 nsew
rlabel locali s 51452 -59649 51631 -59613 8 VDD
port 41 nsew
rlabel locali s 49286 -59649 51397 -59638 8 VDD
port 41 nsew
rlabel locali s 51552 -59613 51631 -59582 8 VDD
port 41 nsew
rlabel locali s 48485 -59638 51397 -59572 8 VDD
port 41 nsew
rlabel locali s 55814 -59473 56432 -59456 8 VDD
port 41 nsew
rlabel locali s 55814 -59456 56257 -59427 8 VDD
port 41 nsew
rlabel locali s 55815 -59427 56257 -59413 8 VDD
port 41 nsew
rlabel locali s 55815 -59413 57104 -59364 8 VDD
port 41 nsew
rlabel locali s 56217 -59364 57104 -59314 8 VDD
port 41 nsew
rlabel locali s 57022 -59314 57056 -59148 8 VDD
port 41 nsew
rlabel locali s 56826 -59314 56860 -59148 8 VDD
port 41 nsew
rlabel locali s 56630 -59314 56664 -59148 8 VDD
port 41 nsew
rlabel locali s 56434 -59314 56468 -59148 8 VDD
port 41 nsew
rlabel locali s 56217 -59314 56251 -58947 8 VDD
port 41 nsew
rlabel locali s 56021 -59364 56055 -58947 8 VDD
port 41 nsew
rlabel locali s 55825 -59364 55859 -58947 8 VDD
port 41 nsew
rlabel locali s 54986 -59473 55158 -59283 8 VDD
port 41 nsew
rlabel locali s 54804 -59283 55522 -59184 8 VDD
port 41 nsew
rlabel locali s 55440 -59184 55474 -58918 8 VDD
port 41 nsew
rlabel locali s 55244 -59184 55278 -58918 8 VDD
port 41 nsew
rlabel locali s 55048 -59184 55082 -58918 8 VDD
port 41 nsew
rlabel locali s 54852 -59184 54886 -58918 8 VDD
port 41 nsew
rlabel locali s 51892 -59567 52014 -58571 8 VDD
port 41 nsew
rlabel locali s 49286 -59572 51397 -59538 8 VDD
port 41 nsew
rlabel locali s 50284 -59538 50902 -59521 8 VDD
port 41 nsew
rlabel locali s 50284 -59521 50727 -59492 8 VDD
port 41 nsew
rlabel locali s 50285 -59492 50727 -59478 8 VDD
port 41 nsew
rlabel locali s 50285 -59478 51574 -59429 8 VDD
port 41 nsew
rlabel locali s 50687 -59429 51574 -59379 8 VDD
port 41 nsew
rlabel locali s 51492 -59379 51526 -59213 8 VDD
port 41 nsew
rlabel locali s 51296 -59379 51330 -59213 8 VDD
port 41 nsew
rlabel locali s 51100 -59379 51134 -59213 8 VDD
port 41 nsew
rlabel locali s 50904 -59379 50938 -59213 8 VDD
port 41 nsew
rlabel locali s 50687 -59379 50721 -59012 8 VDD
port 41 nsew
rlabel locali s 50491 -59429 50525 -59012 8 VDD
port 41 nsew
rlabel locali s 50295 -59429 50329 -59012 8 VDD
port 41 nsew
rlabel locali s 49456 -59538 49628 -59348 8 VDD
port 41 nsew
rlabel locali s 49274 -59348 49992 -59249 8 VDD
port 41 nsew
rlabel locali s 49910 -59249 49944 -58983 8 VDD
port 41 nsew
rlabel locali s 49714 -59249 49748 -58983 8 VDD
port 41 nsew
rlabel locali s 49518 -59249 49552 -58983 8 VDD
port 41 nsew
rlabel locali s 49322 -59249 49356 -58983 8 VDD
port 41 nsew
rlabel locali s 51382 -58571 52014 -58449 8 VDD
port 41 nsew
rlabel locali s 57347 -58208 57749 -58142 8 VDD
port 41 nsew
rlabel locali s 59618 -56471 59652 -56179 8 VDD
port 41 nsew
rlabel locali s 59422 -56471 59456 -56181 8 VDD
port 41 nsew
rlabel locali s 59194 -56671 59228 -56196 8 VDD
port 41 nsew
rlabel locali s 59064 -56671 59098 -56199 8 VDD
port 41 nsew
rlabel locali s 59613 -56179 59656 -56081 8 VDD
port 41 nsew
rlabel locali s 59613 -56081 65928 -56072 8 VDD
port 41 nsew
rlabel locali s 65866 -56072 65928 -56044 8 VDD
port 41 nsew
rlabel locali s 59613 -56072 65793 -56065 8 VDD
port 41 nsew
rlabel locali s 66657 -56027 66774 -56017 8 VDD
port 41 nsew
rlabel locali s 66094 -56027 66192 -56024 8 VDD
port 41 nsew
rlabel locali s 66657 -56017 67062 -55953 8 VDD
port 41 nsew
rlabel locali s 59613 -56065 65689 -56019 8 VDD
port 41 nsew
rlabel locali s 59416 -56181 59459 -56019 8 VDD
port 41 nsew
rlabel locali s 59185 -56196 59235 -56019 8 VDD
port 41 nsew
rlabel locali s 59059 -56199 59109 -56019 8 VDD
port 41 nsew
rlabel locali s 58469 -56671 58503 -56176 8 VDD
port 41 nsew
rlabel locali s 58273 -56671 58307 -56178 8 VDD
port 41 nsew
rlabel locali s 56900 -56913 56934 -56321 8 VDD
port 41 nsew
rlabel locali s 57340 -56216 57438 -56210 8 VDD
port 41 nsew
rlabel locali s 58467 -56176 58505 -56019 8 VDD
port 41 nsew
rlabel locali s 58270 -56178 58308 -56083 8 VDD
port 41 nsew
rlabel locali s 57340 -56210 58020 -56093 8 VDD
port 41 nsew
rlabel locali s 57112 -56204 57174 -56190 8 VDD
port 41 nsew
rlabel locali s 56893 -56321 56938 -56197 8 VDD
port 41 nsew
rlabel locali s 56477 -56913 56511 -56320 8 VDD
port 41 nsew
rlabel locali s 56281 -56913 56315 -56323 8 VDD
port 41 nsew
rlabel locali s 56031 -56501 56065 -56335 8 VDD
port 41 nsew
rlabel locali s 55835 -56501 55869 -56335 8 VDD
port 41 nsew
rlabel locali s 55639 -56501 55673 -56335 8 VDD
port 41 nsew
rlabel locali s 55443 -56501 55477 -56335 8 VDD
port 41 nsew
rlabel locali s 55226 -56702 55260 -56335 8 VDD
port 41 nsew
rlabel locali s 56471 -56320 56516 -56197 8 VDD
port 41 nsew
rlabel locali s 56276 -56323 56321 -56197 8 VDD
port 41 nsew
rlabel locali s 55226 -56335 56113 -56285 8 VDD
port 41 nsew
rlabel locali s 55030 -56702 55064 -56285 8 VDD
port 41 nsew
rlabel locali s 54834 -56702 54868 -56285 8 VDD
port 41 nsew
rlabel locali s 54824 -56285 56113 -56236 8 VDD
port 41 nsew
rlabel locali s 54824 -56236 55266 -56221 8 VDD
port 41 nsew
rlabel locali s 56270 -56197 57039 -56190 8 VDD
port 41 nsew
rlabel locali s 56270 -56190 57174 -56173 8 VDD
port 41 nsew
rlabel locali s 55263 -56187 55452 -56180 8 VDD
port 41 nsew
rlabel locali s 55226 -56180 55452 -56173 8 VDD
port 41 nsew
rlabel locali s 54824 -56173 57174 -56138 8 VDD
port 41 nsew
rlabel locali s 57112 -56138 57174 -56110 8 VDD
port 41 nsew
rlabel locali s 54824 -56138 57039 -56131 8 VDD
port 41 nsew
rlabel locali s 54824 -56131 56935 -56113 8 VDD
port 41 nsew
rlabel locali s 51382 -58449 51504 -56113 8 VDD
port 41 nsew
rlabel locali s 48485 -59572 48551 -58242 8 VDD
port 41 nsew
rlabel locali s 48132 -59656 48216 -59543 8 VDD
port 41 nsew
rlabel locali s 45618 -59660 47833 -59618 8 VDD
port 41 nsew
rlabel locali s 48149 -59543 48215 -58242 8 VDD
port 41 nsew
rlabel locali s 45618 -59618 47729 -59507 8 VDD
port 41 nsew
rlabel locali s 42939 -59667 43151 -59528 8 VDD
port 41 nsew
rlabel locali s 42689 -59682 42768 -59657 8 VDD
port 41 nsew
rlabel locali s 42492 -59800 42537 -59676 8 VDD
port 41 nsew
rlabel locali s 42076 -60392 42110 -59799 8 VDD
port 41 nsew
rlabel locali s 41880 -60392 41914 -59802 8 VDD
port 41 nsew
rlabel locali s 41630 -59980 41664 -59814 8 VDD
port 41 nsew
rlabel locali s 41434 -59980 41468 -59814 8 VDD
port 41 nsew
rlabel locali s 41238 -59980 41272 -59814 8 VDD
port 41 nsew
rlabel locali s 41042 -59980 41076 -59814 8 VDD
port 41 nsew
rlabel locali s 40825 -60181 40859 -59814 8 VDD
port 41 nsew
rlabel locali s 42070 -59799 42115 -59676 8 VDD
port 41 nsew
rlabel locali s 41875 -59802 41920 -59676 8 VDD
port 41 nsew
rlabel locali s 40825 -59814 41712 -59764 8 VDD
port 41 nsew
rlabel locali s 40629 -60181 40663 -59764 8 VDD
port 41 nsew
rlabel locali s 40433 -60181 40467 -59764 8 VDD
port 41 nsew
rlabel locali s 38831 -60361 38865 -59769 8 VDD
port 41 nsew
rlabel locali s 40423 -59764 41712 -59715 8 VDD
port 41 nsew
rlabel locali s 40423 -59715 40865 -59700 8 VDD
port 41 nsew
rlabel locali s 41869 -59676 42638 -59657 8 VDD
port 41 nsew
rlabel locali s 41869 -59657 42768 -59652 8 VDD
port 41 nsew
rlabel locali s 40862 -59666 41051 -59659 8 VDD
port 41 nsew
rlabel locali s 40825 -59659 41051 -59652 8 VDD
port 41 nsew
rlabel locali s 40423 -59652 42768 -59610 8 VDD
port 41 nsew
rlabel locali s 38824 -59769 38869 -59645 8 VDD
port 41 nsew
rlabel locali s 38408 -60361 38442 -59768 8 VDD
port 41 nsew
rlabel locali s 38212 -60361 38246 -59771 8 VDD
port 41 nsew
rlabel locali s 37962 -59949 37996 -59783 8 VDD
port 41 nsew
rlabel locali s 37766 -59949 37800 -59783 8 VDD
port 41 nsew
rlabel locali s 37570 -59949 37604 -59783 8 VDD
port 41 nsew
rlabel locali s 37374 -59949 37408 -59783 8 VDD
port 41 nsew
rlabel locali s 37157 -60150 37191 -59783 8 VDD
port 41 nsew
rlabel locali s 38402 -59768 38447 -59645 8 VDD
port 41 nsew
rlabel locali s 38207 -59771 38252 -59645 8 VDD
port 41 nsew
rlabel locali s 37157 -59783 38044 -59733 8 VDD
port 41 nsew
rlabel locali s 36961 -60150 36995 -59733 8 VDD
port 41 nsew
rlabel locali s 36765 -60150 36799 -59733 8 VDD
port 41 nsew
rlabel locali s 34059 -60381 34093 -59789 8 VDD
port 41 nsew
rlabel locali s 36755 -59733 38044 -59684 8 VDD
port 41 nsew
rlabel locali s 36755 -59684 37197 -59669 8 VDD
port 41 nsew
rlabel locali s 34499 -59684 34638 -59656 8 VDD
port 41 nsew
rlabel locali s 38201 -59645 38970 -59621 8 VDD
port 41 nsew
rlabel locali s 37194 -59635 37383 -59628 8 VDD
port 41 nsew
rlabel locali s 37157 -59628 37383 -59621 8 VDD
port 41 nsew
rlabel locali s 42589 -59610 42768 -59574 8 VDD
port 41 nsew
rlabel locali s 40423 -59610 42534 -59599 8 VDD
port 41 nsew
rlabel locali s 42689 -59574 42768 -59543 8 VDD
port 41 nsew
rlabel locali s 39622 -59599 42534 -59533 8 VDD
port 41 nsew
rlabel locali s 46616 -59507 47234 -59490 8 VDD
port 41 nsew
rlabel locali s 46616 -59490 47059 -59461 8 VDD
port 41 nsew
rlabel locali s 46617 -59461 47059 -59447 8 VDD
port 41 nsew
rlabel locali s 46617 -59447 47906 -59398 8 VDD
port 41 nsew
rlabel locali s 47019 -59398 47906 -59348 8 VDD
port 41 nsew
rlabel locali s 47824 -59348 47858 -59182 8 VDD
port 41 nsew
rlabel locali s 47628 -59348 47662 -59182 8 VDD
port 41 nsew
rlabel locali s 47432 -59348 47466 -59182 8 VDD
port 41 nsew
rlabel locali s 47236 -59348 47270 -59182 8 VDD
port 41 nsew
rlabel locali s 47019 -59348 47053 -58981 8 VDD
port 41 nsew
rlabel locali s 46823 -59398 46857 -58981 8 VDD
port 41 nsew
rlabel locali s 46627 -59398 46661 -58981 8 VDD
port 41 nsew
rlabel locali s 45788 -59507 45960 -59317 8 VDD
port 41 nsew
rlabel locali s 45606 -59317 46324 -59218 8 VDD
port 41 nsew
rlabel locali s 46242 -59218 46276 -58952 8 VDD
port 41 nsew
rlabel locali s 46046 -59218 46080 -58952 8 VDD
port 41 nsew
rlabel locali s 45850 -59218 45884 -58952 8 VDD
port 41 nsew
rlabel locali s 45654 -59218 45688 -58952 8 VDD
port 41 nsew
rlabel locali s 43029 -59528 43151 -58532 8 VDD
port 41 nsew
rlabel locali s 40423 -59533 42534 -59499 8 VDD
port 41 nsew
rlabel locali s 41421 -59499 42039 -59482 8 VDD
port 41 nsew
rlabel locali s 41421 -59482 41864 -59453 8 VDD
port 41 nsew
rlabel locali s 41422 -59453 41864 -59439 8 VDD
port 41 nsew
rlabel locali s 41422 -59439 42711 -59390 8 VDD
port 41 nsew
rlabel locali s 41824 -59390 42711 -59340 8 VDD
port 41 nsew
rlabel locali s 42629 -59340 42663 -59174 8 VDD
port 41 nsew
rlabel locali s 42433 -59340 42467 -59174 8 VDD
port 41 nsew
rlabel locali s 42237 -59340 42271 -59174 8 VDD
port 41 nsew
rlabel locali s 42041 -59340 42075 -59174 8 VDD
port 41 nsew
rlabel locali s 41824 -59340 41858 -58973 8 VDD
port 41 nsew
rlabel locali s 41628 -59390 41662 -58973 8 VDD
port 41 nsew
rlabel locali s 41432 -59390 41466 -58973 8 VDD
port 41 nsew
rlabel locali s 40593 -59499 40765 -59309 8 VDD
port 41 nsew
rlabel locali s 40411 -59309 41129 -59210 8 VDD
port 41 nsew
rlabel locali s 41047 -59210 41081 -58944 8 VDD
port 41 nsew
rlabel locali s 40851 -59210 40885 -58944 8 VDD
port 41 nsew
rlabel locali s 40655 -59210 40689 -58944 8 VDD
port 41 nsew
rlabel locali s 40459 -59210 40493 -58944 8 VDD
port 41 nsew
rlabel locali s 42519 -58532 43151 -58410 8 VDD
port 41 nsew
rlabel locali s 48149 -58242 48551 -58176 8 VDD
port 41 nsew
rlabel locali s 50420 -56505 50454 -56213 8 VDD
port 41 nsew
rlabel locali s 50224 -56505 50258 -56215 8 VDD
port 41 nsew
rlabel locali s 49996 -56705 50030 -56230 8 VDD
port 41 nsew
rlabel locali s 49866 -56705 49900 -56233 8 VDD
port 41 nsew
rlabel locali s 50415 -56213 50458 -56113 8 VDD
port 41 nsew
rlabel locali s 57903 -56093 58020 -56083 8 VDD
port 41 nsew
rlabel locali s 57340 -56093 57438 -56090 8 VDD
port 41 nsew
rlabel locali s 57903 -56083 58308 -56019 8 VDD
port 41 nsew
rlabel locali s 50415 -56113 56935 -56053 8 VDD
port 41 nsew
rlabel locali s 50218 -56215 50261 -56053 8 VDD
port 41 nsew
rlabel locali s 49987 -56230 50037 -56053 8 VDD
port 41 nsew
rlabel locali s 49861 -56233 49911 -56053 8 VDD
port 41 nsew
rlabel locali s 49271 -56705 49305 -56210 8 VDD
port 41 nsew
rlabel locali s 49075 -56705 49109 -56212 8 VDD
port 41 nsew
rlabel locali s 47702 -56947 47736 -56355 8 VDD
port 41 nsew
rlabel locali s 48142 -56250 48240 -56244 8 VDD
port 41 nsew
rlabel locali s 49269 -56210 49307 -56053 8 VDD
port 41 nsew
rlabel locali s 49072 -56212 49110 -56117 8 VDD
port 41 nsew
rlabel locali s 48142 -56244 48822 -56127 8 VDD
port 41 nsew
rlabel locali s 47914 -56238 47976 -56224 8 VDD
port 41 nsew
rlabel locali s 47695 -56355 47740 -56231 8 VDD
port 41 nsew
rlabel locali s 47279 -56947 47313 -56354 8 VDD
port 41 nsew
rlabel locali s 47083 -56947 47117 -56357 8 VDD
port 41 nsew
rlabel locali s 46833 -56535 46867 -56369 8 VDD
port 41 nsew
rlabel locali s 46637 -56535 46671 -56369 8 VDD
port 41 nsew
rlabel locali s 46441 -56535 46475 -56369 8 VDD
port 41 nsew
rlabel locali s 46245 -56535 46279 -56369 8 VDD
port 41 nsew
rlabel locali s 46028 -56736 46062 -56369 8 VDD
port 41 nsew
rlabel locali s 47273 -56354 47318 -56231 8 VDD
port 41 nsew
rlabel locali s 47078 -56357 47123 -56231 8 VDD
port 41 nsew
rlabel locali s 46028 -56369 46915 -56319 8 VDD
port 41 nsew
rlabel locali s 45832 -56736 45866 -56319 8 VDD
port 41 nsew
rlabel locali s 45636 -56736 45670 -56319 8 VDD
port 41 nsew
rlabel locali s 45626 -56319 46915 -56270 8 VDD
port 41 nsew
rlabel locali s 45626 -56270 46068 -56255 8 VDD
port 41 nsew
rlabel locali s 47072 -56231 47841 -56224 8 VDD
port 41 nsew
rlabel locali s 47072 -56224 47976 -56207 8 VDD
port 41 nsew
rlabel locali s 46065 -56221 46254 -56214 8 VDD
port 41 nsew
rlabel locali s 46028 -56214 46254 -56207 8 VDD
port 41 nsew
rlabel locali s 45626 -56207 47976 -56172 8 VDD
port 41 nsew
rlabel locali s 47914 -56172 47976 -56144 8 VDD
port 41 nsew
rlabel locali s 45626 -56172 47841 -56165 8 VDD
port 41 nsew
rlabel locali s 48705 -56127 48822 -56117 8 VDD
port 41 nsew
rlabel locali s 48142 -56127 48240 -56124 8 VDD
port 41 nsew
rlabel locali s 48705 -56117 49110 -56053 8 VDD
port 41 nsew
rlabel locali s 45626 -56165 47737 -56103 8 VDD
port 41 nsew
rlabel locali s 42519 -58410 42641 -56103 8 VDD
port 41 nsew
rlabel locali s 39622 -59533 39688 -58203 8 VDD
port 41 nsew
rlabel locali s 39269 -59617 39353 -59504 8 VDD
port 41 nsew
rlabel locali s 36755 -59621 38970 -59579 8 VDD
port 41 nsew
rlabel locali s 39286 -59504 39352 -58203 8 VDD
port 41 nsew
rlabel locali s 36755 -59579 38866 -59468 8 VDD
port 41 nsew
rlabel locali s 34499 -59656 34711 -59517 8 VDD
port 41 nsew
rlabel locali s 34249 -59671 34328 -59646 8 VDD
port 41 nsew
rlabel locali s 34052 -59789 34097 -59665 8 VDD
port 41 nsew
rlabel locali s 33636 -60381 33670 -59788 8 VDD
port 41 nsew
rlabel locali s 33440 -60381 33474 -59791 8 VDD
port 41 nsew
rlabel locali s 33190 -59969 33224 -59803 8 VDD
port 41 nsew
rlabel locali s 32994 -59969 33028 -59803 8 VDD
port 41 nsew
rlabel locali s 32798 -59969 32832 -59803 8 VDD
port 41 nsew
rlabel locali s 32602 -59969 32636 -59803 8 VDD
port 41 nsew
rlabel locali s 32385 -60170 32419 -59803 8 VDD
port 41 nsew
rlabel locali s 33630 -59788 33675 -59665 8 VDD
port 41 nsew
rlabel locali s 33435 -59791 33480 -59665 8 VDD
port 41 nsew
rlabel locali s 32385 -59803 33272 -59753 8 VDD
port 41 nsew
rlabel locali s 32189 -60170 32223 -59753 8 VDD
port 41 nsew
rlabel locali s 31993 -60170 32027 -59753 8 VDD
port 41 nsew
rlabel locali s 30391 -60350 30425 -59758 8 VDD
port 41 nsew
rlabel locali s 31983 -59753 33272 -59704 8 VDD
port 41 nsew
rlabel locali s 31983 -59704 32425 -59689 8 VDD
port 41 nsew
rlabel locali s 33429 -59665 34198 -59646 8 VDD
port 41 nsew
rlabel locali s 33429 -59646 34328 -59641 8 VDD
port 41 nsew
rlabel locali s 32422 -59655 32611 -59648 8 VDD
port 41 nsew
rlabel locali s 32385 -59648 32611 -59641 8 VDD
port 41 nsew
rlabel locali s 31983 -59641 34328 -59599 8 VDD
port 41 nsew
rlabel locali s 30384 -59758 30429 -59634 8 VDD
port 41 nsew
rlabel locali s 29968 -60350 30002 -59757 8 VDD
port 41 nsew
rlabel locali s 29772 -60350 29806 -59760 8 VDD
port 41 nsew
rlabel locali s 17982 -61967 18071 -60272 8 VDD
port 41 nsew
rlabel locali s 17788 -61967 17822 -61676 8 VDD
port 41 nsew
rlabel locali s 17592 -61967 17626 -61676 8 VDD
port 41 nsew
rlabel locali s 17396 -61967 17430 -61676 8 VDD
port 41 nsew
rlabel locali s 16951 -61967 16985 -61676 8 VDD
port 41 nsew
rlabel locali s 16755 -61967 16789 -61676 8 VDD
port 41 nsew
rlabel locali s 16559 -61967 16593 -61676 8 VDD
port 41 nsew
rlabel locali s 15088 -61967 15122 -61676 8 VDD
port 41 nsew
rlabel locali s 14892 -61967 14926 -61676 8 VDD
port 41 nsew
rlabel locali s 14696 -61967 14730 -61676 8 VDD
port 41 nsew
rlabel locali s 14251 -61967 14285 -61676 8 VDD
port 41 nsew
rlabel locali s 14055 -61967 14089 -61676 8 VDD
port 41 nsew
rlabel locali s 13859 -61967 13893 -61676 8 VDD
port 41 nsew
rlabel locali s 8743 -62029 8777 -61839 8 VDD
port 41 nsew
rlabel locali s 8541 -62151 8587 -62017 8 VDD
port 41 nsew
rlabel locali s 8428 -62151 8474 -62027 8 VDD
port 41 nsew
rlabel locali s 8547 -62017 8581 -61839 8 VDD
port 41 nsew
rlabel locali s 8434 -62027 8468 -61839 8 VDD
port 41 nsew
rlabel locali s 8232 -62151 8278 -62022 8 VDD
port 41 nsew
rlabel locali s 8119 -62151 8165 -62026 8 VDD
port 41 nsew
rlabel locali s 8238 -62022 8272 -61839 8 VDD
port 41 nsew
rlabel locali s 8124 -62026 8158 -61839 8 VDD
port 41 nsew
rlabel locali s 7921 -62151 7967 -62022 8 VDD
port 41 nsew
rlabel locali s 7732 -62151 7772 -62022 8 VDD
port 41 nsew
rlabel locali s 4732 -62220 5784 -62151 8 VDD
port 41 nsew
rlabel locali s 5738 -62151 5784 -62029 8 VDD
port 41 nsew
rlabel locali s 7928 -62022 7962 -61839 8 VDD
port 41 nsew
rlabel locali s 7732 -62022 7766 -61839 8 VDD
port 41 nsew
rlabel locali s 5743 -62029 5777 -61839 8 VDD
port 41 nsew
rlabel locali s 5541 -62151 5587 -62017 8 VDD
port 41 nsew
rlabel locali s 5428 -62151 5474 -62027 8 VDD
port 41 nsew
rlabel locali s 5547 -62017 5581 -61839 8 VDD
port 41 nsew
rlabel locali s 5434 -62027 5468 -61839 8 VDD
port 41 nsew
rlabel locali s 5232 -62151 5278 -62022 8 VDD
port 41 nsew
rlabel locali s 5119 -62151 5165 -62026 8 VDD
port 41 nsew
rlabel locali s 5238 -62022 5272 -61839 8 VDD
port 41 nsew
rlabel locali s 5124 -62026 5158 -61839 8 VDD
port 41 nsew
rlabel locali s 4921 -62151 4967 -62022 8 VDD
port 41 nsew
rlabel locali s 4732 -62151 4772 -62022 8 VDD
port 41 nsew
rlabel locali s 2232 -62220 3284 -62151 8 VDD
port 41 nsew
rlabel locali s 3238 -62151 3284 -62029 8 VDD
port 41 nsew
rlabel locali s 4928 -62022 4962 -61839 8 VDD
port 41 nsew
rlabel locali s 4732 -62022 4766 -61839 8 VDD
port 41 nsew
rlabel locali s 3243 -62029 3277 -61839 8 VDD
port 41 nsew
rlabel locali s 3041 -62151 3087 -62017 8 VDD
port 41 nsew
rlabel locali s 2928 -62151 2974 -62027 8 VDD
port 41 nsew
rlabel locali s 3047 -62017 3081 -61839 8 VDD
port 41 nsew
rlabel locali s 2934 -62027 2968 -61839 8 VDD
port 41 nsew
rlabel locali s 2732 -62151 2778 -62022 8 VDD
port 41 nsew
rlabel locali s 2619 -62151 2665 -62026 8 VDD
port 41 nsew
rlabel locali s 2738 -62022 2772 -61839 8 VDD
port 41 nsew
rlabel locali s 2624 -62026 2658 -61839 8 VDD
port 41 nsew
rlabel locali s 2421 -62151 2467 -62022 8 VDD
port 41 nsew
rlabel locali s 2232 -62151 2272 -62022 8 VDD
port 41 nsew
rlabel locali s 2428 -62022 2462 -61839 8 VDD
port 41 nsew
rlabel locali s 2232 -62022 2266 -61839 8 VDD
port 41 nsew
rlabel locali s 1109 -62258 1224 -61386 8 VDD
port 41 nsew
rlabel locali s 62 -62258 655 -62220 8 VDD
port 41 nsew
rlabel locali s -268 -62220 784 -62151 8 VDD
port 41 nsew
rlabel locali s 738 -62151 784 -62029 8 VDD
port 41 nsew
rlabel locali s 743 -62029 777 -61839 8 VDD
port 41 nsew
rlabel locali s 541 -62151 587 -62017 8 VDD
port 41 nsew
rlabel locali s 428 -62151 474 -62027 8 VDD
port 41 nsew
rlabel locali s 547 -62017 581 -61839 8 VDD
port 41 nsew
rlabel locali s 434 -62027 468 -61839 8 VDD
port 41 nsew
rlabel locali s 232 -62151 278 -62022 8 VDD
port 41 nsew
rlabel locali s 119 -62151 165 -62026 8 VDD
port 41 nsew
rlabel locali s 238 -62022 272 -61839 8 VDD
port 41 nsew
rlabel locali s 124 -62026 158 -61839 8 VDD
port 41 nsew
rlabel locali s -79 -62151 -33 -62022 2 VDD
port 41 nsew
rlabel locali s -268 -62151 -228 -62022 2 VDD
port 41 nsew
rlabel locali s -72 -62022 -38 -61839 2 VDD
port 41 nsew
rlabel locali s -268 -62022 -234 -61839 2 VDD
port 41 nsew
rlabel locali s -1373 -62258 -1259 -61386 2 VDD
port 41 nsew
rlabel locali s -2454 -62258 -1861 -62220 2 VDD
port 41 nsew
rlabel locali s -2768 -62220 -1716 -62151 2 VDD
port 41 nsew
rlabel locali s -1762 -62151 -1716 -62029 2 VDD
port 41 nsew
rlabel locali s -1757 -62029 -1723 -61839 2 VDD
port 41 nsew
rlabel locali s -1959 -62151 -1913 -62017 2 VDD
port 41 nsew
rlabel locali s -2072 -62151 -2026 -62027 2 VDD
port 41 nsew
rlabel locali s -1953 -62017 -1919 -61839 2 VDD
port 41 nsew
rlabel locali s -2066 -62027 -2032 -61839 2 VDD
port 41 nsew
rlabel locali s -2268 -62151 -2222 -62022 2 VDD
port 41 nsew
rlabel locali s -2381 -62151 -2335 -62026 2 VDD
port 41 nsew
rlabel locali s -2262 -62022 -2228 -61839 2 VDD
port 41 nsew
rlabel locali s -2376 -62026 -2342 -61839 2 VDD
port 41 nsew
rlabel locali s -2579 -62151 -2533 -62022 2 VDD
port 41 nsew
rlabel locali s -2768 -62151 -2728 -62022 2 VDD
port 41 nsew
rlabel locali s -2572 -62022 -2538 -61839 2 VDD
port 41 nsew
rlabel locali s -2768 -62022 -2734 -61839 2 VDD
port 41 nsew
rlabel locali s -3941 -62258 -3826 -61421 2 VDD
port 41 nsew
rlabel locali s -5268 -62258 -4216 -62151 2 VDD
port 41 nsew
rlabel locali s -21562 -62284 -18772 -62217 2 VDD
port 41 nsew
rlabel locali s -21374 -62217 -18772 -62201 2 VDD
port 41 nsew
rlabel locali s -4262 -62151 -4216 -62029 2 VDD
port 41 nsew
rlabel locali s -4257 -62029 -4223 -61839 2 VDD
port 41 nsew
rlabel locali s -4459 -62151 -4413 -62017 2 VDD
port 41 nsew
rlabel locali s -4572 -62151 -4526 -62027 2 VDD
port 41 nsew
rlabel locali s -4453 -62017 -4419 -61839 2 VDD
port 41 nsew
rlabel locali s -4566 -62027 -4532 -61839 2 VDD
port 41 nsew
rlabel locali s -4768 -62151 -4722 -62022 2 VDD
port 41 nsew
rlabel locali s -4881 -62151 -4835 -62026 2 VDD
port 41 nsew
rlabel locali s -4762 -62022 -4728 -61839 2 VDD
port 41 nsew
rlabel locali s -4876 -62026 -4842 -61839 2 VDD
port 41 nsew
rlabel locali s -5079 -62151 -5033 -62022 2 VDD
port 41 nsew
rlabel locali s -5268 -62151 -5228 -62022 2 VDD
port 41 nsew
rlabel locali s -5072 -62022 -5038 -61839 2 VDD
port 41 nsew
rlabel locali s -5268 -62022 -5234 -61839 2 VDD
port 41 nsew
rlabel locali s -20226 -62201 -20192 -61925 2 VDD
port 41 nsew
rlabel locali s -20422 -62201 -20388 -61925 2 VDD
port 41 nsew
rlabel locali s -20618 -62201 -20584 -61925 2 VDD
port 41 nsew
rlabel locali s -20814 -62201 -20780 -61925 2 VDD
port 41 nsew
rlabel locali s -21356 -62201 -21322 -61925 2 VDD
port 41 nsew
rlabel locali s -21552 -62217 -21518 -61925 2 VDD
port 41 nsew
rlabel locali s -18948 -61749 -18772 -61662 2 VDD
port 41 nsew
rlabel locali s 1104 -61386 1227 -61250 8 VDD
port 41 nsew
rlabel locali s -1379 -61386 -1256 -61250 2 VDD
port 41 nsew
rlabel locali s -3946 -61421 -3823 -61285 2 VDD
port 41 nsew
rlabel locali s 1103 -60833 1226 -60832 8 VDD
port 41 nsew
rlabel locali s 1103 -60832 1409 -60770 8 VDD
port 41 nsew
rlabel locali s -15506 -60973 -15472 -60807 2 VDD
port 41 nsew
rlabel locali s -15702 -60973 -15668 -60807 2 VDD
port 41 nsew
rlabel locali s -15898 -60973 -15864 -60807 2 VDD
port 41 nsew
rlabel locali s -16094 -60973 -16060 -60807 2 VDD
port 41 nsew
rlabel locali s -16311 -61174 -16277 -60807 2 VDD
port 41 nsew
rlabel locali s 17690 -60566 17724 -60275 8 VDD
port 41 nsew
rlabel locali s 17494 -60566 17528 -60275 8 VDD
port 41 nsew
rlabel locali s 17298 -60566 17332 -60275 8 VDD
port 41 nsew
rlabel locali s 15947 -60566 15981 -60275 8 VDD
port 41 nsew
rlabel locali s 15751 -60566 15785 -60275 8 VDD
port 41 nsew
rlabel locali s 15555 -60566 15589 -60275 8 VDD
port 41 nsew
rlabel locali s 14990 -60566 15024 -60275 8 VDD
port 41 nsew
rlabel locali s 14794 -60566 14828 -60275 8 VDD
port 41 nsew
rlabel locali s 14598 -60566 14632 -60275 8 VDD
port 41 nsew
rlabel locali s 13247 -60566 13281 -60275 8 VDD
port 41 nsew
rlabel locali s 13051 -60566 13085 -60275 8 VDD
port 41 nsew
rlabel locali s 12855 -60566 12889 -60275 8 VDD
port 41 nsew
rlabel locali s 12365 -60566 12399 -60275 8 VDD
port 41 nsew
rlabel locali s 12169 -60566 12203 -60275 8 VDD
port 41 nsew
rlabel locali s 11973 -60566 12007 -60275 8 VDD
port 41 nsew
rlabel locali s 17289 -60275 17784 -60272 8 VDD
port 41 nsew
rlabel locali s 14589 -60275 16042 -60274 8 VDD
port 41 nsew
rlabel locali s 16967 -60272 18071 -60270 8 VDD
port 41 nsew
rlabel locali s 14276 -60274 16042 -60270 8 VDD
port 41 nsew
rlabel locali s 11964 -60275 13342 -60270 8 VDD
port 41 nsew
rlabel locali s 11964 -60270 18071 -60207 8 VDD
port 41 nsew
rlabel locali s 16967 -60207 18071 -60204 8 VDD
port 41 nsew
rlabel locali s 14276 -60207 14749 -60206 8 VDD
port 41 nsew
rlabel locali s 29522 -59938 29556 -59772 8 VDD
port 41 nsew
rlabel locali s 29326 -59938 29360 -59772 8 VDD
port 41 nsew
rlabel locali s 29130 -59938 29164 -59772 8 VDD
port 41 nsew
rlabel locali s 28934 -59938 28968 -59772 8 VDD
port 41 nsew
rlabel locali s 28717 -60139 28751 -59772 8 VDD
port 41 nsew
rlabel locali s 29962 -59757 30007 -59634 8 VDD
port 41 nsew
rlabel locali s 29767 -59760 29812 -59634 8 VDD
port 41 nsew
rlabel locali s 28717 -59772 29604 -59722 8 VDD
port 41 nsew
rlabel locali s 28521 -60139 28555 -59722 8 VDD
port 41 nsew
rlabel locali s 28325 -60139 28359 -59722 8 VDD
port 41 nsew
rlabel locali s 21512 -59756 21575 -59745 8 VDD
port 41 nsew
rlabel locali s 20392 -59749 20478 -59745 8 VDD
port 41 nsew
rlabel locali s 22910 -59740 26199 -59732 8 VDD
port 41 nsew
rlabel locali s 22193 -59745 22267 -59739 8 VDD
port 41 nsew
rlabel locali s 20392 -59745 21575 -59739 8 VDD
port 41 nsew
rlabel locali s 20392 -59739 22267 -59733 8 VDD
port 41 nsew
rlabel locali s 17945 -60204 18071 -59733 8 VDD
port 41 nsew
rlabel locali s 7741 -59996 7864 -59969 8 VDD
port 41 nsew
rlabel locali s 7741 -59969 8794 -59900 8 VDD
port 41 nsew
rlabel locali s 8748 -59900 8794 -59778 8 VDD
port 41 nsew
rlabel locali s 17945 -59733 22267 -59732 8 VDD
port 41 nsew
rlabel locali s 28315 -59722 29604 -59673 8 VDD
port 41 nsew
rlabel locali s 28315 -59673 28757 -59658 8 VDD
port 41 nsew
rlabel locali s 17945 -59732 26199 -59676 8 VDD
port 41 nsew
rlabel locali s 21512 -59676 26199 -59672 8 VDD
port 41 nsew
rlabel locali s 22193 -59672 26199 -59664 8 VDD
port 41 nsew
rlabel locali s 22888 -59664 26199 -59637 8 VDD
port 41 nsew
rlabel locali s 29761 -59634 30530 -59610 8 VDD
port 41 nsew
rlabel locali s 28754 -59624 28943 -59617 8 VDD
port 41 nsew
rlabel locali s 28717 -59617 28943 -59610 8 VDD
port 41 nsew
rlabel locali s 34149 -59599 34328 -59563 8 VDD
port 41 nsew
rlabel locali s 31983 -59599 34094 -59588 8 VDD
port 41 nsew
rlabel locali s 34249 -59563 34328 -59532 8 VDD
port 41 nsew
rlabel locali s 31182 -59588 34094 -59522 8 VDD
port 41 nsew
rlabel locali s 37753 -59468 38371 -59451 8 VDD
port 41 nsew
rlabel locali s 37753 -59451 38196 -59422 8 VDD
port 41 nsew
rlabel locali s 37754 -59422 38196 -59408 8 VDD
port 41 nsew
rlabel locali s 37754 -59408 39043 -59359 8 VDD
port 41 nsew
rlabel locali s 38156 -59359 39043 -59309 8 VDD
port 41 nsew
rlabel locali s 38961 -59309 38995 -59143 8 VDD
port 41 nsew
rlabel locali s 38765 -59309 38799 -59143 8 VDD
port 41 nsew
rlabel locali s 38569 -59309 38603 -59143 8 VDD
port 41 nsew
rlabel locali s 38373 -59309 38407 -59143 8 VDD
port 41 nsew
rlabel locali s 38156 -59309 38190 -58942 8 VDD
port 41 nsew
rlabel locali s 37960 -59359 37994 -58942 8 VDD
port 41 nsew
rlabel locali s 37764 -59359 37798 -58942 8 VDD
port 41 nsew
rlabel locali s 36925 -59468 37097 -59278 8 VDD
port 41 nsew
rlabel locali s 36743 -59278 37461 -59179 8 VDD
port 41 nsew
rlabel locali s 37379 -59179 37413 -58913 8 VDD
port 41 nsew
rlabel locali s 37183 -59179 37217 -58913 8 VDD
port 41 nsew
rlabel locali s 36987 -59179 37021 -58913 8 VDD
port 41 nsew
rlabel locali s 36791 -59179 36825 -58913 8 VDD
port 41 nsew
rlabel locali s 34589 -59517 34711 -58521 8 VDD
port 41 nsew
rlabel locali s 31983 -59522 34094 -59488 8 VDD
port 41 nsew
rlabel locali s 32981 -59488 33599 -59471 8 VDD
port 41 nsew
rlabel locali s 32981 -59471 33424 -59442 8 VDD
port 41 nsew
rlabel locali s 32982 -59442 33424 -59428 8 VDD
port 41 nsew
rlabel locali s 32982 -59428 34271 -59379 8 VDD
port 41 nsew
rlabel locali s 33384 -59379 34271 -59329 8 VDD
port 41 nsew
rlabel locali s 34189 -59329 34223 -59163 8 VDD
port 41 nsew
rlabel locali s 33993 -59329 34027 -59163 8 VDD
port 41 nsew
rlabel locali s 33797 -59329 33831 -59163 8 VDD
port 41 nsew
rlabel locali s 33601 -59329 33635 -59163 8 VDD
port 41 nsew
rlabel locali s 33384 -59329 33418 -58962 8 VDD
port 41 nsew
rlabel locali s 33188 -59379 33222 -58962 8 VDD
port 41 nsew
rlabel locali s 32992 -59379 33026 -58962 8 VDD
port 41 nsew
rlabel locali s 32153 -59488 32325 -59298 8 VDD
port 41 nsew
rlabel locali s 31971 -59298 32689 -59199 8 VDD
port 41 nsew
rlabel locali s 32607 -59199 32641 -58933 8 VDD
port 41 nsew
rlabel locali s 32411 -59199 32445 -58933 8 VDD
port 41 nsew
rlabel locali s 32215 -59199 32249 -58933 8 VDD
port 41 nsew
rlabel locali s 32019 -59199 32053 -58933 8 VDD
port 41 nsew
rlabel locali s 34079 -58521 34711 -58399 8 VDD
port 41 nsew
rlabel locali s 39286 -58203 39688 -58137 8 VDD
port 41 nsew
rlabel locali s 41557 -56466 41591 -56174 8 VDD
port 41 nsew
rlabel locali s 41361 -56466 41395 -56176 8 VDD
port 41 nsew
rlabel locali s 41133 -56666 41167 -56191 8 VDD
port 41 nsew
rlabel locali s 41003 -56666 41037 -56194 8 VDD
port 41 nsew
rlabel locali s 41552 -56174 41595 -56103 8 VDD
port 41 nsew
rlabel locali s 41552 -56103 47737 -56054 8 VDD
port 41 nsew
rlabel locali s 48705 -56053 56935 -56020 8 VDD
port 41 nsew
rlabel locali s 46624 -56054 47242 -56037 8 VDD
port 41 nsew
rlabel locali s 57903 -56019 65689 -55966 8 VDD
port 41 nsew
rlabel locali s 55822 -56020 56440 -56003 8 VDD
port 41 nsew
rlabel locali s 55822 -56003 56265 -55974 8 VDD
port 41 nsew
rlabel locali s 48705 -56020 55166 -56000 8 VDD
port 41 nsew
rlabel locali s 46624 -56037 47067 -56008 8 VDD
port 41 nsew
rlabel locali s 41552 -56054 45968 -56014 8 VDD
port 41 nsew
rlabel locali s 41355 -56176 41398 -56014 8 VDD
port 41 nsew
rlabel locali s 41124 -56191 41174 -56014 8 VDD
port 41 nsew
rlabel locali s 40998 -56194 41048 -56014 8 VDD
port 41 nsew
rlabel locali s 40408 -56666 40442 -56171 8 VDD
port 41 nsew
rlabel locali s 40212 -56666 40246 -56173 8 VDD
port 41 nsew
rlabel locali s 38839 -56908 38873 -56316 8 VDD
port 41 nsew
rlabel locali s 39279 -56211 39377 -56205 8 VDD
port 41 nsew
rlabel locali s 40406 -56171 40444 -56014 8 VDD
port 41 nsew
rlabel locali s 40209 -56173 40247 -56078 8 VDD
port 41 nsew
rlabel locali s 39279 -56205 39959 -56088 8 VDD
port 41 nsew
rlabel locali s 39051 -56199 39113 -56185 8 VDD
port 41 nsew
rlabel locali s 38832 -56316 38877 -56192 8 VDD
port 41 nsew
rlabel locali s 38416 -56908 38450 -56315 8 VDD
port 41 nsew
rlabel locali s 38220 -56908 38254 -56318 8 VDD
port 41 nsew
rlabel locali s 37970 -56496 38004 -56330 8 VDD
port 41 nsew
rlabel locali s 37774 -56496 37808 -56330 8 VDD
port 41 nsew
rlabel locali s 37578 -56496 37612 -56330 8 VDD
port 41 nsew
rlabel locali s 37382 -56496 37416 -56330 8 VDD
port 41 nsew
rlabel locali s 37165 -56697 37199 -56330 8 VDD
port 41 nsew
rlabel locali s 38410 -56315 38455 -56192 8 VDD
port 41 nsew
rlabel locali s 38215 -56318 38260 -56192 8 VDD
port 41 nsew
rlabel locali s 37165 -56330 38052 -56280 8 VDD
port 41 nsew
rlabel locali s 36969 -56697 37003 -56280 8 VDD
port 41 nsew
rlabel locali s 36773 -56697 36807 -56280 8 VDD
port 41 nsew
rlabel locali s 36763 -56280 38052 -56231 8 VDD
port 41 nsew
rlabel locali s 36763 -56231 37205 -56216 8 VDD
port 41 nsew
rlabel locali s 38209 -56192 38978 -56185 8 VDD
port 41 nsew
rlabel locali s 38209 -56185 39113 -56168 8 VDD
port 41 nsew
rlabel locali s 37202 -56182 37391 -56175 8 VDD
port 41 nsew
rlabel locali s 37165 -56175 37391 -56168 8 VDD
port 41 nsew
rlabel locali s 34079 -58399 34201 -56168 8 VDD
port 41 nsew
rlabel locali s 31182 -59522 31248 -58192 8 VDD
port 41 nsew
rlabel locali s 30829 -59606 30913 -59493 8 VDD
port 41 nsew
rlabel locali s 28315 -59610 30530 -59568 8 VDD
port 41 nsew
rlabel locali s 30846 -59493 30912 -58192 8 VDD
port 41 nsew
rlabel locali s 28315 -59568 30426 -59457 8 VDD
port 41 nsew
rlabel locali s 29313 -59457 29931 -59440 8 VDD
port 41 nsew
rlabel locali s 29313 -59440 29756 -59411 8 VDD
port 41 nsew
rlabel locali s 29314 -59411 29756 -59397 8 VDD
port 41 nsew
rlabel locali s 29314 -59397 30603 -59348 8 VDD
port 41 nsew
rlabel locali s 29716 -59348 30603 -59298 8 VDD
port 41 nsew
rlabel locali s 30521 -59298 30555 -59132 8 VDD
port 41 nsew
rlabel locali s 30325 -59298 30359 -59132 8 VDD
port 41 nsew
rlabel locali s 30129 -59298 30163 -59132 8 VDD
port 41 nsew
rlabel locali s 29933 -59298 29967 -59132 8 VDD
port 41 nsew
rlabel locali s 29716 -59298 29750 -58931 8 VDD
port 41 nsew
rlabel locali s 29520 -59348 29554 -58931 8 VDD
port 41 nsew
rlabel locali s 29324 -59348 29358 -58931 8 VDD
port 41 nsew
rlabel locali s 28485 -59457 28657 -59267 8 VDD
port 41 nsew
rlabel locali s 28303 -59267 29021 -59168 8 VDD
port 41 nsew
rlabel locali s 28939 -59168 28973 -58902 8 VDD
port 41 nsew
rlabel locali s 28743 -59168 28777 -58902 8 VDD
port 41 nsew
rlabel locali s 28547 -59168 28581 -58902 8 VDD
port 41 nsew
rlabel locali s 28351 -59168 28385 -58902 8 VDD
port 41 nsew
rlabel locali s 30846 -58192 31248 -58126 8 VDD
port 41 nsew
rlabel locali s 26110 -59637 26199 -57482 8 VDD
port 41 nsew
rlabel locali s 25972 -59637 26006 -58802 8 VDD
port 41 nsew
rlabel locali s 25776 -59637 25810 -58802 8 VDD
port 41 nsew
rlabel locali s 25572 -59637 25606 -58802 8 VDD
port 41 nsew
rlabel locali s 25376 -59637 25410 -58802 8 VDD
port 41 nsew
rlabel locali s 24972 -59637 25006 -58802 8 VDD
port 41 nsew
rlabel locali s 24776 -59637 24810 -58802 8 VDD
port 41 nsew
rlabel locali s 24572 -59637 24606 -58802 8 VDD
port 41 nsew
rlabel locali s 24376 -59637 24410 -58802 8 VDD
port 41 nsew
rlabel locali s 23972 -59637 24006 -58802 8 VDD
port 41 nsew
rlabel locali s 23776 -59637 23810 -58802 8 VDD
port 41 nsew
rlabel locali s 23572 -59637 23606 -58802 8 VDD
port 41 nsew
rlabel locali s 23376 -59637 23410 -58802 8 VDD
port 41 nsew
rlabel locali s 22888 -59637 22922 -59373 8 VDD
port 41 nsew
rlabel locali s 22692 -59664 22726 -59373 8 VDD
port 41 nsew
rlabel locali s 22496 -59664 22530 -59373 8 VDD
port 41 nsew
rlabel locali s 22193 -59664 22267 -59658 8 VDD
port 41 nsew
rlabel locali s 21963 -59672 21997 -59380 8 VDD
port 41 nsew
rlabel locali s 21767 -59672 21801 -59380 8 VDD
port 41 nsew
rlabel locali s 21512 -59672 21575 -59658 8 VDD
port 41 nsew
rlabel locali s 21225 -59676 21259 -59380 8 VDD
port 41 nsew
rlabel locali s 21029 -59676 21063 -59380 8 VDD
port 41 nsew
rlabel locali s 20833 -59676 20867 -59380 8 VDD
port 41 nsew
rlabel locali s 20637 -59676 20671 -59380 8 VDD
port 41 nsew
rlabel locali s 17945 -59676 20478 -59664 8 VDD
port 41 nsew
rlabel locali s 20392 -59664 20478 -59656 8 VDD
port 41 nsew
rlabel locali s 19911 -59664 19959 -59531 8 VDD
port 41 nsew
rlabel locali s 19714 -59664 19762 -59537 8 VDD
port 41 nsew
rlabel locali s 19917 -59531 19951 -59146 8 VDD
port 41 nsew
rlabel locali s 19721 -59537 19755 -59146 8 VDD
port 41 nsew
rlabel locali s 18965 -59664 19013 -59531 8 VDD
port 41 nsew
rlabel locali s 18768 -59664 18816 -59537 8 VDD
port 41 nsew
rlabel locali s 8753 -59778 8787 -59588 8 VDD
port 41 nsew
rlabel locali s 8551 -59900 8597 -59766 8 VDD
port 41 nsew
rlabel locali s 8438 -59900 8484 -59776 8 VDD
port 41 nsew
rlabel locali s 8557 -59766 8591 -59588 8 VDD
port 41 nsew
rlabel locali s 8444 -59776 8478 -59588 8 VDD
port 41 nsew
rlabel locali s 8242 -59900 8288 -59771 8 VDD
port 41 nsew
rlabel locali s 8129 -59900 8175 -59775 8 VDD
port 41 nsew
rlabel locali s 8248 -59771 8282 -59588 8 VDD
port 41 nsew
rlabel locali s 8134 -59775 8168 -59588 8 VDD
port 41 nsew
rlabel locali s 7931 -59900 7977 -59771 8 VDD
port 41 nsew
rlabel locali s 7741 -59900 7864 -59860 8 VDD
port 41 nsew
rlabel locali s 6525 -59997 6648 -59964 8 VDD
port 41 nsew
rlabel locali s 5169 -60002 5292 -59969 8 VDD
port 41 nsew
rlabel locali s 5169 -59969 6065 -59964 8 VDD
port 41 nsew
rlabel locali s 5169 -59964 6648 -59896 8 VDD
port 41 nsew
rlabel locali s 5993 -59896 6648 -59895 8 VDD
port 41 nsew
rlabel locali s 6525 -59895 6648 -59861 8 VDD
port 41 nsew
rlabel locali s 7742 -59860 7782 -59771 8 VDD
port 41 nsew
rlabel locali s 7938 -59771 7972 -59588 8 VDD
port 41 nsew
rlabel locali s 7742 -59771 7776 -59588 8 VDD
port 41 nsew
rlabel locali s 6581 -59861 6615 -59599 8 VDD
port 41 nsew
rlabel locali s 6385 -59895 6419 -59599 8 VDD
port 41 nsew
rlabel locali s 6189 -59895 6223 -59599 8 VDD
port 41 nsew
rlabel locali s 5993 -59895 6027 -59599 8 VDD
port 41 nsew
rlabel locali s 5169 -59896 5490 -59891 8 VDD
port 41 nsew
rlabel locali s 5451 -59891 5485 -59599 8 VDD
port 41 nsew
rlabel locali s 5169 -59891 5292 -59866 8 VDD
port 41 nsew
rlabel locali s 4768 -60000 4891 -59955 8 VDD
port 41 nsew
rlabel locali s 4430 -59955 4891 -59940 8 VDD
port 41 nsew
rlabel locali s 3540 -59977 3663 -59940 8 VDD
port 41 nsew
rlabel locali s 3540 -59940 4891 -59891 8 VDD
port 41 nsew
rlabel locali s 5255 -59866 5289 -59599 8 VDD
port 41 nsew
rlabel locali s 4768 -59891 4891 -59864 8 VDD
port 41 nsew
rlabel locali s 18971 -59531 19005 -59146 8 VDD
port 41 nsew
rlabel locali s 18775 -59537 18809 -59146 8 VDD
port 41 nsew
rlabel locali s 4828 -59864 4862 -59474 8 VDD
port 41 nsew
rlabel locali s 4632 -59891 4666 -59474 8 VDD
port 41 nsew
rlabel locali s 3540 -59891 4470 -59841 8 VDD
port 41 nsew
rlabel locali s 3151 -59976 3274 -59962 8 VDD
port 41 nsew
rlabel locali s 1108 -60770 1223 -59962 8 VDD
port 41 nsew
rlabel locali s -1380 -60798 -1257 -60662 2 VDD
port 41 nsew
rlabel locali s -16311 -60807 -15424 -60757 2 VDD
port 41 nsew
rlabel locali s -16507 -61174 -16473 -60757 2 VDD
port 41 nsew
rlabel locali s -16703 -61174 -16669 -60757 2 VDD
port 41 nsew
rlabel locali s -17088 -61203 -17054 -60937 2 VDD
port 41 nsew
rlabel locali s -17284 -61203 -17250 -60937 2 VDD
port 41 nsew
rlabel locali s -17480 -61203 -17446 -60937 2 VDD
port 41 nsew
rlabel locali s -17676 -61203 -17642 -60937 2 VDD
port 41 nsew
rlabel locali s -17724 -60937 -17006 -60838 2 VDD
port 41 nsew
rlabel locali s -16713 -60757 -15424 -60708 2 VDD
port 41 nsew
rlabel locali s -16713 -60708 -16271 -60694 2 VDD
port 41 nsew
rlabel locali s -16714 -60694 -16271 -60665 2 VDD
port 41 nsew
rlabel locali s 173 -59989 296 -59962 8 VDD
port 41 nsew
rlabel locali s 173 -59962 3274 -59883 8 VDD
port 41 nsew
rlabel locali s 4436 -59841 4470 -59474 8 VDD
port 41 nsew
rlabel locali s 4219 -59841 4253 -59675 8 VDD
port 41 nsew
rlabel locali s 4023 -59841 4057 -59675 8 VDD
port 41 nsew
rlabel locali s 3827 -59841 3861 -59675 8 VDD
port 41 nsew
rlabel locali s 3631 -59841 3665 -59675 8 VDD
port 41 nsew
rlabel locali s 3151 -59883 3274 -59840 8 VDD
port 41 nsew
rlabel locali s 3223 -59840 3257 -59476 8 VDD
port 41 nsew
rlabel locali s 3027 -59883 3061 -59476 8 VDD
port 41 nsew
rlabel locali s 1978 -59883 2865 -59843 8 VDD
port 41 nsew
rlabel locali s 2831 -59843 2865 -59476 8 VDD
port 41 nsew
rlabel locali s 2614 -59843 2648 -59677 8 VDD
port 41 nsew
rlabel locali s 2418 -59843 2452 -59677 8 VDD
port 41 nsew
rlabel locali s 2222 -59843 2256 -59677 8 VDD
port 41 nsew
rlabel locali s 2026 -59843 2060 -59677 8 VDD
port 41 nsew
rlabel locali s 1619 -59883 1653 -59590 8 VDD
port 41 nsew
rlabel locali s 1423 -59883 1457 -59590 8 VDD
port 41 nsew
rlabel locali s 1227 -59883 1261 -59590 8 VDD
port 41 nsew
rlabel locali s 1031 -59883 1065 -59590 8 VDD
port 41 nsew
rlabel locali s 173 -59883 528 -59882 8 VDD
port 41 nsew
rlabel locali s 489 -59882 523 -59590 8 VDD
port 41 nsew
rlabel locali s 173 -59882 327 -59853 8 VDD
port 41 nsew
rlabel locali s -121 -59988 2 -59966 2 VDD
port 41 nsew
rlabel locali s -1376 -60662 -1261 -59966 2 VDD
port 41 nsew
rlabel locali s -3947 -60654 -3824 -60518 2 VDD
port 41 nsew
rlabel locali s -16714 -60665 -16096 -60648 2 VDD
port 41 nsew
rlabel locali s -17542 -60838 -17370 -60667 2 VDD
port 41 nsew
rlabel locali s -18946 -61662 -18774 -60667 2 VDD
port 41 nsew
rlabel locali s -18946 -60667 -17370 -60648 2 VDD
port 41 nsew
rlabel locali s -18946 -60648 -15601 -60537 2 VDD
port 41 nsew
rlabel locali s -2791 -59967 -2318 -59966 2 VDD
port 41 nsew
rlabel locali s -3942 -60518 -3827 -59966 2 VDD
port 41 nsew
rlabel locali s -18946 -60537 -15497 -60495 2 VDD
port 41 nsew
rlabel locali s -16266 -60495 -15497 -60471 2 VDD
port 41 nsew
rlabel locali s -17310 -60495 -17084 -60488 2 VDD
port 41 nsew
rlabel locali s -17273 -60488 -17084 -60481 2 VDD
port 41 nsew
rlabel locali s -15643 -60471 -15598 -60347 2 VDD
port 41 nsew
rlabel locali s -16065 -60471 -16020 -60348 2 VDD
port 41 nsew
rlabel locali s -6113 -59969 -5009 -59966 2 VDD
port 41 nsew
rlabel locali s -6113 -59966 2 -59903 2 VDD
port 41 nsew
rlabel locali s -1384 -59903 2 -59898 2 VDD
port 41 nsew
rlabel locali s -4084 -59903 -2318 -59899 2 VDD
port 41 nsew
rlabel locali s -6113 -59903 -5009 -59901 2 VDD
port 41 nsew
rlabel locali s -4084 -59899 -2631 -59898 2 VDD
port 41 nsew
rlabel locali s -5826 -59901 -5331 -59898 2 VDD
port 41 nsew
rlabel locali s 293 -59853 327 -59590 8 VDD
port 41 nsew
rlabel locali s -121 -59898 2 -59852 2 VDD
port 41 nsew
rlabel locali s -49 -59852 -15 -59607 2 VDD
port 41 nsew
rlabel locali s -245 -59898 -211 -59607 2 VDD
port 41 nsew
rlabel locali s -441 -59898 -407 -59607 2 VDD
port 41 nsew
rlabel locali s -931 -59898 -897 -59607 2 VDD
port 41 nsew
rlabel locali s -1127 -59898 -1093 -59607 2 VDD
port 41 nsew
rlabel locali s -1323 -59898 -1289 -59607 2 VDD
port 41 nsew
rlabel locali s -2674 -59898 -2640 -59607 2 VDD
port 41 nsew
rlabel locali s -2870 -59898 -2836 -59607 2 VDD
port 41 nsew
rlabel locali s -3066 -59898 -3032 -59607 2 VDD
port 41 nsew
rlabel locali s -3631 -59898 -3597 -59607 2 VDD
port 41 nsew
rlabel locali s -3827 -59898 -3793 -59607 2 VDD
port 41 nsew
rlabel locali s -4023 -59898 -3989 -59607 2 VDD
port 41 nsew
rlabel locali s -5374 -59898 -5340 -59607 2 VDD
port 41 nsew
rlabel locali s -5570 -59898 -5536 -59607 2 VDD
port 41 nsew
rlabel locali s -5766 -59898 -5732 -59607 2 VDD
port 41 nsew
rlabel locali s 22938 -58280 22972 -57763 8 VDD
port 41 nsew
rlabel locali s 22742 -58280 22776 -57763 8 VDD
port 41 nsew
rlabel locali s 22546 -58280 22580 -57763 8 VDD
port 41 nsew
rlabel locali s -1935 -58497 -1901 -58206 2 VDD
port 41 nsew
rlabel locali s -2131 -58497 -2097 -58206 2 VDD
port 41 nsew
rlabel locali s -2327 -58497 -2293 -58206 2 VDD
port 41 nsew
rlabel locali s -2772 -58497 -2738 -58206 2 VDD
port 41 nsew
rlabel locali s -2968 -58497 -2934 -58206 2 VDD
port 41 nsew
rlabel locali s -3164 -58497 -3130 -58206 2 VDD
port 41 nsew
rlabel locali s -4635 -58497 -4601 -58206 2 VDD
port 41 nsew
rlabel locali s -4831 -58497 -4797 -58206 2 VDD
port 41 nsew
rlabel locali s -5027 -58497 -4993 -58206 2 VDD
port 41 nsew
rlabel locali s -5472 -58497 -5438 -58206 2 VDD
port 41 nsew
rlabel locali s -5668 -58497 -5634 -58206 2 VDD
port 41 nsew
rlabel locali s -5864 -58497 -5830 -58206 2 VDD
port 41 nsew
rlabel locali s -6113 -59901 -6024 -58206 2 VDD
port 41 nsew
rlabel locali s -15636 -60347 -15602 -59755 2 VDD
port 41 nsew
rlabel locali s -16059 -60348 -16025 -59755 2 VDD
port 41 nsew
rlabel locali s -16260 -60471 -16215 -60345 2 VDD
port 41 nsew
rlabel locali s -17712 -60447 -17270 -60432 2 VDD
port 41 nsew
rlabel locali s -17712 -60432 -16423 -60383 2 VDD
port 41 nsew
rlabel locali s -16255 -60345 -16221 -59755 2 VDD
port 41 nsew
rlabel locali s -17310 -60383 -16423 -60333 2 VDD
port 41 nsew
rlabel locali s -16505 -60333 -16471 -60167 2 VDD
port 41 nsew
rlabel locali s -16701 -60333 -16667 -60167 2 VDD
port 41 nsew
rlabel locali s -16897 -60333 -16863 -60167 2 VDD
port 41 nsew
rlabel locali s -17093 -60333 -17059 -60167 2 VDD
port 41 nsew
rlabel locali s -17310 -60333 -17276 -59966 2 VDD
port 41 nsew
rlabel locali s -17506 -60383 -17472 -59966 2 VDD
port 41 nsew
rlabel locali s -17702 -60383 -17668 -59966 2 VDD
port 41 nsew
rlabel locali s -10665 -59700 -10192 -59699 2 VDD
port 41 nsew
rlabel locali s -13987 -59702 -12883 -59699 2 VDD
port 41 nsew
rlabel locali s -13987 -59699 -7880 -59636 2 VDD
port 41 nsew
rlabel locali s -9258 -59636 -7880 -59631 2 VDD
port 41 nsew
rlabel locali s -11958 -59636 -10192 -59632 2 VDD
port 41 nsew
rlabel locali s -13987 -59636 -12883 -59634 2 VDD
port 41 nsew
rlabel locali s -11958 -59632 -10505 -59631 2 VDD
port 41 nsew
rlabel locali s -13700 -59634 -13205 -59631 2 VDD
port 41 nsew
rlabel locali s -7923 -59631 -7889 -59340 2 VDD
port 41 nsew
rlabel locali s -8119 -59631 -8085 -59340 2 VDD
port 41 nsew
rlabel locali s -8315 -59631 -8281 -59340 2 VDD
port 41 nsew
rlabel locali s -8805 -59631 -8771 -59340 2 VDD
port 41 nsew
rlabel locali s -9001 -59631 -8967 -59340 2 VDD
port 41 nsew
rlabel locali s -9197 -59631 -9163 -59340 2 VDD
port 41 nsew
rlabel locali s -10548 -59631 -10514 -59340 2 VDD
port 41 nsew
rlabel locali s -10744 -59631 -10710 -59340 2 VDD
port 41 nsew
rlabel locali s -10940 -59631 -10906 -59340 2 VDD
port 41 nsew
rlabel locali s -11505 -59631 -11471 -59340 2 VDD
port 41 nsew
rlabel locali s -11701 -59631 -11667 -59340 2 VDD
port 41 nsew
rlabel locali s -11897 -59631 -11863 -59340 2 VDD
port 41 nsew
rlabel locali s -13248 -59631 -13214 -59340 2 VDD
port 41 nsew
rlabel locali s -13444 -59631 -13410 -59340 2 VDD
port 41 nsew
rlabel locali s -13640 -59631 -13606 -59340 2 VDD
port 41 nsew
rlabel locali s -13987 -59634 -13898 -58731 2 VDD
port 41 nsew
rlabel locali s -18908 -59445 -18874 -59060 2 VDD
port 41 nsew
rlabel locali s -18914 -59060 -18866 -58927 2 VDD
port 41 nsew
rlabel locali s -19104 -59445 -19070 -59054 2 VDD
port 41 nsew
rlabel locali s -19813 -59444 -19779 -59059 2 VDD
port 41 nsew
rlabel locali s -19111 -59054 -19063 -58927 2 VDD
port 41 nsew
rlabel locali s -19116 -58927 -18562 -58899 2 VDD
port 41 nsew
rlabel locali s -19819 -59059 -19771 -58926 2 VDD
port 41 nsew
rlabel locali s -20009 -59444 -19975 -59053 2 VDD
port 41 nsew
rlabel locali s -21019 -59715 -20985 -59131 2 VDD
port 41 nsew
rlabel locali s -20016 -59053 -19968 -58926 2 VDD
port 41 nsew
rlabel locali s -21028 -59131 -20975 -59003 2 VDD
port 41 nsew
rlabel locali s -21215 -59715 -21181 -59115 2 VDD
port 41 nsew
rlabel locali s -27269 -59664 -27203 -59463 2 VDD
port 41 nsew
rlabel locali s -27836 -59668 -27341 -59634 2 VDD
port 41 nsew
rlabel locali s -27389 -59634 -27341 -59463 2 VDD
port 41 nsew
rlabel locali s -27389 -59463 -27203 -59432 2 VDD
port 41 nsew
rlabel locali s -27836 -59432 -27203 -59404 2 VDD
port 41 nsew
rlabel locali s -21224 -59115 -21171 -59003 2 VDD
port 41 nsew
rlabel locali s -19117 -58899 -18562 -58858 2 VDD
port 41 nsew
rlabel locali s -19117 -58858 -18564 -58731 2 VDD
port 41 nsew
rlabel locali s -20021 -58926 -19467 -58857 2 VDD
port 41 nsew
rlabel locali s -21224 -59003 -20356 -58870 2 VDD
port 41 nsew
rlabel locali s -27269 -59404 -27203 -58875 2 VDD
port 41 nsew
rlabel locali s -27836 -59404 -27341 -59398 2 VDD
port 41 nsew
rlabel locali s -27389 -59398 -27341 -59196 2 VDD
port 41 nsew
rlabel locali s -27836 -59196 -27341 -59162 2 VDD
port 41 nsew
rlabel locali s -27389 -59162 -27341 -59066 2 VDD
port 41 nsew
rlabel locali s -27836 -59066 -27341 -59032 2 VDD
port 41 nsew
rlabel locali s -27389 -59032 -27341 -58875 2 VDD
port 41 nsew
rlabel locali s -20006 -58857 -19488 -58731 2 VDD
port 41 nsew
rlabel locali s -21164 -58870 -20382 -58731 2 VDD
port 41 nsew
rlabel locali s -27389 -58875 -27203 -58830 2 VDD
port 41 nsew
rlabel locali s -27836 -58830 -27203 -58816 2 VDD
port 41 nsew
rlabel locali s -3642 -58206 -1840 -58201 2 VDD
port 41 nsew
rlabel locali s -6113 -58206 -4540 -58201 2 VDD
port 41 nsew
rlabel locali s -6113 -58201 -888 -58138 2 VDD
port 41 nsew
rlabel locali s 22536 -57763 22978 -57699 8 VDD
port 41 nsew
rlabel locali s 25095 -57482 26199 -57479 8 VDD
port 41 nsew
rlabel locali s 22594 -57699 22826 -57480 8 VDD
port 41 nsew
rlabel locali s 22404 -57480 22877 -57479 8 VDD
port 41 nsew
rlabel locali s 20092 -57479 26199 -57416 8 VDD
port 41 nsew
rlabel locali s 25095 -57416 26199 -57414 8 VDD
port 41 nsew
rlabel locali s 34079 -56168 39113 -56133 8 VDD
port 41 nsew
rlabel locali s 33117 -56455 33151 -56163 8 VDD
port 41 nsew
rlabel locali s 32921 -56455 32955 -56165 8 VDD
port 41 nsew
rlabel locali s 32693 -56655 32727 -56180 8 VDD
port 41 nsew
rlabel locali s 32563 -56655 32597 -56183 8 VDD
port 41 nsew
rlabel locali s 39051 -56133 39113 -56105 8 VDD
port 41 nsew
rlabel locali s 34079 -56133 38978 -56126 8 VDD
port 41 nsew
rlabel locali s 39842 -56088 39959 -56078 8 VDD
port 41 nsew
rlabel locali s 39279 -56088 39377 -56085 8 VDD
port 41 nsew
rlabel locali s 39842 -56078 40247 -56014 8 VDD
port 41 nsew
rlabel locali s 34079 -56126 38874 -56015 8 VDD
port 41 nsew
rlabel locali s 58270 -55966 65689 -55954 8 VDD
port 41 nsew
rlabel locali s 55823 -55974 56265 -55960 8 VDD
port 41 nsew
rlabel locali s 66657 -55953 74842 -55937 8 VDD
port 41 nsew
rlabel locali s 64576 -55954 65194 -55937 8 VDD
port 41 nsew
rlabel locali s 75810 -55936 84206 -55899 8 VDD
port 41 nsew
rlabel locali s 73729 -55937 74347 -55920 8 VDD
port 41 nsew
rlabel locali s 85174 -55898 86927 -55897 8 VDD
port 41 nsew
rlabel locali s 85174 -55897 87973 -55845 8 VDD
port 41 nsew
rlabel locali s 83093 -55899 83711 -55882 8 VDD
port 41 nsew
rlabel locali s 83093 -55882 83536 -55853 8 VDD
port 41 nsew
rlabel locali s 75810 -55899 82437 -55883 8 VDD
port 41 nsew
rlabel locali s 73729 -55920 74172 -55891 8 VDD
port 41 nsew
rlabel locali s 66657 -55937 73073 -55900 8 VDD
port 41 nsew
rlabel locali s 64576 -55937 65019 -55908 8 VDD
port 41 nsew
rlabel locali s 85541 -55845 87973 -55775 8 VDD
port 41 nsew
rlabel locali s 83094 -55853 83536 -55839 8 VDD
port 41 nsew
rlabel locali s 83094 -55839 84383 -55790 8 VDD
port 41 nsew
rlabel locali s 76177 -55883 82437 -55813 8 VDD
port 41 nsew
rlabel locali s 73730 -55891 74172 -55877 8 VDD
port 41 nsew
rlabel locali s 73730 -55877 75019 -55828 8 VDD
port 41 nsew
rlabel locali s 67024 -55900 73073 -55830 8 VDD
port 41 nsew
rlabel locali s 64577 -55908 65019 -55894 8 VDD
port 41 nsew
rlabel locali s 64577 -55894 65866 -55845 8 VDD
port 41 nsew
rlabel locali s 58270 -55954 63920 -55896 8 VDD
port 41 nsew
rlabel locali s 55823 -55960 57112 -55911 8 VDD
port 41 nsew
rlabel locali s 49072 -56000 55166 -55930 8 VDD
port 41 nsew
rlabel locali s 46625 -56008 47067 -55994 8 VDD
port 41 nsew
rlabel locali s 46625 -55994 47914 -55945 8 VDD
port 41 nsew
rlabel locali s 39842 -56014 45968 -55961 8 VDD
port 41 nsew
rlabel locali s 37761 -56015 38379 -55998 8 VDD
port 41 nsew
rlabel locali s 37761 -55998 38204 -55969 8 VDD
port 41 nsew
rlabel locali s 87299 -55775 87774 -51863 8 VDD
port 41 nsew
rlabel locali s 83496 -55790 84383 -55740 8 VDD
port 41 nsew
rlabel locali s 84301 -55740 84335 -55574 8 VDD
port 41 nsew
rlabel locali s 84105 -55740 84139 -55574 8 VDD
port 41 nsew
rlabel locali s 83909 -55740 83943 -55574 8 VDD
port 41 nsew
rlabel locali s 83713 -55740 83747 -55574 8 VDD
port 41 nsew
rlabel locali s 83496 -55740 83530 -55373 8 VDD
port 41 nsew
rlabel locali s 83300 -55790 83334 -55373 8 VDD
port 41 nsew
rlabel locali s 83104 -55790 83138 -55373 8 VDD
port 41 nsew
rlabel locali s 77524 -55813 82437 -55709 8 VDD
port 41 nsew
rlabel locali s 74132 -55828 75019 -55778 8 VDD
port 41 nsew
rlabel locali s 77524 -55709 82801 -55654 8 VDD
port 41 nsew
rlabel locali s 82083 -55654 82801 -55610 8 VDD
port 41 nsew
rlabel locali s 74937 -55778 74971 -55612 8 VDD
port 41 nsew
rlabel locali s 74741 -55778 74775 -55612 8 VDD
port 41 nsew
rlabel locali s 74545 -55778 74579 -55612 8 VDD
port 41 nsew
rlabel locali s 74349 -55778 74383 -55612 8 VDD
port 41 nsew
rlabel locali s 82719 -55610 82753 -55344 8 VDD
port 41 nsew
rlabel locali s 82523 -55610 82557 -55344 8 VDD
port 41 nsew
rlabel locali s 82327 -55610 82361 -55344 8 VDD
port 41 nsew
rlabel locali s 82131 -55610 82165 -55344 8 VDD
port 41 nsew
rlabel locali s 74132 -55778 74166 -55411 8 VDD
port 41 nsew
rlabel locali s 73936 -55828 73970 -55411 8 VDD
port 41 nsew
rlabel locali s 73740 -55828 73774 -55411 8 VDD
port 41 nsew
rlabel locali s 68362 -55830 73073 -55747 8 VDD
port 41 nsew
rlabel locali s 64979 -55845 65866 -55795 8 VDD
port 41 nsew
rlabel locali s 68362 -55747 73437 -55723 8 VDD
port 41 nsew
rlabel locali s 72719 -55723 73437 -55648 8 VDD
port 41 nsew
rlabel locali s 73355 -55648 73389 -55382 8 VDD
port 41 nsew
rlabel locali s 73159 -55648 73193 -55382 8 VDD
port 41 nsew
rlabel locali s 72963 -55648 72997 -55382 8 VDD
port 41 nsew
rlabel locali s 72767 -55648 72801 -55382 8 VDD
port 41 nsew
rlabel locali s 65784 -55795 65818 -55629 8 VDD
port 41 nsew
rlabel locali s 65588 -55795 65622 -55629 8 VDD
port 41 nsew
rlabel locali s 65392 -55795 65426 -55629 8 VDD
port 41 nsew
rlabel locali s 65196 -55795 65230 -55629 8 VDD
port 41 nsew
rlabel locali s 64979 -55795 65013 -55428 8 VDD
port 41 nsew
rlabel locali s 64783 -55845 64817 -55428 8 VDD
port 41 nsew
rlabel locali s 64587 -55845 64621 -55428 8 VDD
port 41 nsew
rlabel locali s 59615 -55896 63920 -55764 8 VDD
port 41 nsew
rlabel locali s 56225 -55911 57112 -55861 8 VDD
port 41 nsew
rlabel locali s 59615 -55764 64284 -55702 8 VDD
port 41 nsew
rlabel locali s 63566 -55702 64284 -55665 8 VDD
port 41 nsew
rlabel locali s 57030 -55861 57064 -55695 8 VDD
port 41 nsew
rlabel locali s 56834 -55861 56868 -55695 8 VDD
port 41 nsew
rlabel locali s 56638 -55861 56672 -55695 8 VDD
port 41 nsew
rlabel locali s 56442 -55861 56476 -55695 8 VDD
port 41 nsew
rlabel locali s 64202 -55665 64236 -55399 8 VDD
port 41 nsew
rlabel locali s 64006 -55665 64040 -55399 8 VDD
port 41 nsew
rlabel locali s 63810 -55665 63844 -55399 8 VDD
port 41 nsew
rlabel locali s 63614 -55665 63648 -55399 8 VDD
port 41 nsew
rlabel locali s 56225 -55861 56259 -55494 8 VDD
port 41 nsew
rlabel locali s 56029 -55911 56063 -55494 8 VDD
port 41 nsew
rlabel locali s 55833 -55911 55867 -55494 8 VDD
port 41 nsew
rlabel locali s 50432 -55930 55166 -55830 8 VDD
port 41 nsew
rlabel locali s 47027 -55945 47914 -55895 8 VDD
port 41 nsew
rlabel locali s 50432 -55830 55530 -55799 8 VDD
port 41 nsew
rlabel locali s 54812 -55799 55530 -55731 8 VDD
port 41 nsew
rlabel locali s 55448 -55731 55482 -55465 8 VDD
port 41 nsew
rlabel locali s 55252 -55731 55286 -55465 8 VDD
port 41 nsew
rlabel locali s 55056 -55731 55090 -55465 8 VDD
port 41 nsew
rlabel locali s 54860 -55731 54894 -55465 8 VDD
port 41 nsew
rlabel locali s 47832 -55895 47866 -55729 8 VDD
port 41 nsew
rlabel locali s 47636 -55895 47670 -55729 8 VDD
port 41 nsew
rlabel locali s 47440 -55895 47474 -55729 8 VDD
port 41 nsew
rlabel locali s 47244 -55895 47278 -55729 8 VDD
port 41 nsew
rlabel locali s 47027 -55895 47061 -55528 8 VDD
port 41 nsew
rlabel locali s 46831 -55945 46865 -55528 8 VDD
port 41 nsew
rlabel locali s 46635 -55945 46669 -55528 8 VDD
port 41 nsew
rlabel locali s 40209 -55961 45968 -55891 8 VDD
port 41 nsew
rlabel locali s 37762 -55969 38204 -55955 8 VDD
port 41 nsew
rlabel locali s 37762 -55955 39051 -55906 8 VDD
port 41 nsew
rlabel locali s 41581 -55891 45968 -55864 8 VDD
port 41 nsew
rlabel locali s 41581 -55864 46332 -55849 8 VDD
port 41 nsew
rlabel locali s 38164 -55906 39051 -55856 8 VDD
port 41 nsew
rlabel locali s 45614 -55849 46332 -55765 8 VDD
port 41 nsew
rlabel locali s 46250 -55765 46284 -55499 8 VDD
port 41 nsew
rlabel locali s 46054 -55765 46088 -55499 8 VDD
port 41 nsew
rlabel locali s 45858 -55765 45892 -55499 8 VDD
port 41 nsew
rlabel locali s 45662 -55765 45696 -55499 8 VDD
port 41 nsew
rlabel locali s 38969 -55856 39003 -55690 8 VDD
port 41 nsew
rlabel locali s 38773 -55856 38807 -55690 8 VDD
port 41 nsew
rlabel locali s 38577 -55856 38611 -55690 8 VDD
port 41 nsew
rlabel locali s 38381 -55856 38415 -55690 8 VDD
port 41 nsew
rlabel locali s 38164 -55856 38198 -55489 8 VDD
port 41 nsew
rlabel locali s 37968 -55906 38002 -55489 8 VDD
port 41 nsew
rlabel locali s 37772 -55906 37806 -55489 8 VDD
port 41 nsew
rlabel locali s 36933 -56015 37105 -55825 8 VDD
port 41 nsew
rlabel locali s 34079 -56015 34201 -56002 8 VDD
port 41 nsew
rlabel locali s 33112 -56163 33155 -56003 8 VDD
port 41 nsew
rlabel locali s 32915 -56165 32958 -56003 8 VDD
port 41 nsew
rlabel locali s 32684 -56180 32734 -56003 8 VDD
port 41 nsew
rlabel locali s 32558 -56183 32608 -56003 8 VDD
port 41 nsew
rlabel locali s 31968 -56655 32002 -56160 8 VDD
port 41 nsew
rlabel locali s 31772 -56655 31806 -56162 8 VDD
port 41 nsew
rlabel locali s 30399 -56897 30433 -56305 8 VDD
port 41 nsew
rlabel locali s 30839 -56200 30937 -56194 8 VDD
port 41 nsew
rlabel locali s 31966 -56160 32004 -56003 8 VDD
port 41 nsew
rlabel locali s 31769 -56162 31807 -56067 8 VDD
port 41 nsew
rlabel locali s 30839 -56194 31519 -56077 8 VDD
port 41 nsew
rlabel locali s 30611 -56188 30673 -56174 8 VDD
port 41 nsew
rlabel locali s 30392 -56305 30437 -56181 8 VDD
port 41 nsew
rlabel locali s 29976 -56897 30010 -56304 8 VDD
port 41 nsew
rlabel locali s 29780 -56897 29814 -56307 8 VDD
port 41 nsew
rlabel locali s 29530 -56485 29564 -56319 8 VDD
port 41 nsew
rlabel locali s 29334 -56485 29368 -56319 8 VDD
port 41 nsew
rlabel locali s 29138 -56485 29172 -56319 8 VDD
port 41 nsew
rlabel locali s 28942 -56485 28976 -56319 8 VDD
port 41 nsew
rlabel locali s 28725 -56686 28759 -56319 8 VDD
port 41 nsew
rlabel locali s 29970 -56304 30015 -56181 8 VDD
port 41 nsew
rlabel locali s 29775 -56307 29820 -56181 8 VDD
port 41 nsew
rlabel locali s 28725 -56319 29612 -56269 8 VDD
port 41 nsew
rlabel locali s 28529 -56686 28563 -56269 8 VDD
port 41 nsew
rlabel locali s 28333 -56686 28367 -56269 8 VDD
port 41 nsew
rlabel locali s 28323 -56269 29612 -56220 8 VDD
port 41 nsew
rlabel locali s 28323 -56220 28765 -56205 8 VDD
port 41 nsew
rlabel locali s 29769 -56181 30538 -56174 8 VDD
port 41 nsew
rlabel locali s 29769 -56174 30673 -56157 8 VDD
port 41 nsew
rlabel locali s 28762 -56171 28951 -56164 8 VDD
port 41 nsew
rlabel locali s 28725 -56164 28951 -56157 8 VDD
port 41 nsew
rlabel locali s 28323 -56157 30673 -56122 8 VDD
port 41 nsew
rlabel locali s 30611 -56122 30673 -56094 8 VDD
port 41 nsew
rlabel locali s 28323 -56122 30538 -56115 8 VDD
port 41 nsew
rlabel locali s 31402 -56077 31519 -56067 8 VDD
port 41 nsew
rlabel locali s 30839 -56077 30937 -56074 8 VDD
port 41 nsew
rlabel locali s 31402 -56067 31807 -56003 8 VDD
port 41 nsew
rlabel locali s 28323 -56115 30434 -56073 8 VDD
port 41 nsew
rlabel locali s 26110 -57414 26199 -56073 8 VDD
port 41 nsew
rlabel locali s 25417 -57414 25912 -57411 8 VDD
port 41 nsew
rlabel locali s 22404 -57416 24170 -57412 8 VDD
port 41 nsew
rlabel locali s 22717 -57412 24170 -57411 8 VDD
port 41 nsew
rlabel locali s 20092 -57416 21470 -57411 8 VDD
port 41 nsew
rlabel locali s 25818 -57411 25852 -57120 8 VDD
port 41 nsew
rlabel locali s 25622 -57411 25656 -57120 8 VDD
port 41 nsew
rlabel locali s 25426 -57411 25460 -57120 8 VDD
port 41 nsew
rlabel locali s 24075 -57411 24109 -57120 8 VDD
port 41 nsew
rlabel locali s 23879 -57411 23913 -57120 8 VDD
port 41 nsew
rlabel locali s 23683 -57411 23717 -57120 8 VDD
port 41 nsew
rlabel locali s 23118 -57411 23152 -57120 8 VDD
port 41 nsew
rlabel locali s 22922 -57411 22956 -57120 8 VDD
port 41 nsew
rlabel locali s 22726 -57411 22760 -57120 8 VDD
port 41 nsew
rlabel locali s 21375 -57411 21409 -57120 8 VDD
port 41 nsew
rlabel locali s 21179 -57411 21213 -57120 8 VDD
port 41 nsew
rlabel locali s 20983 -57411 21017 -57120 8 VDD
port 41 nsew
rlabel locali s 20493 -57411 20527 -57120 8 VDD
port 41 nsew
rlabel locali s 20297 -57411 20331 -57120 8 VDD
port 41 nsew
rlabel locali s 20101 -57411 20135 -57120 8 VDD
port 41 nsew
rlabel locali s 18771 -57445 19639 -57312 8 VDD
port 41 nsew
rlabel locali s 18967 -57312 19020 -57184 8 VDD
port 41 nsew
rlabel locali s 18771 -57312 18824 -57200 8 VDD
port 41 nsew
rlabel locali s -1606 -58138 -1337 -57210 2 VDD
port 41 nsew
rlabel locali s -2637 -58138 -2368 -57210 2 VDD
port 41 nsew
rlabel locali s -3540 -58138 -3271 -57210 2 VDD
port 41 nsew
rlabel locali s -4402 -58138 -4133 -57210 2 VDD
port 41 nsew
rlabel locali s -5279 -58138 -5010 -57210 2 VDD
port 41 nsew
rlabel locali s -5825 -58138 -5556 -57210 2 VDD
port 41 nsew
rlabel locali s -6113 -58138 -6023 -58049 2 VDD
port 41 nsew
rlabel locali s -6730 -58647 -6696 -58057 2 VDD
port 41 nsew
rlabel locali s -6113 -58049 -6024 -57934 2 VDD
port 41 nsew
rlabel locali s -6736 -58057 -6691 -57934 2 VDD
port 41 nsew
rlabel locali s -6926 -58647 -6892 -58054 2 VDD
port 41 nsew
rlabel locali s -7349 -58647 -7315 -58055 2 VDD
port 41 nsew
rlabel locali s -21534 -58731 -13897 -58564 2 VDD
port 41 nsew
rlabel locali s -27269 -58816 -27203 -58604 2 VDD
port 41 nsew
rlabel locali s -27836 -58816 -27341 -58796 2 VDD
port 41 nsew
rlabel locali s -27389 -58796 -27341 -58604 2 VDD
port 41 nsew
rlabel locali s -27389 -58604 -27203 -58594 2 VDD
port 41 nsew
rlabel locali s -6931 -58054 -6886 -57934 2 VDD
port 41 nsew
rlabel locali s -7353 -58055 -7308 -57934 2 VDD
port 41 nsew
rlabel locali s -9809 -58230 -9775 -57939 2 VDD
port 41 nsew
rlabel locali s -10005 -58230 -9971 -57939 2 VDD
port 41 nsew
rlabel locali s -10201 -58230 -10167 -57939 2 VDD
port 41 nsew
rlabel locali s -10646 -58230 -10612 -57939 2 VDD
port 41 nsew
rlabel locali s -10842 -58230 -10808 -57939 2 VDD
port 41 nsew
rlabel locali s -11038 -58230 -11004 -57939 2 VDD
port 41 nsew
rlabel locali s -12509 -58230 -12475 -57939 2 VDD
port 41 nsew
rlabel locali s -12705 -58230 -12671 -57939 2 VDD
port 41 nsew
rlabel locali s -12901 -58230 -12867 -57939 2 VDD
port 41 nsew
rlabel locali s -13346 -58230 -13312 -57939 2 VDD
port 41 nsew
rlabel locali s -13542 -58230 -13508 -57939 2 VDD
port 41 nsew
rlabel locali s -13738 -58230 -13704 -57939 2 VDD
port 41 nsew
rlabel locali s -13987 -58564 -13898 -57939 2 VDD
port 41 nsew
rlabel locali s -11516 -57939 -9714 -57934 2 VDD
port 41 nsew
rlabel locali s -13987 -57939 -12414 -57934 2 VDD
port 41 nsew
rlabel locali s -13987 -57934 -6024 -57871 2 VDD
port 41 nsew
rlabel locali s -27836 -58594 -27203 -58560 2 VDD
port 41 nsew
rlabel locali s -27389 -58560 -27203 -58545 2 VDD
port 41 nsew
rlabel locali s -27269 -58545 -27203 -58363 2 VDD
port 41 nsew
rlabel locali s -27389 -58545 -27341 -58363 2 VDD
port 41 nsew
rlabel locali s -27389 -58363 -27203 -58358 2 VDD
port 41 nsew
rlabel locali s -27836 -58358 -27203 -58324 2 VDD
port 41 nsew
rlabel locali s -27389 -58324 -27203 -58304 2 VDD
port 41 nsew
rlabel locali s -27269 -58304 -27203 -58131 2 VDD
port 41 nsew
rlabel locali s -27389 -58304 -27341 -58131 2 VDD
port 41 nsew
rlabel locali s -27389 -58131 -27203 -58122 2 VDD
port 41 nsew
rlabel locali s -27836 -58122 -27203 -58088 2 VDD
port 41 nsew
rlabel locali s -27389 -58088 -27203 -58072 2 VDD
port 41 nsew
rlabel locali s -9909 -57871 -6024 -57849 2 VDD
port 41 nsew
rlabel locali s -6113 -57849 -6024 -57210 2 VDD
port 41 nsew
rlabel locali s 18976 -57184 19010 -56600 8 VDD
port 41 nsew
rlabel locali s 18780 -57200 18814 -56600 8 VDD
port 41 nsew
rlabel locali s -6113 -57210 -888 -57147 2 VDD
port 41 nsew
rlabel locali s -3642 -57147 -1840 -57142 2 VDD
port 41 nsew
rlabel locali s -6113 -57147 -4540 -57142 2 VDD
port 41 nsew
rlabel locali s -1935 -57142 -1901 -56851 2 VDD
port 41 nsew
rlabel locali s -2131 -57142 -2097 -56851 2 VDD
port 41 nsew
rlabel locali s -2327 -57142 -2293 -56851 2 VDD
port 41 nsew
rlabel locali s -2772 -57142 -2738 -56851 2 VDD
port 41 nsew
rlabel locali s -2968 -57142 -2934 -56851 2 VDD
port 41 nsew
rlabel locali s -3164 -57142 -3130 -56851 2 VDD
port 41 nsew
rlabel locali s -4635 -57142 -4601 -56851 2 VDD
port 41 nsew
rlabel locali s -4831 -57142 -4797 -56851 2 VDD
port 41 nsew
rlabel locali s -5027 -57142 -4993 -56851 2 VDD
port 41 nsew
rlabel locali s -5472 -57142 -5438 -56851 2 VDD
port 41 nsew
rlabel locali s -5668 -57142 -5634 -56851 2 VDD
port 41 nsew
rlabel locali s -5864 -57142 -5830 -56851 2 VDD
port 41 nsew
rlabel locali s 26110 -56073 30434 -56004 8 VDD
port 41 nsew
rlabel locali s 31402 -56003 33155 -56002 8 VDD
port 41 nsew
rlabel locali s 31402 -56002 34201 -55950 8 VDD
port 41 nsew
rlabel locali s 29321 -56004 29939 -55987 8 VDD
port 41 nsew
rlabel locali s 29321 -55987 29764 -55958 8 VDD
port 41 nsew
rlabel locali s 31769 -55950 34201 -55880 8 VDD
port 41 nsew
rlabel locali s 29322 -55958 29764 -55944 8 VDD
port 41 nsew
rlabel locali s 29322 -55944 30611 -55895 8 VDD
port 41 nsew
rlabel locali s 29724 -55895 30611 -55845 8 VDD
port 41 nsew
rlabel locali s 36751 -55825 37469 -55726 8 VDD
port 41 nsew
rlabel locali s 37387 -55726 37421 -55460 8 VDD
port 41 nsew
rlabel locali s 37191 -55726 37225 -55460 8 VDD
port 41 nsew
rlabel locali s 36995 -55726 37029 -55460 8 VDD
port 41 nsew
rlabel locali s 36799 -55726 36833 -55460 8 VDD
port 41 nsew
rlabel locali s 30529 -55845 30563 -55679 8 VDD
port 41 nsew
rlabel locali s 30333 -55845 30367 -55679 8 VDD
port 41 nsew
rlabel locali s 30137 -55845 30171 -55679 8 VDD
port 41 nsew
rlabel locali s 29941 -55845 29975 -55679 8 VDD
port 41 nsew
rlabel locali s 29724 -55845 29758 -55478 8 VDD
port 41 nsew
rlabel locali s 29528 -55895 29562 -55478 8 VDD
port 41 nsew
rlabel locali s 29332 -55895 29366 -55478 8 VDD
port 41 nsew
rlabel locali s 26110 -56004 28665 -55814 8 VDD
port 41 nsew
rlabel locali s 26110 -55814 29029 -55779 8 VDD
port 41 nsew
rlabel locali s 28311 -55779 29029 -55715 8 VDD
port 41 nsew
rlabel locali s 26110 -55779 26199 -55719 8 VDD
port 41 nsew
rlabel locali s 25916 -56010 25950 -55719 8 VDD
port 41 nsew
rlabel locali s 25720 -56010 25754 -55719 8 VDD
port 41 nsew
rlabel locali s 25524 -56010 25558 -55719 8 VDD
port 41 nsew
rlabel locali s 25079 -56010 25113 -55719 8 VDD
port 41 nsew
rlabel locali s 24883 -56010 24917 -55719 8 VDD
port 41 nsew
rlabel locali s 24687 -56010 24721 -55719 8 VDD
port 41 nsew
rlabel locali s 23216 -56010 23250 -55719 8 VDD
port 41 nsew
rlabel locali s 23020 -56010 23054 -55719 8 VDD
port 41 nsew
rlabel locali s 22824 -56010 22858 -55719 8 VDD
port 41 nsew
rlabel locali s 22379 -56010 22413 -55719 8 VDD
port 41 nsew
rlabel locali s 22183 -56010 22217 -55719 8 VDD
port 41 nsew
rlabel locali s 21987 -56010 22021 -55719 8 VDD
port 41 nsew
rlabel locali s 28947 -55715 28981 -55449 8 VDD
port 41 nsew
rlabel locali s 28751 -55715 28785 -55449 8 VDD
port 41 nsew
rlabel locali s 28555 -55715 28589 -55449 8 VDD
port 41 nsew
rlabel locali s 28359 -55715 28393 -55449 8 VDD
port 41 nsew
rlabel locali s 24626 -55719 26199 -55714 8 VDD
port 41 nsew
rlabel locali s 21926 -55719 23728 -55714 8 VDD
port 41 nsew
rlabel locali s 20974 -55714 26199 -55651 8 VDD
port 41 nsew
rlabel locali s 8753 -55760 8787 -55570 8 VDD
port 41 nsew
rlabel locali s 8557 -55760 8591 -55582 8 VDD
port 41 nsew
rlabel locali s 8748 -55570 8794 -55448 8 VDD
port 41 nsew
rlabel locali s 8551 -55582 8597 -55448 8 VDD
port 41 nsew
rlabel locali s 8444 -55760 8478 -55572 8 VDD
port 41 nsew
rlabel locali s 8248 -55760 8282 -55577 8 VDD
port 41 nsew
rlabel locali s 8438 -55572 8484 -55448 8 VDD
port 41 nsew
rlabel locali s 8242 -55577 8288 -55448 8 VDD
port 41 nsew
rlabel locali s 8134 -55760 8168 -55573 8 VDD
port 41 nsew
rlabel locali s 7938 -55760 7972 -55577 8 VDD
port 41 nsew
rlabel locali s 7742 -55760 7776 -55577 8 VDD
port 41 nsew
rlabel locali s 8129 -55573 8175 -55448 8 VDD
port 41 nsew
rlabel locali s 7931 -55577 7977 -55448 8 VDD
port 41 nsew
rlabel locali s 7742 -55577 7782 -55488 8 VDD
port 41 nsew
rlabel locali s 7741 -55488 7864 -55448 8 VDD
port 41 nsew
rlabel locali s 6581 -55749 6615 -55487 8 VDD
port 41 nsew
rlabel locali s 7741 -55448 8794 -55379 8 VDD
port 41 nsew
rlabel locali s 7741 -55379 7864 -55352 8 VDD
port 41 nsew
rlabel locali s 6525 -55487 6648 -55453 8 VDD
port 41 nsew
rlabel locali s 6385 -55749 6419 -55453 8 VDD
port 41 nsew
rlabel locali s 6189 -55749 6223 -55453 8 VDD
port 41 nsew
rlabel locali s 5993 -55749 6027 -55453 8 VDD
port 41 nsew
rlabel locali s 5451 -55749 5485 -55457 8 VDD
port 41 nsew
rlabel locali s 5255 -55749 5289 -55482 8 VDD
port 41 nsew
rlabel locali s 4828 -55874 4862 -55484 8 VDD
port 41 nsew
rlabel locali s 5169 -55482 5292 -55457 8 VDD
port 41 nsew
rlabel locali s 5993 -55453 6648 -55452 8 VDD
port 41 nsew
rlabel locali s 5169 -55457 5490 -55452 8 VDD
port 41 nsew
rlabel locali s 5169 -55452 6648 -55384 8 VDD
port 41 nsew
rlabel locali s 6525 -55384 6648 -55351 8 VDD
port 41 nsew
rlabel locali s 5169 -55384 6065 -55379 8 VDD
port 41 nsew
rlabel locali s 5169 -55379 5292 -55346 8 VDD
port 41 nsew
rlabel locali s 4768 -55484 4891 -55457 8 VDD
port 41 nsew
rlabel locali s 4632 -55874 4666 -55457 8 VDD
port 41 nsew
rlabel locali s 4436 -55874 4470 -55507 8 VDD
port 41 nsew
rlabel locali s 4219 -55673 4253 -55507 8 VDD
port 41 nsew
rlabel locali s 4023 -55673 4057 -55507 8 VDD
port 41 nsew
rlabel locali s 3827 -55673 3861 -55507 8 VDD
port 41 nsew
rlabel locali s 3631 -55673 3665 -55507 8 VDD
port 41 nsew
rlabel locali s 3223 -55872 3257 -55508 8 VDD
port 41 nsew
rlabel locali s 3540 -55507 4470 -55457 8 VDD
port 41 nsew
rlabel locali s 3540 -55457 4891 -55408 8 VDD
port 41 nsew
rlabel locali s 4430 -55408 4891 -55393 8 VDD
port 41 nsew
rlabel locali s 4768 -55393 4891 -55348 8 VDD
port 41 nsew
rlabel locali s 3540 -55408 3663 -55371 8 VDD
port 41 nsew
rlabel locali s 3151 -55508 3274 -55465 8 VDD
port 41 nsew
rlabel locali s 3027 -55872 3061 -55465 8 VDD
port 41 nsew
rlabel locali s 2831 -55872 2865 -55505 8 VDD
port 41 nsew
rlabel locali s 2614 -55671 2648 -55505 8 VDD
port 41 nsew
rlabel locali s 2418 -55671 2452 -55505 8 VDD
port 41 nsew
rlabel locali s 2222 -55671 2256 -55505 8 VDD
port 41 nsew
rlabel locali s 2026 -55671 2060 -55505 8 VDD
port 41 nsew
rlabel locali s 1978 -55505 2865 -55465 8 VDD
port 41 nsew
rlabel locali s 1619 -55758 1653 -55465 8 VDD
port 41 nsew
rlabel locali s 1423 -55758 1457 -55465 8 VDD
port 41 nsew
rlabel locali s 1227 -55758 1261 -55465 8 VDD
port 41 nsew
rlabel locali s 1031 -55758 1065 -55465 8 VDD
port 41 nsew
rlabel locali s 489 -55758 523 -55466 8 VDD
port 41 nsew
rlabel locali s 293 -55758 327 -55495 8 VDD
port 41 nsew
rlabel locali s -49 -55741 -15 -55496 2 VDD
port 41 nsew
rlabel locali s 173 -55495 327 -55466 8 VDD
port 41 nsew
rlabel locali s 173 -55466 528 -55465 8 VDD
port 41 nsew
rlabel locali s 173 -55465 3274 -55386 8 VDD
port 41 nsew
rlabel locali s 3151 -55386 3274 -55372 8 VDD
port 41 nsew
rlabel locali s 1108 -55386 1223 -54578 8 VDD
port 41 nsew
rlabel locali s 173 -55386 296 -55359 8 VDD
port 41 nsew
rlabel locali s -121 -55496 2 -55450 2 VDD
port 41 nsew
rlabel locali s -245 -55741 -211 -55450 2 VDD
port 41 nsew
rlabel locali s -441 -55741 -407 -55450 2 VDD
port 41 nsew
rlabel locali s -931 -55741 -897 -55450 2 VDD
port 41 nsew
rlabel locali s -1127 -55741 -1093 -55450 2 VDD
port 41 nsew
rlabel locali s -1323 -55741 -1289 -55450 2 VDD
port 41 nsew
rlabel locali s -2674 -55741 -2640 -55450 2 VDD
port 41 nsew
rlabel locali s -2870 -55741 -2836 -55450 2 VDD
port 41 nsew
rlabel locali s -3066 -55741 -3032 -55450 2 VDD
port 41 nsew
rlabel locali s -3631 -55741 -3597 -55450 2 VDD
port 41 nsew
rlabel locali s -3827 -55741 -3793 -55450 2 VDD
port 41 nsew
rlabel locali s -4023 -55741 -3989 -55450 2 VDD
port 41 nsew
rlabel locali s -5374 -55741 -5340 -55450 2 VDD
port 41 nsew
rlabel locali s -5570 -55741 -5536 -55450 2 VDD
port 41 nsew
rlabel locali s -5766 -55741 -5732 -55450 2 VDD
port 41 nsew
rlabel locali s -1384 -55450 2 -55445 2 VDD
port 41 nsew
rlabel locali s -4084 -55450 -2631 -55449 2 VDD
port 41 nsew
rlabel locali s -4084 -55449 -2318 -55445 2 VDD
port 41 nsew
rlabel locali s -5826 -55450 -5331 -55447 2 VDD
port 41 nsew
rlabel locali s -6113 -57142 -6024 -55447 2 VDD
port 41 nsew
rlabel locali s -10517 -56949 -10483 -56783 2 VDD
port 41 nsew
rlabel locali s -10713 -56949 -10679 -56783 2 VDD
port 41 nsew
rlabel locali s -10909 -56949 -10875 -56783 2 VDD
port 41 nsew
rlabel locali s -11105 -56949 -11071 -56783 2 VDD
port 41 nsew
rlabel locali s -11322 -57150 -11288 -56783 2 VDD
port 41 nsew
rlabel locali s -11322 -56783 -10435 -56733 2 VDD
port 41 nsew
rlabel locali s -11518 -57150 -11484 -56733 2 VDD
port 41 nsew
rlabel locali s -11714 -57150 -11680 -56733 2 VDD
port 41 nsew
rlabel locali s -12099 -57179 -12065 -56913 2 VDD
port 41 nsew
rlabel locali s -12295 -57179 -12261 -56913 2 VDD
port 41 nsew
rlabel locali s -12491 -57179 -12457 -56913 2 VDD
port 41 nsew
rlabel locali s -12687 -57179 -12653 -56913 2 VDD
port 41 nsew
rlabel locali s -12735 -56913 -12017 -56814 2 VDD
port 41 nsew
rlabel locali s -11724 -56733 -10435 -56684 2 VDD
port 41 nsew
rlabel locali s -11724 -56684 -11282 -56670 2 VDD
port 41 nsew
rlabel locali s -11725 -56670 -11282 -56641 2 VDD
port 41 nsew
rlabel locali s -11725 -56641 -11107 -56624 2 VDD
port 41 nsew
rlabel locali s -12553 -56814 -12381 -56624 2 VDD
port 41 nsew
rlabel locali s -13525 -57871 -13372 -56624 2 VDD
port 41 nsew
rlabel locali s -13525 -56624 -10612 -56513 2 VDD
port 41 nsew
rlabel locali s -13525 -56513 -10508 -56471 2 VDD
port 41 nsew
rlabel locali s -11277 -56471 -10508 -56447 2 VDD
port 41 nsew
rlabel locali s -12321 -56471 -12095 -56464 2 VDD
port 41 nsew
rlabel locali s -12284 -56464 -12095 -56457 2 VDD
port 41 nsew
rlabel locali s -10654 -56447 -10609 -56323 2 VDD
port 41 nsew
rlabel locali s -11076 -56447 -11031 -56324 2 VDD
port 41 nsew
rlabel locali s -10647 -56323 -10613 -55731 2 VDD
port 41 nsew
rlabel locali s -11070 -56324 -11036 -55731 2 VDD
port 41 nsew
rlabel locali s -11271 -56447 -11226 -56321 2 VDD
port 41 nsew
rlabel locali s -12723 -56423 -12281 -56408 2 VDD
port 41 nsew
rlabel locali s -12723 -56408 -11434 -56359 2 VDD
port 41 nsew
rlabel locali s -11266 -56321 -11232 -55731 2 VDD
port 41 nsew
rlabel locali s -12321 -56359 -11434 -56309 2 VDD
port 41 nsew
rlabel locali s -11516 -56309 -11482 -56143 2 VDD
port 41 nsew
rlabel locali s -11712 -56309 -11678 -56143 2 VDD
port 41 nsew
rlabel locali s -11908 -56309 -11874 -56143 2 VDD
port 41 nsew
rlabel locali s -12104 -56309 -12070 -56143 2 VDD
port 41 nsew
rlabel locali s -12321 -56309 -12287 -55942 2 VDD
port 41 nsew
rlabel locali s -12517 -56359 -12483 -55942 2 VDD
port 41 nsew
rlabel locali s -12713 -56359 -12679 -55942 2 VDD
port 41 nsew
rlabel locali s -6113 -55447 -5009 -55445 2 VDD
port 41 nsew
rlabel locali s -6113 -55445 2 -55382 2 VDD
port 41 nsew
rlabel locali s -121 -55382 2 -55360 2 VDD
port 41 nsew
rlabel locali s -1376 -55382 -1261 -54686 2 VDD
port 41 nsew
rlabel locali s -2791 -55382 -2318 -55381 2 VDD
port 41 nsew
rlabel locali s -3942 -55382 -3827 -54830 2 VDD
port 41 nsew
rlabel locali s -6113 -55382 -5009 -55379 2 VDD
port 41 nsew
rlabel locali s -5235 -55379 -5147 -54989 2 VDD
port 41 nsew
rlabel locali s -5417 -55379 -5329 -54989 2 VDD
port 41 nsew
rlabel locali s -5600 -55379 -5512 -54989 2 VDD
port 41 nsew
rlabel locali s -5616 -54989 -5121 -54921 2 VDD
port 41 nsew
rlabel locali s -3947 -54830 -3824 -54694 2 VDD
port 41 nsew
rlabel locali s 1103 -54578 1409 -54516 8 VDD
port 41 nsew
rlabel locali s -1380 -54686 -1257 -54550 2 VDD
port 41 nsew
rlabel locali s -5215 -54921 -5181 -54630 2 VDD
port 41 nsew
rlabel locali s -5411 -54921 -5377 -54630 2 VDD
port 41 nsew
rlabel locali s -5607 -54921 -5573 -54630 2 VDD
port 41 nsew
rlabel locali s -13525 -56471 -13372 -54775 2 VDD
port 41 nsew
rlabel locali s -27269 -58072 -27203 -57525 2 VDD
port 41 nsew
rlabel locali s -27389 -58072 -27341 -57992 2 VDD
port 41 nsew
rlabel locali s -27836 -57992 -27341 -57958 2 VDD
port 41 nsew
rlabel locali s -27389 -57958 -27341 -57756 2 VDD
port 41 nsew
rlabel locali s -27836 -57756 -27341 -57722 2 VDD
port 41 nsew
rlabel locali s -27389 -57722 -27341 -57525 2 VDD
port 41 nsew
rlabel locali s -27389 -57525 -27203 -57520 2 VDD
port 41 nsew
rlabel locali s -27836 -57520 -27203 -57486 2 VDD
port 41 nsew
rlabel locali s -27389 -57486 -27203 -57466 2 VDD
port 41 nsew
rlabel locali s -27269 -57466 -27203 -57296 2 VDD
port 41 nsew
rlabel locali s -27389 -57466 -27341 -57296 2 VDD
port 41 nsew
rlabel locali s -27389 -57296 -27203 -57284 2 VDD
port 41 nsew
rlabel locali s -27836 -57284 -27203 -57250 2 VDD
port 41 nsew
rlabel locali s -27389 -57250 -27203 -57237 2 VDD
port 41 nsew
rlabel locali s -27269 -57237 -27203 -57057 2 VDD
port 41 nsew
rlabel locali s -27389 -57237 -27341 -57057 2 VDD
port 41 nsew
rlabel locali s -27389 -57057 -27203 -57048 2 VDD
port 41 nsew
rlabel locali s -27836 -57048 -27203 -57014 2 VDD
port 41 nsew
rlabel locali s -27389 -57014 -27203 -56998 2 VDD
port 41 nsew
rlabel locali s -27269 -56998 -27203 -56822 2 VDD
port 41 nsew
rlabel locali s -27389 -56998 -27341 -56822 2 VDD
port 41 nsew
rlabel locali s -27389 -56822 -27203 -56812 2 VDD
port 41 nsew
rlabel locali s -27836 -56812 -27203 -56778 2 VDD
port 41 nsew
rlabel locali s -27389 -56778 -27203 -56763 2 VDD
port 41 nsew
rlabel locali s -27269 -56763 -27203 -56586 2 VDD
port 41 nsew
rlabel locali s -27389 -56763 -27341 -56586 2 VDD
port 41 nsew
rlabel locali s -27389 -56586 -27203 -56576 2 VDD
port 41 nsew
rlabel locali s -27836 -56576 -27203 -56542 2 VDD
port 41 nsew
rlabel locali s -27389 -56542 -27203 -56527 2 VDD
port 41 nsew
rlabel locali s -27269 -56527 -27203 -56355 2 VDD
port 41 nsew
rlabel locali s -27389 -56527 -27341 -56355 2 VDD
port 41 nsew
rlabel locali s -27389 -56355 -27203 -56340 2 VDD
port 41 nsew
rlabel locali s -27836 -56340 -27203 -56306 2 VDD
port 41 nsew
rlabel locali s -27389 -56306 -27203 -56296 2 VDD
port 41 nsew
rlabel locali s -15506 -55973 -15472 -55807 2 VDD
port 41 nsew
rlabel locali s -15702 -55973 -15668 -55807 2 VDD
port 41 nsew
rlabel locali s -15898 -55973 -15864 -55807 2 VDD
port 41 nsew
rlabel locali s -16094 -55973 -16060 -55807 2 VDD
port 41 nsew
rlabel locali s -16311 -56174 -16277 -55807 2 VDD
port 41 nsew
rlabel locali s -16311 -55807 -15424 -55757 2 VDD
port 41 nsew
rlabel locali s -16507 -56174 -16473 -55757 2 VDD
port 41 nsew
rlabel locali s -16703 -56174 -16669 -55757 2 VDD
port 41 nsew
rlabel locali s -17088 -56203 -17054 -55937 2 VDD
port 41 nsew
rlabel locali s -17284 -56203 -17250 -55937 2 VDD
port 41 nsew
rlabel locali s -17480 -56203 -17446 -55937 2 VDD
port 41 nsew
rlabel locali s -17676 -56203 -17642 -55937 2 VDD
port 41 nsew
rlabel locali s -17724 -55937 -17006 -55838 2 VDD
port 41 nsew
rlabel locali s -16713 -55757 -15424 -55708 2 VDD
port 41 nsew
rlabel locali s -16713 -55708 -16271 -55694 2 VDD
port 41 nsew
rlabel locali s -16714 -55694 -16271 -55665 2 VDD
port 41 nsew
rlabel locali s -16714 -55665 -16096 -55648 2 VDD
port 41 nsew
rlabel locali s -17542 -55838 -17370 -55648 2 VDD
port 41 nsew
rlabel locali s -18181 -56026 -18147 -55767 2 VDD
port 41 nsew
rlabel locali s -18377 -56026 -18343 -55767 2 VDD
port 41 nsew
rlabel locali s -18919 -56026 -18885 -55767 2 VDD
port 41 nsew
rlabel locali s -19115 -56026 -19081 -55767 2 VDD
port 41 nsew
rlabel locali s -19311 -56026 -19277 -55767 2 VDD
port 41 nsew
rlabel locali s -19507 -56026 -19473 -55767 2 VDD
port 41 nsew
rlabel locali s -20083 -56020 -20049 -55854 2 VDD
port 41 nsew
rlabel locali s -20279 -56020 -20245 -55854 2 VDD
port 41 nsew
rlabel locali s -20475 -56020 -20441 -55854 2 VDD
port 41 nsew
rlabel locali s -20671 -56020 -20637 -55854 2 VDD
port 41 nsew
rlabel locali s -20888 -56221 -20854 -55854 2 VDD
port 41 nsew
rlabel locali s -20888 -55854 -20001 -55804 2 VDD
port 41 nsew
rlabel locali s -21084 -56221 -21050 -55804 2 VDD
port 41 nsew
rlabel locali s -21280 -56221 -21246 -55804 2 VDD
port 41 nsew
rlabel locali s -21290 -55804 -20001 -55767 2 VDD
port 41 nsew
rlabel locali s -22950 -55767 -18147 -55734 2 VDD
port 41 nsew
rlabel locali s -22950 -55734 -18137 -55648 2 VDD
port 41 nsew
rlabel locali s -22950 -55648 -15601 -55600 2 VDD
port 41 nsew
rlabel locali s -27269 -56296 -27203 -55630 2 VDD
port 41 nsew
rlabel locali s -27389 -56296 -27341 -56104 2 VDD
port 41 nsew
rlabel locali s -27836 -56104 -27341 -56070 2 VDD
port 41 nsew
rlabel locali s -27389 -56070 -27341 -55856 2 VDD
port 41 nsew
rlabel locali s -27836 -55856 -27341 -55822 2 VDD
port 41 nsew
rlabel locali s -27389 -55822 -27341 -55630 2 VDD
port 41 nsew
rlabel locali s -27389 -55630 -27203 -55620 2 VDD
port 41 nsew
rlabel locali s -27836 -55620 -27203 -55600 2 VDD
port 41 nsew
rlabel locali s -27836 -55600 -15601 -55586 2 VDD
port 41 nsew
rlabel locali s -27389 -55586 -15601 -55571 2 VDD
port 41 nsew
rlabel locali s -27269 -55571 -15601 -55537 2 VDD
port 41 nsew
rlabel locali s -27269 -55537 -15497 -55535 2 VDD
port 41 nsew
rlabel locali s -17712 -55535 -15497 -55495 2 VDD
port 41 nsew
rlabel locali s -16266 -55495 -15497 -55471 2 VDD
port 41 nsew
rlabel locali s -17310 -55495 -17084 -55488 2 VDD
port 41 nsew
rlabel locali s -17273 -55488 -17084 -55481 2 VDD
port 41 nsew
rlabel locali s -15643 -55471 -15598 -55347 2 VDD
port 41 nsew
rlabel locali s -16065 -55471 -16020 -55348 2 VDD
port 41 nsew
rlabel locali s -10665 -54773 -10192 -54772 2 VDD
port 41 nsew
rlabel locali s -13987 -54775 -12883 -54772 2 VDD
port 41 nsew
rlabel locali s -13987 -54772 -7880 -54709 2 VDD
port 41 nsew
rlabel locali s -15636 -55347 -15602 -54755 2 VDD
port 41 nsew
rlabel locali s -16059 -55348 -16025 -54755 2 VDD
port 41 nsew
rlabel locali s -16260 -55471 -16215 -55345 2 VDD
port 41 nsew
rlabel locali s -17712 -55447 -17270 -55432 2 VDD
port 41 nsew
rlabel locali s -17712 -55432 -16423 -55383 2 VDD
port 41 nsew
rlabel locali s -27269 -55535 -22678 -55396 2 VDD
port 41 nsew
rlabel locali s -27389 -55571 -27341 -55396 2 VDD
port 41 nsew
rlabel locali s -27389 -55396 -22678 -55384 2 VDD
port 41 nsew
rlabel locali s -16255 -55345 -16221 -54755 2 VDD
port 41 nsew
rlabel locali s -17310 -55383 -16423 -55333 2 VDD
port 41 nsew
rlabel locali s -16505 -55333 -16471 -55167 2 VDD
port 41 nsew
rlabel locali s -16701 -55333 -16667 -55167 2 VDD
port 41 nsew
rlabel locali s -16897 -55333 -16863 -55167 2 VDD
port 41 nsew
rlabel locali s -17093 -55333 -17059 -55167 2 VDD
port 41 nsew
rlabel locali s -17310 -55333 -17276 -54966 2 VDD
port 41 nsew
rlabel locali s -17506 -55383 -17472 -54966 2 VDD
port 41 nsew
rlabel locali s -17702 -55383 -17668 -54966 2 VDD
port 41 nsew
rlabel locali s -27836 -55384 -22678 -55350 2 VDD
port 41 nsew
rlabel locali s -27389 -55350 -22678 -55337 2 VDD
port 41 nsew
rlabel locali s -27269 -55337 -22678 -55328 2 VDD
port 41 nsew
rlabel locali s -22950 -55328 -22678 -54866 2 VDD
port 41 nsew
rlabel locali s -27269 -55328 -27203 -55162 2 VDD
port 41 nsew
rlabel locali s -27389 -55337 -27341 -55162 2 VDD
port 41 nsew
rlabel locali s -27389 -55162 -27203 -55148 2 VDD
port 41 nsew
rlabel locali s -27836 -55148 -27203 -55114 2 VDD
port 41 nsew
rlabel locali s -27389 -55114 -27203 -55103 2 VDD
port 41 nsew
rlabel locali s -27269 -55103 -27203 -54925 2 VDD
port 41 nsew
rlabel locali s -27389 -55103 -27341 -54925 2 VDD
port 41 nsew
rlabel locali s -27389 -54925 -27203 -54912 2 VDD
port 41 nsew
rlabel locali s -27836 -54912 -27203 -54878 2 VDD
port 41 nsew
rlabel locali s -27389 -54878 -27203 -54866 2 VDD
port 41 nsew
rlabel locali s -9258 -54709 -7880 -54704 2 VDD
port 41 nsew
rlabel locali s -11958 -54709 -10192 -54705 2 VDD
port 41 nsew
rlabel locali s -13987 -54709 -12883 -54707 2 VDD
port 41 nsew
rlabel locali s -11958 -54705 -10505 -54704 2 VDD
port 41 nsew
rlabel locali s -13700 -54707 -13205 -54704 2 VDD
port 41 nsew
rlabel locali s 1103 -54516 1226 -54515 8 VDD
port 41 nsew
rlabel locali s -7923 -54704 -7889 -54413 2 VDD
port 41 nsew
rlabel locali s -8119 -54704 -8085 -54413 2 VDD
port 41 nsew
rlabel locali s -8315 -54704 -8281 -54413 2 VDD
port 41 nsew
rlabel locali s -8805 -54704 -8771 -54413 2 VDD
port 41 nsew
rlabel locali s -9001 -54704 -8967 -54413 2 VDD
port 41 nsew
rlabel locali s -9197 -54704 -9163 -54413 2 VDD
port 41 nsew
rlabel locali s -10548 -54704 -10514 -54413 2 VDD
port 41 nsew
rlabel locali s -10744 -54704 -10710 -54413 2 VDD
port 41 nsew
rlabel locali s -10940 -54704 -10906 -54413 2 VDD
port 41 nsew
rlabel locali s -11505 -54704 -11471 -54413 2 VDD
port 41 nsew
rlabel locali s -11701 -54704 -11667 -54413 2 VDD
port 41 nsew
rlabel locali s -11897 -54704 -11863 -54413 2 VDD
port 41 nsew
rlabel locali s -13248 -54704 -13214 -54413 2 VDD
port 41 nsew
rlabel locali s -13444 -54704 -13410 -54413 2 VDD
port 41 nsew
rlabel locali s -13640 -54704 -13606 -54413 2 VDD
port 41 nsew
rlabel locali s 1104 -54098 1227 -53962 8 VDD
port 41 nsew
rlabel locali s -1379 -54098 -1256 -53962 2 VDD
port 41 nsew
rlabel locali s 8743 -53509 8777 -53319 8 VDD
port 41 nsew
rlabel locali s 8547 -53509 8581 -53331 8 VDD
port 41 nsew
rlabel locali s 26626 -53252 27729 -51863 8 VDD
port 41 nsew
rlabel locali s 8738 -53319 8784 -53197 8 VDD
port 41 nsew
rlabel locali s 8541 -53331 8587 -53197 8 VDD
port 41 nsew
rlabel locali s 8434 -53509 8468 -53321 8 VDD
port 41 nsew
rlabel locali s 8238 -53509 8272 -53326 8 VDD
port 41 nsew
rlabel locali s 8428 -53321 8474 -53197 8 VDD
port 41 nsew
rlabel locali s 8232 -53326 8278 -53197 8 VDD
port 41 nsew
rlabel locali s 8124 -53509 8158 -53322 8 VDD
port 41 nsew
rlabel locali s 7928 -53509 7962 -53326 8 VDD
port 41 nsew
rlabel locali s 7732 -53509 7766 -53326 8 VDD
port 41 nsew
rlabel locali s 8119 -53322 8165 -53197 8 VDD
port 41 nsew
rlabel locali s 7921 -53326 7967 -53197 8 VDD
port 41 nsew
rlabel locali s 7732 -53326 7772 -53197 8 VDD
port 41 nsew
rlabel locali s 5743 -53509 5777 -53319 8 VDD
port 41 nsew
rlabel locali s 5547 -53509 5581 -53331 8 VDD
port 41 nsew
rlabel locali s 7732 -53197 8784 -53090 8 VDD
port 41 nsew
rlabel locali s 5738 -53319 5784 -53197 8 VDD
port 41 nsew
rlabel locali s 5541 -53331 5587 -53197 8 VDD
port 41 nsew
rlabel locali s 5434 -53509 5468 -53321 8 VDD
port 41 nsew
rlabel locali s 5238 -53509 5272 -53326 8 VDD
port 41 nsew
rlabel locali s 5428 -53321 5474 -53197 8 VDD
port 41 nsew
rlabel locali s 5232 -53326 5278 -53197 8 VDD
port 41 nsew
rlabel locali s 5124 -53509 5158 -53322 8 VDD
port 41 nsew
rlabel locali s 4928 -53509 4962 -53326 8 VDD
port 41 nsew
rlabel locali s 4732 -53509 4766 -53326 8 VDD
port 41 nsew
rlabel locali s 5119 -53322 5165 -53197 8 VDD
port 41 nsew
rlabel locali s 4921 -53326 4967 -53197 8 VDD
port 41 nsew
rlabel locali s 4732 -53326 4772 -53197 8 VDD
port 41 nsew
rlabel locali s 3243 -53509 3277 -53319 8 VDD
port 41 nsew
rlabel locali s 3047 -53509 3081 -53331 8 VDD
port 41 nsew
rlabel locali s 4732 -53197 5784 -53128 8 VDD
port 41 nsew
rlabel locali s 3238 -53319 3284 -53197 8 VDD
port 41 nsew
rlabel locali s 3041 -53331 3087 -53197 8 VDD
port 41 nsew
rlabel locali s 2934 -53509 2968 -53321 8 VDD
port 41 nsew
rlabel locali s 2738 -53509 2772 -53326 8 VDD
port 41 nsew
rlabel locali s 2928 -53321 2974 -53197 8 VDD
port 41 nsew
rlabel locali s 2732 -53326 2778 -53197 8 VDD
port 41 nsew
rlabel locali s 2624 -53509 2658 -53322 8 VDD
port 41 nsew
rlabel locali s 2428 -53509 2462 -53326 8 VDD
port 41 nsew
rlabel locali s 2232 -53509 2266 -53326 8 VDD
port 41 nsew
rlabel locali s 2619 -53322 2665 -53197 8 VDD
port 41 nsew
rlabel locali s 2421 -53326 2467 -53197 8 VDD
port 41 nsew
rlabel locali s 2232 -53326 2272 -53197 8 VDD
port 41 nsew
rlabel locali s 2232 -53197 3284 -53128 8 VDD
port 41 nsew
rlabel locali s 5009 -53128 5602 -53090 8 VDD
port 41 nsew
rlabel locali s 2596 -53128 3189 -53090 8 VDD
port 41 nsew
rlabel locali s 1109 -53962 1224 -53090 8 VDD
port 41 nsew
rlabel locali s 743 -53509 777 -53319 8 VDD
port 41 nsew
rlabel locali s 547 -53509 581 -53331 8 VDD
port 41 nsew
rlabel locali s 738 -53319 784 -53197 8 VDD
port 41 nsew
rlabel locali s 541 -53331 587 -53197 8 VDD
port 41 nsew
rlabel locali s 434 -53509 468 -53321 8 VDD
port 41 nsew
rlabel locali s 238 -53509 272 -53326 8 VDD
port 41 nsew
rlabel locali s 428 -53321 474 -53197 8 VDD
port 41 nsew
rlabel locali s 232 -53326 278 -53197 8 VDD
port 41 nsew
rlabel locali s 124 -53509 158 -53322 8 VDD
port 41 nsew
rlabel locali s -72 -53509 -38 -53326 2 VDD
port 41 nsew
rlabel locali s -268 -53509 -234 -53326 2 VDD
port 41 nsew
rlabel locali s 119 -53322 165 -53197 8 VDD
port 41 nsew
rlabel locali s -79 -53326 -33 -53197 2 VDD
port 41 nsew
rlabel locali s -268 -53326 -228 -53197 2 VDD
port 41 nsew
rlabel locali s -268 -53197 784 -53128 8 VDD
port 41 nsew
rlabel locali s 62 -53128 655 -53090 8 VDD
port 41 nsew
rlabel locali s -1373 -53962 -1259 -53090 2 VDD
port 41 nsew
rlabel locali s -3946 -54063 -3823 -53927 2 VDD
port 41 nsew
rlabel locali s -1757 -53509 -1723 -53319 2 VDD
port 41 nsew
rlabel locali s -1953 -53509 -1919 -53331 2 VDD
port 41 nsew
rlabel locali s -1762 -53319 -1716 -53197 2 VDD
port 41 nsew
rlabel locali s -1959 -53331 -1913 -53197 2 VDD
port 41 nsew
rlabel locali s -2066 -53509 -2032 -53321 2 VDD
port 41 nsew
rlabel locali s -2262 -53509 -2228 -53326 2 VDD
port 41 nsew
rlabel locali s -2072 -53321 -2026 -53197 2 VDD
port 41 nsew
rlabel locali s -2268 -53326 -2222 -53197 2 VDD
port 41 nsew
rlabel locali s -2376 -53509 -2342 -53322 2 VDD
port 41 nsew
rlabel locali s -2572 -53509 -2538 -53326 2 VDD
port 41 nsew
rlabel locali s -2768 -53509 -2734 -53326 2 VDD
port 41 nsew
rlabel locali s -2381 -53322 -2335 -53197 2 VDD
port 41 nsew
rlabel locali s -2579 -53326 -2533 -53197 2 VDD
port 41 nsew
rlabel locali s -2768 -53326 -2728 -53197 2 VDD
port 41 nsew
rlabel locali s -2768 -53197 -1716 -53128 2 VDD
port 41 nsew
rlabel locali s -2454 -53128 -1861 -53090 2 VDD
port 41 nsew
rlabel locali s -3941 -53927 -3826 -53090 2 VDD
port 41 nsew
rlabel locali s -13987 -54707 -13898 -53784 2 VDD
port 41 nsew
rlabel locali s -27269 -54866 -22678 -54695 2 VDD
port 41 nsew
rlabel locali s -27389 -54866 -27341 -54695 2 VDD
port 41 nsew
rlabel locali s -27389 -54695 -22678 -54676 2 VDD
port 41 nsew
rlabel locali s -27836 -54676 -22678 -54642 2 VDD
port 41 nsew
rlabel locali s -27389 -54642 -22678 -54636 2 VDD
port 41 nsew
rlabel locali s -27269 -54636 -22678 -54594 2 VDD
port 41 nsew
rlabel locali s -18141 -54111 -18107 -53945 2 VDD
port 41 nsew
rlabel locali s -18337 -54111 -18303 -53945 2 VDD
port 41 nsew
rlabel locali s -18533 -54111 -18499 -53945 2 VDD
port 41 nsew
rlabel locali s -18729 -54111 -18695 -53945 2 VDD
port 41 nsew
rlabel locali s -18946 -54312 -18912 -53945 2 VDD
port 41 nsew
rlabel locali s -18946 -53945 -18059 -53901 2 VDD
port 41 nsew
rlabel locali s -19142 -54312 -19108 -53901 2 VDD
port 41 nsew
rlabel locali s -19338 -54312 -19304 -53901 2 VDD
port 41 nsew
rlabel locali s -19390 -53901 -18059 -53846 2 VDD
port 41 nsew
rlabel locali s -19390 -53846 -18063 -53784 2 VDD
port 41 nsew
rlabel locali s -20011 -54090 -19977 -53798 2 VDD
port 41 nsew
rlabel locali s -20207 -54090 -20173 -53798 2 VDD
port 41 nsew
rlabel locali s -20212 -53798 -19967 -53784 2 VDD
port 41 nsew
rlabel locali s -20749 -54090 -20715 -53794 2 VDD
port 41 nsew
rlabel locali s -20945 -54090 -20911 -53794 2 VDD
port 41 nsew
rlabel locali s -21141 -54090 -21107 -53794 2 VDD
port 41 nsew
rlabel locali s -21337 -54090 -21303 -53794 2 VDD
port 41 nsew
rlabel locali s -22950 -54594 -22678 -54080 2 VDD
port 41 nsew
rlabel locali s -27269 -54594 -27203 -54455 2 VDD
port 41 nsew
rlabel locali s -27389 -54636 -27341 -54455 2 VDD
port 41 nsew
rlabel locali s -27389 -54455 -27203 -54440 2 VDD
port 41 nsew
rlabel locali s -27836 -54440 -27203 -54406 2 VDD
port 41 nsew
rlabel locali s -27389 -54406 -27203 -54396 2 VDD
port 41 nsew
rlabel locali s -27269 -54396 -27203 -54217 2 VDD
port 41 nsew
rlabel locali s -27389 -54396 -27341 -54217 2 VDD
port 41 nsew
rlabel locali s -27389 -54217 -27203 -54204 2 VDD
port 41 nsew
rlabel locali s -27836 -54204 -27203 -54170 2 VDD
port 41 nsew
rlabel locali s -27389 -54170 -27203 -54158 2 VDD
port 41 nsew
rlabel locali s -27269 -54158 -27203 -54080 2 VDD
port 41 nsew
rlabel locali s -27269 -54080 -22678 -53981 2 VDD
port 41 nsew
rlabel locali s -27389 -54158 -27341 -53981 2 VDD
port 41 nsew
rlabel locali s -27389 -53981 -22678 -53968 2 VDD
port 41 nsew
rlabel locali s -27836 -53968 -22678 -53934 2 VDD
port 41 nsew
rlabel locali s -27389 -53934 -22678 -53922 2 VDD
port 41 nsew
rlabel locali s -27269 -53922 -22678 -53808 2 VDD
port 41 nsew
rlabel locali s -22950 -53808 -22678 -53794 2 VDD
port 41 nsew
rlabel locali s -22950 -53794 -20715 -53784 2 VDD
port 41 nsew
rlabel locali s -4257 -53509 -4223 -53319 2 VDD
port 41 nsew
rlabel locali s -4453 -53509 -4419 -53331 2 VDD
port 41 nsew
rlabel locali s -4262 -53319 -4216 -53197 2 VDD
port 41 nsew
rlabel locali s -4459 -53331 -4413 -53197 2 VDD
port 41 nsew
rlabel locali s -4566 -53509 -4532 -53321 2 VDD
port 41 nsew
rlabel locali s -4762 -53509 -4728 -53326 2 VDD
port 41 nsew
rlabel locali s -4572 -53321 -4526 -53197 2 VDD
port 41 nsew
rlabel locali s -4768 -53326 -4722 -53197 2 VDD
port 41 nsew
rlabel locali s -4876 -53509 -4842 -53322 2 VDD
port 41 nsew
rlabel locali s -5072 -53509 -5038 -53326 2 VDD
port 41 nsew
rlabel locali s -5268 -53509 -5234 -53326 2 VDD
port 41 nsew
rlabel locali s -4881 -53322 -4835 -53197 2 VDD
port 41 nsew
rlabel locali s -5079 -53326 -5033 -53197 2 VDD
port 41 nsew
rlabel locali s -5268 -53326 -5228 -53197 2 VDD
port 41 nsew
rlabel locali s -5268 -53197 -4216 -53090 2 VDD
port 41 nsew
rlabel locali s -6757 -53713 -6723 -53123 2 VDD
port 41 nsew
rlabel locali s -6633 -53090 8829 -52997 8 VDD
port 41 nsew
rlabel locali s -6763 -53123 -6718 -52997 2 VDD
port 41 nsew
rlabel locali s -6953 -53713 -6919 -53120 2 VDD
port 41 nsew
rlabel locali s -7376 -53713 -7342 -53121 2 VDD
port 41 nsew
rlabel locali s -22950 -53784 -13898 -53571 2 VDD
port 41 nsew
rlabel locali s -27269 -53808 -27203 -53750 2 VDD
port 41 nsew
rlabel locali s -27389 -53922 -27341 -53750 2 VDD
port 41 nsew
rlabel locali s -27389 -53750 -27203 -53732 2 VDD
port 41 nsew
rlabel locali s -27836 -53732 -27203 -53698 2 VDD
port 41 nsew
rlabel locali s -27389 -53698 -27203 -53691 2 VDD
port 41 nsew
rlabel locali s -6958 -53120 -6913 -52997 2 VDD
port 41 nsew
rlabel locali s -7380 -53121 -7335 -52997 2 VDD
port 41 nsew
rlabel locali s -9809 -53303 -9775 -53012 2 VDD
port 41 nsew
rlabel locali s -10005 -53303 -9971 -53012 2 VDD
port 41 nsew
rlabel locali s -10201 -53303 -10167 -53012 2 VDD
port 41 nsew
rlabel locali s -10646 -53303 -10612 -53012 2 VDD
port 41 nsew
rlabel locali s -10842 -53303 -10808 -53012 2 VDD
port 41 nsew
rlabel locali s -11038 -53303 -11004 -53012 2 VDD
port 41 nsew
rlabel locali s -12509 -53303 -12475 -53012 2 VDD
port 41 nsew
rlabel locali s -12705 -53303 -12671 -53012 2 VDD
port 41 nsew
rlabel locali s -12901 -53303 -12867 -53012 2 VDD
port 41 nsew
rlabel locali s -13346 -53303 -13312 -53012 2 VDD
port 41 nsew
rlabel locali s -13542 -53303 -13508 -53012 2 VDD
port 41 nsew
rlabel locali s -13738 -53303 -13704 -53012 2 VDD
port 41 nsew
rlabel locali s -13987 -53571 -13898 -53012 2 VDD
port 41 nsew
rlabel locali s -11516 -53012 -9714 -53007 2 VDD
port 41 nsew
rlabel locali s -13987 -53012 -12414 -53007 2 VDD
port 41 nsew
rlabel locali s -13987 -53007 -8762 -52997 2 VDD
port 41 nsew
rlabel locali s -13987 -52997 8829 -52944 2 VDD
port 41 nsew
rlabel locali s -27269 -53691 -27203 -53273 2 VDD
port 41 nsew
rlabel locali s -27389 -53691 -27341 -53496 2 VDD
port 41 nsew
rlabel locali s -27836 -53496 -27341 -53462 2 VDD
port 41 nsew
rlabel locali s -27389 -53462 -27341 -53273 2 VDD
port 41 nsew
rlabel locali s -27389 -53273 -27203 -53260 2 VDD
port 41 nsew
rlabel locali s -27836 -53260 -27203 -53226 2 VDD
port 41 nsew
rlabel locali s -27389 -53226 -27203 -53214 2 VDD
port 41 nsew
rlabel locali s -8962 -52944 8829 -52908 2 VDD
port 41 nsew
rlabel locali s -6631 -52908 8829 -52897 8 VDD
port 41 nsew
rlabel locali s 26626 -51863 87774 -51743 8 VDD
port 41 nsew
rlabel locali s 7598 -52897 8360 -51743 8 VDD
port 41 nsew
rlabel locali s -27269 -53214 -27203 -52226 2 VDD
port 41 nsew
rlabel locali s -27389 -53214 -27341 -53024 2 VDD
port 41 nsew
rlabel locali s -27836 -53024 -27341 -52990 2 VDD
port 41 nsew
rlabel locali s -27389 -52990 -27341 -52788 2 VDD
port 41 nsew
rlabel locali s -27836 -52788 -27341 -52754 2 VDD
port 41 nsew
rlabel locali s -27389 -52754 -27341 -52552 2 VDD
port 41 nsew
rlabel locali s -27836 -52552 -27341 -52518 2 VDD
port 41 nsew
rlabel locali s -27389 -52518 -27341 -52316 2 VDD
port 41 nsew
rlabel locali s -27836 -52316 -27341 -52282 2 VDD
port 41 nsew
rlabel locali s -27389 -52282 -27341 -52116 2 VDD
port 41 nsew
rlabel locali s 7598 -51743 87774 -50981 8 VDD
port 41 nsew
rlabel locali s 26626 -50981 87774 -50760 8 VDD
port 41 nsew
rlabel locali s 83333 -50760 86302 -49082 8 VDD
port 41 nsew
rlabel locali s 83333 -49082 98798 -46113 8 VDD
port 41 nsew
rlabel locali s 95829 -46113 98798 -31308 8 VDD
port 41 nsew
rlabel locali s -6836 -44340 8126 -44147 8 VDD
port 41 nsew
rlabel locali s -22077 -44182 -19475 -44173 2 VDD
port 41 nsew
rlabel locali s 7029 -44147 8081 -44040 8 VDD
port 41 nsew
rlabel locali s 4306 -44147 4899 -44109 8 VDD
port 41 nsew
rlabel locali s 1893 -44147 2486 -44109 8 VDD
port 41 nsew
rlabel locali s 12143 -43924 17368 -43861 8 VDD
port 41 nsew
rlabel locali s 8035 -44040 8081 -43918 8 VDD
port 41 nsew
rlabel locali s 15795 -43861 17368 -43856 8 VDD
port 41 nsew
rlabel locali s 13095 -43861 14897 -43856 8 VDD
port 41 nsew
rlabel locali s 87128 -42165 87162 -41573 8 VDD
port 41 nsew
rlabel locali s 87568 -41468 87707 -41440 8 VDD
port 41 nsew
rlabel locali s 87568 -41440 87780 -41301 8 VDD
port 41 nsew
rlabel locali s 87318 -41455 87397 -41430 8 VDD
port 41 nsew
rlabel locali s 87121 -41573 87166 -41449 8 VDD
port 41 nsew
rlabel locali s 86705 -42165 86739 -41572 8 VDD
port 41 nsew
rlabel locali s 86509 -42165 86543 -41575 8 VDD
port 41 nsew
rlabel locali s 86259 -41753 86293 -41587 8 VDD
port 41 nsew
rlabel locali s 86063 -41753 86097 -41587 8 VDD
port 41 nsew
rlabel locali s 85867 -41753 85901 -41587 8 VDD
port 41 nsew
rlabel locali s 85671 -41753 85705 -41587 8 VDD
port 41 nsew
rlabel locali s 85454 -41954 85488 -41587 8 VDD
port 41 nsew
rlabel locali s 86699 -41572 86744 -41449 8 VDD
port 41 nsew
rlabel locali s 86504 -41575 86549 -41449 8 VDD
port 41 nsew
rlabel locali s 85454 -41587 86341 -41537 8 VDD
port 41 nsew
rlabel locali s 85258 -41954 85292 -41537 8 VDD
port 41 nsew
rlabel locali s 85062 -41954 85096 -41537 8 VDD
port 41 nsew
rlabel locali s 83460 -42134 83494 -41542 8 VDD
port 41 nsew
rlabel locali s 85052 -41537 86341 -41488 8 VDD
port 41 nsew
rlabel locali s 85052 -41488 85494 -41473 8 VDD
port 41 nsew
rlabel locali s 86498 -41449 87267 -41430 8 VDD
port 41 nsew
rlabel locali s 86498 -41430 87397 -41425 8 VDD
port 41 nsew
rlabel locali s 85491 -41439 85680 -41432 8 VDD
port 41 nsew
rlabel locali s 85454 -41432 85680 -41425 8 VDD
port 41 nsew
rlabel locali s 85052 -41425 87397 -41383 8 VDD
port 41 nsew
rlabel locali s 83453 -41542 83498 -41418 8 VDD
port 41 nsew
rlabel locali s 83037 -42134 83071 -41541 8 VDD
port 41 nsew
rlabel locali s 82841 -42134 82875 -41544 8 VDD
port 41 nsew
rlabel locali s 82591 -41722 82625 -41556 8 VDD
port 41 nsew
rlabel locali s 82395 -41722 82429 -41556 8 VDD
port 41 nsew
rlabel locali s 82199 -41722 82233 -41556 8 VDD
port 41 nsew
rlabel locali s 82003 -41722 82037 -41556 8 VDD
port 41 nsew
rlabel locali s 81786 -41923 81820 -41556 8 VDD
port 41 nsew
rlabel locali s 83031 -41541 83076 -41418 8 VDD
port 41 nsew
rlabel locali s 82836 -41544 82881 -41418 8 VDD
port 41 nsew
rlabel locali s 81786 -41556 82673 -41506 8 VDD
port 41 nsew
rlabel locali s 81590 -41923 81624 -41506 8 VDD
port 41 nsew
rlabel locali s 81394 -41923 81428 -41506 8 VDD
port 41 nsew
rlabel locali s 77764 -42203 77798 -41611 8 VDD
port 41 nsew
rlabel locali s 81384 -41506 82673 -41457 8 VDD
port 41 nsew
rlabel locali s 78204 -41506 78343 -41478 8 VDD
port 41 nsew
rlabel locali s 81384 -41457 81826 -41442 8 VDD
port 41 nsew
rlabel locali s 82830 -41418 83599 -41394 8 VDD
port 41 nsew
rlabel locali s 81823 -41408 82012 -41401 8 VDD
port 41 nsew
rlabel locali s 81786 -41401 82012 -41394 8 VDD
port 41 nsew
rlabel locali s 87218 -41383 87397 -41347 8 VDD
port 41 nsew
rlabel locali s 85052 -41383 87163 -41372 8 VDD
port 41 nsew
rlabel locali s 87318 -41347 87397 -41316 8 VDD
port 41 nsew
rlabel locali s 84251 -41372 87163 -41306 8 VDD
port 41 nsew
rlabel locali s 87658 -41301 87780 -40305 8 VDD
port 41 nsew
rlabel locali s 85052 -41306 87163 -41272 8 VDD
port 41 nsew
rlabel locali s 86050 -41272 86668 -41255 8 VDD
port 41 nsew
rlabel locali s 86050 -41255 86493 -41226 8 VDD
port 41 nsew
rlabel locali s 86051 -41226 86493 -41212 8 VDD
port 41 nsew
rlabel locali s 86051 -41212 87340 -41163 8 VDD
port 41 nsew
rlabel locali s 86453 -41163 87340 -41113 8 VDD
port 41 nsew
rlabel locali s 87258 -41113 87292 -40947 8 VDD
port 41 nsew
rlabel locali s 87062 -41113 87096 -40947 8 VDD
port 41 nsew
rlabel locali s 86866 -41113 86900 -40947 8 VDD
port 41 nsew
rlabel locali s 86670 -41113 86704 -40947 8 VDD
port 41 nsew
rlabel locali s 86453 -41113 86487 -40746 8 VDD
port 41 nsew
rlabel locali s 86257 -41163 86291 -40746 8 VDD
port 41 nsew
rlabel locali s 86061 -41163 86095 -40746 8 VDD
port 41 nsew
rlabel locali s 85222 -41272 85394 -41082 8 VDD
port 41 nsew
rlabel locali s 85040 -41082 85758 -40983 8 VDD
port 41 nsew
rlabel locali s 85676 -40983 85710 -40717 8 VDD
port 41 nsew
rlabel locali s 85480 -40983 85514 -40717 8 VDD
port 41 nsew
rlabel locali s 85284 -40983 85318 -40717 8 VDD
port 41 nsew
rlabel locali s 85088 -40983 85122 -40717 8 VDD
port 41 nsew
rlabel locali s 87148 -40305 87780 -40183 8 VDD
port 41 nsew
rlabel locali s 87148 -40183 87270 -37786 8 VDD
port 41 nsew
rlabel locali s 84251 -41306 84317 -39976 8 VDD
port 41 nsew
rlabel locali s 83898 -41390 83982 -41277 8 VDD
port 41 nsew
rlabel locali s 81384 -41394 83599 -41352 8 VDD
port 41 nsew
rlabel locali s 83915 -41277 83981 -39976 8 VDD
port 41 nsew
rlabel locali s 81384 -41352 83495 -41241 8 VDD
port 41 nsew
rlabel locali s 78204 -41478 78416 -41339 8 VDD
port 41 nsew
rlabel locali s 77954 -41493 78033 -41468 8 VDD
port 41 nsew
rlabel locali s 77757 -41611 77802 -41487 8 VDD
port 41 nsew
rlabel locali s 77341 -42203 77375 -41610 8 VDD
port 41 nsew
rlabel locali s 77145 -42203 77179 -41613 8 VDD
port 41 nsew
rlabel locali s 76895 -41791 76929 -41625 8 VDD
port 41 nsew
rlabel locali s 76699 -41791 76733 -41625 8 VDD
port 41 nsew
rlabel locali s 76503 -41791 76537 -41625 8 VDD
port 41 nsew
rlabel locali s 76307 -41791 76341 -41625 8 VDD
port 41 nsew
rlabel locali s 76090 -41992 76124 -41625 8 VDD
port 41 nsew
rlabel locali s 77335 -41610 77380 -41487 8 VDD
port 41 nsew
rlabel locali s 77140 -41613 77185 -41487 8 VDD
port 41 nsew
rlabel locali s 76090 -41625 76977 -41575 8 VDD
port 41 nsew
rlabel locali s 75894 -41992 75928 -41575 8 VDD
port 41 nsew
rlabel locali s 75698 -41992 75732 -41575 8 VDD
port 41 nsew
rlabel locali s 74096 -42172 74130 -41580 8 VDD
port 41 nsew
rlabel locali s 75688 -41575 76977 -41526 8 VDD
port 41 nsew
rlabel locali s 75688 -41526 76130 -41511 8 VDD
port 41 nsew
rlabel locali s 77134 -41487 77903 -41468 8 VDD
port 41 nsew
rlabel locali s 77134 -41468 78033 -41463 8 VDD
port 41 nsew
rlabel locali s 76127 -41477 76316 -41470 8 VDD
port 41 nsew
rlabel locali s 76090 -41470 76316 -41463 8 VDD
port 41 nsew
rlabel locali s 75688 -41463 78033 -41421 8 VDD
port 41 nsew
rlabel locali s 74089 -41580 74134 -41456 8 VDD
port 41 nsew
rlabel locali s 73673 -42172 73707 -41579 8 VDD
port 41 nsew
rlabel locali s 73477 -42172 73511 -41582 8 VDD
port 41 nsew
rlabel locali s 73227 -41760 73261 -41594 8 VDD
port 41 nsew
rlabel locali s 73031 -41760 73065 -41594 8 VDD
port 41 nsew
rlabel locali s 72835 -41760 72869 -41594 8 VDD
port 41 nsew
rlabel locali s 72639 -41760 72673 -41594 8 VDD
port 41 nsew
rlabel locali s 72422 -41961 72456 -41594 8 VDD
port 41 nsew
rlabel locali s 73667 -41579 73712 -41456 8 VDD
port 41 nsew
rlabel locali s 73472 -41582 73517 -41456 8 VDD
port 41 nsew
rlabel locali s 72422 -41594 73309 -41544 8 VDD
port 41 nsew
rlabel locali s 72226 -41961 72260 -41544 8 VDD
port 41 nsew
rlabel locali s 72030 -41961 72064 -41544 8 VDD
port 41 nsew
rlabel locali s 68611 -42220 68645 -41628 8 VDD
port 41 nsew
rlabel locali s 72020 -41544 73309 -41495 8 VDD
port 41 nsew
rlabel locali s 69051 -41523 69190 -41495 8 VDD
port 41 nsew
rlabel locali s 72020 -41495 72462 -41480 8 VDD
port 41 nsew
rlabel locali s 73466 -41456 74235 -41432 8 VDD
port 41 nsew
rlabel locali s 72459 -41446 72648 -41439 8 VDD
port 41 nsew
rlabel locali s 72422 -41439 72648 -41432 8 VDD
port 41 nsew
rlabel locali s 77854 -41421 78033 -41385 8 VDD
port 41 nsew
rlabel locali s 75688 -41421 77799 -41410 8 VDD
port 41 nsew
rlabel locali s 77954 -41385 78033 -41354 8 VDD
port 41 nsew
rlabel locali s 74887 -41410 77799 -41344 8 VDD
port 41 nsew
rlabel locali s 82382 -41241 83000 -41224 8 VDD
port 41 nsew
rlabel locali s 82382 -41224 82825 -41195 8 VDD
port 41 nsew
rlabel locali s 82383 -41195 82825 -41181 8 VDD
port 41 nsew
rlabel locali s 82383 -41181 83672 -41132 8 VDD
port 41 nsew
rlabel locali s 82785 -41132 83672 -41082 8 VDD
port 41 nsew
rlabel locali s 83590 -41082 83624 -40916 8 VDD
port 41 nsew
rlabel locali s 83394 -41082 83428 -40916 8 VDD
port 41 nsew
rlabel locali s 83198 -41082 83232 -40916 8 VDD
port 41 nsew
rlabel locali s 83002 -41082 83036 -40916 8 VDD
port 41 nsew
rlabel locali s 82785 -41082 82819 -40715 8 VDD
port 41 nsew
rlabel locali s 82589 -41132 82623 -40715 8 VDD
port 41 nsew
rlabel locali s 82393 -41132 82427 -40715 8 VDD
port 41 nsew
rlabel locali s 81554 -41241 81726 -41051 8 VDD
port 41 nsew
rlabel locali s 81372 -41051 82090 -40952 8 VDD
port 41 nsew
rlabel locali s 82008 -40952 82042 -40686 8 VDD
port 41 nsew
rlabel locali s 81812 -40952 81846 -40686 8 VDD
port 41 nsew
rlabel locali s 81616 -40952 81650 -40686 8 VDD
port 41 nsew
rlabel locali s 81420 -40952 81454 -40686 8 VDD
port 41 nsew
rlabel locali s 78294 -41339 78416 -40343 8 VDD
port 41 nsew
rlabel locali s 75688 -41344 77799 -41310 8 VDD
port 41 nsew
rlabel locali s 76686 -41310 77304 -41293 8 VDD
port 41 nsew
rlabel locali s 76686 -41293 77129 -41264 8 VDD
port 41 nsew
rlabel locali s 76687 -41264 77129 -41250 8 VDD
port 41 nsew
rlabel locali s 76687 -41250 77976 -41201 8 VDD
port 41 nsew
rlabel locali s 77089 -41201 77976 -41151 8 VDD
port 41 nsew
rlabel locali s 77894 -41151 77928 -40985 8 VDD
port 41 nsew
rlabel locali s 77698 -41151 77732 -40985 8 VDD
port 41 nsew
rlabel locali s 77502 -41151 77536 -40985 8 VDD
port 41 nsew
rlabel locali s 77306 -41151 77340 -40985 8 VDD
port 41 nsew
rlabel locali s 77089 -41151 77123 -40784 8 VDD
port 41 nsew
rlabel locali s 76893 -41201 76927 -40784 8 VDD
port 41 nsew
rlabel locali s 76697 -41201 76731 -40784 8 VDD
port 41 nsew
rlabel locali s 75858 -41310 76030 -41120 8 VDD
port 41 nsew
rlabel locali s 75676 -41120 76394 -41021 8 VDD
port 41 nsew
rlabel locali s 76312 -41021 76346 -40755 8 VDD
port 41 nsew
rlabel locali s 76116 -41021 76150 -40755 8 VDD
port 41 nsew
rlabel locali s 75920 -41021 75954 -40755 8 VDD
port 41 nsew
rlabel locali s 75724 -41021 75758 -40755 8 VDD
port 41 nsew
rlabel locali s 77784 -40343 78416 -40221 8 VDD
port 41 nsew
rlabel locali s 83915 -39976 84317 -39910 8 VDD
port 41 nsew
rlabel locali s 86186 -38239 86220 -37947 8 VDD
port 41 nsew
rlabel locali s 85990 -38239 86024 -37949 8 VDD
port 41 nsew
rlabel locali s 85762 -38439 85796 -37964 8 VDD
port 41 nsew
rlabel locali s 85632 -38439 85666 -37967 8 VDD
port 41 nsew
rlabel locali s 86181 -37947 86224 -37787 8 VDD
port 41 nsew
rlabel locali s 85984 -37949 86027 -37787 8 VDD
port 41 nsew
rlabel locali s 85753 -37964 85803 -37787 8 VDD
port 41 nsew
rlabel locali s 85627 -37967 85677 -37787 8 VDD
port 41 nsew
rlabel locali s 85037 -38439 85071 -37944 8 VDD
port 41 nsew
rlabel locali s 84841 -38439 84875 -37946 8 VDD
port 41 nsew
rlabel locali s 83468 -38681 83502 -38089 8 VDD
port 41 nsew
rlabel locali s 83908 -37984 84006 -37978 8 VDD
port 41 nsew
rlabel locali s 85035 -37944 85073 -37787 8 VDD
port 41 nsew
rlabel locali s 84838 -37946 84876 -37851 8 VDD
port 41 nsew
rlabel locali s 83908 -37978 84588 -37861 8 VDD
port 41 nsew
rlabel locali s 83680 -37972 83742 -37958 8 VDD
port 41 nsew
rlabel locali s 83461 -38089 83506 -37965 8 VDD
port 41 nsew
rlabel locali s 83045 -38681 83079 -38088 8 VDD
port 41 nsew
rlabel locali s 82849 -38681 82883 -38091 8 VDD
port 41 nsew
rlabel locali s 82599 -38269 82633 -38103 8 VDD
port 41 nsew
rlabel locali s 82403 -38269 82437 -38103 8 VDD
port 41 nsew
rlabel locali s 82207 -38269 82241 -38103 8 VDD
port 41 nsew
rlabel locali s 82011 -38269 82045 -38103 8 VDD
port 41 nsew
rlabel locali s 81794 -38470 81828 -38103 8 VDD
port 41 nsew
rlabel locali s 83039 -38088 83084 -37965 8 VDD
port 41 nsew
rlabel locali s 82844 -38091 82889 -37965 8 VDD
port 41 nsew
rlabel locali s 81794 -38103 82681 -38053 8 VDD
port 41 nsew
rlabel locali s 81598 -38470 81632 -38053 8 VDD
port 41 nsew
rlabel locali s 81402 -38470 81436 -38053 8 VDD
port 41 nsew
rlabel locali s 81392 -38053 82681 -38004 8 VDD
port 41 nsew
rlabel locali s 81392 -38004 81834 -37989 8 VDD
port 41 nsew
rlabel locali s 82838 -37965 83607 -37958 8 VDD
port 41 nsew
rlabel locali s 82838 -37958 83742 -37941 8 VDD
port 41 nsew
rlabel locali s 81831 -37955 82020 -37948 8 VDD
port 41 nsew
rlabel locali s 81794 -37948 82020 -37941 8 VDD
port 41 nsew
rlabel locali s 81392 -37941 83742 -37906 8 VDD
port 41 nsew
rlabel locali s 83680 -37906 83742 -37878 8 VDD
port 41 nsew
rlabel locali s 81392 -37906 83607 -37899 8 VDD
port 41 nsew
rlabel locali s 81392 -37899 83503 -37885 8 VDD
port 41 nsew
rlabel locali s 77784 -40221 77906 -37885 8 VDD
port 41 nsew
rlabel locali s 74887 -41344 74953 -40014 8 VDD
port 41 nsew
rlabel locali s 74534 -41428 74618 -41315 8 VDD
port 41 nsew
rlabel locali s 72020 -41432 74235 -41390 8 VDD
port 41 nsew
rlabel locali s 74551 -41315 74617 -40014 8 VDD
port 41 nsew
rlabel locali s 72020 -41390 74131 -41279 8 VDD
port 41 nsew
rlabel locali s 69051 -41495 69263 -41356 8 VDD
port 41 nsew
rlabel locali s 68801 -41510 68880 -41485 8 VDD
port 41 nsew
rlabel locali s 68604 -41628 68649 -41504 8 VDD
port 41 nsew
rlabel locali s 68188 -42220 68222 -41627 8 VDD
port 41 nsew
rlabel locali s 67992 -42220 68026 -41630 8 VDD
port 41 nsew
rlabel locali s 67742 -41808 67776 -41642 8 VDD
port 41 nsew
rlabel locali s 67546 -41808 67580 -41642 8 VDD
port 41 nsew
rlabel locali s 67350 -41808 67384 -41642 8 VDD
port 41 nsew
rlabel locali s 67154 -41808 67188 -41642 8 VDD
port 41 nsew
rlabel locali s 66937 -42009 66971 -41642 8 VDD
port 41 nsew
rlabel locali s 68182 -41627 68227 -41504 8 VDD
port 41 nsew
rlabel locali s 67987 -41630 68032 -41504 8 VDD
port 41 nsew
rlabel locali s 66937 -41642 67824 -41592 8 VDD
port 41 nsew
rlabel locali s 66741 -42009 66775 -41592 8 VDD
port 41 nsew
rlabel locali s 66545 -42009 66579 -41592 8 VDD
port 41 nsew
rlabel locali s 64943 -42189 64977 -41597 8 VDD
port 41 nsew
rlabel locali s 66535 -41592 67824 -41543 8 VDD
port 41 nsew
rlabel locali s 66535 -41543 66977 -41528 8 VDD
port 41 nsew
rlabel locali s 67981 -41504 68750 -41485 8 VDD
port 41 nsew
rlabel locali s 67981 -41485 68880 -41480 8 VDD
port 41 nsew
rlabel locali s 66974 -41494 67163 -41487 8 VDD
port 41 nsew
rlabel locali s 66937 -41487 67163 -41480 8 VDD
port 41 nsew
rlabel locali s 66535 -41480 68880 -41438 8 VDD
port 41 nsew
rlabel locali s 64936 -41597 64981 -41473 8 VDD
port 41 nsew
rlabel locali s 64520 -42189 64554 -41596 8 VDD
port 41 nsew
rlabel locali s 64324 -42189 64358 -41599 8 VDD
port 41 nsew
rlabel locali s 64074 -41777 64108 -41611 8 VDD
port 41 nsew
rlabel locali s 63878 -41777 63912 -41611 8 VDD
port 41 nsew
rlabel locali s 63682 -41777 63716 -41611 8 VDD
port 41 nsew
rlabel locali s 63486 -41777 63520 -41611 8 VDD
port 41 nsew
rlabel locali s 63269 -41978 63303 -41611 8 VDD
port 41 nsew
rlabel locali s 64514 -41596 64559 -41473 8 VDD
port 41 nsew
rlabel locali s 64319 -41599 64364 -41473 8 VDD
port 41 nsew
rlabel locali s 63269 -41611 64156 -41561 8 VDD
port 41 nsew
rlabel locali s 63073 -41978 63107 -41561 8 VDD
port 41 nsew
rlabel locali s 62877 -41978 62911 -41561 8 VDD
port 41 nsew
rlabel locali s 59857 -42286 59891 -41694 8 VDD
port 41 nsew
rlabel locali s 60297 -41589 60436 -41561 8 VDD
port 41 nsew
rlabel locali s 62867 -41561 64156 -41512 8 VDD
port 41 nsew
rlabel locali s 62867 -41512 63309 -41497 8 VDD
port 41 nsew
rlabel locali s 64313 -41473 65082 -41449 8 VDD
port 41 nsew
rlabel locali s 63306 -41463 63495 -41456 8 VDD
port 41 nsew
rlabel locali s 63269 -41456 63495 -41449 8 VDD
port 41 nsew
rlabel locali s 68701 -41438 68880 -41402 8 VDD
port 41 nsew
rlabel locali s 66535 -41438 68646 -41427 8 VDD
port 41 nsew
rlabel locali s 68801 -41402 68880 -41371 8 VDD
port 41 nsew
rlabel locali s 65734 -41427 68646 -41361 8 VDD
port 41 nsew
rlabel locali s 73018 -41279 73636 -41262 8 VDD
port 41 nsew
rlabel locali s 73018 -41262 73461 -41233 8 VDD
port 41 nsew
rlabel locali s 73019 -41233 73461 -41219 8 VDD
port 41 nsew
rlabel locali s 73019 -41219 74308 -41170 8 VDD
port 41 nsew
rlabel locali s 73421 -41170 74308 -41120 8 VDD
port 41 nsew
rlabel locali s 74226 -41120 74260 -40954 8 VDD
port 41 nsew
rlabel locali s 74030 -41120 74064 -40954 8 VDD
port 41 nsew
rlabel locali s 73834 -41120 73868 -40954 8 VDD
port 41 nsew
rlabel locali s 73638 -41120 73672 -40954 8 VDD
port 41 nsew
rlabel locali s 73421 -41120 73455 -40753 8 VDD
port 41 nsew
rlabel locali s 73225 -41170 73259 -40753 8 VDD
port 41 nsew
rlabel locali s 73029 -41170 73063 -40753 8 VDD
port 41 nsew
rlabel locali s 72190 -41279 72362 -41089 8 VDD
port 41 nsew
rlabel locali s 72008 -41089 72726 -40990 8 VDD
port 41 nsew
rlabel locali s 72644 -40990 72678 -40724 8 VDD
port 41 nsew
rlabel locali s 72448 -40990 72482 -40724 8 VDD
port 41 nsew
rlabel locali s 72252 -40990 72286 -40724 8 VDD
port 41 nsew
rlabel locali s 72056 -40990 72090 -40724 8 VDD
port 41 nsew
rlabel locali s 69141 -41356 69263 -40360 8 VDD
port 41 nsew
rlabel locali s 66535 -41361 68646 -41327 8 VDD
port 41 nsew
rlabel locali s 67533 -41327 68151 -41310 8 VDD
port 41 nsew
rlabel locali s 67533 -41310 67976 -41281 8 VDD
port 41 nsew
rlabel locali s 67534 -41281 67976 -41267 8 VDD
port 41 nsew
rlabel locali s 67534 -41267 68823 -41218 8 VDD
port 41 nsew
rlabel locali s 67936 -41218 68823 -41168 8 VDD
port 41 nsew
rlabel locali s 68741 -41168 68775 -41002 8 VDD
port 41 nsew
rlabel locali s 68545 -41168 68579 -41002 8 VDD
port 41 nsew
rlabel locali s 68349 -41168 68383 -41002 8 VDD
port 41 nsew
rlabel locali s 68153 -41168 68187 -41002 8 VDD
port 41 nsew
rlabel locali s 67936 -41168 67970 -40801 8 VDD
port 41 nsew
rlabel locali s 67740 -41218 67774 -40801 8 VDD
port 41 nsew
rlabel locali s 67544 -41218 67578 -40801 8 VDD
port 41 nsew
rlabel locali s 66705 -41327 66877 -41137 8 VDD
port 41 nsew
rlabel locali s 66523 -41137 67241 -41038 8 VDD
port 41 nsew
rlabel locali s 67159 -41038 67193 -40772 8 VDD
port 41 nsew
rlabel locali s 66963 -41038 66997 -40772 8 VDD
port 41 nsew
rlabel locali s 66767 -41038 66801 -40772 8 VDD
port 41 nsew
rlabel locali s 66571 -41038 66605 -40772 8 VDD
port 41 nsew
rlabel locali s 68631 -40360 69263 -40238 8 VDD
port 41 nsew
rlabel locali s 74551 -40014 74953 -39948 8 VDD
port 41 nsew
rlabel locali s 76822 -38277 76856 -37985 8 VDD
port 41 nsew
rlabel locali s 76626 -38277 76660 -37987 8 VDD
port 41 nsew
rlabel locali s 76398 -38477 76432 -38002 8 VDD
port 41 nsew
rlabel locali s 76268 -38477 76302 -38005 8 VDD
port 41 nsew
rlabel locali s 76817 -37985 76860 -37885 8 VDD
port 41 nsew
rlabel locali s 84471 -37861 84588 -37851 8 VDD
port 41 nsew
rlabel locali s 83908 -37861 84006 -37858 8 VDD
port 41 nsew
rlabel locali s 84471 -37851 84876 -37787 8 VDD
port 41 nsew
rlabel locali s 76817 -37885 83503 -37825 8 VDD
port 41 nsew
rlabel locali s 76620 -37987 76663 -37825 8 VDD
port 41 nsew
rlabel locali s 76389 -38002 76439 -37825 8 VDD
port 41 nsew
rlabel locali s 76263 -38005 76313 -37825 8 VDD
port 41 nsew
rlabel locali s 75673 -38477 75707 -37982 8 VDD
port 41 nsew
rlabel locali s 75477 -38477 75511 -37984 8 VDD
port 41 nsew
rlabel locali s 74104 -38719 74138 -38127 8 VDD
port 41 nsew
rlabel locali s 74544 -38022 74642 -38016 8 VDD
port 41 nsew
rlabel locali s 75671 -37982 75709 -37825 8 VDD
port 41 nsew
rlabel locali s 75474 -37984 75512 -37889 8 VDD
port 41 nsew
rlabel locali s 74544 -38016 75224 -37899 8 VDD
port 41 nsew
rlabel locali s 74316 -38010 74378 -37996 8 VDD
port 41 nsew
rlabel locali s 74097 -38127 74142 -38003 8 VDD
port 41 nsew
rlabel locali s 73681 -38719 73715 -38126 8 VDD
port 41 nsew
rlabel locali s 73485 -38719 73519 -38129 8 VDD
port 41 nsew
rlabel locali s 73235 -38307 73269 -38141 8 VDD
port 41 nsew
rlabel locali s 73039 -38307 73073 -38141 8 VDD
port 41 nsew
rlabel locali s 72843 -38307 72877 -38141 8 VDD
port 41 nsew
rlabel locali s 72647 -38307 72681 -38141 8 VDD
port 41 nsew
rlabel locali s 72430 -38508 72464 -38141 8 VDD
port 41 nsew
rlabel locali s 73675 -38126 73720 -38003 8 VDD
port 41 nsew
rlabel locali s 73480 -38129 73525 -38003 8 VDD
port 41 nsew
rlabel locali s 72430 -38141 73317 -38091 8 VDD
port 41 nsew
rlabel locali s 72234 -38508 72268 -38091 8 VDD
port 41 nsew
rlabel locali s 72038 -38508 72072 -38091 8 VDD
port 41 nsew
rlabel locali s 72028 -38091 73317 -38042 8 VDD
port 41 nsew
rlabel locali s 72028 -38042 72470 -38027 8 VDD
port 41 nsew
rlabel locali s 73474 -38003 74243 -37996 8 VDD
port 41 nsew
rlabel locali s 73474 -37996 74378 -37979 8 VDD
port 41 nsew
rlabel locali s 72467 -37993 72656 -37986 8 VDD
port 41 nsew
rlabel locali s 72430 -37986 72656 -37979 8 VDD
port 41 nsew
rlabel locali s 72028 -37979 74378 -37944 8 VDD
port 41 nsew
rlabel locali s 74316 -37944 74378 -37916 8 VDD
port 41 nsew
rlabel locali s 72028 -37944 74243 -37937 8 VDD
port 41 nsew
rlabel locali s 75107 -37899 75224 -37889 8 VDD
port 41 nsew
rlabel locali s 74544 -37899 74642 -37896 8 VDD
port 41 nsew
rlabel locali s 75107 -37889 75512 -37825 8 VDD
port 41 nsew
rlabel locali s 72028 -37937 74139 -37876 8 VDD
port 41 nsew
rlabel locali s 68631 -40238 68753 -37876 8 VDD
port 41 nsew
rlabel locali s 65734 -41361 65800 -40031 8 VDD
port 41 nsew
rlabel locali s 65381 -41445 65465 -41332 8 VDD
port 41 nsew
rlabel locali s 62867 -41449 65082 -41407 8 VDD
port 41 nsew
rlabel locali s 65398 -41332 65464 -40031 8 VDD
port 41 nsew
rlabel locali s 62867 -41407 64978 -41296 8 VDD
port 41 nsew
rlabel locali s 60297 -41561 60509 -41422 8 VDD
port 41 nsew
rlabel locali s 60047 -41576 60126 -41551 8 VDD
port 41 nsew
rlabel locali s 59850 -41694 59895 -41570 8 VDD
port 41 nsew
rlabel locali s 59434 -42286 59468 -41693 8 VDD
port 41 nsew
rlabel locali s 59238 -42286 59272 -41696 8 VDD
port 41 nsew
rlabel locali s 58988 -41874 59022 -41708 8 VDD
port 41 nsew
rlabel locali s 58792 -41874 58826 -41708 8 VDD
port 41 nsew
rlabel locali s 58596 -41874 58630 -41708 8 VDD
port 41 nsew
rlabel locali s 58400 -41874 58434 -41708 8 VDD
port 41 nsew
rlabel locali s 58183 -42075 58217 -41708 8 VDD
port 41 nsew
rlabel locali s 59428 -41693 59473 -41570 8 VDD
port 41 nsew
rlabel locali s 59233 -41696 59278 -41570 8 VDD
port 41 nsew
rlabel locali s 58183 -41708 59070 -41658 8 VDD
port 41 nsew
rlabel locali s 57987 -42075 58021 -41658 8 VDD
port 41 nsew
rlabel locali s 57791 -42075 57825 -41658 8 VDD
port 41 nsew
rlabel locali s 56189 -42255 56223 -41663 8 VDD
port 41 nsew
rlabel locali s 57781 -41658 59070 -41609 8 VDD
port 41 nsew
rlabel locali s 57781 -41609 58223 -41594 8 VDD
port 41 nsew
rlabel locali s 59227 -41570 59996 -41551 8 VDD
port 41 nsew
rlabel locali s 59227 -41551 60126 -41546 8 VDD
port 41 nsew
rlabel locali s 58220 -41560 58409 -41553 8 VDD
port 41 nsew
rlabel locali s 58183 -41553 58409 -41546 8 VDD
port 41 nsew
rlabel locali s 57781 -41546 60126 -41504 8 VDD
port 41 nsew
rlabel locali s 56182 -41663 56227 -41539 8 VDD
port 41 nsew
rlabel locali s 55766 -42255 55800 -41662 8 VDD
port 41 nsew
rlabel locali s 55570 -42255 55604 -41665 8 VDD
port 41 nsew
rlabel locali s 55320 -41843 55354 -41677 8 VDD
port 41 nsew
rlabel locali s 55124 -41843 55158 -41677 8 VDD
port 41 nsew
rlabel locali s 54928 -41843 54962 -41677 8 VDD
port 41 nsew
rlabel locali s 54732 -41843 54766 -41677 8 VDD
port 41 nsew
rlabel locali s 54515 -42044 54549 -41677 8 VDD
port 41 nsew
rlabel locali s 55760 -41662 55805 -41539 8 VDD
port 41 nsew
rlabel locali s 55565 -41665 55610 -41539 8 VDD
port 41 nsew
rlabel locali s 54515 -41677 55402 -41627 8 VDD
port 41 nsew
rlabel locali s 54319 -42044 54353 -41627 8 VDD
port 41 nsew
rlabel locali s 54123 -42044 54157 -41627 8 VDD
port 41 nsew
rlabel locali s 50659 -42320 50693 -41728 8 VDD
port 41 nsew
rlabel locali s 54113 -41627 55402 -41578 8 VDD
port 41 nsew
rlabel locali s 51099 -41623 51238 -41595 8 VDD
port 41 nsew
rlabel locali s 54113 -41578 54555 -41563 8 VDD
port 41 nsew
rlabel locali s 55559 -41539 56328 -41515 8 VDD
port 41 nsew
rlabel locali s 54552 -41529 54741 -41522 8 VDD
port 41 nsew
rlabel locali s 54515 -41522 54741 -41515 8 VDD
port 41 nsew
rlabel locali s 59947 -41504 60126 -41468 8 VDD
port 41 nsew
rlabel locali s 57781 -41504 59892 -41493 8 VDD
port 41 nsew
rlabel locali s 60047 -41468 60126 -41437 8 VDD
port 41 nsew
rlabel locali s 56980 -41493 59892 -41427 8 VDD
port 41 nsew
rlabel locali s 63865 -41296 64483 -41279 8 VDD
port 41 nsew
rlabel locali s 63865 -41279 64308 -41250 8 VDD
port 41 nsew
rlabel locali s 63866 -41250 64308 -41236 8 VDD
port 41 nsew
rlabel locali s 63866 -41236 65155 -41187 8 VDD
port 41 nsew
rlabel locali s 64268 -41187 65155 -41137 8 VDD
port 41 nsew
rlabel locali s 65073 -41137 65107 -40971 8 VDD
port 41 nsew
rlabel locali s 64877 -41137 64911 -40971 8 VDD
port 41 nsew
rlabel locali s 64681 -41137 64715 -40971 8 VDD
port 41 nsew
rlabel locali s 64485 -41137 64519 -40971 8 VDD
port 41 nsew
rlabel locali s 64268 -41137 64302 -40770 8 VDD
port 41 nsew
rlabel locali s 64072 -41187 64106 -40770 8 VDD
port 41 nsew
rlabel locali s 63876 -41187 63910 -40770 8 VDD
port 41 nsew
rlabel locali s 63037 -41296 63209 -41106 8 VDD
port 41 nsew
rlabel locali s 62855 -41106 63573 -41007 8 VDD
port 41 nsew
rlabel locali s 63491 -41007 63525 -40741 8 VDD
port 41 nsew
rlabel locali s 63295 -41007 63329 -40741 8 VDD
port 41 nsew
rlabel locali s 63099 -41007 63133 -40741 8 VDD
port 41 nsew
rlabel locali s 62903 -41007 62937 -40741 8 VDD
port 41 nsew
rlabel locali s 60387 -41422 60509 -40426 8 VDD
port 41 nsew
rlabel locali s 57781 -41427 59892 -41393 8 VDD
port 41 nsew
rlabel locali s 58779 -41393 59397 -41376 8 VDD
port 41 nsew
rlabel locali s 58779 -41376 59222 -41347 8 VDD
port 41 nsew
rlabel locali s 58780 -41347 59222 -41333 8 VDD
port 41 nsew
rlabel locali s 58780 -41333 60069 -41284 8 VDD
port 41 nsew
rlabel locali s 59182 -41284 60069 -41234 8 VDD
port 41 nsew
rlabel locali s 59987 -41234 60021 -41068 8 VDD
port 41 nsew
rlabel locali s 59791 -41234 59825 -41068 8 VDD
port 41 nsew
rlabel locali s 59595 -41234 59629 -41068 8 VDD
port 41 nsew
rlabel locali s 59399 -41234 59433 -41068 8 VDD
port 41 nsew
rlabel locali s 59182 -41234 59216 -40867 8 VDD
port 41 nsew
rlabel locali s 58986 -41284 59020 -40867 8 VDD
port 41 nsew
rlabel locali s 58790 -41284 58824 -40867 8 VDD
port 41 nsew
rlabel locali s 57951 -41393 58123 -41203 8 VDD
port 41 nsew
rlabel locali s 57769 -41203 58487 -41104 8 VDD
port 41 nsew
rlabel locali s 58405 -41104 58439 -40838 8 VDD
port 41 nsew
rlabel locali s 58209 -41104 58243 -40838 8 VDD
port 41 nsew
rlabel locali s 58013 -41104 58047 -40838 8 VDD
port 41 nsew
rlabel locali s 57817 -41104 57851 -40838 8 VDD
port 41 nsew
rlabel locali s 59877 -40426 60509 -40304 8 VDD
port 41 nsew
rlabel locali s 65398 -40031 65800 -39965 8 VDD
port 41 nsew
rlabel locali s 67669 -38294 67703 -38002 8 VDD
port 41 nsew
rlabel locali s 67473 -38294 67507 -38004 8 VDD
port 41 nsew
rlabel locali s 67245 -38494 67279 -38019 8 VDD
port 41 nsew
rlabel locali s 67115 -38494 67149 -38022 8 VDD
port 41 nsew
rlabel locali s 67664 -38002 67707 -37876 8 VDD
port 41 nsew
rlabel locali s 67659 -37876 74139 -37842 8 VDD
port 41 nsew
rlabel locali s 67467 -38004 67510 -37842 8 VDD
port 41 nsew
rlabel locali s 67236 -38019 67286 -37842 8 VDD
port 41 nsew
rlabel locali s 67110 -38022 67160 -37842 8 VDD
port 41 nsew
rlabel locali s 66520 -38494 66554 -37999 8 VDD
port 41 nsew
rlabel locali s 66324 -38494 66358 -38001 8 VDD
port 41 nsew
rlabel locali s 64951 -38736 64985 -38144 8 VDD
port 41 nsew
rlabel locali s 65391 -38039 65489 -38033 8 VDD
port 41 nsew
rlabel locali s 66518 -37999 66556 -37842 8 VDD
port 41 nsew
rlabel locali s 66321 -38001 66359 -37906 8 VDD
port 41 nsew
rlabel locali s 65391 -38033 66071 -37916 8 VDD
port 41 nsew
rlabel locali s 65163 -38027 65225 -38013 8 VDD
port 41 nsew
rlabel locali s 64944 -38144 64989 -38020 8 VDD
port 41 nsew
rlabel locali s 64528 -38736 64562 -38143 8 VDD
port 41 nsew
rlabel locali s 64332 -38736 64366 -38146 8 VDD
port 41 nsew
rlabel locali s 64082 -38324 64116 -38158 8 VDD
port 41 nsew
rlabel locali s 63886 -38324 63920 -38158 8 VDD
port 41 nsew
rlabel locali s 63690 -38324 63724 -38158 8 VDD
port 41 nsew
rlabel locali s 63494 -38324 63528 -38158 8 VDD
port 41 nsew
rlabel locali s 63277 -38525 63311 -38158 8 VDD
port 41 nsew
rlabel locali s 64522 -38143 64567 -38020 8 VDD
port 41 nsew
rlabel locali s 64327 -38146 64372 -38020 8 VDD
port 41 nsew
rlabel locali s 63277 -38158 64164 -38108 8 VDD
port 41 nsew
rlabel locali s 63081 -38525 63115 -38108 8 VDD
port 41 nsew
rlabel locali s 62885 -38525 62919 -38108 8 VDD
port 41 nsew
rlabel locali s 62875 -38108 64164 -38059 8 VDD
port 41 nsew
rlabel locali s 62875 -38059 63317 -38044 8 VDD
port 41 nsew
rlabel locali s 64321 -38020 65090 -38013 8 VDD
port 41 nsew
rlabel locali s 64321 -38013 65225 -37996 8 VDD
port 41 nsew
rlabel locali s 63314 -38010 63503 -38003 8 VDD
port 41 nsew
rlabel locali s 63277 -38003 63503 -37996 8 VDD
port 41 nsew
rlabel locali s 62875 -37996 65225 -37970 8 VDD
port 41 nsew
rlabel locali s 59877 -40304 59999 -37970 8 VDD
port 41 nsew
rlabel locali s 56980 -41427 57046 -40097 8 VDD
port 41 nsew
rlabel locali s 56627 -41511 56711 -41398 8 VDD
port 41 nsew
rlabel locali s 54113 -41515 56328 -41473 8 VDD
port 41 nsew
rlabel locali s 56644 -41398 56710 -40097 8 VDD
port 41 nsew
rlabel locali s 54113 -41473 56224 -41362 8 VDD
port 41 nsew
rlabel locali s 51099 -41595 51311 -41456 8 VDD
port 41 nsew
rlabel locali s 50849 -41610 50928 -41585 8 VDD
port 41 nsew
rlabel locali s 50652 -41728 50697 -41604 8 VDD
port 41 nsew
rlabel locali s 50236 -42320 50270 -41727 8 VDD
port 41 nsew
rlabel locali s 50040 -42320 50074 -41730 8 VDD
port 41 nsew
rlabel locali s 49790 -41908 49824 -41742 8 VDD
port 41 nsew
rlabel locali s 49594 -41908 49628 -41742 8 VDD
port 41 nsew
rlabel locali s 49398 -41908 49432 -41742 8 VDD
port 41 nsew
rlabel locali s 49202 -41908 49236 -41742 8 VDD
port 41 nsew
rlabel locali s 48985 -42109 49019 -41742 8 VDD
port 41 nsew
rlabel locali s 50230 -41727 50275 -41604 8 VDD
port 41 nsew
rlabel locali s 50035 -41730 50080 -41604 8 VDD
port 41 nsew
rlabel locali s 48985 -41742 49872 -41692 8 VDD
port 41 nsew
rlabel locali s 48789 -42109 48823 -41692 8 VDD
port 41 nsew
rlabel locali s 48593 -42109 48627 -41692 8 VDD
port 41 nsew
rlabel locali s 46991 -42289 47025 -41697 8 VDD
port 41 nsew
rlabel locali s 48583 -41692 49872 -41643 8 VDD
port 41 nsew
rlabel locali s 48583 -41643 49025 -41628 8 VDD
port 41 nsew
rlabel locali s 50029 -41604 50798 -41585 8 VDD
port 41 nsew
rlabel locali s 50029 -41585 50928 -41580 8 VDD
port 41 nsew
rlabel locali s 49022 -41594 49211 -41587 8 VDD
port 41 nsew
rlabel locali s 48985 -41587 49211 -41580 8 VDD
port 41 nsew
rlabel locali s 48583 -41580 50928 -41538 8 VDD
port 41 nsew
rlabel locali s 46984 -41697 47029 -41573 8 VDD
port 41 nsew
rlabel locali s 46568 -42289 46602 -41696 8 VDD
port 41 nsew
rlabel locali s 46372 -42289 46406 -41699 8 VDD
port 41 nsew
rlabel locali s 46122 -41877 46156 -41711 8 VDD
port 41 nsew
rlabel locali s 45926 -41877 45960 -41711 8 VDD
port 41 nsew
rlabel locali s 45730 -41877 45764 -41711 8 VDD
port 41 nsew
rlabel locali s 45534 -41877 45568 -41711 8 VDD
port 41 nsew
rlabel locali s 45317 -42078 45351 -41711 8 VDD
port 41 nsew
rlabel locali s 46562 -41696 46607 -41573 8 VDD
port 41 nsew
rlabel locali s 46367 -41699 46412 -41573 8 VDD
port 41 nsew
rlabel locali s 45317 -41711 46204 -41661 8 VDD
port 41 nsew
rlabel locali s 45121 -42078 45155 -41661 8 VDD
port 41 nsew
rlabel locali s 44925 -42078 44959 -41661 8 VDD
port 41 nsew
rlabel locali s 41796 -42281 41830 -41689 8 VDD
port 41 nsew
rlabel locali s 44915 -41661 46204 -41612 8 VDD
port 41 nsew
rlabel locali s 44915 -41612 45357 -41597 8 VDD
port 41 nsew
rlabel locali s 46361 -41573 47130 -41549 8 VDD
port 41 nsew
rlabel locali s 45354 -41563 45543 -41556 8 VDD
port 41 nsew
rlabel locali s 42236 -41584 42375 -41556 8 VDD
port 41 nsew
rlabel locali s 45317 -41556 45543 -41549 8 VDD
port 41 nsew
rlabel locali s 50749 -41538 50928 -41502 8 VDD
port 41 nsew
rlabel locali s 48583 -41538 50694 -41527 8 VDD
port 41 nsew
rlabel locali s 50849 -41502 50928 -41471 8 VDD
port 41 nsew
rlabel locali s 47782 -41527 50694 -41461 8 VDD
port 41 nsew
rlabel locali s 55111 -41362 55729 -41345 8 VDD
port 41 nsew
rlabel locali s 55111 -41345 55554 -41316 8 VDD
port 41 nsew
rlabel locali s 55112 -41316 55554 -41302 8 VDD
port 41 nsew
rlabel locali s 55112 -41302 56401 -41253 8 VDD
port 41 nsew
rlabel locali s 55514 -41253 56401 -41203 8 VDD
port 41 nsew
rlabel locali s 56319 -41203 56353 -41037 8 VDD
port 41 nsew
rlabel locali s 56123 -41203 56157 -41037 8 VDD
port 41 nsew
rlabel locali s 55927 -41203 55961 -41037 8 VDD
port 41 nsew
rlabel locali s 55731 -41203 55765 -41037 8 VDD
port 41 nsew
rlabel locali s 55514 -41203 55548 -40836 8 VDD
port 41 nsew
rlabel locali s 55318 -41253 55352 -40836 8 VDD
port 41 nsew
rlabel locali s 55122 -41253 55156 -40836 8 VDD
port 41 nsew
rlabel locali s 54283 -41362 54455 -41172 8 VDD
port 41 nsew
rlabel locali s 54101 -41172 54819 -41073 8 VDD
port 41 nsew
rlabel locali s 54737 -41073 54771 -40807 8 VDD
port 41 nsew
rlabel locali s 54541 -41073 54575 -40807 8 VDD
port 41 nsew
rlabel locali s 54345 -41073 54379 -40807 8 VDD
port 41 nsew
rlabel locali s 54149 -41073 54183 -40807 8 VDD
port 41 nsew
rlabel locali s 51189 -41456 51311 -40460 8 VDD
port 41 nsew
rlabel locali s 48583 -41461 50694 -41427 8 VDD
port 41 nsew
rlabel locali s 49581 -41427 50199 -41410 8 VDD
port 41 nsew
rlabel locali s 49581 -41410 50024 -41381 8 VDD
port 41 nsew
rlabel locali s 49582 -41381 50024 -41367 8 VDD
port 41 nsew
rlabel locali s 49582 -41367 50871 -41318 8 VDD
port 41 nsew
rlabel locali s 49984 -41318 50871 -41268 8 VDD
port 41 nsew
rlabel locali s 50789 -41268 50823 -41102 8 VDD
port 41 nsew
rlabel locali s 50593 -41268 50627 -41102 8 VDD
port 41 nsew
rlabel locali s 50397 -41268 50431 -41102 8 VDD
port 41 nsew
rlabel locali s 50201 -41268 50235 -41102 8 VDD
port 41 nsew
rlabel locali s 49984 -41268 50018 -40901 8 VDD
port 41 nsew
rlabel locali s 49788 -41318 49822 -40901 8 VDD
port 41 nsew
rlabel locali s 49592 -41318 49626 -40901 8 VDD
port 41 nsew
rlabel locali s 48753 -41427 48925 -41237 8 VDD
port 41 nsew
rlabel locali s 48571 -41237 49289 -41138 8 VDD
port 41 nsew
rlabel locali s 49207 -41138 49241 -40872 8 VDD
port 41 nsew
rlabel locali s 49011 -41138 49045 -40872 8 VDD
port 41 nsew
rlabel locali s 48815 -41138 48849 -40872 8 VDD
port 41 nsew
rlabel locali s 48619 -41138 48653 -40872 8 VDD
port 41 nsew
rlabel locali s 50679 -40460 51311 -40338 8 VDD
port 41 nsew
rlabel locali s 56644 -40097 57046 -40031 8 VDD
port 41 nsew
rlabel locali s 58915 -38360 58949 -38068 8 VDD
port 41 nsew
rlabel locali s 58719 -38360 58753 -38070 8 VDD
port 41 nsew
rlabel locali s 58491 -38560 58525 -38085 8 VDD
port 41 nsew
rlabel locali s 58361 -38560 58395 -38088 8 VDD
port 41 nsew
rlabel locali s 58910 -38068 58953 -37970 8 VDD
port 41 nsew
rlabel locali s 58910 -37970 65225 -37961 8 VDD
port 41 nsew
rlabel locali s 65163 -37961 65225 -37933 8 VDD
port 41 nsew
rlabel locali s 58910 -37961 65090 -37954 8 VDD
port 41 nsew
rlabel locali s 65954 -37916 66071 -37906 8 VDD
port 41 nsew
rlabel locali s 65391 -37916 65489 -37913 8 VDD
port 41 nsew
rlabel locali s 65954 -37906 66359 -37842 8 VDD
port 41 nsew
rlabel locali s 58910 -37954 64986 -37908 8 VDD
port 41 nsew
rlabel locali s 58713 -38070 58756 -37908 8 VDD
port 41 nsew
rlabel locali s 58482 -38085 58532 -37908 8 VDD
port 41 nsew
rlabel locali s 58356 -38088 58406 -37908 8 VDD
port 41 nsew
rlabel locali s 57766 -38560 57800 -38065 8 VDD
port 41 nsew
rlabel locali s 57570 -38560 57604 -38067 8 VDD
port 41 nsew
rlabel locali s 56197 -38802 56231 -38210 8 VDD
port 41 nsew
rlabel locali s 56637 -38105 56735 -38099 8 VDD
port 41 nsew
rlabel locali s 57764 -38065 57802 -37908 8 VDD
port 41 nsew
rlabel locali s 57567 -38067 57605 -37972 8 VDD
port 41 nsew
rlabel locali s 56637 -38099 57317 -37982 8 VDD
port 41 nsew
rlabel locali s 56409 -38093 56471 -38079 8 VDD
port 41 nsew
rlabel locali s 56190 -38210 56235 -38086 8 VDD
port 41 nsew
rlabel locali s 55774 -38802 55808 -38209 8 VDD
port 41 nsew
rlabel locali s 55578 -38802 55612 -38212 8 VDD
port 41 nsew
rlabel locali s 55328 -38390 55362 -38224 8 VDD
port 41 nsew
rlabel locali s 55132 -38390 55166 -38224 8 VDD
port 41 nsew
rlabel locali s 54936 -38390 54970 -38224 8 VDD
port 41 nsew
rlabel locali s 54740 -38390 54774 -38224 8 VDD
port 41 nsew
rlabel locali s 54523 -38591 54557 -38224 8 VDD
port 41 nsew
rlabel locali s 55768 -38209 55813 -38086 8 VDD
port 41 nsew
rlabel locali s 55573 -38212 55618 -38086 8 VDD
port 41 nsew
rlabel locali s 54523 -38224 55410 -38174 8 VDD
port 41 nsew
rlabel locali s 54327 -38591 54361 -38174 8 VDD
port 41 nsew
rlabel locali s 54131 -38591 54165 -38174 8 VDD
port 41 nsew
rlabel locali s 54121 -38174 55410 -38125 8 VDD
port 41 nsew
rlabel locali s 54121 -38125 54563 -38110 8 VDD
port 41 nsew
rlabel locali s 55567 -38086 56336 -38079 8 VDD
port 41 nsew
rlabel locali s 55567 -38079 56471 -38062 8 VDD
port 41 nsew
rlabel locali s 54560 -38076 54749 -38069 8 VDD
port 41 nsew
rlabel locali s 54523 -38069 54749 -38062 8 VDD
port 41 nsew
rlabel locali s 54121 -38062 56471 -38027 8 VDD
port 41 nsew
rlabel locali s 56409 -38027 56471 -37999 8 VDD
port 41 nsew
rlabel locali s 54121 -38027 56336 -38020 8 VDD
port 41 nsew
rlabel locali s 54121 -38020 56232 -38002 8 VDD
port 41 nsew
rlabel locali s 50679 -40338 50801 -38002 8 VDD
port 41 nsew
rlabel locali s 47782 -41461 47848 -40131 8 VDD
port 41 nsew
rlabel locali s 47429 -41545 47513 -41432 8 VDD
port 41 nsew
rlabel locali s 44915 -41549 47130 -41507 8 VDD
port 41 nsew
rlabel locali s 47446 -41432 47512 -40131 8 VDD
port 41 nsew
rlabel locali s 44915 -41507 47026 -41396 8 VDD
port 41 nsew
rlabel locali s 42236 -41556 42448 -41417 8 VDD
port 41 nsew
rlabel locali s 41986 -41571 42065 -41546 8 VDD
port 41 nsew
rlabel locali s 41789 -41689 41834 -41565 8 VDD
port 41 nsew
rlabel locali s 41373 -42281 41407 -41688 8 VDD
port 41 nsew
rlabel locali s 41177 -42281 41211 -41691 8 VDD
port 41 nsew
rlabel locali s 40927 -41869 40961 -41703 8 VDD
port 41 nsew
rlabel locali s 40731 -41869 40765 -41703 8 VDD
port 41 nsew
rlabel locali s 40535 -41869 40569 -41703 8 VDD
port 41 nsew
rlabel locali s 40339 -41869 40373 -41703 8 VDD
port 41 nsew
rlabel locali s 40122 -42070 40156 -41703 8 VDD
port 41 nsew
rlabel locali s 41367 -41688 41412 -41565 8 VDD
port 41 nsew
rlabel locali s 41172 -41691 41217 -41565 8 VDD
port 41 nsew
rlabel locali s 40122 -41703 41009 -41653 8 VDD
port 41 nsew
rlabel locali s 39926 -42070 39960 -41653 8 VDD
port 41 nsew
rlabel locali s 39730 -42070 39764 -41653 8 VDD
port 41 nsew
rlabel locali s 38128 -42250 38162 -41658 8 VDD
port 41 nsew
rlabel locali s 39720 -41653 41009 -41604 8 VDD
port 41 nsew
rlabel locali s 39720 -41604 40162 -41589 8 VDD
port 41 nsew
rlabel locali s 41166 -41565 41935 -41546 8 VDD
port 41 nsew
rlabel locali s 41166 -41546 42065 -41541 8 VDD
port 41 nsew
rlabel locali s 40159 -41555 40348 -41548 8 VDD
port 41 nsew
rlabel locali s 40122 -41548 40348 -41541 8 VDD
port 41 nsew
rlabel locali s 39720 -41541 42065 -41499 8 VDD
port 41 nsew
rlabel locali s 38121 -41658 38166 -41534 8 VDD
port 41 nsew
rlabel locali s 37705 -42250 37739 -41657 8 VDD
port 41 nsew
rlabel locali s 37509 -42250 37543 -41660 8 VDD
port 41 nsew
rlabel locali s 37259 -41838 37293 -41672 8 VDD
port 41 nsew
rlabel locali s 37063 -41838 37097 -41672 8 VDD
port 41 nsew
rlabel locali s 36867 -41838 36901 -41672 8 VDD
port 41 nsew
rlabel locali s 36671 -41838 36705 -41672 8 VDD
port 41 nsew
rlabel locali s 36454 -42039 36488 -41672 8 VDD
port 41 nsew
rlabel locali s 37699 -41657 37744 -41534 8 VDD
port 41 nsew
rlabel locali s 37504 -41660 37549 -41534 8 VDD
port 41 nsew
rlabel locali s 36454 -41672 37341 -41622 8 VDD
port 41 nsew
rlabel locali s 36258 -42039 36292 -41622 8 VDD
port 41 nsew
rlabel locali s 36062 -42039 36096 -41622 8 VDD
port 41 nsew
rlabel locali s 33356 -42270 33390 -41678 8 VDD
port 41 nsew
rlabel locali s 36052 -41622 37341 -41573 8 VDD
port 41 nsew
rlabel locali s 36052 -41573 36494 -41558 8 VDD
port 41 nsew
rlabel locali s 33796 -41573 33935 -41545 8 VDD
port 41 nsew
rlabel locali s 37498 -41534 38267 -41510 8 VDD
port 41 nsew
rlabel locali s 36491 -41524 36680 -41517 8 VDD
port 41 nsew
rlabel locali s 36454 -41517 36680 -41510 8 VDD
port 41 nsew
rlabel locali s 41886 -41499 42065 -41463 8 VDD
port 41 nsew
rlabel locali s 39720 -41499 41831 -41488 8 VDD
port 41 nsew
rlabel locali s 41986 -41463 42065 -41432 8 VDD
port 41 nsew
rlabel locali s 38919 -41488 41831 -41422 8 VDD
port 41 nsew
rlabel locali s 45913 -41396 46531 -41379 8 VDD
port 41 nsew
rlabel locali s 45913 -41379 46356 -41350 8 VDD
port 41 nsew
rlabel locali s 45914 -41350 46356 -41336 8 VDD
port 41 nsew
rlabel locali s 45914 -41336 47203 -41287 8 VDD
port 41 nsew
rlabel locali s 46316 -41287 47203 -41237 8 VDD
port 41 nsew
rlabel locali s 47121 -41237 47155 -41071 8 VDD
port 41 nsew
rlabel locali s 46925 -41237 46959 -41071 8 VDD
port 41 nsew
rlabel locali s 46729 -41237 46763 -41071 8 VDD
port 41 nsew
rlabel locali s 46533 -41237 46567 -41071 8 VDD
port 41 nsew
rlabel locali s 46316 -41237 46350 -40870 8 VDD
port 41 nsew
rlabel locali s 46120 -41287 46154 -40870 8 VDD
port 41 nsew
rlabel locali s 45924 -41287 45958 -40870 8 VDD
port 41 nsew
rlabel locali s 45085 -41396 45257 -41206 8 VDD
port 41 nsew
rlabel locali s 44903 -41206 45621 -41107 8 VDD
port 41 nsew
rlabel locali s 45539 -41107 45573 -40841 8 VDD
port 41 nsew
rlabel locali s 45343 -41107 45377 -40841 8 VDD
port 41 nsew
rlabel locali s 45147 -41107 45181 -40841 8 VDD
port 41 nsew
rlabel locali s 44951 -41107 44985 -40841 8 VDD
port 41 nsew
rlabel locali s 42326 -41417 42448 -40421 8 VDD
port 41 nsew
rlabel locali s 39720 -41422 41831 -41388 8 VDD
port 41 nsew
rlabel locali s 40718 -41388 41336 -41371 8 VDD
port 41 nsew
rlabel locali s 40718 -41371 41161 -41342 8 VDD
port 41 nsew
rlabel locali s 40719 -41342 41161 -41328 8 VDD
port 41 nsew
rlabel locali s 40719 -41328 42008 -41279 8 VDD
port 41 nsew
rlabel locali s 41121 -41279 42008 -41229 8 VDD
port 41 nsew
rlabel locali s 41926 -41229 41960 -41063 8 VDD
port 41 nsew
rlabel locali s 41730 -41229 41764 -41063 8 VDD
port 41 nsew
rlabel locali s 41534 -41229 41568 -41063 8 VDD
port 41 nsew
rlabel locali s 41338 -41229 41372 -41063 8 VDD
port 41 nsew
rlabel locali s 41121 -41229 41155 -40862 8 VDD
port 41 nsew
rlabel locali s 40925 -41279 40959 -40862 8 VDD
port 41 nsew
rlabel locali s 40729 -41279 40763 -40862 8 VDD
port 41 nsew
rlabel locali s 39890 -41388 40062 -41198 8 VDD
port 41 nsew
rlabel locali s 39708 -41198 40426 -41099 8 VDD
port 41 nsew
rlabel locali s 40344 -41099 40378 -40833 8 VDD
port 41 nsew
rlabel locali s 40148 -41099 40182 -40833 8 VDD
port 41 nsew
rlabel locali s 39952 -41099 39986 -40833 8 VDD
port 41 nsew
rlabel locali s 39756 -41099 39790 -40833 8 VDD
port 41 nsew
rlabel locali s 41816 -40421 42448 -40299 8 VDD
port 41 nsew
rlabel locali s 47446 -40131 47848 -40065 8 VDD
port 41 nsew
rlabel locali s 49717 -38394 49751 -38102 8 VDD
port 41 nsew
rlabel locali s 49521 -38394 49555 -38104 8 VDD
port 41 nsew
rlabel locali s 49293 -38594 49327 -38119 8 VDD
port 41 nsew
rlabel locali s 49163 -38594 49197 -38122 8 VDD
port 41 nsew
rlabel locali s 49712 -38102 49755 -38002 8 VDD
port 41 nsew
rlabel locali s 57200 -37982 57317 -37972 8 VDD
port 41 nsew
rlabel locali s 56637 -37982 56735 -37979 8 VDD
port 41 nsew
rlabel locali s 57200 -37972 57605 -37908 8 VDD
port 41 nsew
rlabel locali s 49712 -38002 56232 -37942 8 VDD
port 41 nsew
rlabel locali s 49515 -38104 49558 -37942 8 VDD
port 41 nsew
rlabel locali s 49284 -38119 49334 -37942 8 VDD
port 41 nsew
rlabel locali s 49158 -38122 49208 -37942 8 VDD
port 41 nsew
rlabel locali s 48568 -38594 48602 -38099 8 VDD
port 41 nsew
rlabel locali s 48372 -38594 48406 -38101 8 VDD
port 41 nsew
rlabel locali s 46999 -38836 47033 -38244 8 VDD
port 41 nsew
rlabel locali s 47439 -38139 47537 -38133 8 VDD
port 41 nsew
rlabel locali s 48566 -38099 48604 -37942 8 VDD
port 41 nsew
rlabel locali s 48369 -38101 48407 -38006 8 VDD
port 41 nsew
rlabel locali s 47439 -38133 48119 -38016 8 VDD
port 41 nsew
rlabel locali s 47211 -38127 47273 -38113 8 VDD
port 41 nsew
rlabel locali s 46992 -38244 47037 -38120 8 VDD
port 41 nsew
rlabel locali s 46576 -38836 46610 -38243 8 VDD
port 41 nsew
rlabel locali s 46380 -38836 46414 -38246 8 VDD
port 41 nsew
rlabel locali s 46130 -38424 46164 -38258 8 VDD
port 41 nsew
rlabel locali s 45934 -38424 45968 -38258 8 VDD
port 41 nsew
rlabel locali s 45738 -38424 45772 -38258 8 VDD
port 41 nsew
rlabel locali s 45542 -38424 45576 -38258 8 VDD
port 41 nsew
rlabel locali s 45325 -38625 45359 -38258 8 VDD
port 41 nsew
rlabel locali s 46570 -38243 46615 -38120 8 VDD
port 41 nsew
rlabel locali s 46375 -38246 46420 -38120 8 VDD
port 41 nsew
rlabel locali s 45325 -38258 46212 -38208 8 VDD
port 41 nsew
rlabel locali s 45129 -38625 45163 -38208 8 VDD
port 41 nsew
rlabel locali s 44933 -38625 44967 -38208 8 VDD
port 41 nsew
rlabel locali s 44923 -38208 46212 -38159 8 VDD
port 41 nsew
rlabel locali s 44923 -38159 45365 -38144 8 VDD
port 41 nsew
rlabel locali s 46369 -38120 47138 -38113 8 VDD
port 41 nsew
rlabel locali s 46369 -38113 47273 -38096 8 VDD
port 41 nsew
rlabel locali s 45362 -38110 45551 -38103 8 VDD
port 41 nsew
rlabel locali s 45325 -38103 45551 -38096 8 VDD
port 41 nsew
rlabel locali s 44923 -38096 47273 -38061 8 VDD
port 41 nsew
rlabel locali s 47211 -38061 47273 -38033 8 VDD
port 41 nsew
rlabel locali s 44923 -38061 47138 -38054 8 VDD
port 41 nsew
rlabel locali s 48002 -38016 48119 -38006 8 VDD
port 41 nsew
rlabel locali s 47439 -38016 47537 -38013 8 VDD
port 41 nsew
rlabel locali s 48002 -38006 48407 -37942 8 VDD
port 41 nsew
rlabel locali s 44923 -38054 47034 -37992 8 VDD
port 41 nsew
rlabel locali s 41816 -40299 41938 -37992 8 VDD
port 41 nsew
rlabel locali s 38919 -41422 38985 -40092 8 VDD
port 41 nsew
rlabel locali s 38566 -41506 38650 -41393 8 VDD
port 41 nsew
rlabel locali s 36052 -41510 38267 -41468 8 VDD
port 41 nsew
rlabel locali s 38583 -41393 38649 -40092 8 VDD
port 41 nsew
rlabel locali s 36052 -41468 38163 -41357 8 VDD
port 41 nsew
rlabel locali s 33796 -41545 34008 -41406 8 VDD
port 41 nsew
rlabel locali s 33546 -41560 33625 -41535 8 VDD
port 41 nsew
rlabel locali s 33349 -41678 33394 -41554 8 VDD
port 41 nsew
rlabel locali s 32933 -42270 32967 -41677 8 VDD
port 41 nsew
rlabel locali s 32737 -42270 32771 -41680 8 VDD
port 41 nsew
rlabel locali s 32487 -41858 32521 -41692 8 VDD
port 41 nsew
rlabel locali s 32291 -41858 32325 -41692 8 VDD
port 41 nsew
rlabel locali s 32095 -41858 32129 -41692 8 VDD
port 41 nsew
rlabel locali s 31899 -41858 31933 -41692 8 VDD
port 41 nsew
rlabel locali s 31682 -42059 31716 -41692 8 VDD
port 41 nsew
rlabel locali s 32927 -41677 32972 -41554 8 VDD
port 41 nsew
rlabel locali s 32732 -41680 32777 -41554 8 VDD
port 41 nsew
rlabel locali s 31682 -41692 32569 -41642 8 VDD
port 41 nsew
rlabel locali s 31486 -42059 31520 -41642 8 VDD
port 41 nsew
rlabel locali s 31290 -42059 31324 -41642 8 VDD
port 41 nsew
rlabel locali s 29688 -42239 29722 -41647 8 VDD
port 41 nsew
rlabel locali s 31280 -41642 32569 -41593 8 VDD
port 41 nsew
rlabel locali s 31280 -41593 31722 -41578 8 VDD
port 41 nsew
rlabel locali s 32726 -41554 33495 -41535 8 VDD
port 41 nsew
rlabel locali s 32726 -41535 33625 -41530 8 VDD
port 41 nsew
rlabel locali s 31719 -41544 31908 -41537 8 VDD
port 41 nsew
rlabel locali s 31682 -41537 31908 -41530 8 VDD
port 41 nsew
rlabel locali s 31280 -41530 33625 -41488 8 VDD
port 41 nsew
rlabel locali s 29681 -41647 29726 -41523 8 VDD
port 41 nsew
rlabel locali s 29265 -42239 29299 -41646 8 VDD
port 41 nsew
rlabel locali s 29069 -42239 29103 -41649 8 VDD
port 41 nsew
rlabel locali s 17279 -43856 17368 -42161 8 VDD
port 41 nsew
rlabel locali s 17085 -43856 17119 -43565 8 VDD
port 41 nsew
rlabel locali s 16889 -43856 16923 -43565 8 VDD
port 41 nsew
rlabel locali s 16693 -43856 16727 -43565 8 VDD
port 41 nsew
rlabel locali s 16248 -43856 16282 -43565 8 VDD
port 41 nsew
rlabel locali s 16052 -43856 16086 -43565 8 VDD
port 41 nsew
rlabel locali s 15856 -43856 15890 -43565 8 VDD
port 41 nsew
rlabel locali s 14385 -43856 14419 -43565 8 VDD
port 41 nsew
rlabel locali s 14189 -43856 14223 -43565 8 VDD
port 41 nsew
rlabel locali s 13993 -43856 14027 -43565 8 VDD
port 41 nsew
rlabel locali s 13548 -43856 13582 -43565 8 VDD
port 41 nsew
rlabel locali s 13352 -43856 13386 -43565 8 VDD
port 41 nsew
rlabel locali s 13156 -43856 13190 -43565 8 VDD
port 41 nsew
rlabel locali s 8040 -43918 8074 -43728 8 VDD
port 41 nsew
rlabel locali s 7838 -44040 7884 -43906 8 VDD
port 41 nsew
rlabel locali s 7725 -44040 7771 -43916 8 VDD
port 41 nsew
rlabel locali s 7844 -43906 7878 -43728 8 VDD
port 41 nsew
rlabel locali s 7731 -43916 7765 -43728 8 VDD
port 41 nsew
rlabel locali s 7529 -44040 7575 -43911 8 VDD
port 41 nsew
rlabel locali s 7416 -44040 7462 -43915 8 VDD
port 41 nsew
rlabel locali s 7535 -43911 7569 -43728 8 VDD
port 41 nsew
rlabel locali s 7421 -43915 7455 -43728 8 VDD
port 41 nsew
rlabel locali s 7218 -44040 7264 -43911 8 VDD
port 41 nsew
rlabel locali s 7029 -44040 7069 -43911 8 VDD
port 41 nsew
rlabel locali s 4029 -44109 5081 -44040 8 VDD
port 41 nsew
rlabel locali s 5035 -44040 5081 -43918 8 VDD
port 41 nsew
rlabel locali s 7225 -43911 7259 -43728 8 VDD
port 41 nsew
rlabel locali s 7029 -43911 7063 -43728 8 VDD
port 41 nsew
rlabel locali s 5040 -43918 5074 -43728 8 VDD
port 41 nsew
rlabel locali s 4838 -44040 4884 -43906 8 VDD
port 41 nsew
rlabel locali s 4725 -44040 4771 -43916 8 VDD
port 41 nsew
rlabel locali s 4844 -43906 4878 -43728 8 VDD
port 41 nsew
rlabel locali s 4731 -43916 4765 -43728 8 VDD
port 41 nsew
rlabel locali s 4529 -44040 4575 -43911 8 VDD
port 41 nsew
rlabel locali s 4416 -44040 4462 -43915 8 VDD
port 41 nsew
rlabel locali s 4535 -43911 4569 -43728 8 VDD
port 41 nsew
rlabel locali s 4421 -43915 4455 -43728 8 VDD
port 41 nsew
rlabel locali s 4218 -44040 4264 -43911 8 VDD
port 41 nsew
rlabel locali s 4029 -44040 4069 -43911 8 VDD
port 41 nsew
rlabel locali s 1529 -44109 2581 -44040 8 VDD
port 41 nsew
rlabel locali s 2535 -44040 2581 -43918 8 VDD
port 41 nsew
rlabel locali s 4225 -43911 4259 -43728 8 VDD
port 41 nsew
rlabel locali s 4029 -43911 4063 -43728 8 VDD
port 41 nsew
rlabel locali s 2540 -43918 2574 -43728 8 VDD
port 41 nsew
rlabel locali s 2338 -44040 2384 -43906 8 VDD
port 41 nsew
rlabel locali s 2225 -44040 2271 -43916 8 VDD
port 41 nsew
rlabel locali s 2344 -43906 2378 -43728 8 VDD
port 41 nsew
rlabel locali s 2231 -43916 2265 -43728 8 VDD
port 41 nsew
rlabel locali s 2029 -44040 2075 -43911 8 VDD
port 41 nsew
rlabel locali s 1916 -44040 1962 -43915 8 VDD
port 41 nsew
rlabel locali s 2035 -43911 2069 -43728 8 VDD
port 41 nsew
rlabel locali s 1921 -43915 1955 -43728 8 VDD
port 41 nsew
rlabel locali s 1718 -44040 1764 -43911 8 VDD
port 41 nsew
rlabel locali s 1529 -44040 1569 -43911 8 VDD
port 41 nsew
rlabel locali s 1725 -43911 1759 -43728 8 VDD
port 41 nsew
rlabel locali s 1529 -43911 1563 -43728 8 VDD
port 41 nsew
rlabel locali s 406 -44147 521 -43275 8 VDD
port 41 nsew
rlabel locali s -641 -44147 -48 -44109 2 VDD
port 41 nsew
rlabel locali s -971 -44109 81 -44040 2 VDD
port 41 nsew
rlabel locali s 35 -44040 81 -43918 8 VDD
port 41 nsew
rlabel locali s 40 -43918 74 -43728 8 VDD
port 41 nsew
rlabel locali s -162 -44040 -116 -43906 2 VDD
port 41 nsew
rlabel locali s -275 -44040 -229 -43916 2 VDD
port 41 nsew
rlabel locali s -156 -43906 -122 -43728 2 VDD
port 41 nsew
rlabel locali s -269 -43916 -235 -43728 2 VDD
port 41 nsew
rlabel locali s -471 -44040 -425 -43911 2 VDD
port 41 nsew
rlabel locali s -584 -44040 -538 -43915 2 VDD
port 41 nsew
rlabel locali s -465 -43911 -431 -43728 2 VDD
port 41 nsew
rlabel locali s -579 -43915 -545 -43728 2 VDD
port 41 nsew
rlabel locali s -782 -44040 -736 -43911 2 VDD
port 41 nsew
rlabel locali s -971 -44040 -931 -43911 2 VDD
port 41 nsew
rlabel locali s -775 -43911 -741 -43728 2 VDD
port 41 nsew
rlabel locali s -971 -43911 -937 -43728 2 VDD
port 41 nsew
rlabel locali s -2076 -44147 -1962 -43275 2 VDD
port 41 nsew
rlabel locali s -3157 -44147 -2564 -44109 2 VDD
port 41 nsew
rlabel locali s -3471 -44109 -2419 -44040 2 VDD
port 41 nsew
rlabel locali s -2465 -44040 -2419 -43918 2 VDD
port 41 nsew
rlabel locali s -2460 -43918 -2426 -43728 2 VDD
port 41 nsew
rlabel locali s -2662 -44040 -2616 -43906 2 VDD
port 41 nsew
rlabel locali s -2775 -44040 -2729 -43916 2 VDD
port 41 nsew
rlabel locali s -2656 -43906 -2622 -43728 2 VDD
port 41 nsew
rlabel locali s -2769 -43916 -2735 -43728 2 VDD
port 41 nsew
rlabel locali s -2971 -44040 -2925 -43911 2 VDD
port 41 nsew
rlabel locali s -3084 -44040 -3038 -43915 2 VDD
port 41 nsew
rlabel locali s -2965 -43911 -2931 -43728 2 VDD
port 41 nsew
rlabel locali s -3079 -43915 -3045 -43728 2 VDD
port 41 nsew
rlabel locali s -3282 -44040 -3236 -43911 2 VDD
port 41 nsew
rlabel locali s -3471 -44040 -3431 -43911 2 VDD
port 41 nsew
rlabel locali s -3275 -43911 -3241 -43728 2 VDD
port 41 nsew
rlabel locali s -3471 -43911 -3437 -43728 2 VDD
port 41 nsew
rlabel locali s -4644 -44147 -4529 -43310 2 VDD
port 41 nsew
rlabel locali s -5971 -44147 -4919 -44040 2 VDD
port 41 nsew
rlabel locali s -22265 -44173 -19475 -44106 2 VDD
port 41 nsew
rlabel locali s -22077 -44106 -19475 -44090 2 VDD
port 41 nsew
rlabel locali s -4965 -44040 -4919 -43918 2 VDD
port 41 nsew
rlabel locali s -4960 -43918 -4926 -43728 2 VDD
port 41 nsew
rlabel locali s -5162 -44040 -5116 -43906 2 VDD
port 41 nsew
rlabel locali s -5275 -44040 -5229 -43916 2 VDD
port 41 nsew
rlabel locali s -5156 -43906 -5122 -43728 2 VDD
port 41 nsew
rlabel locali s -5269 -43916 -5235 -43728 2 VDD
port 41 nsew
rlabel locali s -5471 -44040 -5425 -43911 2 VDD
port 41 nsew
rlabel locali s -5584 -44040 -5538 -43915 2 VDD
port 41 nsew
rlabel locali s -5465 -43911 -5431 -43728 2 VDD
port 41 nsew
rlabel locali s -5579 -43915 -5545 -43728 2 VDD
port 41 nsew
rlabel locali s -5782 -44040 -5736 -43911 2 VDD
port 41 nsew
rlabel locali s -5971 -44040 -5931 -43911 2 VDD
port 41 nsew
rlabel locali s -5775 -43911 -5741 -43728 2 VDD
port 41 nsew
rlabel locali s -5971 -43911 -5937 -43728 2 VDD
port 41 nsew
rlabel locali s -20929 -44090 -20895 -43814 2 VDD
port 41 nsew
rlabel locali s -21125 -44090 -21091 -43814 2 VDD
port 41 nsew
rlabel locali s -21321 -44090 -21287 -43814 2 VDD
port 41 nsew
rlabel locali s -21517 -44090 -21483 -43814 2 VDD
port 41 nsew
rlabel locali s -22059 -44090 -22025 -43814 2 VDD
port 41 nsew
rlabel locali s -22255 -44106 -22221 -43814 2 VDD
port 41 nsew
rlabel locali s -19651 -43638 -19475 -43551 2 VDD
port 41 nsew
rlabel locali s 401 -43275 524 -43139 8 VDD
port 41 nsew
rlabel locali s -2082 -43275 -1959 -43139 2 VDD
port 41 nsew
rlabel locali s -4649 -43310 -4526 -43174 2 VDD
port 41 nsew
rlabel locali s 400 -42722 523 -42721 8 VDD
port 41 nsew
rlabel locali s 400 -42721 706 -42659 8 VDD
port 41 nsew
rlabel locali s -16209 -42862 -16175 -42696 2 VDD
port 41 nsew
rlabel locali s -16405 -42862 -16371 -42696 2 VDD
port 41 nsew
rlabel locali s -16601 -42862 -16567 -42696 2 VDD
port 41 nsew
rlabel locali s -16797 -42862 -16763 -42696 2 VDD
port 41 nsew
rlabel locali s -17014 -43063 -16980 -42696 2 VDD
port 41 nsew
rlabel locali s 16987 -42455 17021 -42164 8 VDD
port 41 nsew
rlabel locali s 16791 -42455 16825 -42164 8 VDD
port 41 nsew
rlabel locali s 16595 -42455 16629 -42164 8 VDD
port 41 nsew
rlabel locali s 15244 -42455 15278 -42164 8 VDD
port 41 nsew
rlabel locali s 15048 -42455 15082 -42164 8 VDD
port 41 nsew
rlabel locali s 14852 -42455 14886 -42164 8 VDD
port 41 nsew
rlabel locali s 14287 -42455 14321 -42164 8 VDD
port 41 nsew
rlabel locali s 14091 -42455 14125 -42164 8 VDD
port 41 nsew
rlabel locali s 13895 -42455 13929 -42164 8 VDD
port 41 nsew
rlabel locali s 12544 -42455 12578 -42164 8 VDD
port 41 nsew
rlabel locali s 12348 -42455 12382 -42164 8 VDD
port 41 nsew
rlabel locali s 12152 -42455 12186 -42164 8 VDD
port 41 nsew
rlabel locali s 11662 -42455 11696 -42164 8 VDD
port 41 nsew
rlabel locali s 11466 -42455 11500 -42164 8 VDD
port 41 nsew
rlabel locali s 11270 -42455 11304 -42164 8 VDD
port 41 nsew
rlabel locali s 16586 -42164 17081 -42161 8 VDD
port 41 nsew
rlabel locali s 13886 -42164 15339 -42163 8 VDD
port 41 nsew
rlabel locali s 16264 -42161 17368 -42159 8 VDD
port 41 nsew
rlabel locali s 13573 -42163 15339 -42159 8 VDD
port 41 nsew
rlabel locali s 11261 -42164 12639 -42159 8 VDD
port 41 nsew
rlabel locali s 11261 -42159 17368 -42096 8 VDD
port 41 nsew
rlabel locali s 16264 -42096 17368 -42093 8 VDD
port 41 nsew
rlabel locali s 13573 -42096 14046 -42095 8 VDD
port 41 nsew
rlabel locali s 28819 -41827 28853 -41661 8 VDD
port 41 nsew
rlabel locali s 28623 -41827 28657 -41661 8 VDD
port 41 nsew
rlabel locali s 28427 -41827 28461 -41661 8 VDD
port 41 nsew
rlabel locali s 28231 -41827 28265 -41661 8 VDD
port 41 nsew
rlabel locali s 28014 -42028 28048 -41661 8 VDD
port 41 nsew
rlabel locali s 29259 -41646 29304 -41523 8 VDD
port 41 nsew
rlabel locali s 29064 -41649 29109 -41523 8 VDD
port 41 nsew
rlabel locali s 28014 -41661 28901 -41611 8 VDD
port 41 nsew
rlabel locali s 27818 -42028 27852 -41611 8 VDD
port 41 nsew
rlabel locali s 27622 -42028 27656 -41611 8 VDD
port 41 nsew
rlabel locali s 20809 -41645 20872 -41634 8 VDD
port 41 nsew
rlabel locali s 19689 -41638 19775 -41634 8 VDD
port 41 nsew
rlabel locali s 22207 -41629 25496 -41621 8 VDD
port 41 nsew
rlabel locali s 21490 -41634 21564 -41628 8 VDD
port 41 nsew
rlabel locali s 19689 -41634 20872 -41628 8 VDD
port 41 nsew
rlabel locali s 19689 -41628 21564 -41622 8 VDD
port 41 nsew
rlabel locali s 17242 -42093 17368 -41622 8 VDD
port 41 nsew
rlabel locali s 7038 -41885 7161 -41858 8 VDD
port 41 nsew
rlabel locali s 7038 -41858 8091 -41789 8 VDD
port 41 nsew
rlabel locali s 8045 -41789 8091 -41667 8 VDD
port 41 nsew
rlabel locali s 17242 -41622 21564 -41621 8 VDD
port 41 nsew
rlabel locali s 27612 -41611 28901 -41562 8 VDD
port 41 nsew
rlabel locali s 27612 -41562 28054 -41547 8 VDD
port 41 nsew
rlabel locali s 17242 -41621 25496 -41565 8 VDD
port 41 nsew
rlabel locali s 20809 -41565 25496 -41561 8 VDD
port 41 nsew
rlabel locali s 21490 -41561 25496 -41553 8 VDD
port 41 nsew
rlabel locali s 22185 -41553 25496 -41526 8 VDD
port 41 nsew
rlabel locali s 29058 -41523 29827 -41499 8 VDD
port 41 nsew
rlabel locali s 28051 -41513 28240 -41506 8 VDD
port 41 nsew
rlabel locali s 28014 -41506 28240 -41499 8 VDD
port 41 nsew
rlabel locali s 33446 -41488 33625 -41452 8 VDD
port 41 nsew
rlabel locali s 31280 -41488 33391 -41477 8 VDD
port 41 nsew
rlabel locali s 33546 -41452 33625 -41421 8 VDD
port 41 nsew
rlabel locali s 30479 -41477 33391 -41411 8 VDD
port 41 nsew
rlabel locali s 37050 -41357 37668 -41340 8 VDD
port 41 nsew
rlabel locali s 37050 -41340 37493 -41311 8 VDD
port 41 nsew
rlabel locali s 37051 -41311 37493 -41297 8 VDD
port 41 nsew
rlabel locali s 37051 -41297 38340 -41248 8 VDD
port 41 nsew
rlabel locali s 37453 -41248 38340 -41198 8 VDD
port 41 nsew
rlabel locali s 38258 -41198 38292 -41032 8 VDD
port 41 nsew
rlabel locali s 38062 -41198 38096 -41032 8 VDD
port 41 nsew
rlabel locali s 37866 -41198 37900 -41032 8 VDD
port 41 nsew
rlabel locali s 37670 -41198 37704 -41032 8 VDD
port 41 nsew
rlabel locali s 37453 -41198 37487 -40831 8 VDD
port 41 nsew
rlabel locali s 37257 -41248 37291 -40831 8 VDD
port 41 nsew
rlabel locali s 37061 -41248 37095 -40831 8 VDD
port 41 nsew
rlabel locali s 36222 -41357 36394 -41167 8 VDD
port 41 nsew
rlabel locali s 36040 -41167 36758 -41068 8 VDD
port 41 nsew
rlabel locali s 36676 -41068 36710 -40802 8 VDD
port 41 nsew
rlabel locali s 36480 -41068 36514 -40802 8 VDD
port 41 nsew
rlabel locali s 36284 -41068 36318 -40802 8 VDD
port 41 nsew
rlabel locali s 36088 -41068 36122 -40802 8 VDD
port 41 nsew
rlabel locali s 33886 -41406 34008 -40410 8 VDD
port 41 nsew
rlabel locali s 31280 -41411 33391 -41377 8 VDD
port 41 nsew
rlabel locali s 32278 -41377 32896 -41360 8 VDD
port 41 nsew
rlabel locali s 32278 -41360 32721 -41331 8 VDD
port 41 nsew
rlabel locali s 32279 -41331 32721 -41317 8 VDD
port 41 nsew
rlabel locali s 32279 -41317 33568 -41268 8 VDD
port 41 nsew
rlabel locali s 32681 -41268 33568 -41218 8 VDD
port 41 nsew
rlabel locali s 33486 -41218 33520 -41052 8 VDD
port 41 nsew
rlabel locali s 33290 -41218 33324 -41052 8 VDD
port 41 nsew
rlabel locali s 33094 -41218 33128 -41052 8 VDD
port 41 nsew
rlabel locali s 32898 -41218 32932 -41052 8 VDD
port 41 nsew
rlabel locali s 32681 -41218 32715 -40851 8 VDD
port 41 nsew
rlabel locali s 32485 -41268 32519 -40851 8 VDD
port 41 nsew
rlabel locali s 32289 -41268 32323 -40851 8 VDD
port 41 nsew
rlabel locali s 31450 -41377 31622 -41187 8 VDD
port 41 nsew
rlabel locali s 31268 -41187 31986 -41088 8 VDD
port 41 nsew
rlabel locali s 31904 -41088 31938 -40822 8 VDD
port 41 nsew
rlabel locali s 31708 -41088 31742 -40822 8 VDD
port 41 nsew
rlabel locali s 31512 -41088 31546 -40822 8 VDD
port 41 nsew
rlabel locali s 31316 -41088 31350 -40822 8 VDD
port 41 nsew
rlabel locali s 33376 -40410 34008 -40288 8 VDD
port 41 nsew
rlabel locali s 38583 -40092 38985 -40026 8 VDD
port 41 nsew
rlabel locali s 40854 -38355 40888 -38063 8 VDD
port 41 nsew
rlabel locali s 40658 -38355 40692 -38065 8 VDD
port 41 nsew
rlabel locali s 40430 -38555 40464 -38080 8 VDD
port 41 nsew
rlabel locali s 40300 -38555 40334 -38083 8 VDD
port 41 nsew
rlabel locali s 40849 -38063 40892 -37992 8 VDD
port 41 nsew
rlabel locali s 40849 -37992 47034 -37943 8 VDD
port 41 nsew
rlabel locali s 48002 -37942 56232 -37909 8 VDD
port 41 nsew
rlabel locali s 45921 -37943 46539 -37926 8 VDD
port 41 nsew
rlabel locali s 57200 -37908 64986 -37855 8 VDD
port 41 nsew
rlabel locali s 55119 -37909 55737 -37892 8 VDD
port 41 nsew
rlabel locali s 55119 -37892 55562 -37863 8 VDD
port 41 nsew
rlabel locali s 48002 -37909 54463 -37889 8 VDD
port 41 nsew
rlabel locali s 45921 -37926 46364 -37897 8 VDD
port 41 nsew
rlabel locali s 40849 -37943 45265 -37903 8 VDD
port 41 nsew
rlabel locali s 40652 -38065 40695 -37903 8 VDD
port 41 nsew
rlabel locali s 40421 -38080 40471 -37903 8 VDD
port 41 nsew
rlabel locali s 40295 -38083 40345 -37903 8 VDD
port 41 nsew
rlabel locali s 39705 -38555 39739 -38060 8 VDD
port 41 nsew
rlabel locali s 39509 -38555 39543 -38062 8 VDD
port 41 nsew
rlabel locali s 38136 -38797 38170 -38205 8 VDD
port 41 nsew
rlabel locali s 38576 -38100 38674 -38094 8 VDD
port 41 nsew
rlabel locali s 39703 -38060 39741 -37903 8 VDD
port 41 nsew
rlabel locali s 39506 -38062 39544 -37967 8 VDD
port 41 nsew
rlabel locali s 38576 -38094 39256 -37977 8 VDD
port 41 nsew
rlabel locali s 38348 -38088 38410 -38074 8 VDD
port 41 nsew
rlabel locali s 38129 -38205 38174 -38081 8 VDD
port 41 nsew
rlabel locali s 37713 -38797 37747 -38204 8 VDD
port 41 nsew
rlabel locali s 37517 -38797 37551 -38207 8 VDD
port 41 nsew
rlabel locali s 37267 -38385 37301 -38219 8 VDD
port 41 nsew
rlabel locali s 37071 -38385 37105 -38219 8 VDD
port 41 nsew
rlabel locali s 36875 -38385 36909 -38219 8 VDD
port 41 nsew
rlabel locali s 36679 -38385 36713 -38219 8 VDD
port 41 nsew
rlabel locali s 36462 -38586 36496 -38219 8 VDD
port 41 nsew
rlabel locali s 37707 -38204 37752 -38081 8 VDD
port 41 nsew
rlabel locali s 37512 -38207 37557 -38081 8 VDD
port 41 nsew
rlabel locali s 36462 -38219 37349 -38169 8 VDD
port 41 nsew
rlabel locali s 36266 -38586 36300 -38169 8 VDD
port 41 nsew
rlabel locali s 36070 -38586 36104 -38169 8 VDD
port 41 nsew
rlabel locali s 36060 -38169 37349 -38120 8 VDD
port 41 nsew
rlabel locali s 36060 -38120 36502 -38105 8 VDD
port 41 nsew
rlabel locali s 37506 -38081 38275 -38074 8 VDD
port 41 nsew
rlabel locali s 37506 -38074 38410 -38057 8 VDD
port 41 nsew
rlabel locali s 36499 -38071 36688 -38064 8 VDD
port 41 nsew
rlabel locali s 36462 -38064 36688 -38057 8 VDD
port 41 nsew
rlabel locali s 33376 -40288 33498 -38057 8 VDD
port 41 nsew
rlabel locali s 30479 -41411 30545 -40081 8 VDD
port 41 nsew
rlabel locali s 30126 -41495 30210 -41382 8 VDD
port 41 nsew
rlabel locali s 27612 -41499 29827 -41457 8 VDD
port 41 nsew
rlabel locali s 30143 -41382 30209 -40081 8 VDD
port 41 nsew
rlabel locali s 27612 -41457 29723 -41346 8 VDD
port 41 nsew
rlabel locali s 28610 -41346 29228 -41329 8 VDD
port 41 nsew
rlabel locali s 28610 -41329 29053 -41300 8 VDD
port 41 nsew
rlabel locali s 28611 -41300 29053 -41286 8 VDD
port 41 nsew
rlabel locali s 28611 -41286 29900 -41237 8 VDD
port 41 nsew
rlabel locali s 29013 -41237 29900 -41187 8 VDD
port 41 nsew
rlabel locali s 29818 -41187 29852 -41021 8 VDD
port 41 nsew
rlabel locali s 29622 -41187 29656 -41021 8 VDD
port 41 nsew
rlabel locali s 29426 -41187 29460 -41021 8 VDD
port 41 nsew
rlabel locali s 29230 -41187 29264 -41021 8 VDD
port 41 nsew
rlabel locali s 29013 -41187 29047 -40820 8 VDD
port 41 nsew
rlabel locali s 28817 -41237 28851 -40820 8 VDD
port 41 nsew
rlabel locali s 28621 -41237 28655 -40820 8 VDD
port 41 nsew
rlabel locali s 27782 -41346 27954 -41156 8 VDD
port 41 nsew
rlabel locali s 27600 -41156 28318 -41057 8 VDD
port 41 nsew
rlabel locali s 28236 -41057 28270 -40791 8 VDD
port 41 nsew
rlabel locali s 28040 -41057 28074 -40791 8 VDD
port 41 nsew
rlabel locali s 27844 -41057 27878 -40791 8 VDD
port 41 nsew
rlabel locali s 27648 -41057 27682 -40791 8 VDD
port 41 nsew
rlabel locali s 30143 -40081 30545 -40015 8 VDD
port 41 nsew
rlabel locali s 25407 -41526 25496 -39371 8 VDD
port 41 nsew
rlabel locali s 25269 -41526 25303 -40691 8 VDD
port 41 nsew
rlabel locali s 25073 -41526 25107 -40691 8 VDD
port 41 nsew
rlabel locali s 24869 -41526 24903 -40691 8 VDD
port 41 nsew
rlabel locali s 24673 -41526 24707 -40691 8 VDD
port 41 nsew
rlabel locali s 24269 -41526 24303 -40691 8 VDD
port 41 nsew
rlabel locali s 24073 -41526 24107 -40691 8 VDD
port 41 nsew
rlabel locali s 23869 -41526 23903 -40691 8 VDD
port 41 nsew
rlabel locali s 23673 -41526 23707 -40691 8 VDD
port 41 nsew
rlabel locali s 23269 -41526 23303 -40691 8 VDD
port 41 nsew
rlabel locali s 23073 -41526 23107 -40691 8 VDD
port 41 nsew
rlabel locali s 22869 -41526 22903 -40691 8 VDD
port 41 nsew
rlabel locali s 22673 -41526 22707 -40691 8 VDD
port 41 nsew
rlabel locali s 22185 -41526 22219 -41262 8 VDD
port 41 nsew
rlabel locali s 21989 -41553 22023 -41262 8 VDD
port 41 nsew
rlabel locali s 21793 -41553 21827 -41262 8 VDD
port 41 nsew
rlabel locali s 21490 -41553 21564 -41547 8 VDD
port 41 nsew
rlabel locali s 21260 -41561 21294 -41269 8 VDD
port 41 nsew
rlabel locali s 21064 -41561 21098 -41269 8 VDD
port 41 nsew
rlabel locali s 20809 -41561 20872 -41547 8 VDD
port 41 nsew
rlabel locali s 20522 -41565 20556 -41269 8 VDD
port 41 nsew
rlabel locali s 20326 -41565 20360 -41269 8 VDD
port 41 nsew
rlabel locali s 20130 -41565 20164 -41269 8 VDD
port 41 nsew
rlabel locali s 19934 -41565 19968 -41269 8 VDD
port 41 nsew
rlabel locali s 17242 -41565 19775 -41553 8 VDD
port 41 nsew
rlabel locali s 19689 -41553 19775 -41545 8 VDD
port 41 nsew
rlabel locali s 19208 -41553 19256 -41420 8 VDD
port 41 nsew
rlabel locali s 19011 -41553 19059 -41426 8 VDD
port 41 nsew
rlabel locali s 19214 -41420 19248 -41035 8 VDD
port 41 nsew
rlabel locali s 19018 -41426 19052 -41035 8 VDD
port 41 nsew
rlabel locali s 18262 -41553 18310 -41420 8 VDD
port 41 nsew
rlabel locali s 18065 -41553 18113 -41426 8 VDD
port 41 nsew
rlabel locali s 8050 -41667 8084 -41477 8 VDD
port 41 nsew
rlabel locali s 7848 -41789 7894 -41655 8 VDD
port 41 nsew
rlabel locali s 7735 -41789 7781 -41665 8 VDD
port 41 nsew
rlabel locali s 7854 -41655 7888 -41477 8 VDD
port 41 nsew
rlabel locali s 7741 -41665 7775 -41477 8 VDD
port 41 nsew
rlabel locali s 7539 -41789 7585 -41660 8 VDD
port 41 nsew
rlabel locali s 7426 -41789 7472 -41664 8 VDD
port 41 nsew
rlabel locali s 7545 -41660 7579 -41477 8 VDD
port 41 nsew
rlabel locali s 7431 -41664 7465 -41477 8 VDD
port 41 nsew
rlabel locali s 7228 -41789 7274 -41660 8 VDD
port 41 nsew
rlabel locali s 7038 -41789 7161 -41749 8 VDD
port 41 nsew
rlabel locali s 5822 -41886 5945 -41853 8 VDD
port 41 nsew
rlabel locali s 4466 -41891 4589 -41858 8 VDD
port 41 nsew
rlabel locali s 4466 -41858 5362 -41853 8 VDD
port 41 nsew
rlabel locali s 4466 -41853 5945 -41785 8 VDD
port 41 nsew
rlabel locali s 5290 -41785 5945 -41784 8 VDD
port 41 nsew
rlabel locali s 5822 -41784 5945 -41750 8 VDD
port 41 nsew
rlabel locali s 7039 -41749 7079 -41660 8 VDD
port 41 nsew
rlabel locali s 7235 -41660 7269 -41477 8 VDD
port 41 nsew
rlabel locali s 7039 -41660 7073 -41477 8 VDD
port 41 nsew
rlabel locali s 5878 -41750 5912 -41488 8 VDD
port 41 nsew
rlabel locali s 5682 -41784 5716 -41488 8 VDD
port 41 nsew
rlabel locali s 5486 -41784 5520 -41488 8 VDD
port 41 nsew
rlabel locali s 5290 -41784 5324 -41488 8 VDD
port 41 nsew
rlabel locali s 4466 -41785 4787 -41780 8 VDD
port 41 nsew
rlabel locali s 4748 -41780 4782 -41488 8 VDD
port 41 nsew
rlabel locali s 4466 -41780 4589 -41755 8 VDD
port 41 nsew
rlabel locali s 4065 -41889 4188 -41844 8 VDD
port 41 nsew
rlabel locali s 3727 -41844 4188 -41829 8 VDD
port 41 nsew
rlabel locali s 2837 -41866 2960 -41829 8 VDD
port 41 nsew
rlabel locali s 2837 -41829 4188 -41780 8 VDD
port 41 nsew
rlabel locali s 4552 -41755 4586 -41488 8 VDD
port 41 nsew
rlabel locali s 4065 -41780 4188 -41753 8 VDD
port 41 nsew
rlabel locali s 18268 -41420 18302 -41035 8 VDD
port 41 nsew
rlabel locali s 18072 -41426 18106 -41035 8 VDD
port 41 nsew
rlabel locali s 4125 -41753 4159 -41363 8 VDD
port 41 nsew
rlabel locali s 3929 -41780 3963 -41363 8 VDD
port 41 nsew
rlabel locali s 2837 -41780 3767 -41730 8 VDD
port 41 nsew
rlabel locali s 2448 -41865 2571 -41851 8 VDD
port 41 nsew
rlabel locali s 405 -42659 520 -41851 8 VDD
port 41 nsew
rlabel locali s -2083 -42687 -1960 -42551 2 VDD
port 41 nsew
rlabel locali s -17014 -42696 -16127 -42646 2 VDD
port 41 nsew
rlabel locali s -17210 -43063 -17176 -42646 2 VDD
port 41 nsew
rlabel locali s -17406 -43063 -17372 -42646 2 VDD
port 41 nsew
rlabel locali s -17791 -43092 -17757 -42826 2 VDD
port 41 nsew
rlabel locali s -17987 -43092 -17953 -42826 2 VDD
port 41 nsew
rlabel locali s -18183 -43092 -18149 -42826 2 VDD
port 41 nsew
rlabel locali s -18379 -43092 -18345 -42826 2 VDD
port 41 nsew
rlabel locali s -18427 -42826 -17709 -42727 2 VDD
port 41 nsew
rlabel locali s -17416 -42646 -16127 -42597 2 VDD
port 41 nsew
rlabel locali s -17416 -42597 -16974 -42583 2 VDD
port 41 nsew
rlabel locali s -17417 -42583 -16974 -42554 2 VDD
port 41 nsew
rlabel locali s -530 -41878 -407 -41851 2 VDD
port 41 nsew
rlabel locali s -530 -41851 2571 -41772 8 VDD
port 41 nsew
rlabel locali s 3733 -41730 3767 -41363 8 VDD
port 41 nsew
rlabel locali s 3516 -41730 3550 -41564 8 VDD
port 41 nsew
rlabel locali s 3320 -41730 3354 -41564 8 VDD
port 41 nsew
rlabel locali s 3124 -41730 3158 -41564 8 VDD
port 41 nsew
rlabel locali s 2928 -41730 2962 -41564 8 VDD
port 41 nsew
rlabel locali s 2448 -41772 2571 -41729 8 VDD
port 41 nsew
rlabel locali s 2520 -41729 2554 -41365 8 VDD
port 41 nsew
rlabel locali s 2324 -41772 2358 -41365 8 VDD
port 41 nsew
rlabel locali s 1275 -41772 2162 -41732 8 VDD
port 41 nsew
rlabel locali s 2128 -41732 2162 -41365 8 VDD
port 41 nsew
rlabel locali s 1911 -41732 1945 -41566 8 VDD
port 41 nsew
rlabel locali s 1715 -41732 1749 -41566 8 VDD
port 41 nsew
rlabel locali s 1519 -41732 1553 -41566 8 VDD
port 41 nsew
rlabel locali s 1323 -41732 1357 -41566 8 VDD
port 41 nsew
rlabel locali s 916 -41772 950 -41479 8 VDD
port 41 nsew
rlabel locali s 720 -41772 754 -41479 8 VDD
port 41 nsew
rlabel locali s 524 -41772 558 -41479 8 VDD
port 41 nsew
rlabel locali s 328 -41772 362 -41479 8 VDD
port 41 nsew
rlabel locali s -530 -41772 -175 -41771 2 VDD
port 41 nsew
rlabel locali s -214 -41771 -180 -41479 2 VDD
port 41 nsew
rlabel locali s -530 -41771 -376 -41742 2 VDD
port 41 nsew
rlabel locali s -824 -41877 -701 -41855 2 VDD
port 41 nsew
rlabel locali s -2079 -42551 -1964 -41855 2 VDD
port 41 nsew
rlabel locali s -4650 -42543 -4527 -42407 2 VDD
port 41 nsew
rlabel locali s -17417 -42554 -16799 -42537 2 VDD
port 41 nsew
rlabel locali s -18245 -42727 -18073 -42556 2 VDD
port 41 nsew
rlabel locali s -19649 -43551 -19477 -42556 2 VDD
port 41 nsew
rlabel locali s -19649 -42556 -18073 -42537 2 VDD
port 41 nsew
rlabel locali s -19649 -42537 -16304 -42426 2 VDD
port 41 nsew
rlabel locali s -3494 -41856 -3021 -41855 2 VDD
port 41 nsew
rlabel locali s -4645 -42407 -4530 -41855 2 VDD
port 41 nsew
rlabel locali s -19649 -42426 -16200 -42384 2 VDD
port 41 nsew
rlabel locali s -16969 -42384 -16200 -42360 2 VDD
port 41 nsew
rlabel locali s -18013 -42384 -17787 -42377 2 VDD
port 41 nsew
rlabel locali s -17976 -42377 -17787 -42370 2 VDD
port 41 nsew
rlabel locali s -16346 -42360 -16301 -42236 2 VDD
port 41 nsew
rlabel locali s -16768 -42360 -16723 -42237 2 VDD
port 41 nsew
rlabel locali s -6816 -41858 -5712 -41855 2 VDD
port 41 nsew
rlabel locali s -6816 -41855 -701 -41792 2 VDD
port 41 nsew
rlabel locali s -2087 -41792 -701 -41787 2 VDD
port 41 nsew
rlabel locali s -4787 -41792 -3021 -41788 2 VDD
port 41 nsew
rlabel locali s -6816 -41792 -5712 -41790 2 VDD
port 41 nsew
rlabel locali s -4787 -41788 -3334 -41787 2 VDD
port 41 nsew
rlabel locali s -6529 -41790 -6034 -41787 2 VDD
port 41 nsew
rlabel locali s -410 -41742 -376 -41479 2 VDD
port 41 nsew
rlabel locali s -824 -41787 -701 -41741 2 VDD
port 41 nsew
rlabel locali s -752 -41741 -718 -41496 2 VDD
port 41 nsew
rlabel locali s -948 -41787 -914 -41496 2 VDD
port 41 nsew
rlabel locali s -1144 -41787 -1110 -41496 2 VDD
port 41 nsew
rlabel locali s -1634 -41787 -1600 -41496 2 VDD
port 41 nsew
rlabel locali s -1830 -41787 -1796 -41496 2 VDD
port 41 nsew
rlabel locali s -2026 -41787 -1992 -41496 2 VDD
port 41 nsew
rlabel locali s -3377 -41787 -3343 -41496 2 VDD
port 41 nsew
rlabel locali s -3573 -41787 -3539 -41496 2 VDD
port 41 nsew
rlabel locali s -3769 -41787 -3735 -41496 2 VDD
port 41 nsew
rlabel locali s -4334 -41787 -4300 -41496 2 VDD
port 41 nsew
rlabel locali s -4530 -41787 -4496 -41496 2 VDD
port 41 nsew
rlabel locali s -4726 -41787 -4692 -41496 2 VDD
port 41 nsew
rlabel locali s -6077 -41787 -6043 -41496 2 VDD
port 41 nsew
rlabel locali s -6273 -41787 -6239 -41496 2 VDD
port 41 nsew
rlabel locali s -6469 -41787 -6435 -41496 2 VDD
port 41 nsew
rlabel locali s 22235 -40169 22269 -39652 8 VDD
port 41 nsew
rlabel locali s 22039 -40169 22073 -39652 8 VDD
port 41 nsew
rlabel locali s 21843 -40169 21877 -39652 8 VDD
port 41 nsew
rlabel locali s -2638 -40386 -2604 -40095 2 VDD
port 41 nsew
rlabel locali s -2834 -40386 -2800 -40095 2 VDD
port 41 nsew
rlabel locali s -3030 -40386 -2996 -40095 2 VDD
port 41 nsew
rlabel locali s -3475 -40386 -3441 -40095 2 VDD
port 41 nsew
rlabel locali s -3671 -40386 -3637 -40095 2 VDD
port 41 nsew
rlabel locali s -3867 -40386 -3833 -40095 2 VDD
port 41 nsew
rlabel locali s -5338 -40386 -5304 -40095 2 VDD
port 41 nsew
rlabel locali s -5534 -40386 -5500 -40095 2 VDD
port 41 nsew
rlabel locali s -5730 -40386 -5696 -40095 2 VDD
port 41 nsew
rlabel locali s -6175 -40386 -6141 -40095 2 VDD
port 41 nsew
rlabel locali s -6371 -40386 -6337 -40095 2 VDD
port 41 nsew
rlabel locali s -6567 -40386 -6533 -40095 2 VDD
port 41 nsew
rlabel locali s -6816 -41790 -6727 -40095 2 VDD
port 41 nsew
rlabel locali s -16339 -42236 -16305 -41644 2 VDD
port 41 nsew
rlabel locali s -16762 -42237 -16728 -41644 2 VDD
port 41 nsew
rlabel locali s -16963 -42360 -16918 -42234 2 VDD
port 41 nsew
rlabel locali s -18415 -42336 -17973 -42321 2 VDD
port 41 nsew
rlabel locali s -18415 -42321 -17126 -42272 2 VDD
port 41 nsew
rlabel locali s -16958 -42234 -16924 -41644 2 VDD
port 41 nsew
rlabel locali s -18013 -42272 -17126 -42222 2 VDD
port 41 nsew
rlabel locali s -17208 -42222 -17174 -42056 2 VDD
port 41 nsew
rlabel locali s -17404 -42222 -17370 -42056 2 VDD
port 41 nsew
rlabel locali s -17600 -42222 -17566 -42056 2 VDD
port 41 nsew
rlabel locali s -17796 -42222 -17762 -42056 2 VDD
port 41 nsew
rlabel locali s -18013 -42222 -17979 -41855 2 VDD
port 41 nsew
rlabel locali s -18209 -42272 -18175 -41855 2 VDD
port 41 nsew
rlabel locali s -18405 -42272 -18371 -41855 2 VDD
port 41 nsew
rlabel locali s -11368 -41589 -10895 -41588 2 VDD
port 41 nsew
rlabel locali s -14690 -41591 -13586 -41588 2 VDD
port 41 nsew
rlabel locali s -14690 -41588 -8583 -41525 2 VDD
port 41 nsew
rlabel locali s -9961 -41525 -8583 -41520 2 VDD
port 41 nsew
rlabel locali s -12661 -41525 -10895 -41521 2 VDD
port 41 nsew
rlabel locali s -14690 -41525 -13586 -41523 2 VDD
port 41 nsew
rlabel locali s -12661 -41521 -11208 -41520 2 VDD
port 41 nsew
rlabel locali s -14403 -41523 -13908 -41520 2 VDD
port 41 nsew
rlabel locali s -8626 -41520 -8592 -41229 2 VDD
port 41 nsew
rlabel locali s -8822 -41520 -8788 -41229 2 VDD
port 41 nsew
rlabel locali s -9018 -41520 -8984 -41229 2 VDD
port 41 nsew
rlabel locali s -9508 -41520 -9474 -41229 2 VDD
port 41 nsew
rlabel locali s -9704 -41520 -9670 -41229 2 VDD
port 41 nsew
rlabel locali s -9900 -41520 -9866 -41229 2 VDD
port 41 nsew
rlabel locali s -11251 -41520 -11217 -41229 2 VDD
port 41 nsew
rlabel locali s -11447 -41520 -11413 -41229 2 VDD
port 41 nsew
rlabel locali s -11643 -41520 -11609 -41229 2 VDD
port 41 nsew
rlabel locali s -12208 -41520 -12174 -41229 2 VDD
port 41 nsew
rlabel locali s -12404 -41520 -12370 -41229 2 VDD
port 41 nsew
rlabel locali s -12600 -41520 -12566 -41229 2 VDD
port 41 nsew
rlabel locali s -13951 -41520 -13917 -41229 2 VDD
port 41 nsew
rlabel locali s -14147 -41520 -14113 -41229 2 VDD
port 41 nsew
rlabel locali s -14343 -41520 -14309 -41229 2 VDD
port 41 nsew
rlabel locali s -14690 -41523 -14601 -40620 2 VDD
port 41 nsew
rlabel locali s -19611 -41334 -19577 -40949 2 VDD
port 41 nsew
rlabel locali s -19617 -40949 -19569 -40816 2 VDD
port 41 nsew
rlabel locali s -19807 -41334 -19773 -40943 2 VDD
port 41 nsew
rlabel locali s -20516 -41333 -20482 -40948 2 VDD
port 41 nsew
rlabel locali s -19814 -40943 -19766 -40816 2 VDD
port 41 nsew
rlabel locali s -19819 -40816 -19265 -40788 2 VDD
port 41 nsew
rlabel locali s -20522 -40948 -20474 -40815 2 VDD
port 41 nsew
rlabel locali s -20712 -41333 -20678 -40942 2 VDD
port 41 nsew
rlabel locali s -21722 -41604 -21688 -41020 2 VDD
port 41 nsew
rlabel locali s -20719 -40942 -20671 -40815 2 VDD
port 41 nsew
rlabel locali s -21731 -41020 -21678 -40892 2 VDD
port 41 nsew
rlabel locali s -21918 -41604 -21884 -41004 2 VDD
port 41 nsew
rlabel locali s -25449 -41519 -25383 -41318 2 VDD
port 41 nsew
rlabel locali s -26016 -41523 -25521 -41489 2 VDD
port 41 nsew
rlabel locali s -25569 -41489 -25521 -41318 2 VDD
port 41 nsew
rlabel locali s -25569 -41318 -25383 -41287 2 VDD
port 41 nsew
rlabel locali s -26016 -41287 -25383 -41259 2 VDD
port 41 nsew
rlabel locali s -21927 -41004 -21874 -40892 2 VDD
port 41 nsew
rlabel locali s -19820 -40788 -19265 -40747 2 VDD
port 41 nsew
rlabel locali s -19820 -40747 -19267 -40620 2 VDD
port 41 nsew
rlabel locali s -20724 -40815 -20170 -40746 2 VDD
port 41 nsew
rlabel locali s -21927 -40892 -21059 -40759 2 VDD
port 41 nsew
rlabel locali s -20709 -40746 -20191 -40620 2 VDD
port 41 nsew
rlabel locali s -21867 -40759 -21085 -40620 2 VDD
port 41 nsew
rlabel locali s -25449 -41259 -25383 -40730 2 VDD
port 41 nsew
rlabel locali s -26016 -41259 -25521 -41253 2 VDD
port 41 nsew
rlabel locali s -25569 -41253 -25521 -41051 2 VDD
port 41 nsew
rlabel locali s -26016 -41051 -25521 -41017 2 VDD
port 41 nsew
rlabel locali s -25569 -41017 -25521 -40921 2 VDD
port 41 nsew
rlabel locali s -26016 -40921 -25521 -40887 2 VDD
port 41 nsew
rlabel locali s -25569 -40887 -25521 -40730 2 VDD
port 41 nsew
rlabel locali s -25569 -40730 -25383 -40685 2 VDD
port 41 nsew
rlabel locali s -26016 -40685 -25383 -40671 2 VDD
port 41 nsew
rlabel locali s -4345 -40095 -2543 -40090 2 VDD
port 41 nsew
rlabel locali s -6816 -40095 -5243 -40090 2 VDD
port 41 nsew
rlabel locali s -6816 -40090 -1591 -40027 2 VDD
port 41 nsew
rlabel locali s 21833 -39652 22275 -39588 8 VDD
port 41 nsew
rlabel locali s 24392 -39371 25496 -39368 8 VDD
port 41 nsew
rlabel locali s 21891 -39588 22123 -39369 8 VDD
port 41 nsew
rlabel locali s 21701 -39369 22174 -39368 8 VDD
port 41 nsew
rlabel locali s 19389 -39368 25496 -39305 8 VDD
port 41 nsew
rlabel locali s 24392 -39305 25496 -39303 8 VDD
port 41 nsew
rlabel locali s 33376 -38057 38410 -38022 8 VDD
port 41 nsew
rlabel locali s 32414 -38344 32448 -38052 8 VDD
port 41 nsew
rlabel locali s 32218 -38344 32252 -38054 8 VDD
port 41 nsew
rlabel locali s 31990 -38544 32024 -38069 8 VDD
port 41 nsew
rlabel locali s 31860 -38544 31894 -38072 8 VDD
port 41 nsew
rlabel locali s 38348 -38022 38410 -37994 8 VDD
port 41 nsew
rlabel locali s 33376 -38022 38275 -38015 8 VDD
port 41 nsew
rlabel locali s 39139 -37977 39256 -37967 8 VDD
port 41 nsew
rlabel locali s 38576 -37977 38674 -37974 8 VDD
port 41 nsew
rlabel locali s 39139 -37967 39544 -37903 8 VDD
port 41 nsew
rlabel locali s 33376 -38015 38171 -37904 8 VDD
port 41 nsew
rlabel locali s 57567 -37855 64986 -37843 8 VDD
port 41 nsew
rlabel locali s 55120 -37863 55562 -37849 8 VDD
port 41 nsew
rlabel locali s 65954 -37842 74139 -37826 8 VDD
port 41 nsew
rlabel locali s 63873 -37843 64491 -37826 8 VDD
port 41 nsew
rlabel locali s 75107 -37825 83503 -37788 8 VDD
port 41 nsew
rlabel locali s 73026 -37826 73644 -37809 8 VDD
port 41 nsew
rlabel locali s 84471 -37787 86224 -37786 8 VDD
port 41 nsew
rlabel locali s 84471 -37786 87270 -37734 8 VDD
port 41 nsew
rlabel locali s 82390 -37788 83008 -37771 8 VDD
port 41 nsew
rlabel locali s 82390 -37771 82833 -37742 8 VDD
port 41 nsew
rlabel locali s 75107 -37788 81734 -37772 8 VDD
port 41 nsew
rlabel locali s 73026 -37809 73469 -37780 8 VDD
port 41 nsew
rlabel locali s 65954 -37826 72370 -37789 8 VDD
port 41 nsew
rlabel locali s 63873 -37826 64316 -37797 8 VDD
port 41 nsew
rlabel locali s 84838 -37734 87270 -37664 8 VDD
port 41 nsew
rlabel locali s 82391 -37742 82833 -37728 8 VDD
port 41 nsew
rlabel locali s 82391 -37728 83680 -37679 8 VDD
port 41 nsew
rlabel locali s 75474 -37772 81734 -37702 8 VDD
port 41 nsew
rlabel locali s 73027 -37780 73469 -37766 8 VDD
port 41 nsew
rlabel locali s 73027 -37766 74316 -37717 8 VDD
port 41 nsew
rlabel locali s 66321 -37789 72370 -37719 8 VDD
port 41 nsew
rlabel locali s 63874 -37797 64316 -37783 8 VDD
port 41 nsew
rlabel locali s 63874 -37783 65163 -37734 8 VDD
port 41 nsew
rlabel locali s 57567 -37843 63217 -37785 8 VDD
port 41 nsew
rlabel locali s 55120 -37849 56409 -37800 8 VDD
port 41 nsew
rlabel locali s 48369 -37889 54463 -37819 8 VDD
port 41 nsew
rlabel locali s 45922 -37897 46364 -37883 8 VDD
port 41 nsew
rlabel locali s 45922 -37883 47211 -37834 8 VDD
port 41 nsew
rlabel locali s 39139 -37903 45265 -37850 8 VDD
port 41 nsew
rlabel locali s 37058 -37904 37676 -37887 8 VDD
port 41 nsew
rlabel locali s 37058 -37887 37501 -37858 8 VDD
port 41 nsew
rlabel locali s 86596 -37664 87071 -33752 8 VDD
port 41 nsew
rlabel locali s 82793 -37679 83680 -37629 8 VDD
port 41 nsew
rlabel locali s 83598 -37629 83632 -37463 8 VDD
port 41 nsew
rlabel locali s 83402 -37629 83436 -37463 8 VDD
port 41 nsew
rlabel locali s 83206 -37629 83240 -37463 8 VDD
port 41 nsew
rlabel locali s 83010 -37629 83044 -37463 8 VDD
port 41 nsew
rlabel locali s 82793 -37629 82827 -37262 8 VDD
port 41 nsew
rlabel locali s 82597 -37679 82631 -37262 8 VDD
port 41 nsew
rlabel locali s 82401 -37679 82435 -37262 8 VDD
port 41 nsew
rlabel locali s 76821 -37702 81734 -37598 8 VDD
port 41 nsew
rlabel locali s 73429 -37717 74316 -37667 8 VDD
port 41 nsew
rlabel locali s 76821 -37598 82098 -37543 8 VDD
port 41 nsew
rlabel locali s 81380 -37543 82098 -37499 8 VDD
port 41 nsew
rlabel locali s 74234 -37667 74268 -37501 8 VDD
port 41 nsew
rlabel locali s 74038 -37667 74072 -37501 8 VDD
port 41 nsew
rlabel locali s 73842 -37667 73876 -37501 8 VDD
port 41 nsew
rlabel locali s 73646 -37667 73680 -37501 8 VDD
port 41 nsew
rlabel locali s 82016 -37499 82050 -37233 8 VDD
port 41 nsew
rlabel locali s 81820 -37499 81854 -37233 8 VDD
port 41 nsew
rlabel locali s 81624 -37499 81658 -37233 8 VDD
port 41 nsew
rlabel locali s 81428 -37499 81462 -37233 8 VDD
port 41 nsew
rlabel locali s 73429 -37667 73463 -37300 8 VDD
port 41 nsew
rlabel locali s 73233 -37717 73267 -37300 8 VDD
port 41 nsew
rlabel locali s 73037 -37717 73071 -37300 8 VDD
port 41 nsew
rlabel locali s 67659 -37719 72370 -37636 8 VDD
port 41 nsew
rlabel locali s 64276 -37734 65163 -37684 8 VDD
port 41 nsew
rlabel locali s 67659 -37636 72734 -37612 8 VDD
port 41 nsew
rlabel locali s 72016 -37612 72734 -37537 8 VDD
port 41 nsew
rlabel locali s 72652 -37537 72686 -37271 8 VDD
port 41 nsew
rlabel locali s 72456 -37537 72490 -37271 8 VDD
port 41 nsew
rlabel locali s 72260 -37537 72294 -37271 8 VDD
port 41 nsew
rlabel locali s 72064 -37537 72098 -37271 8 VDD
port 41 nsew
rlabel locali s 65081 -37684 65115 -37518 8 VDD
port 41 nsew
rlabel locali s 64885 -37684 64919 -37518 8 VDD
port 41 nsew
rlabel locali s 64689 -37684 64723 -37518 8 VDD
port 41 nsew
rlabel locali s 64493 -37684 64527 -37518 8 VDD
port 41 nsew
rlabel locali s 64276 -37684 64310 -37317 8 VDD
port 41 nsew
rlabel locali s 64080 -37734 64114 -37317 8 VDD
port 41 nsew
rlabel locali s 63884 -37734 63918 -37317 8 VDD
port 41 nsew
rlabel locali s 58912 -37785 63217 -37653 8 VDD
port 41 nsew
rlabel locali s 55522 -37800 56409 -37750 8 VDD
port 41 nsew
rlabel locali s 58912 -37653 63581 -37591 8 VDD
port 41 nsew
rlabel locali s 62863 -37591 63581 -37554 8 VDD
port 41 nsew
rlabel locali s 56327 -37750 56361 -37584 8 VDD
port 41 nsew
rlabel locali s 56131 -37750 56165 -37584 8 VDD
port 41 nsew
rlabel locali s 55935 -37750 55969 -37584 8 VDD
port 41 nsew
rlabel locali s 55739 -37750 55773 -37584 8 VDD
port 41 nsew
rlabel locali s 63499 -37554 63533 -37288 8 VDD
port 41 nsew
rlabel locali s 63303 -37554 63337 -37288 8 VDD
port 41 nsew
rlabel locali s 63107 -37554 63141 -37288 8 VDD
port 41 nsew
rlabel locali s 62911 -37554 62945 -37288 8 VDD
port 41 nsew
rlabel locali s 55522 -37750 55556 -37383 8 VDD
port 41 nsew
rlabel locali s 55326 -37800 55360 -37383 8 VDD
port 41 nsew
rlabel locali s 55130 -37800 55164 -37383 8 VDD
port 41 nsew
rlabel locali s 49729 -37819 54463 -37719 8 VDD
port 41 nsew
rlabel locali s 46324 -37834 47211 -37784 8 VDD
port 41 nsew
rlabel locali s 49729 -37719 54827 -37688 8 VDD
port 41 nsew
rlabel locali s 54109 -37688 54827 -37620 8 VDD
port 41 nsew
rlabel locali s 54745 -37620 54779 -37354 8 VDD
port 41 nsew
rlabel locali s 54549 -37620 54583 -37354 8 VDD
port 41 nsew
rlabel locali s 54353 -37620 54387 -37354 8 VDD
port 41 nsew
rlabel locali s 54157 -37620 54191 -37354 8 VDD
port 41 nsew
rlabel locali s 47129 -37784 47163 -37618 8 VDD
port 41 nsew
rlabel locali s 46933 -37784 46967 -37618 8 VDD
port 41 nsew
rlabel locali s 46737 -37784 46771 -37618 8 VDD
port 41 nsew
rlabel locali s 46541 -37784 46575 -37618 8 VDD
port 41 nsew
rlabel locali s 46324 -37784 46358 -37417 8 VDD
port 41 nsew
rlabel locali s 46128 -37834 46162 -37417 8 VDD
port 41 nsew
rlabel locali s 45932 -37834 45966 -37417 8 VDD
port 41 nsew
rlabel locali s 39506 -37850 45265 -37780 8 VDD
port 41 nsew
rlabel locali s 37059 -37858 37501 -37844 8 VDD
port 41 nsew
rlabel locali s 37059 -37844 38348 -37795 8 VDD
port 41 nsew
rlabel locali s 40878 -37780 45265 -37753 8 VDD
port 41 nsew
rlabel locali s 40878 -37753 45629 -37738 8 VDD
port 41 nsew
rlabel locali s 37461 -37795 38348 -37745 8 VDD
port 41 nsew
rlabel locali s 44911 -37738 45629 -37654 8 VDD
port 41 nsew
rlabel locali s 45547 -37654 45581 -37388 8 VDD
port 41 nsew
rlabel locali s 45351 -37654 45385 -37388 8 VDD
port 41 nsew
rlabel locali s 45155 -37654 45189 -37388 8 VDD
port 41 nsew
rlabel locali s 44959 -37654 44993 -37388 8 VDD
port 41 nsew
rlabel locali s 38266 -37745 38300 -37579 8 VDD
port 41 nsew
rlabel locali s 38070 -37745 38104 -37579 8 VDD
port 41 nsew
rlabel locali s 37874 -37745 37908 -37579 8 VDD
port 41 nsew
rlabel locali s 37678 -37745 37712 -37579 8 VDD
port 41 nsew
rlabel locali s 37461 -37745 37495 -37378 8 VDD
port 41 nsew
rlabel locali s 37265 -37795 37299 -37378 8 VDD
port 41 nsew
rlabel locali s 37069 -37795 37103 -37378 8 VDD
port 41 nsew
rlabel locali s 36230 -37904 36402 -37714 8 VDD
port 41 nsew
rlabel locali s 33376 -37904 33498 -37891 8 VDD
port 41 nsew
rlabel locali s 32409 -38052 32452 -37892 8 VDD
port 41 nsew
rlabel locali s 32212 -38054 32255 -37892 8 VDD
port 41 nsew
rlabel locali s 31981 -38069 32031 -37892 8 VDD
port 41 nsew
rlabel locali s 31855 -38072 31905 -37892 8 VDD
port 41 nsew
rlabel locali s 31265 -38544 31299 -38049 8 VDD
port 41 nsew
rlabel locali s 31069 -38544 31103 -38051 8 VDD
port 41 nsew
rlabel locali s 29696 -38786 29730 -38194 8 VDD
port 41 nsew
rlabel locali s 30136 -38089 30234 -38083 8 VDD
port 41 nsew
rlabel locali s 31263 -38049 31301 -37892 8 VDD
port 41 nsew
rlabel locali s 31066 -38051 31104 -37956 8 VDD
port 41 nsew
rlabel locali s 30136 -38083 30816 -37966 8 VDD
port 41 nsew
rlabel locali s 29908 -38077 29970 -38063 8 VDD
port 41 nsew
rlabel locali s 29689 -38194 29734 -38070 8 VDD
port 41 nsew
rlabel locali s 29273 -38786 29307 -38193 8 VDD
port 41 nsew
rlabel locali s 29077 -38786 29111 -38196 8 VDD
port 41 nsew
rlabel locali s 28827 -38374 28861 -38208 8 VDD
port 41 nsew
rlabel locali s 28631 -38374 28665 -38208 8 VDD
port 41 nsew
rlabel locali s 28435 -38374 28469 -38208 8 VDD
port 41 nsew
rlabel locali s 28239 -38374 28273 -38208 8 VDD
port 41 nsew
rlabel locali s 28022 -38575 28056 -38208 8 VDD
port 41 nsew
rlabel locali s 29267 -38193 29312 -38070 8 VDD
port 41 nsew
rlabel locali s 29072 -38196 29117 -38070 8 VDD
port 41 nsew
rlabel locali s 28022 -38208 28909 -38158 8 VDD
port 41 nsew
rlabel locali s 27826 -38575 27860 -38158 8 VDD
port 41 nsew
rlabel locali s 27630 -38575 27664 -38158 8 VDD
port 41 nsew
rlabel locali s 27620 -38158 28909 -38109 8 VDD
port 41 nsew
rlabel locali s 27620 -38109 28062 -38094 8 VDD
port 41 nsew
rlabel locali s 29066 -38070 29835 -38063 8 VDD
port 41 nsew
rlabel locali s 29066 -38063 29970 -38046 8 VDD
port 41 nsew
rlabel locali s 28059 -38060 28248 -38053 8 VDD
port 41 nsew
rlabel locali s 28022 -38053 28248 -38046 8 VDD
port 41 nsew
rlabel locali s 27620 -38046 29970 -38011 8 VDD
port 41 nsew
rlabel locali s 29908 -38011 29970 -37983 8 VDD
port 41 nsew
rlabel locali s 27620 -38011 29835 -38004 8 VDD
port 41 nsew
rlabel locali s 30699 -37966 30816 -37956 8 VDD
port 41 nsew
rlabel locali s 30136 -37966 30234 -37963 8 VDD
port 41 nsew
rlabel locali s 30699 -37956 31104 -37892 8 VDD
port 41 nsew
rlabel locali s 27620 -38004 29731 -37962 8 VDD
port 41 nsew
rlabel locali s 25407 -39303 25496 -37962 8 VDD
port 41 nsew
rlabel locali s 24714 -39303 25209 -39300 8 VDD
port 41 nsew
rlabel locali s 21701 -39305 23467 -39301 8 VDD
port 41 nsew
rlabel locali s 22014 -39301 23467 -39300 8 VDD
port 41 nsew
rlabel locali s 19389 -39305 20767 -39300 8 VDD
port 41 nsew
rlabel locali s 25115 -39300 25149 -39009 8 VDD
port 41 nsew
rlabel locali s 24919 -39300 24953 -39009 8 VDD
port 41 nsew
rlabel locali s 24723 -39300 24757 -39009 8 VDD
port 41 nsew
rlabel locali s 23372 -39300 23406 -39009 8 VDD
port 41 nsew
rlabel locali s 23176 -39300 23210 -39009 8 VDD
port 41 nsew
rlabel locali s 22980 -39300 23014 -39009 8 VDD
port 41 nsew
rlabel locali s 22415 -39300 22449 -39009 8 VDD
port 41 nsew
rlabel locali s 22219 -39300 22253 -39009 8 VDD
port 41 nsew
rlabel locali s 22023 -39300 22057 -39009 8 VDD
port 41 nsew
rlabel locali s 20672 -39300 20706 -39009 8 VDD
port 41 nsew
rlabel locali s 20476 -39300 20510 -39009 8 VDD
port 41 nsew
rlabel locali s 20280 -39300 20314 -39009 8 VDD
port 41 nsew
rlabel locali s 19790 -39300 19824 -39009 8 VDD
port 41 nsew
rlabel locali s 19594 -39300 19628 -39009 8 VDD
port 41 nsew
rlabel locali s 19398 -39300 19432 -39009 8 VDD
port 41 nsew
rlabel locali s 18068 -39334 18936 -39201 8 VDD
port 41 nsew
rlabel locali s 18264 -39201 18317 -39073 8 VDD
port 41 nsew
rlabel locali s 18068 -39201 18121 -39089 8 VDD
port 41 nsew
rlabel locali s -2309 -40027 -2040 -39099 2 VDD
port 41 nsew
rlabel locali s -3340 -40027 -3071 -39099 2 VDD
port 41 nsew
rlabel locali s -4243 -40027 -3974 -39099 2 VDD
port 41 nsew
rlabel locali s -5105 -40027 -4836 -39099 2 VDD
port 41 nsew
rlabel locali s -5982 -40027 -5713 -39099 2 VDD
port 41 nsew
rlabel locali s -6528 -40027 -6259 -39099 2 VDD
port 41 nsew
rlabel locali s -6816 -40027 -6726 -39938 2 VDD
port 41 nsew
rlabel locali s -7433 -40536 -7399 -39946 2 VDD
port 41 nsew
rlabel locali s -6816 -39938 -6727 -39823 2 VDD
port 41 nsew
rlabel locali s -7439 -39946 -7394 -39823 2 VDD
port 41 nsew
rlabel locali s -7629 -40536 -7595 -39943 2 VDD
port 41 nsew
rlabel locali s -8052 -40536 -8018 -39944 2 VDD
port 41 nsew
rlabel locali s -22237 -40620 -14600 -40453 2 VDD
port 41 nsew
rlabel locali s -25449 -40671 -25383 -40459 2 VDD
port 41 nsew
rlabel locali s -26016 -40671 -25521 -40651 2 VDD
port 41 nsew
rlabel locali s -25569 -40651 -25521 -40459 2 VDD
port 41 nsew
rlabel locali s -7634 -39943 -7589 -39823 2 VDD
port 41 nsew
rlabel locali s -8056 -39944 -8011 -39823 2 VDD
port 41 nsew
rlabel locali s -10512 -40119 -10478 -39828 2 VDD
port 41 nsew
rlabel locali s -10708 -40119 -10674 -39828 2 VDD
port 41 nsew
rlabel locali s -10904 -40119 -10870 -39828 2 VDD
port 41 nsew
rlabel locali s -11349 -40119 -11315 -39828 2 VDD
port 41 nsew
rlabel locali s -11545 -40119 -11511 -39828 2 VDD
port 41 nsew
rlabel locali s -11741 -40119 -11707 -39828 2 VDD
port 41 nsew
rlabel locali s -13212 -40119 -13178 -39828 2 VDD
port 41 nsew
rlabel locali s -13408 -40119 -13374 -39828 2 VDD
port 41 nsew
rlabel locali s -13604 -40119 -13570 -39828 2 VDD
port 41 nsew
rlabel locali s -14049 -40119 -14015 -39828 2 VDD
port 41 nsew
rlabel locali s -14245 -40119 -14211 -39828 2 VDD
port 41 nsew
rlabel locali s -14441 -40119 -14407 -39828 2 VDD
port 41 nsew
rlabel locali s -14690 -40453 -14601 -39828 2 VDD
port 41 nsew
rlabel locali s -12219 -39828 -10417 -39823 2 VDD
port 41 nsew
rlabel locali s -14690 -39828 -13117 -39823 2 VDD
port 41 nsew
rlabel locali s -14690 -39823 -6727 -39760 2 VDD
port 41 nsew
rlabel locali s -25569 -40459 -25383 -40449 2 VDD
port 41 nsew
rlabel locali s -26016 -40449 -25383 -40415 2 VDD
port 41 nsew
rlabel locali s -25569 -40415 -25383 -40400 2 VDD
port 41 nsew
rlabel locali s -25449 -40400 -25383 -40218 2 VDD
port 41 nsew
rlabel locali s -25569 -40400 -25521 -40218 2 VDD
port 41 nsew
rlabel locali s -25569 -40218 -25383 -40213 2 VDD
port 41 nsew
rlabel locali s -26016 -40213 -25383 -40179 2 VDD
port 41 nsew
rlabel locali s -25569 -40179 -25383 -40159 2 VDD
port 41 nsew
rlabel locali s -25449 -40159 -25383 -39986 2 VDD
port 41 nsew
rlabel locali s -25569 -40159 -25521 -39986 2 VDD
port 41 nsew
rlabel locali s -25569 -39986 -25383 -39977 2 VDD
port 41 nsew
rlabel locali s -26016 -39977 -25383 -39943 2 VDD
port 41 nsew
rlabel locali s -25569 -39943 -25383 -39927 2 VDD
port 41 nsew
rlabel locali s -10612 -39760 -6727 -39738 2 VDD
port 41 nsew
rlabel locali s -6816 -39738 -6727 -39099 2 VDD
port 41 nsew
rlabel locali s 18273 -39073 18307 -38489 8 VDD
port 41 nsew
rlabel locali s 18077 -39089 18111 -38489 8 VDD
port 41 nsew
rlabel locali s -6816 -39099 -1591 -39036 2 VDD
port 41 nsew
rlabel locali s -4345 -39036 -2543 -39031 2 VDD
port 41 nsew
rlabel locali s -6816 -39036 -5243 -39031 2 VDD
port 41 nsew
rlabel locali s -2638 -39031 -2604 -38740 2 VDD
port 41 nsew
rlabel locali s -2834 -39031 -2800 -38740 2 VDD
port 41 nsew
rlabel locali s -3030 -39031 -2996 -38740 2 VDD
port 41 nsew
rlabel locali s -3475 -39031 -3441 -38740 2 VDD
port 41 nsew
rlabel locali s -3671 -39031 -3637 -38740 2 VDD
port 41 nsew
rlabel locali s -3867 -39031 -3833 -38740 2 VDD
port 41 nsew
rlabel locali s -5338 -39031 -5304 -38740 2 VDD
port 41 nsew
rlabel locali s -5534 -39031 -5500 -38740 2 VDD
port 41 nsew
rlabel locali s -5730 -39031 -5696 -38740 2 VDD
port 41 nsew
rlabel locali s -6175 -39031 -6141 -38740 2 VDD
port 41 nsew
rlabel locali s -6371 -39031 -6337 -38740 2 VDD
port 41 nsew
rlabel locali s -6567 -39031 -6533 -38740 2 VDD
port 41 nsew
rlabel locali s 25407 -37962 29731 -37893 8 VDD
port 41 nsew
rlabel locali s 30699 -37892 32452 -37891 8 VDD
port 41 nsew
rlabel locali s 30699 -37891 33498 -37839 8 VDD
port 41 nsew
rlabel locali s 28618 -37893 29236 -37876 8 VDD
port 41 nsew
rlabel locali s 28618 -37876 29061 -37847 8 VDD
port 41 nsew
rlabel locali s 31066 -37839 33498 -37769 8 VDD
port 41 nsew
rlabel locali s 28619 -37847 29061 -37833 8 VDD
port 41 nsew
rlabel locali s 28619 -37833 29908 -37784 8 VDD
port 41 nsew
rlabel locali s 29021 -37784 29908 -37734 8 VDD
port 41 nsew
rlabel locali s 36048 -37714 36766 -37615 8 VDD
port 41 nsew
rlabel locali s 36684 -37615 36718 -37349 8 VDD
port 41 nsew
rlabel locali s 36488 -37615 36522 -37349 8 VDD
port 41 nsew
rlabel locali s 36292 -37615 36326 -37349 8 VDD
port 41 nsew
rlabel locali s 36096 -37615 36130 -37349 8 VDD
port 41 nsew
rlabel locali s 29826 -37734 29860 -37568 8 VDD
port 41 nsew
rlabel locali s 29630 -37734 29664 -37568 8 VDD
port 41 nsew
rlabel locali s 29434 -37734 29468 -37568 8 VDD
port 41 nsew
rlabel locali s 29238 -37734 29272 -37568 8 VDD
port 41 nsew
rlabel locali s 29021 -37734 29055 -37367 8 VDD
port 41 nsew
rlabel locali s 28825 -37784 28859 -37367 8 VDD
port 41 nsew
rlabel locali s 28629 -37784 28663 -37367 8 VDD
port 41 nsew
rlabel locali s 25407 -37893 27962 -37703 8 VDD
port 41 nsew
rlabel locali s 25407 -37703 28326 -37668 8 VDD
port 41 nsew
rlabel locali s 27608 -37668 28326 -37604 8 VDD
port 41 nsew
rlabel locali s 25407 -37668 25496 -37608 8 VDD
port 41 nsew
rlabel locali s 25213 -37899 25247 -37608 8 VDD
port 41 nsew
rlabel locali s 25017 -37899 25051 -37608 8 VDD
port 41 nsew
rlabel locali s 24821 -37899 24855 -37608 8 VDD
port 41 nsew
rlabel locali s 24376 -37899 24410 -37608 8 VDD
port 41 nsew
rlabel locali s 24180 -37899 24214 -37608 8 VDD
port 41 nsew
rlabel locali s 23984 -37899 24018 -37608 8 VDD
port 41 nsew
rlabel locali s 22513 -37899 22547 -37608 8 VDD
port 41 nsew
rlabel locali s 22317 -37899 22351 -37608 8 VDD
port 41 nsew
rlabel locali s 22121 -37899 22155 -37608 8 VDD
port 41 nsew
rlabel locali s 21676 -37899 21710 -37608 8 VDD
port 41 nsew
rlabel locali s 21480 -37899 21514 -37608 8 VDD
port 41 nsew
rlabel locali s 21284 -37899 21318 -37608 8 VDD
port 41 nsew
rlabel locali s 28244 -37604 28278 -37338 8 VDD
port 41 nsew
rlabel locali s 28048 -37604 28082 -37338 8 VDD
port 41 nsew
rlabel locali s 27852 -37604 27886 -37338 8 VDD
port 41 nsew
rlabel locali s 27656 -37604 27690 -37338 8 VDD
port 41 nsew
rlabel locali s 23923 -37608 25496 -37603 8 VDD
port 41 nsew
rlabel locali s 21223 -37608 23025 -37603 8 VDD
port 41 nsew
rlabel locali s 20271 -37603 25496 -37540 8 VDD
port 41 nsew
rlabel locali s 8050 -37649 8084 -37459 8 VDD
port 41 nsew
rlabel locali s 7854 -37649 7888 -37471 8 VDD
port 41 nsew
rlabel locali s 8045 -37459 8091 -37337 8 VDD
port 41 nsew
rlabel locali s 7848 -37471 7894 -37337 8 VDD
port 41 nsew
rlabel locali s 7741 -37649 7775 -37461 8 VDD
port 41 nsew
rlabel locali s 7545 -37649 7579 -37466 8 VDD
port 41 nsew
rlabel locali s 7735 -37461 7781 -37337 8 VDD
port 41 nsew
rlabel locali s 7539 -37466 7585 -37337 8 VDD
port 41 nsew
rlabel locali s 7431 -37649 7465 -37462 8 VDD
port 41 nsew
rlabel locali s 7235 -37649 7269 -37466 8 VDD
port 41 nsew
rlabel locali s 7039 -37649 7073 -37466 8 VDD
port 41 nsew
rlabel locali s 7426 -37462 7472 -37337 8 VDD
port 41 nsew
rlabel locali s 7228 -37466 7274 -37337 8 VDD
port 41 nsew
rlabel locali s 7039 -37466 7079 -37377 8 VDD
port 41 nsew
rlabel locali s 7038 -37377 7161 -37337 8 VDD
port 41 nsew
rlabel locali s 5878 -37638 5912 -37376 8 VDD
port 41 nsew
rlabel locali s 7038 -37337 8091 -37268 8 VDD
port 41 nsew
rlabel locali s 7038 -37268 7161 -37241 8 VDD
port 41 nsew
rlabel locali s 5822 -37376 5945 -37342 8 VDD
port 41 nsew
rlabel locali s 5682 -37638 5716 -37342 8 VDD
port 41 nsew
rlabel locali s 5486 -37638 5520 -37342 8 VDD
port 41 nsew
rlabel locali s 5290 -37638 5324 -37342 8 VDD
port 41 nsew
rlabel locali s 4748 -37638 4782 -37346 8 VDD
port 41 nsew
rlabel locali s 4552 -37638 4586 -37371 8 VDD
port 41 nsew
rlabel locali s 4125 -37763 4159 -37373 8 VDD
port 41 nsew
rlabel locali s 4466 -37371 4589 -37346 8 VDD
port 41 nsew
rlabel locali s 5290 -37342 5945 -37341 8 VDD
port 41 nsew
rlabel locali s 4466 -37346 4787 -37341 8 VDD
port 41 nsew
rlabel locali s 4466 -37341 5945 -37273 8 VDD
port 41 nsew
rlabel locali s 5822 -37273 5945 -37240 8 VDD
port 41 nsew
rlabel locali s 4466 -37273 5362 -37268 8 VDD
port 41 nsew
rlabel locali s 4466 -37268 4589 -37235 8 VDD
port 41 nsew
rlabel locali s 4065 -37373 4188 -37346 8 VDD
port 41 nsew
rlabel locali s 3929 -37763 3963 -37346 8 VDD
port 41 nsew
rlabel locali s 3733 -37763 3767 -37396 8 VDD
port 41 nsew
rlabel locali s 3516 -37562 3550 -37396 8 VDD
port 41 nsew
rlabel locali s 3320 -37562 3354 -37396 8 VDD
port 41 nsew
rlabel locali s 3124 -37562 3158 -37396 8 VDD
port 41 nsew
rlabel locali s 2928 -37562 2962 -37396 8 VDD
port 41 nsew
rlabel locali s 2520 -37761 2554 -37397 8 VDD
port 41 nsew
rlabel locali s 2837 -37396 3767 -37346 8 VDD
port 41 nsew
rlabel locali s 2837 -37346 4188 -37297 8 VDD
port 41 nsew
rlabel locali s 3727 -37297 4188 -37282 8 VDD
port 41 nsew
rlabel locali s 4065 -37282 4188 -37237 8 VDD
port 41 nsew
rlabel locali s 2837 -37297 2960 -37260 8 VDD
port 41 nsew
rlabel locali s 2448 -37397 2571 -37354 8 VDD
port 41 nsew
rlabel locali s 2324 -37761 2358 -37354 8 VDD
port 41 nsew
rlabel locali s 2128 -37761 2162 -37394 8 VDD
port 41 nsew
rlabel locali s 1911 -37560 1945 -37394 8 VDD
port 41 nsew
rlabel locali s 1715 -37560 1749 -37394 8 VDD
port 41 nsew
rlabel locali s 1519 -37560 1553 -37394 8 VDD
port 41 nsew
rlabel locali s 1323 -37560 1357 -37394 8 VDD
port 41 nsew
rlabel locali s 1275 -37394 2162 -37354 8 VDD
port 41 nsew
rlabel locali s 916 -37647 950 -37354 8 VDD
port 41 nsew
rlabel locali s 720 -37647 754 -37354 8 VDD
port 41 nsew
rlabel locali s 524 -37647 558 -37354 8 VDD
port 41 nsew
rlabel locali s 328 -37647 362 -37354 8 VDD
port 41 nsew
rlabel locali s -214 -37647 -180 -37355 2 VDD
port 41 nsew
rlabel locali s -410 -37647 -376 -37384 2 VDD
port 41 nsew
rlabel locali s -752 -37630 -718 -37385 2 VDD
port 41 nsew
rlabel locali s -530 -37384 -376 -37355 2 VDD
port 41 nsew
rlabel locali s -530 -37355 -175 -37354 2 VDD
port 41 nsew
rlabel locali s -530 -37354 2571 -37275 8 VDD
port 41 nsew
rlabel locali s 2448 -37275 2571 -37261 8 VDD
port 41 nsew
rlabel locali s 405 -37275 520 -36467 8 VDD
port 41 nsew
rlabel locali s -530 -37275 -407 -37248 2 VDD
port 41 nsew
rlabel locali s -824 -37385 -701 -37339 2 VDD
port 41 nsew
rlabel locali s -948 -37630 -914 -37339 2 VDD
port 41 nsew
rlabel locali s -1144 -37630 -1110 -37339 2 VDD
port 41 nsew
rlabel locali s -1634 -37630 -1600 -37339 2 VDD
port 41 nsew
rlabel locali s -1830 -37630 -1796 -37339 2 VDD
port 41 nsew
rlabel locali s -2026 -37630 -1992 -37339 2 VDD
port 41 nsew
rlabel locali s -3377 -37630 -3343 -37339 2 VDD
port 41 nsew
rlabel locali s -3573 -37630 -3539 -37339 2 VDD
port 41 nsew
rlabel locali s -3769 -37630 -3735 -37339 2 VDD
port 41 nsew
rlabel locali s -4334 -37630 -4300 -37339 2 VDD
port 41 nsew
rlabel locali s -4530 -37630 -4496 -37339 2 VDD
port 41 nsew
rlabel locali s -4726 -37630 -4692 -37339 2 VDD
port 41 nsew
rlabel locali s -6077 -37630 -6043 -37339 2 VDD
port 41 nsew
rlabel locali s -6273 -37630 -6239 -37339 2 VDD
port 41 nsew
rlabel locali s -6469 -37630 -6435 -37339 2 VDD
port 41 nsew
rlabel locali s -2087 -37339 -701 -37334 2 VDD
port 41 nsew
rlabel locali s -4787 -37339 -3334 -37338 2 VDD
port 41 nsew
rlabel locali s -4787 -37338 -3021 -37334 2 VDD
port 41 nsew
rlabel locali s -6529 -37339 -6034 -37336 2 VDD
port 41 nsew
rlabel locali s -6816 -39031 -6727 -37336 2 VDD
port 41 nsew
rlabel locali s -11220 -38838 -11186 -38672 2 VDD
port 41 nsew
rlabel locali s -11416 -38838 -11382 -38672 2 VDD
port 41 nsew
rlabel locali s -11612 -38838 -11578 -38672 2 VDD
port 41 nsew
rlabel locali s -11808 -38838 -11774 -38672 2 VDD
port 41 nsew
rlabel locali s -12025 -39039 -11991 -38672 2 VDD
port 41 nsew
rlabel locali s -12025 -38672 -11138 -38622 2 VDD
port 41 nsew
rlabel locali s -12221 -39039 -12187 -38622 2 VDD
port 41 nsew
rlabel locali s -12417 -39039 -12383 -38622 2 VDD
port 41 nsew
rlabel locali s -12802 -39068 -12768 -38802 2 VDD
port 41 nsew
rlabel locali s -12998 -39068 -12964 -38802 2 VDD
port 41 nsew
rlabel locali s -13194 -39068 -13160 -38802 2 VDD
port 41 nsew
rlabel locali s -13390 -39068 -13356 -38802 2 VDD
port 41 nsew
rlabel locali s -13438 -38802 -12720 -38703 2 VDD
port 41 nsew
rlabel locali s -12427 -38622 -11138 -38573 2 VDD
port 41 nsew
rlabel locali s -12427 -38573 -11985 -38559 2 VDD
port 41 nsew
rlabel locali s -12428 -38559 -11985 -38530 2 VDD
port 41 nsew
rlabel locali s -12428 -38530 -11810 -38513 2 VDD
port 41 nsew
rlabel locali s -13256 -38703 -13084 -38513 2 VDD
port 41 nsew
rlabel locali s -14228 -39760 -14075 -38513 2 VDD
port 41 nsew
rlabel locali s -14228 -38513 -11315 -38402 2 VDD
port 41 nsew
rlabel locali s -14228 -38402 -11211 -38360 2 VDD
port 41 nsew
rlabel locali s -11980 -38360 -11211 -38336 2 VDD
port 41 nsew
rlabel locali s -13024 -38360 -12798 -38353 2 VDD
port 41 nsew
rlabel locali s -12987 -38353 -12798 -38346 2 VDD
port 41 nsew
rlabel locali s -11357 -38336 -11312 -38212 2 VDD
port 41 nsew
rlabel locali s -11779 -38336 -11734 -38213 2 VDD
port 41 nsew
rlabel locali s -11350 -38212 -11316 -37620 2 VDD
port 41 nsew
rlabel locali s -11773 -38213 -11739 -37620 2 VDD
port 41 nsew
rlabel locali s -11974 -38336 -11929 -38210 2 VDD
port 41 nsew
rlabel locali s -13426 -38312 -12984 -38297 2 VDD
port 41 nsew
rlabel locali s -13426 -38297 -12137 -38248 2 VDD
port 41 nsew
rlabel locali s -11969 -38210 -11935 -37620 2 VDD
port 41 nsew
rlabel locali s -13024 -38248 -12137 -38198 2 VDD
port 41 nsew
rlabel locali s -12219 -38198 -12185 -38032 2 VDD
port 41 nsew
rlabel locali s -12415 -38198 -12381 -38032 2 VDD
port 41 nsew
rlabel locali s -12611 -38198 -12577 -38032 2 VDD
port 41 nsew
rlabel locali s -12807 -38198 -12773 -38032 2 VDD
port 41 nsew
rlabel locali s -13024 -38198 -12990 -37831 2 VDD
port 41 nsew
rlabel locali s -13220 -38248 -13186 -37831 2 VDD
port 41 nsew
rlabel locali s -13416 -38248 -13382 -37831 2 VDD
port 41 nsew
rlabel locali s -6816 -37336 -5712 -37334 2 VDD
port 41 nsew
rlabel locali s -6816 -37334 -701 -37271 2 VDD
port 41 nsew
rlabel locali s -824 -37271 -701 -37249 2 VDD
port 41 nsew
rlabel locali s -2079 -37271 -1964 -36575 2 VDD
port 41 nsew
rlabel locali s -3494 -37271 -3021 -37270 2 VDD
port 41 nsew
rlabel locali s -4645 -37271 -4530 -36719 2 VDD
port 41 nsew
rlabel locali s -6816 -37271 -5712 -37268 2 VDD
port 41 nsew
rlabel locali s -5938 -37268 -5850 -36878 2 VDD
port 41 nsew
rlabel locali s -6120 -37268 -6032 -36878 2 VDD
port 41 nsew
rlabel locali s -6303 -37268 -6215 -36878 2 VDD
port 41 nsew
rlabel locali s -6319 -36878 -5824 -36810 2 VDD
port 41 nsew
rlabel locali s -4650 -36719 -4527 -36583 2 VDD
port 41 nsew
rlabel locali s 400 -36467 706 -36405 8 VDD
port 41 nsew
rlabel locali s -2083 -36575 -1960 -36439 2 VDD
port 41 nsew
rlabel locali s -5918 -36810 -5884 -36519 2 VDD
port 41 nsew
rlabel locali s -6114 -36810 -6080 -36519 2 VDD
port 41 nsew
rlabel locali s -6310 -36810 -6276 -36519 2 VDD
port 41 nsew
rlabel locali s -14228 -38360 -14075 -36664 2 VDD
port 41 nsew
rlabel locali s -25449 -39927 -25383 -39380 2 VDD
port 41 nsew
rlabel locali s -25569 -39927 -25521 -39847 2 VDD
port 41 nsew
rlabel locali s -26016 -39847 -25521 -39813 2 VDD
port 41 nsew
rlabel locali s -25569 -39813 -25521 -39611 2 VDD
port 41 nsew
rlabel locali s -26016 -39611 -25521 -39577 2 VDD
port 41 nsew
rlabel locali s -25569 -39577 -25521 -39380 2 VDD
port 41 nsew
rlabel locali s -25569 -39380 -25383 -39375 2 VDD
port 41 nsew
rlabel locali s -26016 -39375 -25383 -39341 2 VDD
port 41 nsew
rlabel locali s -25569 -39341 -25383 -39321 2 VDD
port 41 nsew
rlabel locali s -25449 -39321 -25383 -39151 2 VDD
port 41 nsew
rlabel locali s -25569 -39321 -25521 -39151 2 VDD
port 41 nsew
rlabel locali s -25569 -39151 -25383 -39139 2 VDD
port 41 nsew
rlabel locali s -26016 -39139 -25383 -39105 2 VDD
port 41 nsew
rlabel locali s -25569 -39105 -25383 -39092 2 VDD
port 41 nsew
rlabel locali s -25449 -39092 -25383 -38912 2 VDD
port 41 nsew
rlabel locali s -25569 -39092 -25521 -38912 2 VDD
port 41 nsew
rlabel locali s -25569 -38912 -25383 -38903 2 VDD
port 41 nsew
rlabel locali s -26016 -38903 -25383 -38869 2 VDD
port 41 nsew
rlabel locali s -25569 -38869 -25383 -38853 2 VDD
port 41 nsew
rlabel locali s -25449 -38853 -25383 -38677 2 VDD
port 41 nsew
rlabel locali s -25569 -38853 -25521 -38677 2 VDD
port 41 nsew
rlabel locali s -25569 -38677 -25383 -38667 2 VDD
port 41 nsew
rlabel locali s -26016 -38667 -25383 -38633 2 VDD
port 41 nsew
rlabel locali s -25569 -38633 -25383 -38618 2 VDD
port 41 nsew
rlabel locali s -25449 -38618 -25383 -38441 2 VDD
port 41 nsew
rlabel locali s -25569 -38618 -25521 -38441 2 VDD
port 41 nsew
rlabel locali s -25569 -38441 -25383 -38431 2 VDD
port 41 nsew
rlabel locali s -26016 -38431 -25383 -38397 2 VDD
port 41 nsew
rlabel locali s -25569 -38397 -25383 -38382 2 VDD
port 41 nsew
rlabel locali s -25449 -38382 -25383 -38210 2 VDD
port 41 nsew
rlabel locali s -25569 -38382 -25521 -38210 2 VDD
port 41 nsew
rlabel locali s -25569 -38210 -25383 -38195 2 VDD
port 41 nsew
rlabel locali s -26016 -38195 -25383 -38161 2 VDD
port 41 nsew
rlabel locali s -25569 -38161 -25383 -38151 2 VDD
port 41 nsew
rlabel locali s -16209 -37862 -16175 -37696 2 VDD
port 41 nsew
rlabel locali s -16405 -37862 -16371 -37696 2 VDD
port 41 nsew
rlabel locali s -16601 -37862 -16567 -37696 2 VDD
port 41 nsew
rlabel locali s -16797 -37862 -16763 -37696 2 VDD
port 41 nsew
rlabel locali s -17014 -38063 -16980 -37696 2 VDD
port 41 nsew
rlabel locali s -17014 -37696 -16127 -37646 2 VDD
port 41 nsew
rlabel locali s -17210 -38063 -17176 -37646 2 VDD
port 41 nsew
rlabel locali s -17406 -38063 -17372 -37646 2 VDD
port 41 nsew
rlabel locali s -17791 -38092 -17757 -37826 2 VDD
port 41 nsew
rlabel locali s -17987 -38092 -17953 -37826 2 VDD
port 41 nsew
rlabel locali s -18183 -38092 -18149 -37826 2 VDD
port 41 nsew
rlabel locali s -18379 -38092 -18345 -37826 2 VDD
port 41 nsew
rlabel locali s -18427 -37826 -17709 -37727 2 VDD
port 41 nsew
rlabel locali s -17416 -37646 -16127 -37597 2 VDD
port 41 nsew
rlabel locali s -17416 -37597 -16974 -37583 2 VDD
port 41 nsew
rlabel locali s -17417 -37583 -16974 -37554 2 VDD
port 41 nsew
rlabel locali s -17417 -37554 -16799 -37537 2 VDD
port 41 nsew
rlabel locali s -18245 -37727 -18073 -37537 2 VDD
port 41 nsew
rlabel locali s -18884 -37915 -18850 -37656 2 VDD
port 41 nsew
rlabel locali s -19080 -37915 -19046 -37656 2 VDD
port 41 nsew
rlabel locali s -19622 -37915 -19588 -37656 2 VDD
port 41 nsew
rlabel locali s -19818 -37915 -19784 -37656 2 VDD
port 41 nsew
rlabel locali s -20014 -37915 -19980 -37656 2 VDD
port 41 nsew
rlabel locali s -20210 -37915 -20176 -37656 2 VDD
port 41 nsew
rlabel locali s -20786 -37909 -20752 -37743 2 VDD
port 41 nsew
rlabel locali s -20982 -37909 -20948 -37743 2 VDD
port 41 nsew
rlabel locali s -21178 -37909 -21144 -37743 2 VDD
port 41 nsew
rlabel locali s -21374 -37909 -21340 -37743 2 VDD
port 41 nsew
rlabel locali s -21591 -38110 -21557 -37743 2 VDD
port 41 nsew
rlabel locali s -21591 -37743 -20704 -37693 2 VDD
port 41 nsew
rlabel locali s -21787 -38110 -21753 -37693 2 VDD
port 41 nsew
rlabel locali s -21983 -38110 -21949 -37693 2 VDD
port 41 nsew
rlabel locali s -21993 -37693 -20704 -37656 2 VDD
port 41 nsew
rlabel locali s -23653 -37656 -18850 -37623 2 VDD
port 41 nsew
rlabel locali s -23653 -37623 -18840 -37593 2 VDD
port 41 nsew
rlabel locali s -25449 -38151 -25383 -37593 2 VDD
port 41 nsew
rlabel locali s -25449 -37593 -18840 -37537 2 VDD
port 41 nsew
rlabel locali s -25449 -37537 -16304 -37485 2 VDD
port 41 nsew
rlabel locali s -25569 -38151 -25521 -37959 2 VDD
port 41 nsew
rlabel locali s -26016 -37959 -25521 -37925 2 VDD
port 41 nsew
rlabel locali s -25569 -37925 -25521 -37711 2 VDD
port 41 nsew
rlabel locali s -26016 -37711 -25521 -37677 2 VDD
port 41 nsew
rlabel locali s -25569 -37677 -25521 -37485 2 VDD
port 41 nsew
rlabel locali s -25569 -37485 -16304 -37475 2 VDD
port 41 nsew
rlabel locali s -26016 -37475 -16304 -37441 2 VDD
port 41 nsew
rlabel locali s -25569 -37441 -16304 -37426 2 VDD
port 41 nsew
rlabel locali s -25449 -37426 -16200 -37424 2 VDD
port 41 nsew
rlabel locali s -18415 -37424 -16200 -37384 2 VDD
port 41 nsew
rlabel locali s -16969 -37384 -16200 -37360 2 VDD
port 41 nsew
rlabel locali s -18013 -37384 -17787 -37377 2 VDD
port 41 nsew
rlabel locali s -17976 -37377 -17787 -37370 2 VDD
port 41 nsew
rlabel locali s -16346 -37360 -16301 -37236 2 VDD
port 41 nsew
rlabel locali s -16768 -37360 -16723 -37237 2 VDD
port 41 nsew
rlabel locali s -11368 -36662 -10895 -36661 2 VDD
port 41 nsew
rlabel locali s -14690 -36664 -13586 -36661 2 VDD
port 41 nsew
rlabel locali s -14690 -36661 -8583 -36598 2 VDD
port 41 nsew
rlabel locali s -16339 -37236 -16305 -36644 2 VDD
port 41 nsew
rlabel locali s -16762 -37237 -16728 -36644 2 VDD
port 41 nsew
rlabel locali s -16963 -37360 -16918 -37234 2 VDD
port 41 nsew
rlabel locali s -18415 -37336 -17973 -37321 2 VDD
port 41 nsew
rlabel locali s -18415 -37321 -17126 -37272 2 VDD
port 41 nsew
rlabel locali s -25449 -37424 -23381 -37321 2 VDD
port 41 nsew
rlabel locali s -16958 -37234 -16924 -36644 2 VDD
port 41 nsew
rlabel locali s -18013 -37272 -17126 -37222 2 VDD
port 41 nsew
rlabel locali s -17208 -37222 -17174 -37056 2 VDD
port 41 nsew
rlabel locali s -17404 -37222 -17370 -37056 2 VDD
port 41 nsew
rlabel locali s -17600 -37222 -17566 -37056 2 VDD
port 41 nsew
rlabel locali s -17796 -37222 -17762 -37056 2 VDD
port 41 nsew
rlabel locali s -18013 -37222 -17979 -36855 2 VDD
port 41 nsew
rlabel locali s -18209 -37272 -18175 -36855 2 VDD
port 41 nsew
rlabel locali s -18405 -37272 -18371 -36855 2 VDD
port 41 nsew
rlabel locali s -9961 -36598 -8583 -36593 2 VDD
port 41 nsew
rlabel locali s -12661 -36598 -10895 -36594 2 VDD
port 41 nsew
rlabel locali s -14690 -36598 -13586 -36596 2 VDD
port 41 nsew
rlabel locali s -12661 -36594 -11208 -36593 2 VDD
port 41 nsew
rlabel locali s -14403 -36596 -13908 -36593 2 VDD
port 41 nsew
rlabel locali s 400 -36405 523 -36404 8 VDD
port 41 nsew
rlabel locali s -8626 -36593 -8592 -36302 2 VDD
port 41 nsew
rlabel locali s -8822 -36593 -8788 -36302 2 VDD
port 41 nsew
rlabel locali s -9018 -36593 -8984 -36302 2 VDD
port 41 nsew
rlabel locali s -9508 -36593 -9474 -36302 2 VDD
port 41 nsew
rlabel locali s -9704 -36593 -9670 -36302 2 VDD
port 41 nsew
rlabel locali s -9900 -36593 -9866 -36302 2 VDD
port 41 nsew
rlabel locali s -11251 -36593 -11217 -36302 2 VDD
port 41 nsew
rlabel locali s -11447 -36593 -11413 -36302 2 VDD
port 41 nsew
rlabel locali s -11643 -36593 -11609 -36302 2 VDD
port 41 nsew
rlabel locali s -12208 -36593 -12174 -36302 2 VDD
port 41 nsew
rlabel locali s -12404 -36593 -12370 -36302 2 VDD
port 41 nsew
rlabel locali s -12600 -36593 -12566 -36302 2 VDD
port 41 nsew
rlabel locali s -13951 -36593 -13917 -36302 2 VDD
port 41 nsew
rlabel locali s -14147 -36593 -14113 -36302 2 VDD
port 41 nsew
rlabel locali s -14343 -36593 -14309 -36302 2 VDD
port 41 nsew
rlabel locali s 401 -35987 524 -35851 8 VDD
port 41 nsew
rlabel locali s -2082 -35987 -1959 -35851 2 VDD
port 41 nsew
rlabel locali s 8040 -35398 8074 -35208 8 VDD
port 41 nsew
rlabel locali s 7844 -35398 7878 -35220 8 VDD
port 41 nsew
rlabel locali s 25923 -35141 27026 -33752 8 VDD
port 41 nsew
rlabel locali s 8035 -35208 8081 -35086 8 VDD
port 41 nsew
rlabel locali s 7838 -35220 7884 -35086 8 VDD
port 41 nsew
rlabel locali s 7731 -35398 7765 -35210 8 VDD
port 41 nsew
rlabel locali s 7535 -35398 7569 -35215 8 VDD
port 41 nsew
rlabel locali s 7725 -35210 7771 -35086 8 VDD
port 41 nsew
rlabel locali s 7529 -35215 7575 -35086 8 VDD
port 41 nsew
rlabel locali s 7421 -35398 7455 -35211 8 VDD
port 41 nsew
rlabel locali s 7225 -35398 7259 -35215 8 VDD
port 41 nsew
rlabel locali s 7029 -35398 7063 -35215 8 VDD
port 41 nsew
rlabel locali s 7416 -35211 7462 -35086 8 VDD
port 41 nsew
rlabel locali s 7218 -35215 7264 -35086 8 VDD
port 41 nsew
rlabel locali s 7029 -35215 7069 -35086 8 VDD
port 41 nsew
rlabel locali s 5040 -35398 5074 -35208 8 VDD
port 41 nsew
rlabel locali s 4844 -35398 4878 -35220 8 VDD
port 41 nsew
rlabel locali s 7029 -35086 8081 -34979 8 VDD
port 41 nsew
rlabel locali s 5035 -35208 5081 -35086 8 VDD
port 41 nsew
rlabel locali s 4838 -35220 4884 -35086 8 VDD
port 41 nsew
rlabel locali s 4731 -35398 4765 -35210 8 VDD
port 41 nsew
rlabel locali s 4535 -35398 4569 -35215 8 VDD
port 41 nsew
rlabel locali s 4725 -35210 4771 -35086 8 VDD
port 41 nsew
rlabel locali s 4529 -35215 4575 -35086 8 VDD
port 41 nsew
rlabel locali s 4421 -35398 4455 -35211 8 VDD
port 41 nsew
rlabel locali s 4225 -35398 4259 -35215 8 VDD
port 41 nsew
rlabel locali s 4029 -35398 4063 -35215 8 VDD
port 41 nsew
rlabel locali s 4416 -35211 4462 -35086 8 VDD
port 41 nsew
rlabel locali s 4218 -35215 4264 -35086 8 VDD
port 41 nsew
rlabel locali s 4029 -35215 4069 -35086 8 VDD
port 41 nsew
rlabel locali s 2540 -35398 2574 -35208 8 VDD
port 41 nsew
rlabel locali s 2344 -35398 2378 -35220 8 VDD
port 41 nsew
rlabel locali s 4029 -35086 5081 -35017 8 VDD
port 41 nsew
rlabel locali s 2535 -35208 2581 -35086 8 VDD
port 41 nsew
rlabel locali s 2338 -35220 2384 -35086 8 VDD
port 41 nsew
rlabel locali s 2231 -35398 2265 -35210 8 VDD
port 41 nsew
rlabel locali s 2035 -35398 2069 -35215 8 VDD
port 41 nsew
rlabel locali s 2225 -35210 2271 -35086 8 VDD
port 41 nsew
rlabel locali s 2029 -35215 2075 -35086 8 VDD
port 41 nsew
rlabel locali s 1921 -35398 1955 -35211 8 VDD
port 41 nsew
rlabel locali s 1725 -35398 1759 -35215 8 VDD
port 41 nsew
rlabel locali s 1529 -35398 1563 -35215 8 VDD
port 41 nsew
rlabel locali s 1916 -35211 1962 -35086 8 VDD
port 41 nsew
rlabel locali s 1718 -35215 1764 -35086 8 VDD
port 41 nsew
rlabel locali s 1529 -35215 1569 -35086 8 VDD
port 41 nsew
rlabel locali s 1529 -35086 2581 -35017 8 VDD
port 41 nsew
rlabel locali s 4306 -35017 4899 -34979 8 VDD
port 41 nsew
rlabel locali s 1893 -35017 2486 -34979 8 VDD
port 41 nsew
rlabel locali s 406 -35851 521 -34979 8 VDD
port 41 nsew
rlabel locali s 40 -35398 74 -35208 8 VDD
port 41 nsew
rlabel locali s -156 -35398 -122 -35220 2 VDD
port 41 nsew
rlabel locali s 35 -35208 81 -35086 8 VDD
port 41 nsew
rlabel locali s -162 -35220 -116 -35086 2 VDD
port 41 nsew
rlabel locali s -269 -35398 -235 -35210 2 VDD
port 41 nsew
rlabel locali s -465 -35398 -431 -35215 2 VDD
port 41 nsew
rlabel locali s -275 -35210 -229 -35086 2 VDD
port 41 nsew
rlabel locali s -471 -35215 -425 -35086 2 VDD
port 41 nsew
rlabel locali s -579 -35398 -545 -35211 2 VDD
port 41 nsew
rlabel locali s -775 -35398 -741 -35215 2 VDD
port 41 nsew
rlabel locali s -971 -35398 -937 -35215 2 VDD
port 41 nsew
rlabel locali s -584 -35211 -538 -35086 2 VDD
port 41 nsew
rlabel locali s -782 -35215 -736 -35086 2 VDD
port 41 nsew
rlabel locali s -971 -35215 -931 -35086 2 VDD
port 41 nsew
rlabel locali s -971 -35086 81 -35017 2 VDD
port 41 nsew
rlabel locali s -641 -35017 -48 -34979 2 VDD
port 41 nsew
rlabel locali s -2076 -35851 -1962 -34979 2 VDD
port 41 nsew
rlabel locali s -4649 -35952 -4526 -35816 2 VDD
port 41 nsew
rlabel locali s -2460 -35398 -2426 -35208 2 VDD
port 41 nsew
rlabel locali s -2656 -35398 -2622 -35220 2 VDD
port 41 nsew
rlabel locali s -2465 -35208 -2419 -35086 2 VDD
port 41 nsew
rlabel locali s -2662 -35220 -2616 -35086 2 VDD
port 41 nsew
rlabel locali s -2769 -35398 -2735 -35210 2 VDD
port 41 nsew
rlabel locali s -2965 -35398 -2931 -35215 2 VDD
port 41 nsew
rlabel locali s -2775 -35210 -2729 -35086 2 VDD
port 41 nsew
rlabel locali s -2971 -35215 -2925 -35086 2 VDD
port 41 nsew
rlabel locali s -3079 -35398 -3045 -35211 2 VDD
port 41 nsew
rlabel locali s -3275 -35398 -3241 -35215 2 VDD
port 41 nsew
rlabel locali s -3471 -35398 -3437 -35215 2 VDD
port 41 nsew
rlabel locali s -3084 -35211 -3038 -35086 2 VDD
port 41 nsew
rlabel locali s -3282 -35215 -3236 -35086 2 VDD
port 41 nsew
rlabel locali s -3471 -35215 -3431 -35086 2 VDD
port 41 nsew
rlabel locali s -3471 -35086 -2419 -35017 2 VDD
port 41 nsew
rlabel locali s -3157 -35017 -2564 -34979 2 VDD
port 41 nsew
rlabel locali s -4644 -35816 -4529 -34979 2 VDD
port 41 nsew
rlabel locali s -14690 -36596 -14601 -35673 2 VDD
port 41 nsew
rlabel locali s -23653 -37321 -23381 -36532 2 VDD
port 41 nsew
rlabel locali s -25449 -37321 -25383 -37251 2 VDD
port 41 nsew
rlabel locali s -25569 -37426 -25521 -37251 2 VDD
port 41 nsew
rlabel locali s -25569 -37251 -25383 -37239 2 VDD
port 41 nsew
rlabel locali s -26016 -37239 -25383 -37205 2 VDD
port 41 nsew
rlabel locali s -25569 -37205 -25383 -37192 2 VDD
port 41 nsew
rlabel locali s -25449 -37192 -25383 -37017 2 VDD
port 41 nsew
rlabel locali s -25569 -37192 -25521 -37017 2 VDD
port 41 nsew
rlabel locali s -25569 -37017 -25383 -37003 2 VDD
port 41 nsew
rlabel locali s -26016 -37003 -25383 -36969 2 VDD
port 41 nsew
rlabel locali s -25569 -36969 -25383 -36958 2 VDD
port 41 nsew
rlabel locali s -25449 -36958 -25383 -36780 2 VDD
port 41 nsew
rlabel locali s -25569 -36958 -25521 -36780 2 VDD
port 41 nsew
rlabel locali s -25569 -36780 -25383 -36767 2 VDD
port 41 nsew
rlabel locali s -26016 -36767 -25383 -36733 2 VDD
port 41 nsew
rlabel locali s -25569 -36733 -25383 -36721 2 VDD
port 41 nsew
rlabel locali s -25449 -36721 -25383 -36550 2 VDD
port 41 nsew
rlabel locali s -25569 -36721 -25521 -36550 2 VDD
port 41 nsew
rlabel locali s -25569 -36550 -25383 -36532 2 VDD
port 41 nsew
rlabel locali s -25569 -36532 -23381 -36531 2 VDD
port 41 nsew
rlabel locali s -26016 -36531 -23381 -36497 2 VDD
port 41 nsew
rlabel locali s -25569 -36497 -23381 -36491 2 VDD
port 41 nsew
rlabel locali s -25449 -36491 -23381 -36310 2 VDD
port 41 nsew
rlabel locali s -25569 -36491 -25521 -36310 2 VDD
port 41 nsew
rlabel locali s -25569 -36310 -23381 -36295 2 VDD
port 41 nsew
rlabel locali s -26016 -36295 -23381 -36261 2 VDD
port 41 nsew
rlabel locali s -25569 -36261 -23381 -36260 2 VDD
port 41 nsew
rlabel locali s -18844 -36000 -18810 -35834 2 VDD
port 41 nsew
rlabel locali s -19040 -36000 -19006 -35834 2 VDD
port 41 nsew
rlabel locali s -19236 -36000 -19202 -35834 2 VDD
port 41 nsew
rlabel locali s -19432 -36000 -19398 -35834 2 VDD
port 41 nsew
rlabel locali s -19649 -36201 -19615 -35834 2 VDD
port 41 nsew
rlabel locali s -19649 -35834 -18762 -35790 2 VDD
port 41 nsew
rlabel locali s -19845 -36201 -19811 -35790 2 VDD
port 41 nsew
rlabel locali s -20041 -36201 -20007 -35790 2 VDD
port 41 nsew
rlabel locali s -20093 -35790 -18762 -35735 2 VDD
port 41 nsew
rlabel locali s -20093 -35735 -18766 -35673 2 VDD
port 41 nsew
rlabel locali s -20714 -35979 -20680 -35687 2 VDD
port 41 nsew
rlabel locali s -20910 -35979 -20876 -35687 2 VDD
port 41 nsew
rlabel locali s -20915 -35687 -20670 -35673 2 VDD
port 41 nsew
rlabel locali s -21452 -35979 -21418 -35683 2 VDD
port 41 nsew
rlabel locali s -21648 -35979 -21614 -35683 2 VDD
port 41 nsew
rlabel locali s -21844 -35979 -21810 -35683 2 VDD
port 41 nsew
rlabel locali s -22040 -35979 -22006 -35683 2 VDD
port 41 nsew
rlabel locali s -23653 -36260 -23381 -35732 2 VDD
port 41 nsew
rlabel locali s -25569 -36260 -25383 -36251 2 VDD
port 41 nsew
rlabel locali s -25449 -36251 -25383 -36072 2 VDD
port 41 nsew
rlabel locali s -25569 -36251 -25521 -36072 2 VDD
port 41 nsew
rlabel locali s -25569 -36072 -25383 -36059 2 VDD
port 41 nsew
rlabel locali s -26016 -36059 -25383 -36025 2 VDD
port 41 nsew
rlabel locali s -25569 -36025 -25383 -36013 2 VDD
port 41 nsew
rlabel locali s -25449 -36013 -25383 -35836 2 VDD
port 41 nsew
rlabel locali s -25569 -36013 -25521 -35836 2 VDD
port 41 nsew
rlabel locali s -25569 -35836 -25383 -35823 2 VDD
port 41 nsew
rlabel locali s -26016 -35823 -25383 -35789 2 VDD
port 41 nsew
rlabel locali s -25569 -35789 -25383 -35777 2 VDD
port 41 nsew
rlabel locali s -25449 -35777 -25383 -35732 2 VDD
port 41 nsew
rlabel locali s -25449 -35732 -23381 -35683 2 VDD
port 41 nsew
rlabel locali s -25449 -35683 -21418 -35673 2 VDD
port 41 nsew
rlabel locali s -25449 -35673 -14601 -35605 2 VDD
port 41 nsew
rlabel locali s -25569 -35777 -25521 -35605 2 VDD
port 41 nsew
rlabel locali s -4960 -35398 -4926 -35208 2 VDD
port 41 nsew
rlabel locali s -5156 -35398 -5122 -35220 2 VDD
port 41 nsew
rlabel locali s -4965 -35208 -4919 -35086 2 VDD
port 41 nsew
rlabel locali s -5162 -35220 -5116 -35086 2 VDD
port 41 nsew
rlabel locali s -5269 -35398 -5235 -35210 2 VDD
port 41 nsew
rlabel locali s -5465 -35398 -5431 -35215 2 VDD
port 41 nsew
rlabel locali s -5275 -35210 -5229 -35086 2 VDD
port 41 nsew
rlabel locali s -5471 -35215 -5425 -35086 2 VDD
port 41 nsew
rlabel locali s -5579 -35398 -5545 -35211 2 VDD
port 41 nsew
rlabel locali s -5775 -35398 -5741 -35215 2 VDD
port 41 nsew
rlabel locali s -5971 -35398 -5937 -35215 2 VDD
port 41 nsew
rlabel locali s -5584 -35211 -5538 -35086 2 VDD
port 41 nsew
rlabel locali s -5782 -35215 -5736 -35086 2 VDD
port 41 nsew
rlabel locali s -5971 -35215 -5931 -35086 2 VDD
port 41 nsew
rlabel locali s -5971 -35086 -4919 -34979 2 VDD
port 41 nsew
rlabel locali s -7460 -35602 -7426 -35012 2 VDD
port 41 nsew
rlabel locali s -7336 -34979 8126 -34886 8 VDD
port 41 nsew
rlabel locali s -7466 -35012 -7421 -34886 2 VDD
port 41 nsew
rlabel locali s -7656 -35602 -7622 -35009 2 VDD
port 41 nsew
rlabel locali s -8079 -35602 -8045 -35010 2 VDD
port 41 nsew
rlabel locali s -25569 -35605 -14601 -35587 2 VDD
port 41 nsew
rlabel locali s -26016 -35587 -14601 -35553 2 VDD
port 41 nsew
rlabel locali s -25569 -35553 -14601 -35546 2 VDD
port 41 nsew
rlabel locali s -25449 -35546 -14601 -35460 2 VDD
port 41 nsew
rlabel locali s -7661 -35009 -7616 -34886 2 VDD
port 41 nsew
rlabel locali s -8083 -35010 -8038 -34886 2 VDD
port 41 nsew
rlabel locali s -10512 -35192 -10478 -34901 2 VDD
port 41 nsew
rlabel locali s -10708 -35192 -10674 -34901 2 VDD
port 41 nsew
rlabel locali s -10904 -35192 -10870 -34901 2 VDD
port 41 nsew
rlabel locali s -11349 -35192 -11315 -34901 2 VDD
port 41 nsew
rlabel locali s -11545 -35192 -11511 -34901 2 VDD
port 41 nsew
rlabel locali s -11741 -35192 -11707 -34901 2 VDD
port 41 nsew
rlabel locali s -13212 -35192 -13178 -34901 2 VDD
port 41 nsew
rlabel locali s -13408 -35192 -13374 -34901 2 VDD
port 41 nsew
rlabel locali s -13604 -35192 -13570 -34901 2 VDD
port 41 nsew
rlabel locali s -14049 -35192 -14015 -34901 2 VDD
port 41 nsew
rlabel locali s -14245 -35192 -14211 -34901 2 VDD
port 41 nsew
rlabel locali s -14441 -35192 -14407 -34901 2 VDD
port 41 nsew
rlabel locali s -14690 -35460 -14601 -34901 2 VDD
port 41 nsew
rlabel locali s -12219 -34901 -10417 -34896 2 VDD
port 41 nsew
rlabel locali s -14690 -34901 -13117 -34896 2 VDD
port 41 nsew
rlabel locali s -14690 -34896 -9465 -34886 2 VDD
port 41 nsew
rlabel locali s -14690 -34886 8126 -34833 2 VDD
port 41 nsew
rlabel locali s -25449 -35460 -25383 -35128 2 VDD
port 41 nsew
rlabel locali s -25569 -35546 -25521 -35351 2 VDD
port 41 nsew
rlabel locali s -26016 -35351 -25521 -35317 2 VDD
port 41 nsew
rlabel locali s -25569 -35317 -25521 -35128 2 VDD
port 41 nsew
rlabel locali s -25569 -35128 -25383 -35115 2 VDD
port 41 nsew
rlabel locali s -26016 -35115 -25383 -35081 2 VDD
port 41 nsew
rlabel locali s -25569 -35081 -25383 -35069 2 VDD
port 41 nsew
rlabel locali s -9665 -34833 8126 -34797 2 VDD
port 41 nsew
rlabel locali s -7334 -34797 8126 -34786 8 VDD
port 41 nsew
rlabel locali s 25923 -33752 87071 -33632 8 VDD
port 41 nsew
rlabel locali s 6895 -34786 7657 -33632 8 VDD
port 41 nsew
rlabel locali s -25449 -35069 -25383 -34081 2 VDD
port 41 nsew
rlabel locali s -25569 -35069 -25521 -34879 2 VDD
port 41 nsew
rlabel locali s -26016 -34879 -25521 -34845 2 VDD
port 41 nsew
rlabel locali s -25569 -34845 -25521 -34643 2 VDD
port 41 nsew
rlabel locali s -26016 -34643 -25521 -34609 2 VDD
port 41 nsew
rlabel locali s -25569 -34609 -25521 -34407 2 VDD
port 41 nsew
rlabel locali s -26016 -34407 -25521 -34373 2 VDD
port 41 nsew
rlabel locali s -25569 -34373 -25521 -34171 2 VDD
port 41 nsew
rlabel locali s -26016 -34171 -25521 -34137 2 VDD
port 41 nsew
rlabel locali s -25569 -34137 -25521 -33971 2 VDD
port 41 nsew
rlabel locali s 6895 -33632 87071 -32870 8 VDD
port 41 nsew
rlabel locali s 25923 -32870 87071 -32649 8 VDD
port 41 nsew
rlabel locali s 83333 -32649 86302 -31308 8 VDD
port 41 nsew
rlabel locali s 83333 -31308 98798 -28339 8 VDD
port 41 nsew
rlabel locali s 95829 -28339 98798 -15816 8 VDD
port 41 nsew
rlabel locali s -7534 -27749 7428 -27556 2 VDD
port 41 nsew
rlabel locali s -22775 -27591 -20173 -27582 2 VDD
port 41 nsew
rlabel locali s 6331 -27556 7383 -27449 8 VDD
port 41 nsew
rlabel locali s 3608 -27556 4201 -27518 8 VDD
port 41 nsew
rlabel locali s 1195 -27556 1788 -27518 8 VDD
port 41 nsew
rlabel locali s 11445 -27333 16670 -27270 8 VDD
port 41 nsew
rlabel locali s 7337 -27449 7383 -27327 8 VDD
port 41 nsew
rlabel locali s 15097 -27270 16670 -27265 8 VDD
port 41 nsew
rlabel locali s 12397 -27270 14199 -27265 8 VDD
port 41 nsew
rlabel locali s 86430 -25574 86464 -24982 8 VDD
port 41 nsew
rlabel locali s 86870 -24877 87009 -24849 8 VDD
port 41 nsew
rlabel locali s 86870 -24849 87082 -24710 8 VDD
port 41 nsew
rlabel locali s 86620 -24864 86699 -24839 8 VDD
port 41 nsew
rlabel locali s 86423 -24982 86468 -24858 8 VDD
port 41 nsew
rlabel locali s 86007 -25574 86041 -24981 8 VDD
port 41 nsew
rlabel locali s 85811 -25574 85845 -24984 8 VDD
port 41 nsew
rlabel locali s 85561 -25162 85595 -24996 8 VDD
port 41 nsew
rlabel locali s 85365 -25162 85399 -24996 8 VDD
port 41 nsew
rlabel locali s 85169 -25162 85203 -24996 8 VDD
port 41 nsew
rlabel locali s 84973 -25162 85007 -24996 8 VDD
port 41 nsew
rlabel locali s 84756 -25363 84790 -24996 8 VDD
port 41 nsew
rlabel locali s 86001 -24981 86046 -24858 8 VDD
port 41 nsew
rlabel locali s 85806 -24984 85851 -24858 8 VDD
port 41 nsew
rlabel locali s 84756 -24996 85643 -24946 8 VDD
port 41 nsew
rlabel locali s 84560 -25363 84594 -24946 8 VDD
port 41 nsew
rlabel locali s 84364 -25363 84398 -24946 8 VDD
port 41 nsew
rlabel locali s 82762 -25543 82796 -24951 8 VDD
port 41 nsew
rlabel locali s 84354 -24946 85643 -24897 8 VDD
port 41 nsew
rlabel locali s 84354 -24897 84796 -24882 8 VDD
port 41 nsew
rlabel locali s 85800 -24858 86569 -24839 8 VDD
port 41 nsew
rlabel locali s 85800 -24839 86699 -24834 8 VDD
port 41 nsew
rlabel locali s 84793 -24848 84982 -24841 8 VDD
port 41 nsew
rlabel locali s 84756 -24841 84982 -24834 8 VDD
port 41 nsew
rlabel locali s 84354 -24834 86699 -24792 8 VDD
port 41 nsew
rlabel locali s 82755 -24951 82800 -24827 8 VDD
port 41 nsew
rlabel locali s 82339 -25543 82373 -24950 8 VDD
port 41 nsew
rlabel locali s 82143 -25543 82177 -24953 8 VDD
port 41 nsew
rlabel locali s 81893 -25131 81927 -24965 8 VDD
port 41 nsew
rlabel locali s 81697 -25131 81731 -24965 8 VDD
port 41 nsew
rlabel locali s 81501 -25131 81535 -24965 8 VDD
port 41 nsew
rlabel locali s 81305 -25131 81339 -24965 8 VDD
port 41 nsew
rlabel locali s 81088 -25332 81122 -24965 8 VDD
port 41 nsew
rlabel locali s 82333 -24950 82378 -24827 8 VDD
port 41 nsew
rlabel locali s 82138 -24953 82183 -24827 8 VDD
port 41 nsew
rlabel locali s 81088 -24965 81975 -24915 8 VDD
port 41 nsew
rlabel locali s 80892 -25332 80926 -24915 8 VDD
port 41 nsew
rlabel locali s 80696 -25332 80730 -24915 8 VDD
port 41 nsew
rlabel locali s 77066 -25612 77100 -25020 8 VDD
port 41 nsew
rlabel locali s 80686 -24915 81975 -24866 8 VDD
port 41 nsew
rlabel locali s 77506 -24915 77645 -24887 8 VDD
port 41 nsew
rlabel locali s 80686 -24866 81128 -24851 8 VDD
port 41 nsew
rlabel locali s 82132 -24827 82901 -24803 8 VDD
port 41 nsew
rlabel locali s 81125 -24817 81314 -24810 8 VDD
port 41 nsew
rlabel locali s 81088 -24810 81314 -24803 8 VDD
port 41 nsew
rlabel locali s 86520 -24792 86699 -24756 8 VDD
port 41 nsew
rlabel locali s 84354 -24792 86465 -24781 8 VDD
port 41 nsew
rlabel locali s 86620 -24756 86699 -24725 8 VDD
port 41 nsew
rlabel locali s 83553 -24781 86465 -24715 8 VDD
port 41 nsew
rlabel locali s 86960 -24710 87082 -23714 8 VDD
port 41 nsew
rlabel locali s 84354 -24715 86465 -24681 8 VDD
port 41 nsew
rlabel locali s 85352 -24681 85970 -24664 8 VDD
port 41 nsew
rlabel locali s 85352 -24664 85795 -24635 8 VDD
port 41 nsew
rlabel locali s 85353 -24635 85795 -24621 8 VDD
port 41 nsew
rlabel locali s 85353 -24621 86642 -24572 8 VDD
port 41 nsew
rlabel locali s 85755 -24572 86642 -24522 8 VDD
port 41 nsew
rlabel locali s 86560 -24522 86594 -24356 8 VDD
port 41 nsew
rlabel locali s 86364 -24522 86398 -24356 8 VDD
port 41 nsew
rlabel locali s 86168 -24522 86202 -24356 8 VDD
port 41 nsew
rlabel locali s 85972 -24522 86006 -24356 8 VDD
port 41 nsew
rlabel locali s 85755 -24522 85789 -24155 8 VDD
port 41 nsew
rlabel locali s 85559 -24572 85593 -24155 8 VDD
port 41 nsew
rlabel locali s 85363 -24572 85397 -24155 8 VDD
port 41 nsew
rlabel locali s 84524 -24681 84696 -24491 8 VDD
port 41 nsew
rlabel locali s 84342 -24491 85060 -24392 8 VDD
port 41 nsew
rlabel locali s 84978 -24392 85012 -24126 8 VDD
port 41 nsew
rlabel locali s 84782 -24392 84816 -24126 8 VDD
port 41 nsew
rlabel locali s 84586 -24392 84620 -24126 8 VDD
port 41 nsew
rlabel locali s 84390 -24392 84424 -24126 8 VDD
port 41 nsew
rlabel locali s 86450 -23714 87082 -23592 8 VDD
port 41 nsew
rlabel locali s 86450 -23592 86572 -21195 8 VDD
port 41 nsew
rlabel locali s 83553 -24715 83619 -23385 8 VDD
port 41 nsew
rlabel locali s 83200 -24799 83284 -24686 8 VDD
port 41 nsew
rlabel locali s 80686 -24803 82901 -24761 8 VDD
port 41 nsew
rlabel locali s 83217 -24686 83283 -23385 8 VDD
port 41 nsew
rlabel locali s 80686 -24761 82797 -24650 8 VDD
port 41 nsew
rlabel locali s 77506 -24887 77718 -24748 8 VDD
port 41 nsew
rlabel locali s 77256 -24902 77335 -24877 8 VDD
port 41 nsew
rlabel locali s 77059 -25020 77104 -24896 8 VDD
port 41 nsew
rlabel locali s 76643 -25612 76677 -25019 8 VDD
port 41 nsew
rlabel locali s 76447 -25612 76481 -25022 8 VDD
port 41 nsew
rlabel locali s 76197 -25200 76231 -25034 8 VDD
port 41 nsew
rlabel locali s 76001 -25200 76035 -25034 8 VDD
port 41 nsew
rlabel locali s 75805 -25200 75839 -25034 8 VDD
port 41 nsew
rlabel locali s 75609 -25200 75643 -25034 8 VDD
port 41 nsew
rlabel locali s 75392 -25401 75426 -25034 8 VDD
port 41 nsew
rlabel locali s 76637 -25019 76682 -24896 8 VDD
port 41 nsew
rlabel locali s 76442 -25022 76487 -24896 8 VDD
port 41 nsew
rlabel locali s 75392 -25034 76279 -24984 8 VDD
port 41 nsew
rlabel locali s 75196 -25401 75230 -24984 8 VDD
port 41 nsew
rlabel locali s 75000 -25401 75034 -24984 8 VDD
port 41 nsew
rlabel locali s 73398 -25581 73432 -24989 8 VDD
port 41 nsew
rlabel locali s 74990 -24984 76279 -24935 8 VDD
port 41 nsew
rlabel locali s 74990 -24935 75432 -24920 8 VDD
port 41 nsew
rlabel locali s 76436 -24896 77205 -24877 8 VDD
port 41 nsew
rlabel locali s 76436 -24877 77335 -24872 8 VDD
port 41 nsew
rlabel locali s 75429 -24886 75618 -24879 8 VDD
port 41 nsew
rlabel locali s 75392 -24879 75618 -24872 8 VDD
port 41 nsew
rlabel locali s 74990 -24872 77335 -24830 8 VDD
port 41 nsew
rlabel locali s 73391 -24989 73436 -24865 8 VDD
port 41 nsew
rlabel locali s 72975 -25581 73009 -24988 8 VDD
port 41 nsew
rlabel locali s 72779 -25581 72813 -24991 8 VDD
port 41 nsew
rlabel locali s 72529 -25169 72563 -25003 8 VDD
port 41 nsew
rlabel locali s 72333 -25169 72367 -25003 8 VDD
port 41 nsew
rlabel locali s 72137 -25169 72171 -25003 8 VDD
port 41 nsew
rlabel locali s 71941 -25169 71975 -25003 8 VDD
port 41 nsew
rlabel locali s 71724 -25370 71758 -25003 8 VDD
port 41 nsew
rlabel locali s 72969 -24988 73014 -24865 8 VDD
port 41 nsew
rlabel locali s 72774 -24991 72819 -24865 8 VDD
port 41 nsew
rlabel locali s 71724 -25003 72611 -24953 8 VDD
port 41 nsew
rlabel locali s 71528 -25370 71562 -24953 8 VDD
port 41 nsew
rlabel locali s 71332 -25370 71366 -24953 8 VDD
port 41 nsew
rlabel locali s 67913 -25629 67947 -25037 8 VDD
port 41 nsew
rlabel locali s 71322 -24953 72611 -24904 8 VDD
port 41 nsew
rlabel locali s 68353 -24932 68492 -24904 8 VDD
port 41 nsew
rlabel locali s 71322 -24904 71764 -24889 8 VDD
port 41 nsew
rlabel locali s 72768 -24865 73537 -24841 8 VDD
port 41 nsew
rlabel locali s 71761 -24855 71950 -24848 8 VDD
port 41 nsew
rlabel locali s 71724 -24848 71950 -24841 8 VDD
port 41 nsew
rlabel locali s 77156 -24830 77335 -24794 8 VDD
port 41 nsew
rlabel locali s 74990 -24830 77101 -24819 8 VDD
port 41 nsew
rlabel locali s 77256 -24794 77335 -24763 8 VDD
port 41 nsew
rlabel locali s 74189 -24819 77101 -24753 8 VDD
port 41 nsew
rlabel locali s 81684 -24650 82302 -24633 8 VDD
port 41 nsew
rlabel locali s 81684 -24633 82127 -24604 8 VDD
port 41 nsew
rlabel locali s 81685 -24604 82127 -24590 8 VDD
port 41 nsew
rlabel locali s 81685 -24590 82974 -24541 8 VDD
port 41 nsew
rlabel locali s 82087 -24541 82974 -24491 8 VDD
port 41 nsew
rlabel locali s 82892 -24491 82926 -24325 8 VDD
port 41 nsew
rlabel locali s 82696 -24491 82730 -24325 8 VDD
port 41 nsew
rlabel locali s 82500 -24491 82534 -24325 8 VDD
port 41 nsew
rlabel locali s 82304 -24491 82338 -24325 8 VDD
port 41 nsew
rlabel locali s 82087 -24491 82121 -24124 8 VDD
port 41 nsew
rlabel locali s 81891 -24541 81925 -24124 8 VDD
port 41 nsew
rlabel locali s 81695 -24541 81729 -24124 8 VDD
port 41 nsew
rlabel locali s 80856 -24650 81028 -24460 8 VDD
port 41 nsew
rlabel locali s 80674 -24460 81392 -24361 8 VDD
port 41 nsew
rlabel locali s 81310 -24361 81344 -24095 8 VDD
port 41 nsew
rlabel locali s 81114 -24361 81148 -24095 8 VDD
port 41 nsew
rlabel locali s 80918 -24361 80952 -24095 8 VDD
port 41 nsew
rlabel locali s 80722 -24361 80756 -24095 8 VDD
port 41 nsew
rlabel locali s 77596 -24748 77718 -23752 8 VDD
port 41 nsew
rlabel locali s 74990 -24753 77101 -24719 8 VDD
port 41 nsew
rlabel locali s 75988 -24719 76606 -24702 8 VDD
port 41 nsew
rlabel locali s 75988 -24702 76431 -24673 8 VDD
port 41 nsew
rlabel locali s 75989 -24673 76431 -24659 8 VDD
port 41 nsew
rlabel locali s 75989 -24659 77278 -24610 8 VDD
port 41 nsew
rlabel locali s 76391 -24610 77278 -24560 8 VDD
port 41 nsew
rlabel locali s 77196 -24560 77230 -24394 8 VDD
port 41 nsew
rlabel locali s 77000 -24560 77034 -24394 8 VDD
port 41 nsew
rlabel locali s 76804 -24560 76838 -24394 8 VDD
port 41 nsew
rlabel locali s 76608 -24560 76642 -24394 8 VDD
port 41 nsew
rlabel locali s 76391 -24560 76425 -24193 8 VDD
port 41 nsew
rlabel locali s 76195 -24610 76229 -24193 8 VDD
port 41 nsew
rlabel locali s 75999 -24610 76033 -24193 8 VDD
port 41 nsew
rlabel locali s 75160 -24719 75332 -24529 8 VDD
port 41 nsew
rlabel locali s 74978 -24529 75696 -24430 8 VDD
port 41 nsew
rlabel locali s 75614 -24430 75648 -24164 8 VDD
port 41 nsew
rlabel locali s 75418 -24430 75452 -24164 8 VDD
port 41 nsew
rlabel locali s 75222 -24430 75256 -24164 8 VDD
port 41 nsew
rlabel locali s 75026 -24430 75060 -24164 8 VDD
port 41 nsew
rlabel locali s 77086 -23752 77718 -23630 8 VDD
port 41 nsew
rlabel locali s 83217 -23385 83619 -23319 8 VDD
port 41 nsew
rlabel locali s 85488 -21648 85522 -21356 8 VDD
port 41 nsew
rlabel locali s 85292 -21648 85326 -21358 8 VDD
port 41 nsew
rlabel locali s 85064 -21848 85098 -21373 8 VDD
port 41 nsew
rlabel locali s 84934 -21848 84968 -21376 8 VDD
port 41 nsew
rlabel locali s 85483 -21356 85526 -21196 8 VDD
port 41 nsew
rlabel locali s 85286 -21358 85329 -21196 8 VDD
port 41 nsew
rlabel locali s 85055 -21373 85105 -21196 8 VDD
port 41 nsew
rlabel locali s 84929 -21376 84979 -21196 8 VDD
port 41 nsew
rlabel locali s 84339 -21848 84373 -21353 8 VDD
port 41 nsew
rlabel locali s 84143 -21848 84177 -21355 8 VDD
port 41 nsew
rlabel locali s 82770 -22090 82804 -21498 8 VDD
port 41 nsew
rlabel locali s 83210 -21393 83308 -21387 8 VDD
port 41 nsew
rlabel locali s 84337 -21353 84375 -21196 8 VDD
port 41 nsew
rlabel locali s 84140 -21355 84178 -21260 8 VDD
port 41 nsew
rlabel locali s 83210 -21387 83890 -21270 8 VDD
port 41 nsew
rlabel locali s 82982 -21381 83044 -21367 8 VDD
port 41 nsew
rlabel locali s 82763 -21498 82808 -21374 8 VDD
port 41 nsew
rlabel locali s 82347 -22090 82381 -21497 8 VDD
port 41 nsew
rlabel locali s 82151 -22090 82185 -21500 8 VDD
port 41 nsew
rlabel locali s 81901 -21678 81935 -21512 8 VDD
port 41 nsew
rlabel locali s 81705 -21678 81739 -21512 8 VDD
port 41 nsew
rlabel locali s 81509 -21678 81543 -21512 8 VDD
port 41 nsew
rlabel locali s 81313 -21678 81347 -21512 8 VDD
port 41 nsew
rlabel locali s 81096 -21879 81130 -21512 8 VDD
port 41 nsew
rlabel locali s 82341 -21497 82386 -21374 8 VDD
port 41 nsew
rlabel locali s 82146 -21500 82191 -21374 8 VDD
port 41 nsew
rlabel locali s 81096 -21512 81983 -21462 8 VDD
port 41 nsew
rlabel locali s 80900 -21879 80934 -21462 8 VDD
port 41 nsew
rlabel locali s 80704 -21879 80738 -21462 8 VDD
port 41 nsew
rlabel locali s 80694 -21462 81983 -21413 8 VDD
port 41 nsew
rlabel locali s 80694 -21413 81136 -21398 8 VDD
port 41 nsew
rlabel locali s 82140 -21374 82909 -21367 8 VDD
port 41 nsew
rlabel locali s 82140 -21367 83044 -21350 8 VDD
port 41 nsew
rlabel locali s 81133 -21364 81322 -21357 8 VDD
port 41 nsew
rlabel locali s 81096 -21357 81322 -21350 8 VDD
port 41 nsew
rlabel locali s 80694 -21350 83044 -21315 8 VDD
port 41 nsew
rlabel locali s 82982 -21315 83044 -21287 8 VDD
port 41 nsew
rlabel locali s 80694 -21315 82909 -21308 8 VDD
port 41 nsew
rlabel locali s 80694 -21308 82805 -21294 8 VDD
port 41 nsew
rlabel locali s 77086 -23630 77208 -21294 8 VDD
port 41 nsew
rlabel locali s 74189 -24753 74255 -23423 8 VDD
port 41 nsew
rlabel locali s 73836 -24837 73920 -24724 8 VDD
port 41 nsew
rlabel locali s 71322 -24841 73537 -24799 8 VDD
port 41 nsew
rlabel locali s 73853 -24724 73919 -23423 8 VDD
port 41 nsew
rlabel locali s 71322 -24799 73433 -24688 8 VDD
port 41 nsew
rlabel locali s 68353 -24904 68565 -24765 8 VDD
port 41 nsew
rlabel locali s 68103 -24919 68182 -24894 8 VDD
port 41 nsew
rlabel locali s 67906 -25037 67951 -24913 8 VDD
port 41 nsew
rlabel locali s 67490 -25629 67524 -25036 8 VDD
port 41 nsew
rlabel locali s 67294 -25629 67328 -25039 8 VDD
port 41 nsew
rlabel locali s 67044 -25217 67078 -25051 8 VDD
port 41 nsew
rlabel locali s 66848 -25217 66882 -25051 8 VDD
port 41 nsew
rlabel locali s 66652 -25217 66686 -25051 8 VDD
port 41 nsew
rlabel locali s 66456 -25217 66490 -25051 8 VDD
port 41 nsew
rlabel locali s 66239 -25418 66273 -25051 8 VDD
port 41 nsew
rlabel locali s 67484 -25036 67529 -24913 8 VDD
port 41 nsew
rlabel locali s 67289 -25039 67334 -24913 8 VDD
port 41 nsew
rlabel locali s 66239 -25051 67126 -25001 8 VDD
port 41 nsew
rlabel locali s 66043 -25418 66077 -25001 8 VDD
port 41 nsew
rlabel locali s 65847 -25418 65881 -25001 8 VDD
port 41 nsew
rlabel locali s 64245 -25598 64279 -25006 8 VDD
port 41 nsew
rlabel locali s 65837 -25001 67126 -24952 8 VDD
port 41 nsew
rlabel locali s 65837 -24952 66279 -24937 8 VDD
port 41 nsew
rlabel locali s 67283 -24913 68052 -24894 8 VDD
port 41 nsew
rlabel locali s 67283 -24894 68182 -24889 8 VDD
port 41 nsew
rlabel locali s 66276 -24903 66465 -24896 8 VDD
port 41 nsew
rlabel locali s 66239 -24896 66465 -24889 8 VDD
port 41 nsew
rlabel locali s 65837 -24889 68182 -24847 8 VDD
port 41 nsew
rlabel locali s 64238 -25006 64283 -24882 8 VDD
port 41 nsew
rlabel locali s 63822 -25598 63856 -25005 8 VDD
port 41 nsew
rlabel locali s 63626 -25598 63660 -25008 8 VDD
port 41 nsew
rlabel locali s 63376 -25186 63410 -25020 8 VDD
port 41 nsew
rlabel locali s 63180 -25186 63214 -25020 8 VDD
port 41 nsew
rlabel locali s 62984 -25186 63018 -25020 8 VDD
port 41 nsew
rlabel locali s 62788 -25186 62822 -25020 8 VDD
port 41 nsew
rlabel locali s 62571 -25387 62605 -25020 8 VDD
port 41 nsew
rlabel locali s 63816 -25005 63861 -24882 8 VDD
port 41 nsew
rlabel locali s 63621 -25008 63666 -24882 8 VDD
port 41 nsew
rlabel locali s 62571 -25020 63458 -24970 8 VDD
port 41 nsew
rlabel locali s 62375 -25387 62409 -24970 8 VDD
port 41 nsew
rlabel locali s 62179 -25387 62213 -24970 8 VDD
port 41 nsew
rlabel locali s 59159 -25695 59193 -25103 8 VDD
port 41 nsew
rlabel locali s 59599 -24998 59738 -24970 8 VDD
port 41 nsew
rlabel locali s 62169 -24970 63458 -24921 8 VDD
port 41 nsew
rlabel locali s 62169 -24921 62611 -24906 8 VDD
port 41 nsew
rlabel locali s 63615 -24882 64384 -24858 8 VDD
port 41 nsew
rlabel locali s 62608 -24872 62797 -24865 8 VDD
port 41 nsew
rlabel locali s 62571 -24865 62797 -24858 8 VDD
port 41 nsew
rlabel locali s 68003 -24847 68182 -24811 8 VDD
port 41 nsew
rlabel locali s 65837 -24847 67948 -24836 8 VDD
port 41 nsew
rlabel locali s 68103 -24811 68182 -24780 8 VDD
port 41 nsew
rlabel locali s 65036 -24836 67948 -24770 8 VDD
port 41 nsew
rlabel locali s 72320 -24688 72938 -24671 8 VDD
port 41 nsew
rlabel locali s 72320 -24671 72763 -24642 8 VDD
port 41 nsew
rlabel locali s 72321 -24642 72763 -24628 8 VDD
port 41 nsew
rlabel locali s 72321 -24628 73610 -24579 8 VDD
port 41 nsew
rlabel locali s 72723 -24579 73610 -24529 8 VDD
port 41 nsew
rlabel locali s 73528 -24529 73562 -24363 8 VDD
port 41 nsew
rlabel locali s 73332 -24529 73366 -24363 8 VDD
port 41 nsew
rlabel locali s 73136 -24529 73170 -24363 8 VDD
port 41 nsew
rlabel locali s 72940 -24529 72974 -24363 8 VDD
port 41 nsew
rlabel locali s 72723 -24529 72757 -24162 8 VDD
port 41 nsew
rlabel locali s 72527 -24579 72561 -24162 8 VDD
port 41 nsew
rlabel locali s 72331 -24579 72365 -24162 8 VDD
port 41 nsew
rlabel locali s 71492 -24688 71664 -24498 8 VDD
port 41 nsew
rlabel locali s 71310 -24498 72028 -24399 8 VDD
port 41 nsew
rlabel locali s 71946 -24399 71980 -24133 8 VDD
port 41 nsew
rlabel locali s 71750 -24399 71784 -24133 8 VDD
port 41 nsew
rlabel locali s 71554 -24399 71588 -24133 8 VDD
port 41 nsew
rlabel locali s 71358 -24399 71392 -24133 8 VDD
port 41 nsew
rlabel locali s 68443 -24765 68565 -23769 8 VDD
port 41 nsew
rlabel locali s 65837 -24770 67948 -24736 8 VDD
port 41 nsew
rlabel locali s 66835 -24736 67453 -24719 8 VDD
port 41 nsew
rlabel locali s 66835 -24719 67278 -24690 8 VDD
port 41 nsew
rlabel locali s 66836 -24690 67278 -24676 8 VDD
port 41 nsew
rlabel locali s 66836 -24676 68125 -24627 8 VDD
port 41 nsew
rlabel locali s 67238 -24627 68125 -24577 8 VDD
port 41 nsew
rlabel locali s 68043 -24577 68077 -24411 8 VDD
port 41 nsew
rlabel locali s 67847 -24577 67881 -24411 8 VDD
port 41 nsew
rlabel locali s 67651 -24577 67685 -24411 8 VDD
port 41 nsew
rlabel locali s 67455 -24577 67489 -24411 8 VDD
port 41 nsew
rlabel locali s 67238 -24577 67272 -24210 8 VDD
port 41 nsew
rlabel locali s 67042 -24627 67076 -24210 8 VDD
port 41 nsew
rlabel locali s 66846 -24627 66880 -24210 8 VDD
port 41 nsew
rlabel locali s 66007 -24736 66179 -24546 8 VDD
port 41 nsew
rlabel locali s 65825 -24546 66543 -24447 8 VDD
port 41 nsew
rlabel locali s 66461 -24447 66495 -24181 8 VDD
port 41 nsew
rlabel locali s 66265 -24447 66299 -24181 8 VDD
port 41 nsew
rlabel locali s 66069 -24447 66103 -24181 8 VDD
port 41 nsew
rlabel locali s 65873 -24447 65907 -24181 8 VDD
port 41 nsew
rlabel locali s 67933 -23769 68565 -23647 8 VDD
port 41 nsew
rlabel locali s 73853 -23423 74255 -23357 8 VDD
port 41 nsew
rlabel locali s 76124 -21686 76158 -21394 8 VDD
port 41 nsew
rlabel locali s 75928 -21686 75962 -21396 8 VDD
port 41 nsew
rlabel locali s 75700 -21886 75734 -21411 8 VDD
port 41 nsew
rlabel locali s 75570 -21886 75604 -21414 8 VDD
port 41 nsew
rlabel locali s 76119 -21394 76162 -21294 8 VDD
port 41 nsew
rlabel locali s 83773 -21270 83890 -21260 8 VDD
port 41 nsew
rlabel locali s 83210 -21270 83308 -21267 8 VDD
port 41 nsew
rlabel locali s 83773 -21260 84178 -21196 8 VDD
port 41 nsew
rlabel locali s 76119 -21294 82805 -21234 8 VDD
port 41 nsew
rlabel locali s 75922 -21396 75965 -21234 8 VDD
port 41 nsew
rlabel locali s 75691 -21411 75741 -21234 8 VDD
port 41 nsew
rlabel locali s 75565 -21414 75615 -21234 8 VDD
port 41 nsew
rlabel locali s 74975 -21886 75009 -21391 8 VDD
port 41 nsew
rlabel locali s 74779 -21886 74813 -21393 8 VDD
port 41 nsew
rlabel locali s 73406 -22128 73440 -21536 8 VDD
port 41 nsew
rlabel locali s 73846 -21431 73944 -21425 8 VDD
port 41 nsew
rlabel locali s 74973 -21391 75011 -21234 8 VDD
port 41 nsew
rlabel locali s 74776 -21393 74814 -21298 8 VDD
port 41 nsew
rlabel locali s 73846 -21425 74526 -21308 8 VDD
port 41 nsew
rlabel locali s 73618 -21419 73680 -21405 8 VDD
port 41 nsew
rlabel locali s 73399 -21536 73444 -21412 8 VDD
port 41 nsew
rlabel locali s 72983 -22128 73017 -21535 8 VDD
port 41 nsew
rlabel locali s 72787 -22128 72821 -21538 8 VDD
port 41 nsew
rlabel locali s 72537 -21716 72571 -21550 8 VDD
port 41 nsew
rlabel locali s 72341 -21716 72375 -21550 8 VDD
port 41 nsew
rlabel locali s 72145 -21716 72179 -21550 8 VDD
port 41 nsew
rlabel locali s 71949 -21716 71983 -21550 8 VDD
port 41 nsew
rlabel locali s 71732 -21917 71766 -21550 8 VDD
port 41 nsew
rlabel locali s 72977 -21535 73022 -21412 8 VDD
port 41 nsew
rlabel locali s 72782 -21538 72827 -21412 8 VDD
port 41 nsew
rlabel locali s 71732 -21550 72619 -21500 8 VDD
port 41 nsew
rlabel locali s 71536 -21917 71570 -21500 8 VDD
port 41 nsew
rlabel locali s 71340 -21917 71374 -21500 8 VDD
port 41 nsew
rlabel locali s 71330 -21500 72619 -21451 8 VDD
port 41 nsew
rlabel locali s 71330 -21451 71772 -21436 8 VDD
port 41 nsew
rlabel locali s 72776 -21412 73545 -21405 8 VDD
port 41 nsew
rlabel locali s 72776 -21405 73680 -21388 8 VDD
port 41 nsew
rlabel locali s 71769 -21402 71958 -21395 8 VDD
port 41 nsew
rlabel locali s 71732 -21395 71958 -21388 8 VDD
port 41 nsew
rlabel locali s 71330 -21388 73680 -21353 8 VDD
port 41 nsew
rlabel locali s 73618 -21353 73680 -21325 8 VDD
port 41 nsew
rlabel locali s 71330 -21353 73545 -21346 8 VDD
port 41 nsew
rlabel locali s 74409 -21308 74526 -21298 8 VDD
port 41 nsew
rlabel locali s 73846 -21308 73944 -21305 8 VDD
port 41 nsew
rlabel locali s 74409 -21298 74814 -21234 8 VDD
port 41 nsew
rlabel locali s 71330 -21346 73441 -21285 8 VDD
port 41 nsew
rlabel locali s 67933 -23647 68055 -21285 8 VDD
port 41 nsew
rlabel locali s 65036 -24770 65102 -23440 8 VDD
port 41 nsew
rlabel locali s 64683 -24854 64767 -24741 8 VDD
port 41 nsew
rlabel locali s 62169 -24858 64384 -24816 8 VDD
port 41 nsew
rlabel locali s 64700 -24741 64766 -23440 8 VDD
port 41 nsew
rlabel locali s 62169 -24816 64280 -24705 8 VDD
port 41 nsew
rlabel locali s 59599 -24970 59811 -24831 8 VDD
port 41 nsew
rlabel locali s 59349 -24985 59428 -24960 8 VDD
port 41 nsew
rlabel locali s 59152 -25103 59197 -24979 8 VDD
port 41 nsew
rlabel locali s 58736 -25695 58770 -25102 8 VDD
port 41 nsew
rlabel locali s 58540 -25695 58574 -25105 8 VDD
port 41 nsew
rlabel locali s 58290 -25283 58324 -25117 8 VDD
port 41 nsew
rlabel locali s 58094 -25283 58128 -25117 8 VDD
port 41 nsew
rlabel locali s 57898 -25283 57932 -25117 8 VDD
port 41 nsew
rlabel locali s 57702 -25283 57736 -25117 8 VDD
port 41 nsew
rlabel locali s 57485 -25484 57519 -25117 8 VDD
port 41 nsew
rlabel locali s 58730 -25102 58775 -24979 8 VDD
port 41 nsew
rlabel locali s 58535 -25105 58580 -24979 8 VDD
port 41 nsew
rlabel locali s 57485 -25117 58372 -25067 8 VDD
port 41 nsew
rlabel locali s 57289 -25484 57323 -25067 8 VDD
port 41 nsew
rlabel locali s 57093 -25484 57127 -25067 8 VDD
port 41 nsew
rlabel locali s 55491 -25664 55525 -25072 8 VDD
port 41 nsew
rlabel locali s 57083 -25067 58372 -25018 8 VDD
port 41 nsew
rlabel locali s 57083 -25018 57525 -25003 8 VDD
port 41 nsew
rlabel locali s 58529 -24979 59298 -24960 8 VDD
port 41 nsew
rlabel locali s 58529 -24960 59428 -24955 8 VDD
port 41 nsew
rlabel locali s 57522 -24969 57711 -24962 8 VDD
port 41 nsew
rlabel locali s 57485 -24962 57711 -24955 8 VDD
port 41 nsew
rlabel locali s 57083 -24955 59428 -24913 8 VDD
port 41 nsew
rlabel locali s 55484 -25072 55529 -24948 8 VDD
port 41 nsew
rlabel locali s 55068 -25664 55102 -25071 8 VDD
port 41 nsew
rlabel locali s 54872 -25664 54906 -25074 8 VDD
port 41 nsew
rlabel locali s 54622 -25252 54656 -25086 8 VDD
port 41 nsew
rlabel locali s 54426 -25252 54460 -25086 8 VDD
port 41 nsew
rlabel locali s 54230 -25252 54264 -25086 8 VDD
port 41 nsew
rlabel locali s 54034 -25252 54068 -25086 8 VDD
port 41 nsew
rlabel locali s 53817 -25453 53851 -25086 8 VDD
port 41 nsew
rlabel locali s 55062 -25071 55107 -24948 8 VDD
port 41 nsew
rlabel locali s 54867 -25074 54912 -24948 8 VDD
port 41 nsew
rlabel locali s 53817 -25086 54704 -25036 8 VDD
port 41 nsew
rlabel locali s 53621 -25453 53655 -25036 8 VDD
port 41 nsew
rlabel locali s 53425 -25453 53459 -25036 8 VDD
port 41 nsew
rlabel locali s 49961 -25729 49995 -25137 8 VDD
port 41 nsew
rlabel locali s 53415 -25036 54704 -24987 8 VDD
port 41 nsew
rlabel locali s 50401 -25032 50540 -25004 8 VDD
port 41 nsew
rlabel locali s 53415 -24987 53857 -24972 8 VDD
port 41 nsew
rlabel locali s 54861 -24948 55630 -24924 8 VDD
port 41 nsew
rlabel locali s 53854 -24938 54043 -24931 8 VDD
port 41 nsew
rlabel locali s 53817 -24931 54043 -24924 8 VDD
port 41 nsew
rlabel locali s 59249 -24913 59428 -24877 8 VDD
port 41 nsew
rlabel locali s 57083 -24913 59194 -24902 8 VDD
port 41 nsew
rlabel locali s 59349 -24877 59428 -24846 8 VDD
port 41 nsew
rlabel locali s 56282 -24902 59194 -24836 8 VDD
port 41 nsew
rlabel locali s 63167 -24705 63785 -24688 8 VDD
port 41 nsew
rlabel locali s 63167 -24688 63610 -24659 8 VDD
port 41 nsew
rlabel locali s 63168 -24659 63610 -24645 8 VDD
port 41 nsew
rlabel locali s 63168 -24645 64457 -24596 8 VDD
port 41 nsew
rlabel locali s 63570 -24596 64457 -24546 8 VDD
port 41 nsew
rlabel locali s 64375 -24546 64409 -24380 8 VDD
port 41 nsew
rlabel locali s 64179 -24546 64213 -24380 8 VDD
port 41 nsew
rlabel locali s 63983 -24546 64017 -24380 8 VDD
port 41 nsew
rlabel locali s 63787 -24546 63821 -24380 8 VDD
port 41 nsew
rlabel locali s 63570 -24546 63604 -24179 8 VDD
port 41 nsew
rlabel locali s 63374 -24596 63408 -24179 8 VDD
port 41 nsew
rlabel locali s 63178 -24596 63212 -24179 8 VDD
port 41 nsew
rlabel locali s 62339 -24705 62511 -24515 8 VDD
port 41 nsew
rlabel locali s 62157 -24515 62875 -24416 8 VDD
port 41 nsew
rlabel locali s 62793 -24416 62827 -24150 8 VDD
port 41 nsew
rlabel locali s 62597 -24416 62631 -24150 8 VDD
port 41 nsew
rlabel locali s 62401 -24416 62435 -24150 8 VDD
port 41 nsew
rlabel locali s 62205 -24416 62239 -24150 8 VDD
port 41 nsew
rlabel locali s 59689 -24831 59811 -23835 8 VDD
port 41 nsew
rlabel locali s 57083 -24836 59194 -24802 8 VDD
port 41 nsew
rlabel locali s 58081 -24802 58699 -24785 8 VDD
port 41 nsew
rlabel locali s 58081 -24785 58524 -24756 8 VDD
port 41 nsew
rlabel locali s 58082 -24756 58524 -24742 8 VDD
port 41 nsew
rlabel locali s 58082 -24742 59371 -24693 8 VDD
port 41 nsew
rlabel locali s 58484 -24693 59371 -24643 8 VDD
port 41 nsew
rlabel locali s 59289 -24643 59323 -24477 8 VDD
port 41 nsew
rlabel locali s 59093 -24643 59127 -24477 8 VDD
port 41 nsew
rlabel locali s 58897 -24643 58931 -24477 8 VDD
port 41 nsew
rlabel locali s 58701 -24643 58735 -24477 8 VDD
port 41 nsew
rlabel locali s 58484 -24643 58518 -24276 8 VDD
port 41 nsew
rlabel locali s 58288 -24693 58322 -24276 8 VDD
port 41 nsew
rlabel locali s 58092 -24693 58126 -24276 8 VDD
port 41 nsew
rlabel locali s 57253 -24802 57425 -24612 8 VDD
port 41 nsew
rlabel locali s 57071 -24612 57789 -24513 8 VDD
port 41 nsew
rlabel locali s 57707 -24513 57741 -24247 8 VDD
port 41 nsew
rlabel locali s 57511 -24513 57545 -24247 8 VDD
port 41 nsew
rlabel locali s 57315 -24513 57349 -24247 8 VDD
port 41 nsew
rlabel locali s 57119 -24513 57153 -24247 8 VDD
port 41 nsew
rlabel locali s 59179 -23835 59811 -23713 8 VDD
port 41 nsew
rlabel locali s 64700 -23440 65102 -23374 8 VDD
port 41 nsew
rlabel locali s 66971 -21703 67005 -21411 8 VDD
port 41 nsew
rlabel locali s 66775 -21703 66809 -21413 8 VDD
port 41 nsew
rlabel locali s 66547 -21903 66581 -21428 8 VDD
port 41 nsew
rlabel locali s 66417 -21903 66451 -21431 8 VDD
port 41 nsew
rlabel locali s 66966 -21411 67009 -21285 8 VDD
port 41 nsew
rlabel locali s 66961 -21285 73441 -21251 8 VDD
port 41 nsew
rlabel locali s 66769 -21413 66812 -21251 8 VDD
port 41 nsew
rlabel locali s 66538 -21428 66588 -21251 8 VDD
port 41 nsew
rlabel locali s 66412 -21431 66462 -21251 8 VDD
port 41 nsew
rlabel locali s 65822 -21903 65856 -21408 8 VDD
port 41 nsew
rlabel locali s 65626 -21903 65660 -21410 8 VDD
port 41 nsew
rlabel locali s 64253 -22145 64287 -21553 8 VDD
port 41 nsew
rlabel locali s 64693 -21448 64791 -21442 8 VDD
port 41 nsew
rlabel locali s 65820 -21408 65858 -21251 8 VDD
port 41 nsew
rlabel locali s 65623 -21410 65661 -21315 8 VDD
port 41 nsew
rlabel locali s 64693 -21442 65373 -21325 8 VDD
port 41 nsew
rlabel locali s 64465 -21436 64527 -21422 8 VDD
port 41 nsew
rlabel locali s 64246 -21553 64291 -21429 8 VDD
port 41 nsew
rlabel locali s 63830 -22145 63864 -21552 8 VDD
port 41 nsew
rlabel locali s 63634 -22145 63668 -21555 8 VDD
port 41 nsew
rlabel locali s 63384 -21733 63418 -21567 8 VDD
port 41 nsew
rlabel locali s 63188 -21733 63222 -21567 8 VDD
port 41 nsew
rlabel locali s 62992 -21733 63026 -21567 8 VDD
port 41 nsew
rlabel locali s 62796 -21733 62830 -21567 8 VDD
port 41 nsew
rlabel locali s 62579 -21934 62613 -21567 8 VDD
port 41 nsew
rlabel locali s 63824 -21552 63869 -21429 8 VDD
port 41 nsew
rlabel locali s 63629 -21555 63674 -21429 8 VDD
port 41 nsew
rlabel locali s 62579 -21567 63466 -21517 8 VDD
port 41 nsew
rlabel locali s 62383 -21934 62417 -21517 8 VDD
port 41 nsew
rlabel locali s 62187 -21934 62221 -21517 8 VDD
port 41 nsew
rlabel locali s 62177 -21517 63466 -21468 8 VDD
port 41 nsew
rlabel locali s 62177 -21468 62619 -21453 8 VDD
port 41 nsew
rlabel locali s 63623 -21429 64392 -21422 8 VDD
port 41 nsew
rlabel locali s 63623 -21422 64527 -21405 8 VDD
port 41 nsew
rlabel locali s 62616 -21419 62805 -21412 8 VDD
port 41 nsew
rlabel locali s 62579 -21412 62805 -21405 8 VDD
port 41 nsew
rlabel locali s 62177 -21405 64527 -21379 8 VDD
port 41 nsew
rlabel locali s 59179 -23713 59301 -21379 8 VDD
port 41 nsew
rlabel locali s 56282 -24836 56348 -23506 8 VDD
port 41 nsew
rlabel locali s 55929 -24920 56013 -24807 8 VDD
port 41 nsew
rlabel locali s 53415 -24924 55630 -24882 8 VDD
port 41 nsew
rlabel locali s 55946 -24807 56012 -23506 8 VDD
port 41 nsew
rlabel locali s 53415 -24882 55526 -24771 8 VDD
port 41 nsew
rlabel locali s 50401 -25004 50613 -24865 8 VDD
port 41 nsew
rlabel locali s 50151 -25019 50230 -24994 8 VDD
port 41 nsew
rlabel locali s 49954 -25137 49999 -25013 8 VDD
port 41 nsew
rlabel locali s 49538 -25729 49572 -25136 8 VDD
port 41 nsew
rlabel locali s 49342 -25729 49376 -25139 8 VDD
port 41 nsew
rlabel locali s 49092 -25317 49126 -25151 8 VDD
port 41 nsew
rlabel locali s 48896 -25317 48930 -25151 8 VDD
port 41 nsew
rlabel locali s 48700 -25317 48734 -25151 8 VDD
port 41 nsew
rlabel locali s 48504 -25317 48538 -25151 8 VDD
port 41 nsew
rlabel locali s 48287 -25518 48321 -25151 8 VDD
port 41 nsew
rlabel locali s 49532 -25136 49577 -25013 8 VDD
port 41 nsew
rlabel locali s 49337 -25139 49382 -25013 8 VDD
port 41 nsew
rlabel locali s 48287 -25151 49174 -25101 8 VDD
port 41 nsew
rlabel locali s 48091 -25518 48125 -25101 8 VDD
port 41 nsew
rlabel locali s 47895 -25518 47929 -25101 8 VDD
port 41 nsew
rlabel locali s 46293 -25698 46327 -25106 8 VDD
port 41 nsew
rlabel locali s 47885 -25101 49174 -25052 8 VDD
port 41 nsew
rlabel locali s 47885 -25052 48327 -25037 8 VDD
port 41 nsew
rlabel locali s 49331 -25013 50100 -24994 8 VDD
port 41 nsew
rlabel locali s 49331 -24994 50230 -24989 8 VDD
port 41 nsew
rlabel locali s 48324 -25003 48513 -24996 8 VDD
port 41 nsew
rlabel locali s 48287 -24996 48513 -24989 8 VDD
port 41 nsew
rlabel locali s 47885 -24989 50230 -24947 8 VDD
port 41 nsew
rlabel locali s 46286 -25106 46331 -24982 8 VDD
port 41 nsew
rlabel locali s 45870 -25698 45904 -25105 8 VDD
port 41 nsew
rlabel locali s 45674 -25698 45708 -25108 8 VDD
port 41 nsew
rlabel locali s 45424 -25286 45458 -25120 8 VDD
port 41 nsew
rlabel locali s 45228 -25286 45262 -25120 8 VDD
port 41 nsew
rlabel locali s 45032 -25286 45066 -25120 8 VDD
port 41 nsew
rlabel locali s 44836 -25286 44870 -25120 8 VDD
port 41 nsew
rlabel locali s 44619 -25487 44653 -25120 8 VDD
port 41 nsew
rlabel locali s 45864 -25105 45909 -24982 8 VDD
port 41 nsew
rlabel locali s 45669 -25108 45714 -24982 8 VDD
port 41 nsew
rlabel locali s 44619 -25120 45506 -25070 8 VDD
port 41 nsew
rlabel locali s 44423 -25487 44457 -25070 8 VDD
port 41 nsew
rlabel locali s 44227 -25487 44261 -25070 8 VDD
port 41 nsew
rlabel locali s 41098 -25690 41132 -25098 8 VDD
port 41 nsew
rlabel locali s 44217 -25070 45506 -25021 8 VDD
port 41 nsew
rlabel locali s 44217 -25021 44659 -25006 8 VDD
port 41 nsew
rlabel locali s 45663 -24982 46432 -24958 8 VDD
port 41 nsew
rlabel locali s 44656 -24972 44845 -24965 8 VDD
port 41 nsew
rlabel locali s 41538 -24993 41677 -24965 8 VDD
port 41 nsew
rlabel locali s 44619 -24965 44845 -24958 8 VDD
port 41 nsew
rlabel locali s 50051 -24947 50230 -24911 8 VDD
port 41 nsew
rlabel locali s 47885 -24947 49996 -24936 8 VDD
port 41 nsew
rlabel locali s 50151 -24911 50230 -24880 8 VDD
port 41 nsew
rlabel locali s 47084 -24936 49996 -24870 8 VDD
port 41 nsew
rlabel locali s 54413 -24771 55031 -24754 8 VDD
port 41 nsew
rlabel locali s 54413 -24754 54856 -24725 8 VDD
port 41 nsew
rlabel locali s 54414 -24725 54856 -24711 8 VDD
port 41 nsew
rlabel locali s 54414 -24711 55703 -24662 8 VDD
port 41 nsew
rlabel locali s 54816 -24662 55703 -24612 8 VDD
port 41 nsew
rlabel locali s 55621 -24612 55655 -24446 8 VDD
port 41 nsew
rlabel locali s 55425 -24612 55459 -24446 8 VDD
port 41 nsew
rlabel locali s 55229 -24612 55263 -24446 8 VDD
port 41 nsew
rlabel locali s 55033 -24612 55067 -24446 8 VDD
port 41 nsew
rlabel locali s 54816 -24612 54850 -24245 8 VDD
port 41 nsew
rlabel locali s 54620 -24662 54654 -24245 8 VDD
port 41 nsew
rlabel locali s 54424 -24662 54458 -24245 8 VDD
port 41 nsew
rlabel locali s 53585 -24771 53757 -24581 8 VDD
port 41 nsew
rlabel locali s 53403 -24581 54121 -24482 8 VDD
port 41 nsew
rlabel locali s 54039 -24482 54073 -24216 8 VDD
port 41 nsew
rlabel locali s 53843 -24482 53877 -24216 8 VDD
port 41 nsew
rlabel locali s 53647 -24482 53681 -24216 8 VDD
port 41 nsew
rlabel locali s 53451 -24482 53485 -24216 8 VDD
port 41 nsew
rlabel locali s 50491 -24865 50613 -23869 8 VDD
port 41 nsew
rlabel locali s 47885 -24870 49996 -24836 8 VDD
port 41 nsew
rlabel locali s 48883 -24836 49501 -24819 8 VDD
port 41 nsew
rlabel locali s 48883 -24819 49326 -24790 8 VDD
port 41 nsew
rlabel locali s 48884 -24790 49326 -24776 8 VDD
port 41 nsew
rlabel locali s 48884 -24776 50173 -24727 8 VDD
port 41 nsew
rlabel locali s 49286 -24727 50173 -24677 8 VDD
port 41 nsew
rlabel locali s 50091 -24677 50125 -24511 8 VDD
port 41 nsew
rlabel locali s 49895 -24677 49929 -24511 8 VDD
port 41 nsew
rlabel locali s 49699 -24677 49733 -24511 8 VDD
port 41 nsew
rlabel locali s 49503 -24677 49537 -24511 8 VDD
port 41 nsew
rlabel locali s 49286 -24677 49320 -24310 8 VDD
port 41 nsew
rlabel locali s 49090 -24727 49124 -24310 8 VDD
port 41 nsew
rlabel locali s 48894 -24727 48928 -24310 8 VDD
port 41 nsew
rlabel locali s 48055 -24836 48227 -24646 8 VDD
port 41 nsew
rlabel locali s 47873 -24646 48591 -24547 8 VDD
port 41 nsew
rlabel locali s 48509 -24547 48543 -24281 8 VDD
port 41 nsew
rlabel locali s 48313 -24547 48347 -24281 8 VDD
port 41 nsew
rlabel locali s 48117 -24547 48151 -24281 8 VDD
port 41 nsew
rlabel locali s 47921 -24547 47955 -24281 8 VDD
port 41 nsew
rlabel locali s 49981 -23869 50613 -23747 8 VDD
port 41 nsew
rlabel locali s 55946 -23506 56348 -23440 8 VDD
port 41 nsew
rlabel locali s 58217 -21769 58251 -21477 8 VDD
port 41 nsew
rlabel locali s 58021 -21769 58055 -21479 8 VDD
port 41 nsew
rlabel locali s 57793 -21969 57827 -21494 8 VDD
port 41 nsew
rlabel locali s 57663 -21969 57697 -21497 8 VDD
port 41 nsew
rlabel locali s 58212 -21477 58255 -21379 8 VDD
port 41 nsew
rlabel locali s 58212 -21379 64527 -21370 8 VDD
port 41 nsew
rlabel locali s 64465 -21370 64527 -21342 8 VDD
port 41 nsew
rlabel locali s 58212 -21370 64392 -21363 8 VDD
port 41 nsew
rlabel locali s 65256 -21325 65373 -21315 8 VDD
port 41 nsew
rlabel locali s 64693 -21325 64791 -21322 8 VDD
port 41 nsew
rlabel locali s 65256 -21315 65661 -21251 8 VDD
port 41 nsew
rlabel locali s 58212 -21363 64288 -21317 8 VDD
port 41 nsew
rlabel locali s 58015 -21479 58058 -21317 8 VDD
port 41 nsew
rlabel locali s 57784 -21494 57834 -21317 8 VDD
port 41 nsew
rlabel locali s 57658 -21497 57708 -21317 8 VDD
port 41 nsew
rlabel locali s 57068 -21969 57102 -21474 8 VDD
port 41 nsew
rlabel locali s 56872 -21969 56906 -21476 8 VDD
port 41 nsew
rlabel locali s 55499 -22211 55533 -21619 8 VDD
port 41 nsew
rlabel locali s 55939 -21514 56037 -21508 8 VDD
port 41 nsew
rlabel locali s 57066 -21474 57104 -21317 8 VDD
port 41 nsew
rlabel locali s 56869 -21476 56907 -21381 8 VDD
port 41 nsew
rlabel locali s 55939 -21508 56619 -21391 8 VDD
port 41 nsew
rlabel locali s 55711 -21502 55773 -21488 8 VDD
port 41 nsew
rlabel locali s 55492 -21619 55537 -21495 8 VDD
port 41 nsew
rlabel locali s 55076 -22211 55110 -21618 8 VDD
port 41 nsew
rlabel locali s 54880 -22211 54914 -21621 8 VDD
port 41 nsew
rlabel locali s 54630 -21799 54664 -21633 8 VDD
port 41 nsew
rlabel locali s 54434 -21799 54468 -21633 8 VDD
port 41 nsew
rlabel locali s 54238 -21799 54272 -21633 8 VDD
port 41 nsew
rlabel locali s 54042 -21799 54076 -21633 8 VDD
port 41 nsew
rlabel locali s 53825 -22000 53859 -21633 8 VDD
port 41 nsew
rlabel locali s 55070 -21618 55115 -21495 8 VDD
port 41 nsew
rlabel locali s 54875 -21621 54920 -21495 8 VDD
port 41 nsew
rlabel locali s 53825 -21633 54712 -21583 8 VDD
port 41 nsew
rlabel locali s 53629 -22000 53663 -21583 8 VDD
port 41 nsew
rlabel locali s 53433 -22000 53467 -21583 8 VDD
port 41 nsew
rlabel locali s 53423 -21583 54712 -21534 8 VDD
port 41 nsew
rlabel locali s 53423 -21534 53865 -21519 8 VDD
port 41 nsew
rlabel locali s 54869 -21495 55638 -21488 8 VDD
port 41 nsew
rlabel locali s 54869 -21488 55773 -21471 8 VDD
port 41 nsew
rlabel locali s 53862 -21485 54051 -21478 8 VDD
port 41 nsew
rlabel locali s 53825 -21478 54051 -21471 8 VDD
port 41 nsew
rlabel locali s 53423 -21471 55773 -21436 8 VDD
port 41 nsew
rlabel locali s 55711 -21436 55773 -21408 8 VDD
port 41 nsew
rlabel locali s 53423 -21436 55638 -21429 8 VDD
port 41 nsew
rlabel locali s 53423 -21429 55534 -21411 8 VDD
port 41 nsew
rlabel locali s 49981 -23747 50103 -21411 8 VDD
port 41 nsew
rlabel locali s 47084 -24870 47150 -23540 8 VDD
port 41 nsew
rlabel locali s 46731 -24954 46815 -24841 8 VDD
port 41 nsew
rlabel locali s 44217 -24958 46432 -24916 8 VDD
port 41 nsew
rlabel locali s 46748 -24841 46814 -23540 8 VDD
port 41 nsew
rlabel locali s 44217 -24916 46328 -24805 8 VDD
port 41 nsew
rlabel locali s 41538 -24965 41750 -24826 8 VDD
port 41 nsew
rlabel locali s 41288 -24980 41367 -24955 8 VDD
port 41 nsew
rlabel locali s 41091 -25098 41136 -24974 8 VDD
port 41 nsew
rlabel locali s 40675 -25690 40709 -25097 8 VDD
port 41 nsew
rlabel locali s 40479 -25690 40513 -25100 8 VDD
port 41 nsew
rlabel locali s 40229 -25278 40263 -25112 8 VDD
port 41 nsew
rlabel locali s 40033 -25278 40067 -25112 8 VDD
port 41 nsew
rlabel locali s 39837 -25278 39871 -25112 8 VDD
port 41 nsew
rlabel locali s 39641 -25278 39675 -25112 8 VDD
port 41 nsew
rlabel locali s 39424 -25479 39458 -25112 8 VDD
port 41 nsew
rlabel locali s 40669 -25097 40714 -24974 8 VDD
port 41 nsew
rlabel locali s 40474 -25100 40519 -24974 8 VDD
port 41 nsew
rlabel locali s 39424 -25112 40311 -25062 8 VDD
port 41 nsew
rlabel locali s 39228 -25479 39262 -25062 8 VDD
port 41 nsew
rlabel locali s 39032 -25479 39066 -25062 8 VDD
port 41 nsew
rlabel locali s 37430 -25659 37464 -25067 8 VDD
port 41 nsew
rlabel locali s 39022 -25062 40311 -25013 8 VDD
port 41 nsew
rlabel locali s 39022 -25013 39464 -24998 8 VDD
port 41 nsew
rlabel locali s 40468 -24974 41237 -24955 8 VDD
port 41 nsew
rlabel locali s 40468 -24955 41367 -24950 8 VDD
port 41 nsew
rlabel locali s 39461 -24964 39650 -24957 8 VDD
port 41 nsew
rlabel locali s 39424 -24957 39650 -24950 8 VDD
port 41 nsew
rlabel locali s 39022 -24950 41367 -24908 8 VDD
port 41 nsew
rlabel locali s 37423 -25067 37468 -24943 8 VDD
port 41 nsew
rlabel locali s 37007 -25659 37041 -25066 8 VDD
port 41 nsew
rlabel locali s 36811 -25659 36845 -25069 8 VDD
port 41 nsew
rlabel locali s 36561 -25247 36595 -25081 8 VDD
port 41 nsew
rlabel locali s 36365 -25247 36399 -25081 8 VDD
port 41 nsew
rlabel locali s 36169 -25247 36203 -25081 8 VDD
port 41 nsew
rlabel locali s 35973 -25247 36007 -25081 8 VDD
port 41 nsew
rlabel locali s 35756 -25448 35790 -25081 8 VDD
port 41 nsew
rlabel locali s 37001 -25066 37046 -24943 8 VDD
port 41 nsew
rlabel locali s 36806 -25069 36851 -24943 8 VDD
port 41 nsew
rlabel locali s 35756 -25081 36643 -25031 8 VDD
port 41 nsew
rlabel locali s 35560 -25448 35594 -25031 8 VDD
port 41 nsew
rlabel locali s 35364 -25448 35398 -25031 8 VDD
port 41 nsew
rlabel locali s 32658 -25679 32692 -25087 8 VDD
port 41 nsew
rlabel locali s 35354 -25031 36643 -24982 8 VDD
port 41 nsew
rlabel locali s 35354 -24982 35796 -24967 8 VDD
port 41 nsew
rlabel locali s 33098 -24982 33237 -24954 8 VDD
port 41 nsew
rlabel locali s 36800 -24943 37569 -24919 8 VDD
port 41 nsew
rlabel locali s 35793 -24933 35982 -24926 8 VDD
port 41 nsew
rlabel locali s 35756 -24926 35982 -24919 8 VDD
port 41 nsew
rlabel locali s 41188 -24908 41367 -24872 8 VDD
port 41 nsew
rlabel locali s 39022 -24908 41133 -24897 8 VDD
port 41 nsew
rlabel locali s 41288 -24872 41367 -24841 8 VDD
port 41 nsew
rlabel locali s 38221 -24897 41133 -24831 8 VDD
port 41 nsew
rlabel locali s 45215 -24805 45833 -24788 8 VDD
port 41 nsew
rlabel locali s 45215 -24788 45658 -24759 8 VDD
port 41 nsew
rlabel locali s 45216 -24759 45658 -24745 8 VDD
port 41 nsew
rlabel locali s 45216 -24745 46505 -24696 8 VDD
port 41 nsew
rlabel locali s 45618 -24696 46505 -24646 8 VDD
port 41 nsew
rlabel locali s 46423 -24646 46457 -24480 8 VDD
port 41 nsew
rlabel locali s 46227 -24646 46261 -24480 8 VDD
port 41 nsew
rlabel locali s 46031 -24646 46065 -24480 8 VDD
port 41 nsew
rlabel locali s 45835 -24646 45869 -24480 8 VDD
port 41 nsew
rlabel locali s 45618 -24646 45652 -24279 8 VDD
port 41 nsew
rlabel locali s 45422 -24696 45456 -24279 8 VDD
port 41 nsew
rlabel locali s 45226 -24696 45260 -24279 8 VDD
port 41 nsew
rlabel locali s 44387 -24805 44559 -24615 8 VDD
port 41 nsew
rlabel locali s 44205 -24615 44923 -24516 8 VDD
port 41 nsew
rlabel locali s 44841 -24516 44875 -24250 8 VDD
port 41 nsew
rlabel locali s 44645 -24516 44679 -24250 8 VDD
port 41 nsew
rlabel locali s 44449 -24516 44483 -24250 8 VDD
port 41 nsew
rlabel locali s 44253 -24516 44287 -24250 8 VDD
port 41 nsew
rlabel locali s 41628 -24826 41750 -23830 8 VDD
port 41 nsew
rlabel locali s 39022 -24831 41133 -24797 8 VDD
port 41 nsew
rlabel locali s 40020 -24797 40638 -24780 8 VDD
port 41 nsew
rlabel locali s 40020 -24780 40463 -24751 8 VDD
port 41 nsew
rlabel locali s 40021 -24751 40463 -24737 8 VDD
port 41 nsew
rlabel locali s 40021 -24737 41310 -24688 8 VDD
port 41 nsew
rlabel locali s 40423 -24688 41310 -24638 8 VDD
port 41 nsew
rlabel locali s 41228 -24638 41262 -24472 8 VDD
port 41 nsew
rlabel locali s 41032 -24638 41066 -24472 8 VDD
port 41 nsew
rlabel locali s 40836 -24638 40870 -24472 8 VDD
port 41 nsew
rlabel locali s 40640 -24638 40674 -24472 8 VDD
port 41 nsew
rlabel locali s 40423 -24638 40457 -24271 8 VDD
port 41 nsew
rlabel locali s 40227 -24688 40261 -24271 8 VDD
port 41 nsew
rlabel locali s 40031 -24688 40065 -24271 8 VDD
port 41 nsew
rlabel locali s 39192 -24797 39364 -24607 8 VDD
port 41 nsew
rlabel locali s 39010 -24607 39728 -24508 8 VDD
port 41 nsew
rlabel locali s 39646 -24508 39680 -24242 8 VDD
port 41 nsew
rlabel locali s 39450 -24508 39484 -24242 8 VDD
port 41 nsew
rlabel locali s 39254 -24508 39288 -24242 8 VDD
port 41 nsew
rlabel locali s 39058 -24508 39092 -24242 8 VDD
port 41 nsew
rlabel locali s 41118 -23830 41750 -23708 8 VDD
port 41 nsew
rlabel locali s 46748 -23540 47150 -23474 8 VDD
port 41 nsew
rlabel locali s 49019 -21803 49053 -21511 8 VDD
port 41 nsew
rlabel locali s 48823 -21803 48857 -21513 8 VDD
port 41 nsew
rlabel locali s 48595 -22003 48629 -21528 8 VDD
port 41 nsew
rlabel locali s 48465 -22003 48499 -21531 8 VDD
port 41 nsew
rlabel locali s 49014 -21511 49057 -21411 8 VDD
port 41 nsew
rlabel locali s 56502 -21391 56619 -21381 8 VDD
port 41 nsew
rlabel locali s 55939 -21391 56037 -21388 8 VDD
port 41 nsew
rlabel locali s 56502 -21381 56907 -21317 8 VDD
port 41 nsew
rlabel locali s 49014 -21411 55534 -21351 8 VDD
port 41 nsew
rlabel locali s 48817 -21513 48860 -21351 8 VDD
port 41 nsew
rlabel locali s 48586 -21528 48636 -21351 8 VDD
port 41 nsew
rlabel locali s 48460 -21531 48510 -21351 8 VDD
port 41 nsew
rlabel locali s 47870 -22003 47904 -21508 8 VDD
port 41 nsew
rlabel locali s 47674 -22003 47708 -21510 8 VDD
port 41 nsew
rlabel locali s 46301 -22245 46335 -21653 8 VDD
port 41 nsew
rlabel locali s 46741 -21548 46839 -21542 8 VDD
port 41 nsew
rlabel locali s 47868 -21508 47906 -21351 8 VDD
port 41 nsew
rlabel locali s 47671 -21510 47709 -21415 8 VDD
port 41 nsew
rlabel locali s 46741 -21542 47421 -21425 8 VDD
port 41 nsew
rlabel locali s 46513 -21536 46575 -21522 8 VDD
port 41 nsew
rlabel locali s 46294 -21653 46339 -21529 8 VDD
port 41 nsew
rlabel locali s 45878 -22245 45912 -21652 8 VDD
port 41 nsew
rlabel locali s 45682 -22245 45716 -21655 8 VDD
port 41 nsew
rlabel locali s 45432 -21833 45466 -21667 8 VDD
port 41 nsew
rlabel locali s 45236 -21833 45270 -21667 8 VDD
port 41 nsew
rlabel locali s 45040 -21833 45074 -21667 8 VDD
port 41 nsew
rlabel locali s 44844 -21833 44878 -21667 8 VDD
port 41 nsew
rlabel locali s 44627 -22034 44661 -21667 8 VDD
port 41 nsew
rlabel locali s 45872 -21652 45917 -21529 8 VDD
port 41 nsew
rlabel locali s 45677 -21655 45722 -21529 8 VDD
port 41 nsew
rlabel locali s 44627 -21667 45514 -21617 8 VDD
port 41 nsew
rlabel locali s 44431 -22034 44465 -21617 8 VDD
port 41 nsew
rlabel locali s 44235 -22034 44269 -21617 8 VDD
port 41 nsew
rlabel locali s 44225 -21617 45514 -21568 8 VDD
port 41 nsew
rlabel locali s 44225 -21568 44667 -21553 8 VDD
port 41 nsew
rlabel locali s 45671 -21529 46440 -21522 8 VDD
port 41 nsew
rlabel locali s 45671 -21522 46575 -21505 8 VDD
port 41 nsew
rlabel locali s 44664 -21519 44853 -21512 8 VDD
port 41 nsew
rlabel locali s 44627 -21512 44853 -21505 8 VDD
port 41 nsew
rlabel locali s 44225 -21505 46575 -21470 8 VDD
port 41 nsew
rlabel locali s 46513 -21470 46575 -21442 8 VDD
port 41 nsew
rlabel locali s 44225 -21470 46440 -21463 8 VDD
port 41 nsew
rlabel locali s 47304 -21425 47421 -21415 8 VDD
port 41 nsew
rlabel locali s 46741 -21425 46839 -21422 8 VDD
port 41 nsew
rlabel locali s 47304 -21415 47709 -21351 8 VDD
port 41 nsew
rlabel locali s 44225 -21463 46336 -21401 8 VDD
port 41 nsew
rlabel locali s 41118 -23708 41240 -21401 8 VDD
port 41 nsew
rlabel locali s 38221 -24831 38287 -23501 8 VDD
port 41 nsew
rlabel locali s 37868 -24915 37952 -24802 8 VDD
port 41 nsew
rlabel locali s 35354 -24919 37569 -24877 8 VDD
port 41 nsew
rlabel locali s 37885 -24802 37951 -23501 8 VDD
port 41 nsew
rlabel locali s 35354 -24877 37465 -24766 8 VDD
port 41 nsew
rlabel locali s 33098 -24954 33310 -24815 8 VDD
port 41 nsew
rlabel locali s 32848 -24969 32927 -24944 8 VDD
port 41 nsew
rlabel locali s 32651 -25087 32696 -24963 8 VDD
port 41 nsew
rlabel locali s 32235 -25679 32269 -25086 8 VDD
port 41 nsew
rlabel locali s 32039 -25679 32073 -25089 8 VDD
port 41 nsew
rlabel locali s 31789 -25267 31823 -25101 8 VDD
port 41 nsew
rlabel locali s 31593 -25267 31627 -25101 8 VDD
port 41 nsew
rlabel locali s 31397 -25267 31431 -25101 8 VDD
port 41 nsew
rlabel locali s 31201 -25267 31235 -25101 8 VDD
port 41 nsew
rlabel locali s 30984 -25468 31018 -25101 8 VDD
port 41 nsew
rlabel locali s 32229 -25086 32274 -24963 8 VDD
port 41 nsew
rlabel locali s 32034 -25089 32079 -24963 8 VDD
port 41 nsew
rlabel locali s 30984 -25101 31871 -25051 8 VDD
port 41 nsew
rlabel locali s 30788 -25468 30822 -25051 8 VDD
port 41 nsew
rlabel locali s 30592 -25468 30626 -25051 8 VDD
port 41 nsew
rlabel locali s 28990 -25648 29024 -25056 8 VDD
port 41 nsew
rlabel locali s 30582 -25051 31871 -25002 8 VDD
port 41 nsew
rlabel locali s 30582 -25002 31024 -24987 8 VDD
port 41 nsew
rlabel locali s 32028 -24963 32797 -24944 8 VDD
port 41 nsew
rlabel locali s 32028 -24944 32927 -24939 8 VDD
port 41 nsew
rlabel locali s 31021 -24953 31210 -24946 8 VDD
port 41 nsew
rlabel locali s 30984 -24946 31210 -24939 8 VDD
port 41 nsew
rlabel locali s 30582 -24939 32927 -24897 8 VDD
port 41 nsew
rlabel locali s 28983 -25056 29028 -24932 8 VDD
port 41 nsew
rlabel locali s 28567 -25648 28601 -25055 8 VDD
port 41 nsew
rlabel locali s 28371 -25648 28405 -25058 8 VDD
port 41 nsew
rlabel locali s 16581 -27265 16670 -25570 8 VDD
port 41 nsew
rlabel locali s 16387 -27265 16421 -26974 8 VDD
port 41 nsew
rlabel locali s 16191 -27265 16225 -26974 8 VDD
port 41 nsew
rlabel locali s 15995 -27265 16029 -26974 8 VDD
port 41 nsew
rlabel locali s 15550 -27265 15584 -26974 8 VDD
port 41 nsew
rlabel locali s 15354 -27265 15388 -26974 8 VDD
port 41 nsew
rlabel locali s 15158 -27265 15192 -26974 8 VDD
port 41 nsew
rlabel locali s 13687 -27265 13721 -26974 8 VDD
port 41 nsew
rlabel locali s 13491 -27265 13525 -26974 8 VDD
port 41 nsew
rlabel locali s 13295 -27265 13329 -26974 8 VDD
port 41 nsew
rlabel locali s 12850 -27265 12884 -26974 8 VDD
port 41 nsew
rlabel locali s 12654 -27265 12688 -26974 8 VDD
port 41 nsew
rlabel locali s 12458 -27265 12492 -26974 8 VDD
port 41 nsew
rlabel locali s 7342 -27327 7376 -27137 8 VDD
port 41 nsew
rlabel locali s 7140 -27449 7186 -27315 8 VDD
port 41 nsew
rlabel locali s 7027 -27449 7073 -27325 8 VDD
port 41 nsew
rlabel locali s 7146 -27315 7180 -27137 8 VDD
port 41 nsew
rlabel locali s 7033 -27325 7067 -27137 8 VDD
port 41 nsew
rlabel locali s 6831 -27449 6877 -27320 8 VDD
port 41 nsew
rlabel locali s 6718 -27449 6764 -27324 8 VDD
port 41 nsew
rlabel locali s 6837 -27320 6871 -27137 8 VDD
port 41 nsew
rlabel locali s 6723 -27324 6757 -27137 8 VDD
port 41 nsew
rlabel locali s 6520 -27449 6566 -27320 8 VDD
port 41 nsew
rlabel locali s 6331 -27449 6371 -27320 8 VDD
port 41 nsew
rlabel locali s 3331 -27518 4383 -27449 8 VDD
port 41 nsew
rlabel locali s 4337 -27449 4383 -27327 8 VDD
port 41 nsew
rlabel locali s 6527 -27320 6561 -27137 8 VDD
port 41 nsew
rlabel locali s 6331 -27320 6365 -27137 8 VDD
port 41 nsew
rlabel locali s 4342 -27327 4376 -27137 8 VDD
port 41 nsew
rlabel locali s 4140 -27449 4186 -27315 8 VDD
port 41 nsew
rlabel locali s 4027 -27449 4073 -27325 8 VDD
port 41 nsew
rlabel locali s 4146 -27315 4180 -27137 8 VDD
port 41 nsew
rlabel locali s 4033 -27325 4067 -27137 8 VDD
port 41 nsew
rlabel locali s 3831 -27449 3877 -27320 8 VDD
port 41 nsew
rlabel locali s 3718 -27449 3764 -27324 8 VDD
port 41 nsew
rlabel locali s 3837 -27320 3871 -27137 8 VDD
port 41 nsew
rlabel locali s 3723 -27324 3757 -27137 8 VDD
port 41 nsew
rlabel locali s 3520 -27449 3566 -27320 8 VDD
port 41 nsew
rlabel locali s 3331 -27449 3371 -27320 8 VDD
port 41 nsew
rlabel locali s 831 -27518 1883 -27449 8 VDD
port 41 nsew
rlabel locali s 1837 -27449 1883 -27327 8 VDD
port 41 nsew
rlabel locali s 3527 -27320 3561 -27137 8 VDD
port 41 nsew
rlabel locali s 3331 -27320 3365 -27137 8 VDD
port 41 nsew
rlabel locali s 1842 -27327 1876 -27137 8 VDD
port 41 nsew
rlabel locali s 1640 -27449 1686 -27315 8 VDD
port 41 nsew
rlabel locali s 1527 -27449 1573 -27325 8 VDD
port 41 nsew
rlabel locali s 1646 -27315 1680 -27137 8 VDD
port 41 nsew
rlabel locali s 1533 -27325 1567 -27137 8 VDD
port 41 nsew
rlabel locali s 1331 -27449 1377 -27320 8 VDD
port 41 nsew
rlabel locali s 1218 -27449 1264 -27324 8 VDD
port 41 nsew
rlabel locali s 1337 -27320 1371 -27137 8 VDD
port 41 nsew
rlabel locali s 1223 -27324 1257 -27137 8 VDD
port 41 nsew
rlabel locali s 1020 -27449 1066 -27320 8 VDD
port 41 nsew
rlabel locali s 831 -27449 871 -27320 8 VDD
port 41 nsew
rlabel locali s 1027 -27320 1061 -27137 8 VDD
port 41 nsew
rlabel locali s 831 -27320 865 -27137 8 VDD
port 41 nsew
rlabel locali s -292 -27556 -177 -26684 2 VDD
port 41 nsew
rlabel locali s -1339 -27556 -746 -27518 2 VDD
port 41 nsew
rlabel locali s -1669 -27518 -617 -27449 2 VDD
port 41 nsew
rlabel locali s -663 -27449 -617 -27327 2 VDD
port 41 nsew
rlabel locali s -658 -27327 -624 -27137 2 VDD
port 41 nsew
rlabel locali s -860 -27449 -814 -27315 2 VDD
port 41 nsew
rlabel locali s -973 -27449 -927 -27325 2 VDD
port 41 nsew
rlabel locali s -854 -27315 -820 -27137 2 VDD
port 41 nsew
rlabel locali s -967 -27325 -933 -27137 2 VDD
port 41 nsew
rlabel locali s -1169 -27449 -1123 -27320 2 VDD
port 41 nsew
rlabel locali s -1282 -27449 -1236 -27324 2 VDD
port 41 nsew
rlabel locali s -1163 -27320 -1129 -27137 2 VDD
port 41 nsew
rlabel locali s -1277 -27324 -1243 -27137 2 VDD
port 41 nsew
rlabel locali s -1480 -27449 -1434 -27320 2 VDD
port 41 nsew
rlabel locali s -1669 -27449 -1629 -27320 2 VDD
port 41 nsew
rlabel locali s -1473 -27320 -1439 -27137 2 VDD
port 41 nsew
rlabel locali s -1669 -27320 -1635 -27137 2 VDD
port 41 nsew
rlabel locali s -2774 -27556 -2660 -26684 2 VDD
port 41 nsew
rlabel locali s -3855 -27556 -3262 -27518 2 VDD
port 41 nsew
rlabel locali s -4169 -27518 -3117 -27449 2 VDD
port 41 nsew
rlabel locali s -3163 -27449 -3117 -27327 2 VDD
port 41 nsew
rlabel locali s -3158 -27327 -3124 -27137 2 VDD
port 41 nsew
rlabel locali s -3360 -27449 -3314 -27315 2 VDD
port 41 nsew
rlabel locali s -3473 -27449 -3427 -27325 2 VDD
port 41 nsew
rlabel locali s -3354 -27315 -3320 -27137 2 VDD
port 41 nsew
rlabel locali s -3467 -27325 -3433 -27137 2 VDD
port 41 nsew
rlabel locali s -3669 -27449 -3623 -27320 2 VDD
port 41 nsew
rlabel locali s -3782 -27449 -3736 -27324 2 VDD
port 41 nsew
rlabel locali s -3663 -27320 -3629 -27137 2 VDD
port 41 nsew
rlabel locali s -3777 -27324 -3743 -27137 2 VDD
port 41 nsew
rlabel locali s -3980 -27449 -3934 -27320 2 VDD
port 41 nsew
rlabel locali s -4169 -27449 -4129 -27320 2 VDD
port 41 nsew
rlabel locali s -3973 -27320 -3939 -27137 2 VDD
port 41 nsew
rlabel locali s -4169 -27320 -4135 -27137 2 VDD
port 41 nsew
rlabel locali s -5342 -27556 -5227 -26719 2 VDD
port 41 nsew
rlabel locali s -6669 -27556 -5617 -27449 2 VDD
port 41 nsew
rlabel locali s -22963 -27582 -20173 -27515 2 VDD
port 41 nsew
rlabel locali s -22775 -27515 -20173 -27499 2 VDD
port 41 nsew
rlabel locali s -5663 -27449 -5617 -27327 2 VDD
port 41 nsew
rlabel locali s -5658 -27327 -5624 -27137 2 VDD
port 41 nsew
rlabel locali s -5860 -27449 -5814 -27315 2 VDD
port 41 nsew
rlabel locali s -5973 -27449 -5927 -27325 2 VDD
port 41 nsew
rlabel locali s -5854 -27315 -5820 -27137 2 VDD
port 41 nsew
rlabel locali s -5967 -27325 -5933 -27137 2 VDD
port 41 nsew
rlabel locali s -6169 -27449 -6123 -27320 2 VDD
port 41 nsew
rlabel locali s -6282 -27449 -6236 -27324 2 VDD
port 41 nsew
rlabel locali s -6163 -27320 -6129 -27137 2 VDD
port 41 nsew
rlabel locali s -6277 -27324 -6243 -27137 2 VDD
port 41 nsew
rlabel locali s -6480 -27449 -6434 -27320 2 VDD
port 41 nsew
rlabel locali s -6669 -27449 -6629 -27320 2 VDD
port 41 nsew
rlabel locali s -6473 -27320 -6439 -27137 2 VDD
port 41 nsew
rlabel locali s -6669 -27320 -6635 -27137 2 VDD
port 41 nsew
rlabel locali s -21627 -27499 -21593 -27223 2 VDD
port 41 nsew
rlabel locali s -21823 -27499 -21789 -27223 2 VDD
port 41 nsew
rlabel locali s -22019 -27499 -21985 -27223 2 VDD
port 41 nsew
rlabel locali s -22215 -27499 -22181 -27223 2 VDD
port 41 nsew
rlabel locali s -22757 -27499 -22723 -27223 2 VDD
port 41 nsew
rlabel locali s -22953 -27515 -22919 -27223 2 VDD
port 41 nsew
rlabel locali s -20349 -27047 -20173 -26960 2 VDD
port 41 nsew
rlabel locali s -297 -26684 -174 -26548 2 VDD
port 41 nsew
rlabel locali s -2780 -26684 -2657 -26548 2 VDD
port 41 nsew
rlabel locali s -5347 -26719 -5224 -26583 2 VDD
port 41 nsew
rlabel locali s -298 -26131 -175 -26130 2 VDD
port 41 nsew
rlabel locali s -298 -26130 8 -26068 2 VDD
port 41 nsew
rlabel locali s -16907 -26271 -16873 -26105 2 VDD
port 41 nsew
rlabel locali s -17103 -26271 -17069 -26105 2 VDD
port 41 nsew
rlabel locali s -17299 -26271 -17265 -26105 2 VDD
port 41 nsew
rlabel locali s -17495 -26271 -17461 -26105 2 VDD
port 41 nsew
rlabel locali s -17712 -26472 -17678 -26105 2 VDD
port 41 nsew
rlabel locali s 16289 -25864 16323 -25573 8 VDD
port 41 nsew
rlabel locali s 16093 -25864 16127 -25573 8 VDD
port 41 nsew
rlabel locali s 15897 -25864 15931 -25573 8 VDD
port 41 nsew
rlabel locali s 14546 -25864 14580 -25573 8 VDD
port 41 nsew
rlabel locali s 14350 -25864 14384 -25573 8 VDD
port 41 nsew
rlabel locali s 14154 -25864 14188 -25573 8 VDD
port 41 nsew
rlabel locali s 13589 -25864 13623 -25573 8 VDD
port 41 nsew
rlabel locali s 13393 -25864 13427 -25573 8 VDD
port 41 nsew
rlabel locali s 13197 -25864 13231 -25573 8 VDD
port 41 nsew
rlabel locali s 11846 -25864 11880 -25573 8 VDD
port 41 nsew
rlabel locali s 11650 -25864 11684 -25573 8 VDD
port 41 nsew
rlabel locali s 11454 -25864 11488 -25573 8 VDD
port 41 nsew
rlabel locali s 10964 -25864 10998 -25573 8 VDD
port 41 nsew
rlabel locali s 10768 -25864 10802 -25573 8 VDD
port 41 nsew
rlabel locali s 10572 -25864 10606 -25573 8 VDD
port 41 nsew
rlabel locali s 15888 -25573 16383 -25570 8 VDD
port 41 nsew
rlabel locali s 13188 -25573 14641 -25572 8 VDD
port 41 nsew
rlabel locali s 15566 -25570 16670 -25568 8 VDD
port 41 nsew
rlabel locali s 12875 -25572 14641 -25568 8 VDD
port 41 nsew
rlabel locali s 10563 -25573 11941 -25568 8 VDD
port 41 nsew
rlabel locali s 10563 -25568 16670 -25505 8 VDD
port 41 nsew
rlabel locali s 15566 -25505 16670 -25502 8 VDD
port 41 nsew
rlabel locali s 12875 -25505 13348 -25504 8 VDD
port 41 nsew
rlabel locali s 28121 -25236 28155 -25070 8 VDD
port 41 nsew
rlabel locali s 27925 -25236 27959 -25070 8 VDD
port 41 nsew
rlabel locali s 27729 -25236 27763 -25070 8 VDD
port 41 nsew
rlabel locali s 27533 -25236 27567 -25070 8 VDD
port 41 nsew
rlabel locali s 27316 -25437 27350 -25070 8 VDD
port 41 nsew
rlabel locali s 28561 -25055 28606 -24932 8 VDD
port 41 nsew
rlabel locali s 28366 -25058 28411 -24932 8 VDD
port 41 nsew
rlabel locali s 27316 -25070 28203 -25020 8 VDD
port 41 nsew
rlabel locali s 27120 -25437 27154 -25020 8 VDD
port 41 nsew
rlabel locali s 26924 -25437 26958 -25020 8 VDD
port 41 nsew
rlabel locali s 20111 -25054 20174 -25043 8 VDD
port 41 nsew
rlabel locali s 18991 -25047 19077 -25043 8 VDD
port 41 nsew
rlabel locali s 21509 -25038 24798 -25030 8 VDD
port 41 nsew
rlabel locali s 20792 -25043 20866 -25037 8 VDD
port 41 nsew
rlabel locali s 18991 -25043 20174 -25037 8 VDD
port 41 nsew
rlabel locali s 18991 -25037 20866 -25031 8 VDD
port 41 nsew
rlabel locali s 16544 -25502 16670 -25031 8 VDD
port 41 nsew
rlabel locali s 6340 -25294 6463 -25267 8 VDD
port 41 nsew
rlabel locali s 6340 -25267 7393 -25198 8 VDD
port 41 nsew
rlabel locali s 7347 -25198 7393 -25076 8 VDD
port 41 nsew
rlabel locali s 16544 -25031 20866 -25030 8 VDD
port 41 nsew
rlabel locali s 26914 -25020 28203 -24971 8 VDD
port 41 nsew
rlabel locali s 26914 -24971 27356 -24956 8 VDD
port 41 nsew
rlabel locali s 16544 -25030 24798 -24974 8 VDD
port 41 nsew
rlabel locali s 20111 -24974 24798 -24970 8 VDD
port 41 nsew
rlabel locali s 20792 -24970 24798 -24962 8 VDD
port 41 nsew
rlabel locali s 21487 -24962 24798 -24935 8 VDD
port 41 nsew
rlabel locali s 28360 -24932 29129 -24908 8 VDD
port 41 nsew
rlabel locali s 27353 -24922 27542 -24915 8 VDD
port 41 nsew
rlabel locali s 27316 -24915 27542 -24908 8 VDD
port 41 nsew
rlabel locali s 32748 -24897 32927 -24861 8 VDD
port 41 nsew
rlabel locali s 30582 -24897 32693 -24886 8 VDD
port 41 nsew
rlabel locali s 32848 -24861 32927 -24830 8 VDD
port 41 nsew
rlabel locali s 29781 -24886 32693 -24820 8 VDD
port 41 nsew
rlabel locali s 36352 -24766 36970 -24749 8 VDD
port 41 nsew
rlabel locali s 36352 -24749 36795 -24720 8 VDD
port 41 nsew
rlabel locali s 36353 -24720 36795 -24706 8 VDD
port 41 nsew
rlabel locali s 36353 -24706 37642 -24657 8 VDD
port 41 nsew
rlabel locali s 36755 -24657 37642 -24607 8 VDD
port 41 nsew
rlabel locali s 37560 -24607 37594 -24441 8 VDD
port 41 nsew
rlabel locali s 37364 -24607 37398 -24441 8 VDD
port 41 nsew
rlabel locali s 37168 -24607 37202 -24441 8 VDD
port 41 nsew
rlabel locali s 36972 -24607 37006 -24441 8 VDD
port 41 nsew
rlabel locali s 36755 -24607 36789 -24240 8 VDD
port 41 nsew
rlabel locali s 36559 -24657 36593 -24240 8 VDD
port 41 nsew
rlabel locali s 36363 -24657 36397 -24240 8 VDD
port 41 nsew
rlabel locali s 35524 -24766 35696 -24576 8 VDD
port 41 nsew
rlabel locali s 35342 -24576 36060 -24477 8 VDD
port 41 nsew
rlabel locali s 35978 -24477 36012 -24211 8 VDD
port 41 nsew
rlabel locali s 35782 -24477 35816 -24211 8 VDD
port 41 nsew
rlabel locali s 35586 -24477 35620 -24211 8 VDD
port 41 nsew
rlabel locali s 35390 -24477 35424 -24211 8 VDD
port 41 nsew
rlabel locali s 33188 -24815 33310 -23819 8 VDD
port 41 nsew
rlabel locali s 30582 -24820 32693 -24786 8 VDD
port 41 nsew
rlabel locali s 31580 -24786 32198 -24769 8 VDD
port 41 nsew
rlabel locali s 31580 -24769 32023 -24740 8 VDD
port 41 nsew
rlabel locali s 31581 -24740 32023 -24726 8 VDD
port 41 nsew
rlabel locali s 31581 -24726 32870 -24677 8 VDD
port 41 nsew
rlabel locali s 31983 -24677 32870 -24627 8 VDD
port 41 nsew
rlabel locali s 32788 -24627 32822 -24461 8 VDD
port 41 nsew
rlabel locali s 32592 -24627 32626 -24461 8 VDD
port 41 nsew
rlabel locali s 32396 -24627 32430 -24461 8 VDD
port 41 nsew
rlabel locali s 32200 -24627 32234 -24461 8 VDD
port 41 nsew
rlabel locali s 31983 -24627 32017 -24260 8 VDD
port 41 nsew
rlabel locali s 31787 -24677 31821 -24260 8 VDD
port 41 nsew
rlabel locali s 31591 -24677 31625 -24260 8 VDD
port 41 nsew
rlabel locali s 30752 -24786 30924 -24596 8 VDD
port 41 nsew
rlabel locali s 30570 -24596 31288 -24497 8 VDD
port 41 nsew
rlabel locali s 31206 -24497 31240 -24231 8 VDD
port 41 nsew
rlabel locali s 31010 -24497 31044 -24231 8 VDD
port 41 nsew
rlabel locali s 30814 -24497 30848 -24231 8 VDD
port 41 nsew
rlabel locali s 30618 -24497 30652 -24231 8 VDD
port 41 nsew
rlabel locali s 32678 -23819 33310 -23697 8 VDD
port 41 nsew
rlabel locali s 37885 -23501 38287 -23435 8 VDD
port 41 nsew
rlabel locali s 40156 -21764 40190 -21472 8 VDD
port 41 nsew
rlabel locali s 39960 -21764 39994 -21474 8 VDD
port 41 nsew
rlabel locali s 39732 -21964 39766 -21489 8 VDD
port 41 nsew
rlabel locali s 39602 -21964 39636 -21492 8 VDD
port 41 nsew
rlabel locali s 40151 -21472 40194 -21401 8 VDD
port 41 nsew
rlabel locali s 40151 -21401 46336 -21352 8 VDD
port 41 nsew
rlabel locali s 47304 -21351 55534 -21318 8 VDD
port 41 nsew
rlabel locali s 45223 -21352 45841 -21335 8 VDD
port 41 nsew
rlabel locali s 56502 -21317 64288 -21264 8 VDD
port 41 nsew
rlabel locali s 54421 -21318 55039 -21301 8 VDD
port 41 nsew
rlabel locali s 54421 -21301 54864 -21272 8 VDD
port 41 nsew
rlabel locali s 47304 -21318 53765 -21298 8 VDD
port 41 nsew
rlabel locali s 45223 -21335 45666 -21306 8 VDD
port 41 nsew
rlabel locali s 40151 -21352 44567 -21312 8 VDD
port 41 nsew
rlabel locali s 39954 -21474 39997 -21312 8 VDD
port 41 nsew
rlabel locali s 39723 -21489 39773 -21312 8 VDD
port 41 nsew
rlabel locali s 39597 -21492 39647 -21312 8 VDD
port 41 nsew
rlabel locali s 39007 -21964 39041 -21469 8 VDD
port 41 nsew
rlabel locali s 38811 -21964 38845 -21471 8 VDD
port 41 nsew
rlabel locali s 37438 -22206 37472 -21614 8 VDD
port 41 nsew
rlabel locali s 37878 -21509 37976 -21503 8 VDD
port 41 nsew
rlabel locali s 39005 -21469 39043 -21312 8 VDD
port 41 nsew
rlabel locali s 38808 -21471 38846 -21376 8 VDD
port 41 nsew
rlabel locali s 37878 -21503 38558 -21386 8 VDD
port 41 nsew
rlabel locali s 37650 -21497 37712 -21483 8 VDD
port 41 nsew
rlabel locali s 37431 -21614 37476 -21490 8 VDD
port 41 nsew
rlabel locali s 37015 -22206 37049 -21613 8 VDD
port 41 nsew
rlabel locali s 36819 -22206 36853 -21616 8 VDD
port 41 nsew
rlabel locali s 36569 -21794 36603 -21628 8 VDD
port 41 nsew
rlabel locali s 36373 -21794 36407 -21628 8 VDD
port 41 nsew
rlabel locali s 36177 -21794 36211 -21628 8 VDD
port 41 nsew
rlabel locali s 35981 -21794 36015 -21628 8 VDD
port 41 nsew
rlabel locali s 35764 -21995 35798 -21628 8 VDD
port 41 nsew
rlabel locali s 37009 -21613 37054 -21490 8 VDD
port 41 nsew
rlabel locali s 36814 -21616 36859 -21490 8 VDD
port 41 nsew
rlabel locali s 35764 -21628 36651 -21578 8 VDD
port 41 nsew
rlabel locali s 35568 -21995 35602 -21578 8 VDD
port 41 nsew
rlabel locali s 35372 -21995 35406 -21578 8 VDD
port 41 nsew
rlabel locali s 35362 -21578 36651 -21529 8 VDD
port 41 nsew
rlabel locali s 35362 -21529 35804 -21514 8 VDD
port 41 nsew
rlabel locali s 36808 -21490 37577 -21483 8 VDD
port 41 nsew
rlabel locali s 36808 -21483 37712 -21466 8 VDD
port 41 nsew
rlabel locali s 35801 -21480 35990 -21473 8 VDD
port 41 nsew
rlabel locali s 35764 -21473 35990 -21466 8 VDD
port 41 nsew
rlabel locali s 32678 -23697 32800 -21466 8 VDD
port 41 nsew
rlabel locali s 29781 -24820 29847 -23490 8 VDD
port 41 nsew
rlabel locali s 29428 -24904 29512 -24791 8 VDD
port 41 nsew
rlabel locali s 26914 -24908 29129 -24866 8 VDD
port 41 nsew
rlabel locali s 29445 -24791 29511 -23490 8 VDD
port 41 nsew
rlabel locali s 26914 -24866 29025 -24755 8 VDD
port 41 nsew
rlabel locali s 27912 -24755 28530 -24738 8 VDD
port 41 nsew
rlabel locali s 27912 -24738 28355 -24709 8 VDD
port 41 nsew
rlabel locali s 27913 -24709 28355 -24695 8 VDD
port 41 nsew
rlabel locali s 27913 -24695 29202 -24646 8 VDD
port 41 nsew
rlabel locali s 28315 -24646 29202 -24596 8 VDD
port 41 nsew
rlabel locali s 29120 -24596 29154 -24430 8 VDD
port 41 nsew
rlabel locali s 28924 -24596 28958 -24430 8 VDD
port 41 nsew
rlabel locali s 28728 -24596 28762 -24430 8 VDD
port 41 nsew
rlabel locali s 28532 -24596 28566 -24430 8 VDD
port 41 nsew
rlabel locali s 28315 -24596 28349 -24229 8 VDD
port 41 nsew
rlabel locali s 28119 -24646 28153 -24229 8 VDD
port 41 nsew
rlabel locali s 27923 -24646 27957 -24229 8 VDD
port 41 nsew
rlabel locali s 27084 -24755 27256 -24565 8 VDD
port 41 nsew
rlabel locali s 26902 -24565 27620 -24466 8 VDD
port 41 nsew
rlabel locali s 27538 -24466 27572 -24200 8 VDD
port 41 nsew
rlabel locali s 27342 -24466 27376 -24200 8 VDD
port 41 nsew
rlabel locali s 27146 -24466 27180 -24200 8 VDD
port 41 nsew
rlabel locali s 26950 -24466 26984 -24200 8 VDD
port 41 nsew
rlabel locali s 29445 -23490 29847 -23424 8 VDD
port 41 nsew
rlabel locali s 24709 -24935 24798 -22780 8 VDD
port 41 nsew
rlabel locali s 24571 -24935 24605 -24100 8 VDD
port 41 nsew
rlabel locali s 24375 -24935 24409 -24100 8 VDD
port 41 nsew
rlabel locali s 24171 -24935 24205 -24100 8 VDD
port 41 nsew
rlabel locali s 23975 -24935 24009 -24100 8 VDD
port 41 nsew
rlabel locali s 23571 -24935 23605 -24100 8 VDD
port 41 nsew
rlabel locali s 23375 -24935 23409 -24100 8 VDD
port 41 nsew
rlabel locali s 23171 -24935 23205 -24100 8 VDD
port 41 nsew
rlabel locali s 22975 -24935 23009 -24100 8 VDD
port 41 nsew
rlabel locali s 22571 -24935 22605 -24100 8 VDD
port 41 nsew
rlabel locali s 22375 -24935 22409 -24100 8 VDD
port 41 nsew
rlabel locali s 22171 -24935 22205 -24100 8 VDD
port 41 nsew
rlabel locali s 21975 -24935 22009 -24100 8 VDD
port 41 nsew
rlabel locali s 21487 -24935 21521 -24671 8 VDD
port 41 nsew
rlabel locali s 21291 -24962 21325 -24671 8 VDD
port 41 nsew
rlabel locali s 21095 -24962 21129 -24671 8 VDD
port 41 nsew
rlabel locali s 20792 -24962 20866 -24956 8 VDD
port 41 nsew
rlabel locali s 20562 -24970 20596 -24678 8 VDD
port 41 nsew
rlabel locali s 20366 -24970 20400 -24678 8 VDD
port 41 nsew
rlabel locali s 20111 -24970 20174 -24956 8 VDD
port 41 nsew
rlabel locali s 19824 -24974 19858 -24678 8 VDD
port 41 nsew
rlabel locali s 19628 -24974 19662 -24678 8 VDD
port 41 nsew
rlabel locali s 19432 -24974 19466 -24678 8 VDD
port 41 nsew
rlabel locali s 19236 -24974 19270 -24678 8 VDD
port 41 nsew
rlabel locali s 16544 -24974 19077 -24962 8 VDD
port 41 nsew
rlabel locali s 18991 -24962 19077 -24954 8 VDD
port 41 nsew
rlabel locali s 18510 -24962 18558 -24829 8 VDD
port 41 nsew
rlabel locali s 18313 -24962 18361 -24835 8 VDD
port 41 nsew
rlabel locali s 18516 -24829 18550 -24444 8 VDD
port 41 nsew
rlabel locali s 18320 -24835 18354 -24444 8 VDD
port 41 nsew
rlabel locali s 17564 -24962 17612 -24829 8 VDD
port 41 nsew
rlabel locali s 17367 -24962 17415 -24835 8 VDD
port 41 nsew
rlabel locali s 7352 -25076 7386 -24886 8 VDD
port 41 nsew
rlabel locali s 7150 -25198 7196 -25064 8 VDD
port 41 nsew
rlabel locali s 7037 -25198 7083 -25074 8 VDD
port 41 nsew
rlabel locali s 7156 -25064 7190 -24886 8 VDD
port 41 nsew
rlabel locali s 7043 -25074 7077 -24886 8 VDD
port 41 nsew
rlabel locali s 6841 -25198 6887 -25069 8 VDD
port 41 nsew
rlabel locali s 6728 -25198 6774 -25073 8 VDD
port 41 nsew
rlabel locali s 6847 -25069 6881 -24886 8 VDD
port 41 nsew
rlabel locali s 6733 -25073 6767 -24886 8 VDD
port 41 nsew
rlabel locali s 6530 -25198 6576 -25069 8 VDD
port 41 nsew
rlabel locali s 6340 -25198 6463 -25158 8 VDD
port 41 nsew
rlabel locali s 5124 -25295 5247 -25262 8 VDD
port 41 nsew
rlabel locali s 3768 -25300 3891 -25267 8 VDD
port 41 nsew
rlabel locali s 3768 -25267 4664 -25262 8 VDD
port 41 nsew
rlabel locali s 3768 -25262 5247 -25194 8 VDD
port 41 nsew
rlabel locali s 4592 -25194 5247 -25193 8 VDD
port 41 nsew
rlabel locali s 5124 -25193 5247 -25159 8 VDD
port 41 nsew
rlabel locali s 6341 -25158 6381 -25069 8 VDD
port 41 nsew
rlabel locali s 6537 -25069 6571 -24886 8 VDD
port 41 nsew
rlabel locali s 6341 -25069 6375 -24886 8 VDD
port 41 nsew
rlabel locali s 5180 -25159 5214 -24897 8 VDD
port 41 nsew
rlabel locali s 4984 -25193 5018 -24897 8 VDD
port 41 nsew
rlabel locali s 4788 -25193 4822 -24897 8 VDD
port 41 nsew
rlabel locali s 4592 -25193 4626 -24897 8 VDD
port 41 nsew
rlabel locali s 3768 -25194 4089 -25189 8 VDD
port 41 nsew
rlabel locali s 4050 -25189 4084 -24897 8 VDD
port 41 nsew
rlabel locali s 3768 -25189 3891 -25164 8 VDD
port 41 nsew
rlabel locali s 3367 -25298 3490 -25253 8 VDD
port 41 nsew
rlabel locali s 3029 -25253 3490 -25238 8 VDD
port 41 nsew
rlabel locali s 2139 -25275 2262 -25238 8 VDD
port 41 nsew
rlabel locali s 2139 -25238 3490 -25189 8 VDD
port 41 nsew
rlabel locali s 3854 -25164 3888 -24897 8 VDD
port 41 nsew
rlabel locali s 3367 -25189 3490 -25162 8 VDD
port 41 nsew
rlabel locali s 17570 -24829 17604 -24444 8 VDD
port 41 nsew
rlabel locali s 17374 -24835 17408 -24444 8 VDD
port 41 nsew
rlabel locali s 3427 -25162 3461 -24772 8 VDD
port 41 nsew
rlabel locali s 3231 -25189 3265 -24772 8 VDD
port 41 nsew
rlabel locali s 2139 -25189 3069 -25139 8 VDD
port 41 nsew
rlabel locali s 1750 -25274 1873 -25260 8 VDD
port 41 nsew
rlabel locali s -293 -26068 -178 -25260 2 VDD
port 41 nsew
rlabel locali s -2781 -26096 -2658 -25960 2 VDD
port 41 nsew
rlabel locali s -17712 -26105 -16825 -26055 2 VDD
port 41 nsew
rlabel locali s -17908 -26472 -17874 -26055 2 VDD
port 41 nsew
rlabel locali s -18104 -26472 -18070 -26055 2 VDD
port 41 nsew
rlabel locali s -18489 -26501 -18455 -26235 2 VDD
port 41 nsew
rlabel locali s -18685 -26501 -18651 -26235 2 VDD
port 41 nsew
rlabel locali s -18881 -26501 -18847 -26235 2 VDD
port 41 nsew
rlabel locali s -19077 -26501 -19043 -26235 2 VDD
port 41 nsew
rlabel locali s -19125 -26235 -18407 -26136 2 VDD
port 41 nsew
rlabel locali s -18114 -26055 -16825 -26006 2 VDD
port 41 nsew
rlabel locali s -18114 -26006 -17672 -25992 2 VDD
port 41 nsew
rlabel locali s -18115 -25992 -17672 -25963 2 VDD
port 41 nsew
rlabel locali s -1228 -25287 -1105 -25260 2 VDD
port 41 nsew
rlabel locali s -1228 -25260 1873 -25181 8 VDD
port 41 nsew
rlabel locali s 3035 -25139 3069 -24772 8 VDD
port 41 nsew
rlabel locali s 2818 -25139 2852 -24973 8 VDD
port 41 nsew
rlabel locali s 2622 -25139 2656 -24973 8 VDD
port 41 nsew
rlabel locali s 2426 -25139 2460 -24973 8 VDD
port 41 nsew
rlabel locali s 2230 -25139 2264 -24973 8 VDD
port 41 nsew
rlabel locali s 1750 -25181 1873 -25138 8 VDD
port 41 nsew
rlabel locali s 1822 -25138 1856 -24774 8 VDD
port 41 nsew
rlabel locali s 1626 -25181 1660 -24774 8 VDD
port 41 nsew
rlabel locali s 577 -25181 1464 -25141 8 VDD
port 41 nsew
rlabel locali s 1430 -25141 1464 -24774 8 VDD
port 41 nsew
rlabel locali s 1213 -25141 1247 -24975 8 VDD
port 41 nsew
rlabel locali s 1017 -25141 1051 -24975 8 VDD
port 41 nsew
rlabel locali s 821 -25141 855 -24975 8 VDD
port 41 nsew
rlabel locali s 625 -25141 659 -24975 8 VDD
port 41 nsew
rlabel locali s 218 -25181 252 -24888 8 VDD
port 41 nsew
rlabel locali s 22 -25181 56 -24888 8 VDD
port 41 nsew
rlabel locali s -174 -25181 -140 -24888 2 VDD
port 41 nsew
rlabel locali s -370 -25181 -336 -24888 2 VDD
port 41 nsew
rlabel locali s -1228 -25181 -873 -25180 2 VDD
port 41 nsew
rlabel locali s -912 -25180 -878 -24888 2 VDD
port 41 nsew
rlabel locali s -1228 -25180 -1074 -25151 2 VDD
port 41 nsew
rlabel locali s -1522 -25286 -1399 -25264 2 VDD
port 41 nsew
rlabel locali s -2777 -25960 -2662 -25264 2 VDD
port 41 nsew
rlabel locali s -5348 -25952 -5225 -25816 2 VDD
port 41 nsew
rlabel locali s -18115 -25963 -17497 -25946 2 VDD
port 41 nsew
rlabel locali s -18943 -26136 -18771 -25965 2 VDD
port 41 nsew
rlabel locali s -20347 -26960 -20175 -25965 2 VDD
port 41 nsew
rlabel locali s -20347 -25965 -18771 -25946 2 VDD
port 41 nsew
rlabel locali s -20347 -25946 -17002 -25835 2 VDD
port 41 nsew
rlabel locali s -4192 -25265 -3719 -25264 2 VDD
port 41 nsew
rlabel locali s -5343 -25816 -5228 -25264 2 VDD
port 41 nsew
rlabel locali s -20347 -25835 -16898 -25793 2 VDD
port 41 nsew
rlabel locali s -17667 -25793 -16898 -25769 2 VDD
port 41 nsew
rlabel locali s -18711 -25793 -18485 -25786 2 VDD
port 41 nsew
rlabel locali s -18674 -25786 -18485 -25779 2 VDD
port 41 nsew
rlabel locali s -17044 -25769 -16999 -25645 2 VDD
port 41 nsew
rlabel locali s -17466 -25769 -17421 -25646 2 VDD
port 41 nsew
rlabel locali s -7514 -25267 -6410 -25264 2 VDD
port 41 nsew
rlabel locali s -7514 -25264 -1399 -25201 2 VDD
port 41 nsew
rlabel locali s -2785 -25201 -1399 -25196 2 VDD
port 41 nsew
rlabel locali s -5485 -25201 -3719 -25197 2 VDD
port 41 nsew
rlabel locali s -7514 -25201 -6410 -25199 2 VDD
port 41 nsew
rlabel locali s -5485 -25197 -4032 -25196 2 VDD
port 41 nsew
rlabel locali s -7227 -25199 -6732 -25196 2 VDD
port 41 nsew
rlabel locali s -1108 -25151 -1074 -24888 2 VDD
port 41 nsew
rlabel locali s -1522 -25196 -1399 -25150 2 VDD
port 41 nsew
rlabel locali s -1450 -25150 -1416 -24905 2 VDD
port 41 nsew
rlabel locali s -1646 -25196 -1612 -24905 2 VDD
port 41 nsew
rlabel locali s -1842 -25196 -1808 -24905 2 VDD
port 41 nsew
rlabel locali s -2332 -25196 -2298 -24905 2 VDD
port 41 nsew
rlabel locali s -2528 -25196 -2494 -24905 2 VDD
port 41 nsew
rlabel locali s -2724 -25196 -2690 -24905 2 VDD
port 41 nsew
rlabel locali s -4075 -25196 -4041 -24905 2 VDD
port 41 nsew
rlabel locali s -4271 -25196 -4237 -24905 2 VDD
port 41 nsew
rlabel locali s -4467 -25196 -4433 -24905 2 VDD
port 41 nsew
rlabel locali s -5032 -25196 -4998 -24905 2 VDD
port 41 nsew
rlabel locali s -5228 -25196 -5194 -24905 2 VDD
port 41 nsew
rlabel locali s -5424 -25196 -5390 -24905 2 VDD
port 41 nsew
rlabel locali s -6775 -25196 -6741 -24905 2 VDD
port 41 nsew
rlabel locali s -6971 -25196 -6937 -24905 2 VDD
port 41 nsew
rlabel locali s -7167 -25196 -7133 -24905 2 VDD
port 41 nsew
rlabel locali s 21537 -23578 21571 -23061 8 VDD
port 41 nsew
rlabel locali s 21341 -23578 21375 -23061 8 VDD
port 41 nsew
rlabel locali s 21145 -23578 21179 -23061 8 VDD
port 41 nsew
rlabel locali s -3336 -23795 -3302 -23504 2 VDD
port 41 nsew
rlabel locali s -3532 -23795 -3498 -23504 2 VDD
port 41 nsew
rlabel locali s -3728 -23795 -3694 -23504 2 VDD
port 41 nsew
rlabel locali s -4173 -23795 -4139 -23504 2 VDD
port 41 nsew
rlabel locali s -4369 -23795 -4335 -23504 2 VDD
port 41 nsew
rlabel locali s -4565 -23795 -4531 -23504 2 VDD
port 41 nsew
rlabel locali s -6036 -23795 -6002 -23504 2 VDD
port 41 nsew
rlabel locali s -6232 -23795 -6198 -23504 2 VDD
port 41 nsew
rlabel locali s -6428 -23795 -6394 -23504 2 VDD
port 41 nsew
rlabel locali s -6873 -23795 -6839 -23504 2 VDD
port 41 nsew
rlabel locali s -7069 -23795 -7035 -23504 2 VDD
port 41 nsew
rlabel locali s -7265 -23795 -7231 -23504 2 VDD
port 41 nsew
rlabel locali s -7514 -25199 -7425 -23504 2 VDD
port 41 nsew
rlabel locali s -17037 -25645 -17003 -25053 2 VDD
port 41 nsew
rlabel locali s -17460 -25646 -17426 -25053 2 VDD
port 41 nsew
rlabel locali s -17661 -25769 -17616 -25643 2 VDD
port 41 nsew
rlabel locali s -19113 -25745 -18671 -25730 2 VDD
port 41 nsew
rlabel locali s -19113 -25730 -17824 -25681 2 VDD
port 41 nsew
rlabel locali s -17656 -25643 -17622 -25053 2 VDD
port 41 nsew
rlabel locali s -18711 -25681 -17824 -25631 2 VDD
port 41 nsew
rlabel locali s -17906 -25631 -17872 -25465 2 VDD
port 41 nsew
rlabel locali s -18102 -25631 -18068 -25465 2 VDD
port 41 nsew
rlabel locali s -18298 -25631 -18264 -25465 2 VDD
port 41 nsew
rlabel locali s -18494 -25631 -18460 -25465 2 VDD
port 41 nsew
rlabel locali s -18711 -25631 -18677 -25264 2 VDD
port 41 nsew
rlabel locali s -18907 -25681 -18873 -25264 2 VDD
port 41 nsew
rlabel locali s -19103 -25681 -19069 -25264 2 VDD
port 41 nsew
rlabel locali s -12066 -24998 -11593 -24997 2 VDD
port 41 nsew
rlabel locali s -15388 -25000 -14284 -24997 2 VDD
port 41 nsew
rlabel locali s -15388 -24997 -9281 -24934 2 VDD
port 41 nsew
rlabel locali s -10659 -24934 -9281 -24929 2 VDD
port 41 nsew
rlabel locali s -13359 -24934 -11593 -24930 2 VDD
port 41 nsew
rlabel locali s -15388 -24934 -14284 -24932 2 VDD
port 41 nsew
rlabel locali s -13359 -24930 -11906 -24929 2 VDD
port 41 nsew
rlabel locali s -15101 -24932 -14606 -24929 2 VDD
port 41 nsew
rlabel locali s -9324 -24929 -9290 -24638 2 VDD
port 41 nsew
rlabel locali s -9520 -24929 -9486 -24638 2 VDD
port 41 nsew
rlabel locali s -9716 -24929 -9682 -24638 2 VDD
port 41 nsew
rlabel locali s -10206 -24929 -10172 -24638 2 VDD
port 41 nsew
rlabel locali s -10402 -24929 -10368 -24638 2 VDD
port 41 nsew
rlabel locali s -10598 -24929 -10564 -24638 2 VDD
port 41 nsew
rlabel locali s -11949 -24929 -11915 -24638 2 VDD
port 41 nsew
rlabel locali s -12145 -24929 -12111 -24638 2 VDD
port 41 nsew
rlabel locali s -12341 -24929 -12307 -24638 2 VDD
port 41 nsew
rlabel locali s -12906 -24929 -12872 -24638 2 VDD
port 41 nsew
rlabel locali s -13102 -24929 -13068 -24638 2 VDD
port 41 nsew
rlabel locali s -13298 -24929 -13264 -24638 2 VDD
port 41 nsew
rlabel locali s -14649 -24929 -14615 -24638 2 VDD
port 41 nsew
rlabel locali s -14845 -24929 -14811 -24638 2 VDD
port 41 nsew
rlabel locali s -15041 -24929 -15007 -24638 2 VDD
port 41 nsew
rlabel locali s -15388 -24932 -15299 -24029 2 VDD
port 41 nsew
rlabel locali s -20309 -24743 -20275 -24358 2 VDD
port 41 nsew
rlabel locali s -20315 -24358 -20267 -24225 2 VDD
port 41 nsew
rlabel locali s -20505 -24743 -20471 -24352 2 VDD
port 41 nsew
rlabel locali s -21214 -24742 -21180 -24357 2 VDD
port 41 nsew
rlabel locali s -20512 -24352 -20464 -24225 2 VDD
port 41 nsew
rlabel locali s -20517 -24225 -19963 -24197 2 VDD
port 41 nsew
rlabel locali s -21220 -24357 -21172 -24224 2 VDD
port 41 nsew
rlabel locali s -21410 -24742 -21376 -24351 2 VDD
port 41 nsew
rlabel locali s -22420 -25013 -22386 -24429 2 VDD
port 41 nsew
rlabel locali s -21417 -24351 -21369 -24224 2 VDD
port 41 nsew
rlabel locali s -22429 -24429 -22376 -24301 2 VDD
port 41 nsew
rlabel locali s -22616 -25013 -22582 -24413 2 VDD
port 41 nsew
rlabel locali s -22625 -24413 -22572 -24301 2 VDD
port 41 nsew
rlabel locali s -20518 -24197 -19963 -24156 2 VDD
port 41 nsew
rlabel locali s -20518 -24156 -19965 -24029 2 VDD
port 41 nsew
rlabel locali s -21422 -24224 -20868 -24155 2 VDD
port 41 nsew
rlabel locali s -22625 -24301 -21757 -24168 2 VDD
port 41 nsew
rlabel locali s -21407 -24155 -20889 -24029 2 VDD
port 41 nsew
rlabel locali s -22565 -24168 -21783 -24029 2 VDD
port 41 nsew
rlabel locali s -5043 -23504 -3241 -23499 2 VDD
port 41 nsew
rlabel locali s -7514 -23504 -5941 -23499 2 VDD
port 41 nsew
rlabel locali s -7514 -23499 -2289 -23436 2 VDD
port 41 nsew
rlabel locali s 21135 -23061 21577 -22997 8 VDD
port 41 nsew
rlabel locali s 23694 -22780 24798 -22777 8 VDD
port 41 nsew
rlabel locali s 21193 -22997 21425 -22778 8 VDD
port 41 nsew
rlabel locali s 21003 -22778 21476 -22777 8 VDD
port 41 nsew
rlabel locali s 18691 -22777 24798 -22714 8 VDD
port 41 nsew
rlabel locali s 23694 -22714 24798 -22712 8 VDD
port 41 nsew
rlabel locali s 32678 -21466 37712 -21431 8 VDD
port 41 nsew
rlabel locali s 31716 -21753 31750 -21461 8 VDD
port 41 nsew
rlabel locali s 31520 -21753 31554 -21463 8 VDD
port 41 nsew
rlabel locali s 31292 -21953 31326 -21478 8 VDD
port 41 nsew
rlabel locali s 31162 -21953 31196 -21481 8 VDD
port 41 nsew
rlabel locali s 37650 -21431 37712 -21403 8 VDD
port 41 nsew
rlabel locali s 32678 -21431 37577 -21424 8 VDD
port 41 nsew
rlabel locali s 38441 -21386 38558 -21376 8 VDD
port 41 nsew
rlabel locali s 37878 -21386 37976 -21383 8 VDD
port 41 nsew
rlabel locali s 38441 -21376 38846 -21312 8 VDD
port 41 nsew
rlabel locali s 32678 -21424 37473 -21313 8 VDD
port 41 nsew
rlabel locali s 56869 -21264 64288 -21252 8 VDD
port 41 nsew
rlabel locali s 54422 -21272 54864 -21258 8 VDD
port 41 nsew
rlabel locali s 65256 -21251 73441 -21235 8 VDD
port 41 nsew
rlabel locali s 63175 -21252 63793 -21235 8 VDD
port 41 nsew
rlabel locali s 74409 -21234 82805 -21197 8 VDD
port 41 nsew
rlabel locali s 72328 -21235 72946 -21218 8 VDD
port 41 nsew
rlabel locali s 83773 -21196 85526 -21195 8 VDD
port 41 nsew
rlabel locali s 83773 -21195 86572 -21143 8 VDD
port 41 nsew
rlabel locali s 81692 -21197 82310 -21180 8 VDD
port 41 nsew
rlabel locali s 81692 -21180 82135 -21151 8 VDD
port 41 nsew
rlabel locali s 74409 -21197 81036 -21181 8 VDD
port 41 nsew
rlabel locali s 72328 -21218 72771 -21189 8 VDD
port 41 nsew
rlabel locali s 65256 -21235 71672 -21198 8 VDD
port 41 nsew
rlabel locali s 63175 -21235 63618 -21206 8 VDD
port 41 nsew
rlabel locali s 84140 -21143 86572 -21073 8 VDD
port 41 nsew
rlabel locali s 81693 -21151 82135 -21137 8 VDD
port 41 nsew
rlabel locali s 81693 -21137 82982 -21088 8 VDD
port 41 nsew
rlabel locali s 74776 -21181 81036 -21111 8 VDD
port 41 nsew
rlabel locali s 72329 -21189 72771 -21175 8 VDD
port 41 nsew
rlabel locali s 72329 -21175 73618 -21126 8 VDD
port 41 nsew
rlabel locali s 65623 -21198 71672 -21128 8 VDD
port 41 nsew
rlabel locali s 63176 -21206 63618 -21192 8 VDD
port 41 nsew
rlabel locali s 63176 -21192 64465 -21143 8 VDD
port 41 nsew
rlabel locali s 56869 -21252 62519 -21194 8 VDD
port 41 nsew
rlabel locali s 54422 -21258 55711 -21209 8 VDD
port 41 nsew
rlabel locali s 47671 -21298 53765 -21228 8 VDD
port 41 nsew
rlabel locali s 45224 -21306 45666 -21292 8 VDD
port 41 nsew
rlabel locali s 45224 -21292 46513 -21243 8 VDD
port 41 nsew
rlabel locali s 38441 -21312 44567 -21259 8 VDD
port 41 nsew
rlabel locali s 36360 -21313 36978 -21296 8 VDD
port 41 nsew
rlabel locali s 36360 -21296 36803 -21267 8 VDD
port 41 nsew
rlabel locali s 85898 -21073 86373 -17161 8 VDD
port 41 nsew
rlabel locali s 82095 -21088 82982 -21038 8 VDD
port 41 nsew
rlabel locali s 82900 -21038 82934 -20872 8 VDD
port 41 nsew
rlabel locali s 82704 -21038 82738 -20872 8 VDD
port 41 nsew
rlabel locali s 82508 -21038 82542 -20872 8 VDD
port 41 nsew
rlabel locali s 82312 -21038 82346 -20872 8 VDD
port 41 nsew
rlabel locali s 82095 -21038 82129 -20671 8 VDD
port 41 nsew
rlabel locali s 81899 -21088 81933 -20671 8 VDD
port 41 nsew
rlabel locali s 81703 -21088 81737 -20671 8 VDD
port 41 nsew
rlabel locali s 76123 -21111 81036 -21007 8 VDD
port 41 nsew
rlabel locali s 72731 -21126 73618 -21076 8 VDD
port 41 nsew
rlabel locali s 76123 -21007 81400 -20952 8 VDD
port 41 nsew
rlabel locali s 80682 -20952 81400 -20908 8 VDD
port 41 nsew
rlabel locali s 73536 -21076 73570 -20910 8 VDD
port 41 nsew
rlabel locali s 73340 -21076 73374 -20910 8 VDD
port 41 nsew
rlabel locali s 73144 -21076 73178 -20910 8 VDD
port 41 nsew
rlabel locali s 72948 -21076 72982 -20910 8 VDD
port 41 nsew
rlabel locali s 81318 -20908 81352 -20642 8 VDD
port 41 nsew
rlabel locali s 81122 -20908 81156 -20642 8 VDD
port 41 nsew
rlabel locali s 80926 -20908 80960 -20642 8 VDD
port 41 nsew
rlabel locali s 80730 -20908 80764 -20642 8 VDD
port 41 nsew
rlabel locali s 72731 -21076 72765 -20709 8 VDD
port 41 nsew
rlabel locali s 72535 -21126 72569 -20709 8 VDD
port 41 nsew
rlabel locali s 72339 -21126 72373 -20709 8 VDD
port 41 nsew
rlabel locali s 66961 -21128 71672 -21045 8 VDD
port 41 nsew
rlabel locali s 63578 -21143 64465 -21093 8 VDD
port 41 nsew
rlabel locali s 66961 -21045 72036 -21021 8 VDD
port 41 nsew
rlabel locali s 71318 -21021 72036 -20946 8 VDD
port 41 nsew
rlabel locali s 71954 -20946 71988 -20680 8 VDD
port 41 nsew
rlabel locali s 71758 -20946 71792 -20680 8 VDD
port 41 nsew
rlabel locali s 71562 -20946 71596 -20680 8 VDD
port 41 nsew
rlabel locali s 71366 -20946 71400 -20680 8 VDD
port 41 nsew
rlabel locali s 64383 -21093 64417 -20927 8 VDD
port 41 nsew
rlabel locali s 64187 -21093 64221 -20927 8 VDD
port 41 nsew
rlabel locali s 63991 -21093 64025 -20927 8 VDD
port 41 nsew
rlabel locali s 63795 -21093 63829 -20927 8 VDD
port 41 nsew
rlabel locali s 63578 -21093 63612 -20726 8 VDD
port 41 nsew
rlabel locali s 63382 -21143 63416 -20726 8 VDD
port 41 nsew
rlabel locali s 63186 -21143 63220 -20726 8 VDD
port 41 nsew
rlabel locali s 58214 -21194 62519 -21062 8 VDD
port 41 nsew
rlabel locali s 54824 -21209 55711 -21159 8 VDD
port 41 nsew
rlabel locali s 58214 -21062 62883 -21000 8 VDD
port 41 nsew
rlabel locali s 62165 -21000 62883 -20963 8 VDD
port 41 nsew
rlabel locali s 55629 -21159 55663 -20993 8 VDD
port 41 nsew
rlabel locali s 55433 -21159 55467 -20993 8 VDD
port 41 nsew
rlabel locali s 55237 -21159 55271 -20993 8 VDD
port 41 nsew
rlabel locali s 55041 -21159 55075 -20993 8 VDD
port 41 nsew
rlabel locali s 62801 -20963 62835 -20697 8 VDD
port 41 nsew
rlabel locali s 62605 -20963 62639 -20697 8 VDD
port 41 nsew
rlabel locali s 62409 -20963 62443 -20697 8 VDD
port 41 nsew
rlabel locali s 62213 -20963 62247 -20697 8 VDD
port 41 nsew
rlabel locali s 54824 -21159 54858 -20792 8 VDD
port 41 nsew
rlabel locali s 54628 -21209 54662 -20792 8 VDD
port 41 nsew
rlabel locali s 54432 -21209 54466 -20792 8 VDD
port 41 nsew
rlabel locali s 49031 -21228 53765 -21128 8 VDD
port 41 nsew
rlabel locali s 45626 -21243 46513 -21193 8 VDD
port 41 nsew
rlabel locali s 49031 -21128 54129 -21097 8 VDD
port 41 nsew
rlabel locali s 53411 -21097 54129 -21029 8 VDD
port 41 nsew
rlabel locali s 54047 -21029 54081 -20763 8 VDD
port 41 nsew
rlabel locali s 53851 -21029 53885 -20763 8 VDD
port 41 nsew
rlabel locali s 53655 -21029 53689 -20763 8 VDD
port 41 nsew
rlabel locali s 53459 -21029 53493 -20763 8 VDD
port 41 nsew
rlabel locali s 46431 -21193 46465 -21027 8 VDD
port 41 nsew
rlabel locali s 46235 -21193 46269 -21027 8 VDD
port 41 nsew
rlabel locali s 46039 -21193 46073 -21027 8 VDD
port 41 nsew
rlabel locali s 45843 -21193 45877 -21027 8 VDD
port 41 nsew
rlabel locali s 45626 -21193 45660 -20826 8 VDD
port 41 nsew
rlabel locali s 45430 -21243 45464 -20826 8 VDD
port 41 nsew
rlabel locali s 45234 -21243 45268 -20826 8 VDD
port 41 nsew
rlabel locali s 38808 -21259 44567 -21189 8 VDD
port 41 nsew
rlabel locali s 36361 -21267 36803 -21253 8 VDD
port 41 nsew
rlabel locali s 36361 -21253 37650 -21204 8 VDD
port 41 nsew
rlabel locali s 40180 -21189 44567 -21162 8 VDD
port 41 nsew
rlabel locali s 40180 -21162 44931 -21147 8 VDD
port 41 nsew
rlabel locali s 36763 -21204 37650 -21154 8 VDD
port 41 nsew
rlabel locali s 44213 -21147 44931 -21063 8 VDD
port 41 nsew
rlabel locali s 44849 -21063 44883 -20797 8 VDD
port 41 nsew
rlabel locali s 44653 -21063 44687 -20797 8 VDD
port 41 nsew
rlabel locali s 44457 -21063 44491 -20797 8 VDD
port 41 nsew
rlabel locali s 44261 -21063 44295 -20797 8 VDD
port 41 nsew
rlabel locali s 37568 -21154 37602 -20988 8 VDD
port 41 nsew
rlabel locali s 37372 -21154 37406 -20988 8 VDD
port 41 nsew
rlabel locali s 37176 -21154 37210 -20988 8 VDD
port 41 nsew
rlabel locali s 36980 -21154 37014 -20988 8 VDD
port 41 nsew
rlabel locali s 36763 -21154 36797 -20787 8 VDD
port 41 nsew
rlabel locali s 36567 -21204 36601 -20787 8 VDD
port 41 nsew
rlabel locali s 36371 -21204 36405 -20787 8 VDD
port 41 nsew
rlabel locali s 35532 -21313 35704 -21123 8 VDD
port 41 nsew
rlabel locali s 32678 -21313 32800 -21300 8 VDD
port 41 nsew
rlabel locali s 31711 -21461 31754 -21301 8 VDD
port 41 nsew
rlabel locali s 31514 -21463 31557 -21301 8 VDD
port 41 nsew
rlabel locali s 31283 -21478 31333 -21301 8 VDD
port 41 nsew
rlabel locali s 31157 -21481 31207 -21301 8 VDD
port 41 nsew
rlabel locali s 30567 -21953 30601 -21458 8 VDD
port 41 nsew
rlabel locali s 30371 -21953 30405 -21460 8 VDD
port 41 nsew
rlabel locali s 28998 -22195 29032 -21603 8 VDD
port 41 nsew
rlabel locali s 29438 -21498 29536 -21492 8 VDD
port 41 nsew
rlabel locali s 30565 -21458 30603 -21301 8 VDD
port 41 nsew
rlabel locali s 30368 -21460 30406 -21365 8 VDD
port 41 nsew
rlabel locali s 29438 -21492 30118 -21375 8 VDD
port 41 nsew
rlabel locali s 29210 -21486 29272 -21472 8 VDD
port 41 nsew
rlabel locali s 28991 -21603 29036 -21479 8 VDD
port 41 nsew
rlabel locali s 28575 -22195 28609 -21602 8 VDD
port 41 nsew
rlabel locali s 28379 -22195 28413 -21605 8 VDD
port 41 nsew
rlabel locali s 28129 -21783 28163 -21617 8 VDD
port 41 nsew
rlabel locali s 27933 -21783 27967 -21617 8 VDD
port 41 nsew
rlabel locali s 27737 -21783 27771 -21617 8 VDD
port 41 nsew
rlabel locali s 27541 -21783 27575 -21617 8 VDD
port 41 nsew
rlabel locali s 27324 -21984 27358 -21617 8 VDD
port 41 nsew
rlabel locali s 28569 -21602 28614 -21479 8 VDD
port 41 nsew
rlabel locali s 28374 -21605 28419 -21479 8 VDD
port 41 nsew
rlabel locali s 27324 -21617 28211 -21567 8 VDD
port 41 nsew
rlabel locali s 27128 -21984 27162 -21567 8 VDD
port 41 nsew
rlabel locali s 26932 -21984 26966 -21567 8 VDD
port 41 nsew
rlabel locali s 26922 -21567 28211 -21518 8 VDD
port 41 nsew
rlabel locali s 26922 -21518 27364 -21503 8 VDD
port 41 nsew
rlabel locali s 28368 -21479 29137 -21472 8 VDD
port 41 nsew
rlabel locali s 28368 -21472 29272 -21455 8 VDD
port 41 nsew
rlabel locali s 27361 -21469 27550 -21462 8 VDD
port 41 nsew
rlabel locali s 27324 -21462 27550 -21455 8 VDD
port 41 nsew
rlabel locali s 26922 -21455 29272 -21420 8 VDD
port 41 nsew
rlabel locali s 29210 -21420 29272 -21392 8 VDD
port 41 nsew
rlabel locali s 26922 -21420 29137 -21413 8 VDD
port 41 nsew
rlabel locali s 30001 -21375 30118 -21365 8 VDD
port 41 nsew
rlabel locali s 29438 -21375 29536 -21372 8 VDD
port 41 nsew
rlabel locali s 30001 -21365 30406 -21301 8 VDD
port 41 nsew
rlabel locali s 26922 -21413 29033 -21371 8 VDD
port 41 nsew
rlabel locali s 24709 -22712 24798 -21371 8 VDD
port 41 nsew
rlabel locali s 24016 -22712 24511 -22709 8 VDD
port 41 nsew
rlabel locali s 21003 -22714 22769 -22710 8 VDD
port 41 nsew
rlabel locali s 21316 -22710 22769 -22709 8 VDD
port 41 nsew
rlabel locali s 18691 -22714 20069 -22709 8 VDD
port 41 nsew
rlabel locali s 24417 -22709 24451 -22418 8 VDD
port 41 nsew
rlabel locali s 24221 -22709 24255 -22418 8 VDD
port 41 nsew
rlabel locali s 24025 -22709 24059 -22418 8 VDD
port 41 nsew
rlabel locali s 22674 -22709 22708 -22418 8 VDD
port 41 nsew
rlabel locali s 22478 -22709 22512 -22418 8 VDD
port 41 nsew
rlabel locali s 22282 -22709 22316 -22418 8 VDD
port 41 nsew
rlabel locali s 21717 -22709 21751 -22418 8 VDD
port 41 nsew
rlabel locali s 21521 -22709 21555 -22418 8 VDD
port 41 nsew
rlabel locali s 21325 -22709 21359 -22418 8 VDD
port 41 nsew
rlabel locali s 19974 -22709 20008 -22418 8 VDD
port 41 nsew
rlabel locali s 19778 -22709 19812 -22418 8 VDD
port 41 nsew
rlabel locali s 19582 -22709 19616 -22418 8 VDD
port 41 nsew
rlabel locali s 19092 -22709 19126 -22418 8 VDD
port 41 nsew
rlabel locali s 18896 -22709 18930 -22418 8 VDD
port 41 nsew
rlabel locali s 18700 -22709 18734 -22418 8 VDD
port 41 nsew
rlabel locali s 17370 -22743 18238 -22610 8 VDD
port 41 nsew
rlabel locali s 17566 -22610 17619 -22482 8 VDD
port 41 nsew
rlabel locali s 17370 -22610 17423 -22498 8 VDD
port 41 nsew
rlabel locali s -3007 -23436 -2738 -22508 2 VDD
port 41 nsew
rlabel locali s -4038 -23436 -3769 -22508 2 VDD
port 41 nsew
rlabel locali s -4941 -23436 -4672 -22508 2 VDD
port 41 nsew
rlabel locali s -5803 -23436 -5534 -22508 2 VDD
port 41 nsew
rlabel locali s -6680 -23436 -6411 -22508 2 VDD
port 41 nsew
rlabel locali s -7226 -23436 -6957 -22508 2 VDD
port 41 nsew
rlabel locali s -7514 -23436 -7424 -23347 2 VDD
port 41 nsew
rlabel locali s -8131 -23945 -8097 -23355 2 VDD
port 41 nsew
rlabel locali s -7514 -23347 -7425 -23232 2 VDD
port 41 nsew
rlabel locali s -8137 -23355 -8092 -23232 2 VDD
port 41 nsew
rlabel locali s -8327 -23945 -8293 -23352 2 VDD
port 41 nsew
rlabel locali s -8750 -23945 -8716 -23353 2 VDD
port 41 nsew
rlabel locali s -22935 -24029 -15298 -23862 2 VDD
port 41 nsew
rlabel locali s -8332 -23352 -8287 -23232 2 VDD
port 41 nsew
rlabel locali s -8754 -23353 -8709 -23232 2 VDD
port 41 nsew
rlabel locali s -11210 -23528 -11176 -23237 2 VDD
port 41 nsew
rlabel locali s -11406 -23528 -11372 -23237 2 VDD
port 41 nsew
rlabel locali s -11602 -23528 -11568 -23237 2 VDD
port 41 nsew
rlabel locali s -12047 -23528 -12013 -23237 2 VDD
port 41 nsew
rlabel locali s -12243 -23528 -12209 -23237 2 VDD
port 41 nsew
rlabel locali s -12439 -23528 -12405 -23237 2 VDD
port 41 nsew
rlabel locali s -13910 -23528 -13876 -23237 2 VDD
port 41 nsew
rlabel locali s -14106 -23528 -14072 -23237 2 VDD
port 41 nsew
rlabel locali s -14302 -23528 -14268 -23237 2 VDD
port 41 nsew
rlabel locali s -14747 -23528 -14713 -23237 2 VDD
port 41 nsew
rlabel locali s -14943 -23528 -14909 -23237 2 VDD
port 41 nsew
rlabel locali s -15139 -23528 -15105 -23237 2 VDD
port 41 nsew
rlabel locali s -15388 -23862 -15299 -23237 2 VDD
port 41 nsew
rlabel locali s -12917 -23237 -11115 -23232 2 VDD
port 41 nsew
rlabel locali s -15388 -23237 -13815 -23232 2 VDD
port 41 nsew
rlabel locali s -15388 -23232 -7425 -23169 2 VDD
port 41 nsew
rlabel locali s -11310 -23169 -7425 -23147 2 VDD
port 41 nsew
rlabel locali s -7514 -23147 -7425 -22508 2 VDD
port 41 nsew
rlabel locali s 17575 -22482 17609 -21898 8 VDD
port 41 nsew
rlabel locali s 17379 -22498 17413 -21898 8 VDD
port 41 nsew
rlabel locali s -7514 -22508 -2289 -22445 2 VDD
port 41 nsew
rlabel locali s -5043 -22445 -3241 -22440 2 VDD
port 41 nsew
rlabel locali s -7514 -22445 -5941 -22440 2 VDD
port 41 nsew
rlabel locali s -3336 -22440 -3302 -22149 2 VDD
port 41 nsew
rlabel locali s -3532 -22440 -3498 -22149 2 VDD
port 41 nsew
rlabel locali s -3728 -22440 -3694 -22149 2 VDD
port 41 nsew
rlabel locali s -4173 -22440 -4139 -22149 2 VDD
port 41 nsew
rlabel locali s -4369 -22440 -4335 -22149 2 VDD
port 41 nsew
rlabel locali s -4565 -22440 -4531 -22149 2 VDD
port 41 nsew
rlabel locali s -6036 -22440 -6002 -22149 2 VDD
port 41 nsew
rlabel locali s -6232 -22440 -6198 -22149 2 VDD
port 41 nsew
rlabel locali s -6428 -22440 -6394 -22149 2 VDD
port 41 nsew
rlabel locali s -6873 -22440 -6839 -22149 2 VDD
port 41 nsew
rlabel locali s -7069 -22440 -7035 -22149 2 VDD
port 41 nsew
rlabel locali s -7265 -22440 -7231 -22149 2 VDD
port 41 nsew
rlabel locali s 24709 -21371 29033 -21302 8 VDD
port 41 nsew
rlabel locali s 30001 -21301 31754 -21300 8 VDD
port 41 nsew
rlabel locali s 30001 -21300 32800 -21248 8 VDD
port 41 nsew
rlabel locali s 27920 -21302 28538 -21285 8 VDD
port 41 nsew
rlabel locali s 27920 -21285 28363 -21256 8 VDD
port 41 nsew
rlabel locali s 30368 -21248 32800 -21178 8 VDD
port 41 nsew
rlabel locali s 27921 -21256 28363 -21242 8 VDD
port 41 nsew
rlabel locali s 27921 -21242 29210 -21193 8 VDD
port 41 nsew
rlabel locali s 28323 -21193 29210 -21143 8 VDD
port 41 nsew
rlabel locali s 35350 -21123 36068 -21024 8 VDD
port 41 nsew
rlabel locali s 35986 -21024 36020 -20758 8 VDD
port 41 nsew
rlabel locali s 35790 -21024 35824 -20758 8 VDD
port 41 nsew
rlabel locali s 35594 -21024 35628 -20758 8 VDD
port 41 nsew
rlabel locali s 35398 -21024 35432 -20758 8 VDD
port 41 nsew
rlabel locali s 29128 -21143 29162 -20977 8 VDD
port 41 nsew
rlabel locali s 28932 -21143 28966 -20977 8 VDD
port 41 nsew
rlabel locali s 28736 -21143 28770 -20977 8 VDD
port 41 nsew
rlabel locali s 28540 -21143 28574 -20977 8 VDD
port 41 nsew
rlabel locali s 28323 -21143 28357 -20776 8 VDD
port 41 nsew
rlabel locali s 28127 -21193 28161 -20776 8 VDD
port 41 nsew
rlabel locali s 27931 -21193 27965 -20776 8 VDD
port 41 nsew
rlabel locali s 24709 -21302 27264 -21112 8 VDD
port 41 nsew
rlabel locali s 24709 -21112 27628 -21077 8 VDD
port 41 nsew
rlabel locali s 26910 -21077 27628 -21013 8 VDD
port 41 nsew
rlabel locali s 24709 -21077 24798 -21017 8 VDD
port 41 nsew
rlabel locali s 24515 -21308 24549 -21017 8 VDD
port 41 nsew
rlabel locali s 24319 -21308 24353 -21017 8 VDD
port 41 nsew
rlabel locali s 24123 -21308 24157 -21017 8 VDD
port 41 nsew
rlabel locali s 23678 -21308 23712 -21017 8 VDD
port 41 nsew
rlabel locali s 23482 -21308 23516 -21017 8 VDD
port 41 nsew
rlabel locali s 23286 -21308 23320 -21017 8 VDD
port 41 nsew
rlabel locali s 21815 -21308 21849 -21017 8 VDD
port 41 nsew
rlabel locali s 21619 -21308 21653 -21017 8 VDD
port 41 nsew
rlabel locali s 21423 -21308 21457 -21017 8 VDD
port 41 nsew
rlabel locali s 20978 -21308 21012 -21017 8 VDD
port 41 nsew
rlabel locali s 20782 -21308 20816 -21017 8 VDD
port 41 nsew
rlabel locali s 20586 -21308 20620 -21017 8 VDD
port 41 nsew
rlabel locali s 27546 -21013 27580 -20747 8 VDD
port 41 nsew
rlabel locali s 27350 -21013 27384 -20747 8 VDD
port 41 nsew
rlabel locali s 27154 -21013 27188 -20747 8 VDD
port 41 nsew
rlabel locali s 26958 -21013 26992 -20747 8 VDD
port 41 nsew
rlabel locali s 23225 -21017 24798 -21012 8 VDD
port 41 nsew
rlabel locali s 20525 -21017 22327 -21012 8 VDD
port 41 nsew
rlabel locali s 19573 -21012 24798 -20949 8 VDD
port 41 nsew
rlabel locali s 7352 -21058 7386 -20868 8 VDD
port 41 nsew
rlabel locali s 7156 -21058 7190 -20880 8 VDD
port 41 nsew
rlabel locali s 7347 -20868 7393 -20746 8 VDD
port 41 nsew
rlabel locali s 7150 -20880 7196 -20746 8 VDD
port 41 nsew
rlabel locali s 7043 -21058 7077 -20870 8 VDD
port 41 nsew
rlabel locali s 6847 -21058 6881 -20875 8 VDD
port 41 nsew
rlabel locali s 7037 -20870 7083 -20746 8 VDD
port 41 nsew
rlabel locali s 6841 -20875 6887 -20746 8 VDD
port 41 nsew
rlabel locali s 6733 -21058 6767 -20871 8 VDD
port 41 nsew
rlabel locali s 6537 -21058 6571 -20875 8 VDD
port 41 nsew
rlabel locali s 6341 -21058 6375 -20875 8 VDD
port 41 nsew
rlabel locali s 6728 -20871 6774 -20746 8 VDD
port 41 nsew
rlabel locali s 6530 -20875 6576 -20746 8 VDD
port 41 nsew
rlabel locali s 6341 -20875 6381 -20786 8 VDD
port 41 nsew
rlabel locali s 6340 -20786 6463 -20746 8 VDD
port 41 nsew
rlabel locali s 5180 -21047 5214 -20785 8 VDD
port 41 nsew
rlabel locali s 6340 -20746 7393 -20677 8 VDD
port 41 nsew
rlabel locali s 6340 -20677 6463 -20650 8 VDD
port 41 nsew
rlabel locali s 5124 -20785 5247 -20751 8 VDD
port 41 nsew
rlabel locali s 4984 -21047 5018 -20751 8 VDD
port 41 nsew
rlabel locali s 4788 -21047 4822 -20751 8 VDD
port 41 nsew
rlabel locali s 4592 -21047 4626 -20751 8 VDD
port 41 nsew
rlabel locali s 4050 -21047 4084 -20755 8 VDD
port 41 nsew
rlabel locali s 3854 -21047 3888 -20780 8 VDD
port 41 nsew
rlabel locali s 3427 -21172 3461 -20782 8 VDD
port 41 nsew
rlabel locali s 3768 -20780 3891 -20755 8 VDD
port 41 nsew
rlabel locali s 4592 -20751 5247 -20750 8 VDD
port 41 nsew
rlabel locali s 3768 -20755 4089 -20750 8 VDD
port 41 nsew
rlabel locali s 3768 -20750 5247 -20682 8 VDD
port 41 nsew
rlabel locali s 5124 -20682 5247 -20649 8 VDD
port 41 nsew
rlabel locali s 3768 -20682 4664 -20677 8 VDD
port 41 nsew
rlabel locali s 3768 -20677 3891 -20644 8 VDD
port 41 nsew
rlabel locali s 3367 -20782 3490 -20755 8 VDD
port 41 nsew
rlabel locali s 3231 -21172 3265 -20755 8 VDD
port 41 nsew
rlabel locali s 3035 -21172 3069 -20805 8 VDD
port 41 nsew
rlabel locali s 2818 -20971 2852 -20805 8 VDD
port 41 nsew
rlabel locali s 2622 -20971 2656 -20805 8 VDD
port 41 nsew
rlabel locali s 2426 -20971 2460 -20805 8 VDD
port 41 nsew
rlabel locali s 2230 -20971 2264 -20805 8 VDD
port 41 nsew
rlabel locali s 1822 -21170 1856 -20806 8 VDD
port 41 nsew
rlabel locali s 2139 -20805 3069 -20755 8 VDD
port 41 nsew
rlabel locali s 2139 -20755 3490 -20706 8 VDD
port 41 nsew
rlabel locali s 3029 -20706 3490 -20691 8 VDD
port 41 nsew
rlabel locali s 3367 -20691 3490 -20646 8 VDD
port 41 nsew
rlabel locali s 2139 -20706 2262 -20669 8 VDD
port 41 nsew
rlabel locali s 1750 -20806 1873 -20763 8 VDD
port 41 nsew
rlabel locali s 1626 -21170 1660 -20763 8 VDD
port 41 nsew
rlabel locali s 1430 -21170 1464 -20803 8 VDD
port 41 nsew
rlabel locali s 1213 -20969 1247 -20803 8 VDD
port 41 nsew
rlabel locali s 1017 -20969 1051 -20803 8 VDD
port 41 nsew
rlabel locali s 821 -20969 855 -20803 8 VDD
port 41 nsew
rlabel locali s 625 -20969 659 -20803 8 VDD
port 41 nsew
rlabel locali s 577 -20803 1464 -20763 8 VDD
port 41 nsew
rlabel locali s 218 -21056 252 -20763 8 VDD
port 41 nsew
rlabel locali s 22 -21056 56 -20763 8 VDD
port 41 nsew
rlabel locali s -174 -21056 -140 -20763 2 VDD
port 41 nsew
rlabel locali s -370 -21056 -336 -20763 2 VDD
port 41 nsew
rlabel locali s -912 -21056 -878 -20764 2 VDD
port 41 nsew
rlabel locali s -1108 -21056 -1074 -20793 2 VDD
port 41 nsew
rlabel locali s -1450 -21039 -1416 -20794 2 VDD
port 41 nsew
rlabel locali s -1228 -20793 -1074 -20764 2 VDD
port 41 nsew
rlabel locali s -1228 -20764 -873 -20763 2 VDD
port 41 nsew
rlabel locali s -1228 -20763 1873 -20684 8 VDD
port 41 nsew
rlabel locali s 1750 -20684 1873 -20670 8 VDD
port 41 nsew
rlabel locali s -293 -20684 -178 -19876 2 VDD
port 41 nsew
rlabel locali s -1228 -20684 -1105 -20657 2 VDD
port 41 nsew
rlabel locali s -1522 -20794 -1399 -20748 2 VDD
port 41 nsew
rlabel locali s -1646 -21039 -1612 -20748 2 VDD
port 41 nsew
rlabel locali s -1842 -21039 -1808 -20748 2 VDD
port 41 nsew
rlabel locali s -2332 -21039 -2298 -20748 2 VDD
port 41 nsew
rlabel locali s -2528 -21039 -2494 -20748 2 VDD
port 41 nsew
rlabel locali s -2724 -21039 -2690 -20748 2 VDD
port 41 nsew
rlabel locali s -4075 -21039 -4041 -20748 2 VDD
port 41 nsew
rlabel locali s -4271 -21039 -4237 -20748 2 VDD
port 41 nsew
rlabel locali s -4467 -21039 -4433 -20748 2 VDD
port 41 nsew
rlabel locali s -5032 -21039 -4998 -20748 2 VDD
port 41 nsew
rlabel locali s -5228 -21039 -5194 -20748 2 VDD
port 41 nsew
rlabel locali s -5424 -21039 -5390 -20748 2 VDD
port 41 nsew
rlabel locali s -6775 -21039 -6741 -20748 2 VDD
port 41 nsew
rlabel locali s -6971 -21039 -6937 -20748 2 VDD
port 41 nsew
rlabel locali s -7167 -21039 -7133 -20748 2 VDD
port 41 nsew
rlabel locali s -2785 -20748 -1399 -20743 2 VDD
port 41 nsew
rlabel locali s -5485 -20748 -4032 -20747 2 VDD
port 41 nsew
rlabel locali s -5485 -20747 -3719 -20743 2 VDD
port 41 nsew
rlabel locali s -7227 -20748 -6732 -20745 2 VDD
port 41 nsew
rlabel locali s -7514 -22440 -7425 -20745 2 VDD
port 41 nsew
rlabel locali s -11918 -22247 -11884 -22081 2 VDD
port 41 nsew
rlabel locali s -12114 -22247 -12080 -22081 2 VDD
port 41 nsew
rlabel locali s -12310 -22247 -12276 -22081 2 VDD
port 41 nsew
rlabel locali s -12506 -22247 -12472 -22081 2 VDD
port 41 nsew
rlabel locali s -12723 -22448 -12689 -22081 2 VDD
port 41 nsew
rlabel locali s -12723 -22081 -11836 -22031 2 VDD
port 41 nsew
rlabel locali s -12919 -22448 -12885 -22031 2 VDD
port 41 nsew
rlabel locali s -13115 -22448 -13081 -22031 2 VDD
port 41 nsew
rlabel locali s -13500 -22477 -13466 -22211 2 VDD
port 41 nsew
rlabel locali s -13696 -22477 -13662 -22211 2 VDD
port 41 nsew
rlabel locali s -13892 -22477 -13858 -22211 2 VDD
port 41 nsew
rlabel locali s -14088 -22477 -14054 -22211 2 VDD
port 41 nsew
rlabel locali s -14136 -22211 -13418 -22112 2 VDD
port 41 nsew
rlabel locali s -13125 -22031 -11836 -21982 2 VDD
port 41 nsew
rlabel locali s -13125 -21982 -12683 -21968 2 VDD
port 41 nsew
rlabel locali s -13126 -21968 -12683 -21939 2 VDD
port 41 nsew
rlabel locali s -13126 -21939 -12508 -21922 2 VDD
port 41 nsew
rlabel locali s -13954 -22112 -13782 -21922 2 VDD
port 41 nsew
rlabel locali s -14926 -23169 -14773 -21922 2 VDD
port 41 nsew
rlabel locali s -14926 -21922 -12013 -21811 2 VDD
port 41 nsew
rlabel locali s -14926 -21811 -11909 -21769 2 VDD
port 41 nsew
rlabel locali s -12678 -21769 -11909 -21745 2 VDD
port 41 nsew
rlabel locali s -13722 -21769 -13496 -21762 2 VDD
port 41 nsew
rlabel locali s -13685 -21762 -13496 -21755 2 VDD
port 41 nsew
rlabel locali s -12055 -21745 -12010 -21621 2 VDD
port 41 nsew
rlabel locali s -12477 -21745 -12432 -21622 2 VDD
port 41 nsew
rlabel locali s -12048 -21621 -12014 -21029 2 VDD
port 41 nsew
rlabel locali s -12471 -21622 -12437 -21029 2 VDD
port 41 nsew
rlabel locali s -12672 -21745 -12627 -21619 2 VDD
port 41 nsew
rlabel locali s -14124 -21721 -13682 -21706 2 VDD
port 41 nsew
rlabel locali s -14124 -21706 -12835 -21657 2 VDD
port 41 nsew
rlabel locali s -12667 -21619 -12633 -21029 2 VDD
port 41 nsew
rlabel locali s -13722 -21657 -12835 -21607 2 VDD
port 41 nsew
rlabel locali s -12917 -21607 -12883 -21441 2 VDD
port 41 nsew
rlabel locali s -13113 -21607 -13079 -21441 2 VDD
port 41 nsew
rlabel locali s -13309 -21607 -13275 -21441 2 VDD
port 41 nsew
rlabel locali s -13505 -21607 -13471 -21441 2 VDD
port 41 nsew
rlabel locali s -13722 -21607 -13688 -21240 2 VDD
port 41 nsew
rlabel locali s -13918 -21657 -13884 -21240 2 VDD
port 41 nsew
rlabel locali s -14114 -21657 -14080 -21240 2 VDD
port 41 nsew
rlabel locali s -7514 -20745 -6410 -20743 2 VDD
port 41 nsew
rlabel locali s -7514 -20743 -1399 -20680 2 VDD
port 41 nsew
rlabel locali s -1522 -20680 -1399 -20658 2 VDD
port 41 nsew
rlabel locali s -2777 -20680 -2662 -19984 2 VDD
port 41 nsew
rlabel locali s -4192 -20680 -3719 -20679 2 VDD
port 41 nsew
rlabel locali s -5343 -20680 -5228 -20128 2 VDD
port 41 nsew
rlabel locali s -7514 -20680 -6410 -20677 2 VDD
port 41 nsew
rlabel locali s -6636 -20677 -6548 -20287 2 VDD
port 41 nsew
rlabel locali s -6818 -20677 -6730 -20287 2 VDD
port 41 nsew
rlabel locali s -7001 -20677 -6913 -20287 2 VDD
port 41 nsew
rlabel locali s -7017 -20287 -6522 -20219 2 VDD
port 41 nsew
rlabel locali s -5348 -20128 -5225 -19992 2 VDD
port 41 nsew
rlabel locali s -298 -19876 8 -19814 2 VDD
port 41 nsew
rlabel locali s -2781 -19984 -2658 -19848 2 VDD
port 41 nsew
rlabel locali s -6616 -20219 -6582 -19928 2 VDD
port 41 nsew
rlabel locali s -6812 -20219 -6778 -19928 2 VDD
port 41 nsew
rlabel locali s -7008 -20219 -6974 -19928 2 VDD
port 41 nsew
rlabel locali s -14926 -21769 -14773 -20073 2 VDD
port 41 nsew
rlabel locali s -16907 -21271 -16873 -21105 2 VDD
port 41 nsew
rlabel locali s -17103 -21271 -17069 -21105 2 VDD
port 41 nsew
rlabel locali s -17299 -21271 -17265 -21105 2 VDD
port 41 nsew
rlabel locali s -17495 -21271 -17461 -21105 2 VDD
port 41 nsew
rlabel locali s -17712 -21472 -17678 -21105 2 VDD
port 41 nsew
rlabel locali s -17712 -21105 -16825 -21055 2 VDD
port 41 nsew
rlabel locali s -17908 -21472 -17874 -21055 2 VDD
port 41 nsew
rlabel locali s -18104 -21472 -18070 -21055 2 VDD
port 41 nsew
rlabel locali s -18489 -21501 -18455 -21235 2 VDD
port 41 nsew
rlabel locali s -18685 -21501 -18651 -21235 2 VDD
port 41 nsew
rlabel locali s -18881 -21501 -18847 -21235 2 VDD
port 41 nsew
rlabel locali s -19077 -21501 -19043 -21235 2 VDD
port 41 nsew
rlabel locali s -19125 -21235 -18407 -21136 2 VDD
port 41 nsew
rlabel locali s -18114 -21055 -16825 -21006 2 VDD
port 41 nsew
rlabel locali s -18114 -21006 -17672 -20992 2 VDD
port 41 nsew
rlabel locali s -18115 -20992 -17672 -20963 2 VDD
port 41 nsew
rlabel locali s -18115 -20963 -17497 -20946 2 VDD
port 41 nsew
rlabel locali s -18943 -21136 -18771 -20946 2 VDD
port 41 nsew
rlabel locali s -19582 -21324 -19548 -21065 2 VDD
port 41 nsew
rlabel locali s -19778 -21324 -19744 -21065 2 VDD
port 41 nsew
rlabel locali s -20320 -21324 -20286 -21065 2 VDD
port 41 nsew
rlabel locali s -20516 -21324 -20482 -21065 2 VDD
port 41 nsew
rlabel locali s -20712 -21324 -20678 -21065 2 VDD
port 41 nsew
rlabel locali s -20908 -21324 -20874 -21065 2 VDD
port 41 nsew
rlabel locali s -21484 -21318 -21450 -21152 2 VDD
port 41 nsew
rlabel locali s -21680 -21318 -21646 -21152 2 VDD
port 41 nsew
rlabel locali s -21876 -21318 -21842 -21152 2 VDD
port 41 nsew
rlabel locali s -22072 -21318 -22038 -21152 2 VDD
port 41 nsew
rlabel locali s -22289 -21519 -22255 -21152 2 VDD
port 41 nsew
rlabel locali s -22289 -21152 -21402 -21102 2 VDD
port 41 nsew
rlabel locali s -22485 -21519 -22451 -21102 2 VDD
port 41 nsew
rlabel locali s -22681 -21519 -22647 -21102 2 VDD
port 41 nsew
rlabel locali s -22691 -21102 -21402 -21065 2 VDD
port 41 nsew
rlabel locali s -24351 -21065 -19548 -21032 2 VDD
port 41 nsew
rlabel locali s -24351 -21032 -19538 -20946 2 VDD
port 41 nsew
rlabel locali s -24351 -20946 -17002 -20835 2 VDD
port 41 nsew
rlabel locali s -24351 -20835 -16898 -20833 2 VDD
port 41 nsew
rlabel locali s -19113 -20833 -16898 -20793 2 VDD
port 41 nsew
rlabel locali s -17667 -20793 -16898 -20769 2 VDD
port 41 nsew
rlabel locali s -18711 -20793 -18485 -20786 2 VDD
port 41 nsew
rlabel locali s -18674 -20786 -18485 -20779 2 VDD
port 41 nsew
rlabel locali s -17044 -20769 -16999 -20645 2 VDD
port 41 nsew
rlabel locali s -17466 -20769 -17421 -20646 2 VDD
port 41 nsew
rlabel locali s -12066 -20071 -11593 -20070 2 VDD
port 41 nsew
rlabel locali s -15388 -20073 -14284 -20070 2 VDD
port 41 nsew
rlabel locali s -15388 -20070 -9281 -20007 2 VDD
port 41 nsew
rlabel locali s -17037 -20645 -17003 -20053 2 VDD
port 41 nsew
rlabel locali s -17460 -20646 -17426 -20053 2 VDD
port 41 nsew
rlabel locali s -17661 -20769 -17616 -20643 2 VDD
port 41 nsew
rlabel locali s -19113 -20745 -18671 -20730 2 VDD
port 41 nsew
rlabel locali s -19113 -20730 -17824 -20681 2 VDD
port 41 nsew
rlabel locali s -17656 -20643 -17622 -20053 2 VDD
port 41 nsew
rlabel locali s -18711 -20681 -17824 -20631 2 VDD
port 41 nsew
rlabel locali s -17906 -20631 -17872 -20465 2 VDD
port 41 nsew
rlabel locali s -18102 -20631 -18068 -20465 2 VDD
port 41 nsew
rlabel locali s -18298 -20631 -18264 -20465 2 VDD
port 41 nsew
rlabel locali s -18494 -20631 -18460 -20465 2 VDD
port 41 nsew
rlabel locali s -18711 -20631 -18677 -20264 2 VDD
port 41 nsew
rlabel locali s -18907 -20681 -18873 -20264 2 VDD
port 41 nsew
rlabel locali s -19103 -20681 -19069 -20264 2 VDD
port 41 nsew
rlabel locali s -10659 -20007 -9281 -20002 2 VDD
port 41 nsew
rlabel locali s -13359 -20007 -11593 -20003 2 VDD
port 41 nsew
rlabel locali s -15388 -20007 -14284 -20005 2 VDD
port 41 nsew
rlabel locali s -13359 -20003 -11906 -20002 2 VDD
port 41 nsew
rlabel locali s -15101 -20005 -14606 -20002 2 VDD
port 41 nsew
rlabel locali s -298 -19814 -175 -19813 2 VDD
port 41 nsew
rlabel locali s -9324 -20002 -9290 -19711 2 VDD
port 41 nsew
rlabel locali s -9520 -20002 -9486 -19711 2 VDD
port 41 nsew
rlabel locali s -9716 -20002 -9682 -19711 2 VDD
port 41 nsew
rlabel locali s -10206 -20002 -10172 -19711 2 VDD
port 41 nsew
rlabel locali s -10402 -20002 -10368 -19711 2 VDD
port 41 nsew
rlabel locali s -10598 -20002 -10564 -19711 2 VDD
port 41 nsew
rlabel locali s -11949 -20002 -11915 -19711 2 VDD
port 41 nsew
rlabel locali s -12145 -20002 -12111 -19711 2 VDD
port 41 nsew
rlabel locali s -12341 -20002 -12307 -19711 2 VDD
port 41 nsew
rlabel locali s -12906 -20002 -12872 -19711 2 VDD
port 41 nsew
rlabel locali s -13102 -20002 -13068 -19711 2 VDD
port 41 nsew
rlabel locali s -13298 -20002 -13264 -19711 2 VDD
port 41 nsew
rlabel locali s -14649 -20002 -14615 -19711 2 VDD
port 41 nsew
rlabel locali s -14845 -20002 -14811 -19711 2 VDD
port 41 nsew
rlabel locali s -15041 -20002 -15007 -19711 2 VDD
port 41 nsew
rlabel locali s -297 -19396 -174 -19260 2 VDD
port 41 nsew
rlabel locali s -2780 -19396 -2657 -19260 2 VDD
port 41 nsew
rlabel locali s 7342 -18807 7376 -18617 8 VDD
port 41 nsew
rlabel locali s 7146 -18807 7180 -18629 8 VDD
port 41 nsew
rlabel locali s 25225 -18550 26328 -17161 8 VDD
port 41 nsew
rlabel locali s 7337 -18617 7383 -18495 8 VDD
port 41 nsew
rlabel locali s 7140 -18629 7186 -18495 8 VDD
port 41 nsew
rlabel locali s 7033 -18807 7067 -18619 8 VDD
port 41 nsew
rlabel locali s 6837 -18807 6871 -18624 8 VDD
port 41 nsew
rlabel locali s 7027 -18619 7073 -18495 8 VDD
port 41 nsew
rlabel locali s 6831 -18624 6877 -18495 8 VDD
port 41 nsew
rlabel locali s 6723 -18807 6757 -18620 8 VDD
port 41 nsew
rlabel locali s 6527 -18807 6561 -18624 8 VDD
port 41 nsew
rlabel locali s 6331 -18807 6365 -18624 8 VDD
port 41 nsew
rlabel locali s 6718 -18620 6764 -18495 8 VDD
port 41 nsew
rlabel locali s 6520 -18624 6566 -18495 8 VDD
port 41 nsew
rlabel locali s 6331 -18624 6371 -18495 8 VDD
port 41 nsew
rlabel locali s 4342 -18807 4376 -18617 8 VDD
port 41 nsew
rlabel locali s 4146 -18807 4180 -18629 8 VDD
port 41 nsew
rlabel locali s 6331 -18495 7383 -18388 8 VDD
port 41 nsew
rlabel locali s 4337 -18617 4383 -18495 8 VDD
port 41 nsew
rlabel locali s 4140 -18629 4186 -18495 8 VDD
port 41 nsew
rlabel locali s 4033 -18807 4067 -18619 8 VDD
port 41 nsew
rlabel locali s 3837 -18807 3871 -18624 8 VDD
port 41 nsew
rlabel locali s 4027 -18619 4073 -18495 8 VDD
port 41 nsew
rlabel locali s 3831 -18624 3877 -18495 8 VDD
port 41 nsew
rlabel locali s 3723 -18807 3757 -18620 8 VDD
port 41 nsew
rlabel locali s 3527 -18807 3561 -18624 8 VDD
port 41 nsew
rlabel locali s 3331 -18807 3365 -18624 8 VDD
port 41 nsew
rlabel locali s 3718 -18620 3764 -18495 8 VDD
port 41 nsew
rlabel locali s 3520 -18624 3566 -18495 8 VDD
port 41 nsew
rlabel locali s 3331 -18624 3371 -18495 8 VDD
port 41 nsew
rlabel locali s 1842 -18807 1876 -18617 8 VDD
port 41 nsew
rlabel locali s 1646 -18807 1680 -18629 8 VDD
port 41 nsew
rlabel locali s 3331 -18495 4383 -18426 8 VDD
port 41 nsew
rlabel locali s 1837 -18617 1883 -18495 8 VDD
port 41 nsew
rlabel locali s 1640 -18629 1686 -18495 8 VDD
port 41 nsew
rlabel locali s 1533 -18807 1567 -18619 8 VDD
port 41 nsew
rlabel locali s 1337 -18807 1371 -18624 8 VDD
port 41 nsew
rlabel locali s 1527 -18619 1573 -18495 8 VDD
port 41 nsew
rlabel locali s 1331 -18624 1377 -18495 8 VDD
port 41 nsew
rlabel locali s 1223 -18807 1257 -18620 8 VDD
port 41 nsew
rlabel locali s 1027 -18807 1061 -18624 8 VDD
port 41 nsew
rlabel locali s 831 -18807 865 -18624 8 VDD
port 41 nsew
rlabel locali s 1218 -18620 1264 -18495 8 VDD
port 41 nsew
rlabel locali s 1020 -18624 1066 -18495 8 VDD
port 41 nsew
rlabel locali s 831 -18624 871 -18495 8 VDD
port 41 nsew
rlabel locali s 831 -18495 1883 -18426 8 VDD
port 41 nsew
rlabel locali s 3608 -18426 4201 -18388 8 VDD
port 41 nsew
rlabel locali s 1195 -18426 1788 -18388 8 VDD
port 41 nsew
rlabel locali s -292 -19260 -177 -18388 2 VDD
port 41 nsew
rlabel locali s -658 -18807 -624 -18617 2 VDD
port 41 nsew
rlabel locali s -854 -18807 -820 -18629 2 VDD
port 41 nsew
rlabel locali s -663 -18617 -617 -18495 2 VDD
port 41 nsew
rlabel locali s -860 -18629 -814 -18495 2 VDD
port 41 nsew
rlabel locali s -967 -18807 -933 -18619 2 VDD
port 41 nsew
rlabel locali s -1163 -18807 -1129 -18624 2 VDD
port 41 nsew
rlabel locali s -973 -18619 -927 -18495 2 VDD
port 41 nsew
rlabel locali s -1169 -18624 -1123 -18495 2 VDD
port 41 nsew
rlabel locali s -1277 -18807 -1243 -18620 2 VDD
port 41 nsew
rlabel locali s -1473 -18807 -1439 -18624 2 VDD
port 41 nsew
rlabel locali s -1669 -18807 -1635 -18624 2 VDD
port 41 nsew
rlabel locali s -1282 -18620 -1236 -18495 2 VDD
port 41 nsew
rlabel locali s -1480 -18624 -1434 -18495 2 VDD
port 41 nsew
rlabel locali s -1669 -18624 -1629 -18495 2 VDD
port 41 nsew
rlabel locali s -1669 -18495 -617 -18426 2 VDD
port 41 nsew
rlabel locali s -1339 -18426 -746 -18388 2 VDD
port 41 nsew
rlabel locali s -2774 -19260 -2660 -18388 2 VDD
port 41 nsew
rlabel locali s -5347 -19361 -5224 -19225 2 VDD
port 41 nsew
rlabel locali s -3158 -18807 -3124 -18617 2 VDD
port 41 nsew
rlabel locali s -3354 -18807 -3320 -18629 2 VDD
port 41 nsew
rlabel locali s -3163 -18617 -3117 -18495 2 VDD
port 41 nsew
rlabel locali s -3360 -18629 -3314 -18495 2 VDD
port 41 nsew
rlabel locali s -3467 -18807 -3433 -18619 2 VDD
port 41 nsew
rlabel locali s -3663 -18807 -3629 -18624 2 VDD
port 41 nsew
rlabel locali s -3473 -18619 -3427 -18495 2 VDD
port 41 nsew
rlabel locali s -3669 -18624 -3623 -18495 2 VDD
port 41 nsew
rlabel locali s -3777 -18807 -3743 -18620 2 VDD
port 41 nsew
rlabel locali s -3973 -18807 -3939 -18624 2 VDD
port 41 nsew
rlabel locali s -4169 -18807 -4135 -18624 2 VDD
port 41 nsew
rlabel locali s -3782 -18620 -3736 -18495 2 VDD
port 41 nsew
rlabel locali s -3980 -18624 -3934 -18495 2 VDD
port 41 nsew
rlabel locali s -4169 -18624 -4129 -18495 2 VDD
port 41 nsew
rlabel locali s -4169 -18495 -3117 -18426 2 VDD
port 41 nsew
rlabel locali s -3855 -18426 -3262 -18388 2 VDD
port 41 nsew
rlabel locali s -5342 -19225 -5227 -18388 2 VDD
port 41 nsew
rlabel locali s -15388 -20005 -15299 -19082 2 VDD
port 41 nsew
rlabel locali s -19542 -19409 -19508 -19243 2 VDD
port 41 nsew
rlabel locali s -19738 -19409 -19704 -19243 2 VDD
port 41 nsew
rlabel locali s -19934 -19409 -19900 -19243 2 VDD
port 41 nsew
rlabel locali s -20130 -19409 -20096 -19243 2 VDD
port 41 nsew
rlabel locali s -20347 -19610 -20313 -19243 2 VDD
port 41 nsew
rlabel locali s -20347 -19243 -19460 -19199 2 VDD
port 41 nsew
rlabel locali s -20543 -19610 -20509 -19199 2 VDD
port 41 nsew
rlabel locali s -20739 -19610 -20705 -19199 2 VDD
port 41 nsew
rlabel locali s -20791 -19199 -19460 -19144 2 VDD
port 41 nsew
rlabel locali s -20791 -19144 -19464 -19082 2 VDD
port 41 nsew
rlabel locali s -21412 -19388 -21378 -19096 2 VDD
port 41 nsew
rlabel locali s -21608 -19388 -21574 -19096 2 VDD
port 41 nsew
rlabel locali s -21613 -19096 -21368 -19082 2 VDD
port 41 nsew
rlabel locali s -22150 -19388 -22116 -19092 2 VDD
port 41 nsew
rlabel locali s -22346 -19388 -22312 -19092 2 VDD
port 41 nsew
rlabel locali s -22542 -19388 -22508 -19092 2 VDD
port 41 nsew
rlabel locali s -22738 -19388 -22704 -19092 2 VDD
port 41 nsew
rlabel locali s -24351 -20833 -24079 -19092 2 VDD
port 41 nsew
rlabel locali s -24351 -19092 -22116 -19082 2 VDD
port 41 nsew
rlabel locali s -5658 -18807 -5624 -18617 2 VDD
port 41 nsew
rlabel locali s -5854 -18807 -5820 -18629 2 VDD
port 41 nsew
rlabel locali s -5663 -18617 -5617 -18495 2 VDD
port 41 nsew
rlabel locali s -5860 -18629 -5814 -18495 2 VDD
port 41 nsew
rlabel locali s -5967 -18807 -5933 -18619 2 VDD
port 41 nsew
rlabel locali s -6163 -18807 -6129 -18624 2 VDD
port 41 nsew
rlabel locali s -5973 -18619 -5927 -18495 2 VDD
port 41 nsew
rlabel locali s -6169 -18624 -6123 -18495 2 VDD
port 41 nsew
rlabel locali s -6277 -18807 -6243 -18620 2 VDD
port 41 nsew
rlabel locali s -6473 -18807 -6439 -18624 2 VDD
port 41 nsew
rlabel locali s -6669 -18807 -6635 -18624 2 VDD
port 41 nsew
rlabel locali s -6282 -18620 -6236 -18495 2 VDD
port 41 nsew
rlabel locali s -6480 -18624 -6434 -18495 2 VDD
port 41 nsew
rlabel locali s -6669 -18624 -6629 -18495 2 VDD
port 41 nsew
rlabel locali s -6669 -18495 -5617 -18388 2 VDD
port 41 nsew
rlabel locali s -8158 -19011 -8124 -18421 2 VDD
port 41 nsew
rlabel locali s -8034 -18388 7428 -18295 2 VDD
port 41 nsew
rlabel locali s -8164 -18421 -8119 -18295 2 VDD
port 41 nsew
rlabel locali s -8354 -19011 -8320 -18418 2 VDD
port 41 nsew
rlabel locali s -8777 -19011 -8743 -18419 2 VDD
port 41 nsew
rlabel locali s -24351 -19082 -15299 -18869 2 VDD
port 41 nsew
rlabel locali s -8359 -18418 -8314 -18295 2 VDD
port 41 nsew
rlabel locali s -8781 -18419 -8736 -18295 2 VDD
port 41 nsew
rlabel locali s -11210 -18601 -11176 -18310 2 VDD
port 41 nsew
rlabel locali s -11406 -18601 -11372 -18310 2 VDD
port 41 nsew
rlabel locali s -11602 -18601 -11568 -18310 2 VDD
port 41 nsew
rlabel locali s -12047 -18601 -12013 -18310 2 VDD
port 41 nsew
rlabel locali s -12243 -18601 -12209 -18310 2 VDD
port 41 nsew
rlabel locali s -12439 -18601 -12405 -18310 2 VDD
port 41 nsew
rlabel locali s -13910 -18601 -13876 -18310 2 VDD
port 41 nsew
rlabel locali s -14106 -18601 -14072 -18310 2 VDD
port 41 nsew
rlabel locali s -14302 -18601 -14268 -18310 2 VDD
port 41 nsew
rlabel locali s -14747 -18601 -14713 -18310 2 VDD
port 41 nsew
rlabel locali s -14943 -18601 -14909 -18310 2 VDD
port 41 nsew
rlabel locali s -15139 -18601 -15105 -18310 2 VDD
port 41 nsew
rlabel locali s -15388 -18869 -15299 -18310 2 VDD
port 41 nsew
rlabel locali s -12917 -18310 -11115 -18305 2 VDD
port 41 nsew
rlabel locali s -15388 -18310 -13815 -18305 2 VDD
port 41 nsew
rlabel locali s -15388 -18305 -10163 -18295 2 VDD
port 41 nsew
rlabel locali s -15388 -18295 7428 -18242 2 VDD
port 41 nsew
rlabel locali s -10363 -18242 7428 -18206 2 VDD
port 41 nsew
rlabel locali s -8032 -18206 7428 -18195 2 VDD
port 41 nsew
rlabel locali s 25225 -17161 86373 -17041 8 VDD
port 41 nsew
rlabel locali s 6197 -18195 6959 -17041 8 VDD
port 41 nsew
rlabel locali s 6197 -17041 86373 -16279 8 VDD
port 41 nsew
rlabel locali s -9810 -18206 -9410 -16765 2 VDD
port 41 nsew
rlabel locali s -11883 -18242 -11533 -16765 2 VDD
port 41 nsew
rlabel locali s -14106 -18242 -13756 -16765 2 VDD
port 41 nsew
rlabel locali s -14987 -16765 -7549 -16699 2 VDD
port 41 nsew
rlabel locali s -7809 -16699 -7750 -16627 2 VDD
port 41 nsew
rlabel locali s -8397 -16699 -8338 -16627 2 VDD
port 41 nsew
rlabel locali s -8668 -16699 -8609 -16627 2 VDD
port 41 nsew
rlabel locali s -8909 -16699 -8850 -16627 2 VDD
port 41 nsew
rlabel locali s -9141 -16699 -9082 -16627 2 VDD
port 41 nsew
rlabel locali s -9747 -16699 -9688 -16627 2 VDD
port 41 nsew
rlabel locali s -9976 -16699 -9917 -16627 2 VDD
port 41 nsew
rlabel locali s -10215 -16699 -10156 -16627 2 VDD
port 41 nsew
rlabel locali s -10450 -16699 -10391 -16627 2 VDD
port 41 nsew
rlabel locali s -10686 -16699 -10627 -16627 2 VDD
port 41 nsew
rlabel locali s -10917 -16699 -10858 -16627 2 VDD
port 41 nsew
rlabel locali s -11642 -16699 -11583 -16627 2 VDD
port 41 nsew
rlabel locali s -11876 -16699 -11817 -16627 2 VDD
port 41 nsew
rlabel locali s -12110 -16699 -12051 -16627 2 VDD
port 41 nsew
rlabel locali s -12347 -16699 -12288 -16627 2 VDD
port 41 nsew
rlabel locali s -12577 -16699 -12518 -16627 2 VDD
port 41 nsew
rlabel locali s -12817 -16699 -12758 -16627 2 VDD
port 41 nsew
rlabel locali s -13055 -16699 -12996 -16627 2 VDD
port 41 nsew
rlabel locali s -13291 -16699 -13232 -16627 2 VDD
port 41 nsew
rlabel locali s -13522 -16699 -13463 -16627 2 VDD
port 41 nsew
rlabel locali s -13999 -16699 -13940 -16627 2 VDD
port 41 nsew
rlabel locali s -15097 -16627 -7545 -16579 2 VDD
port 41 nsew
rlabel locali s 25225 -16279 86373 -16058 8 VDD
port 41 nsew
rlabel locali s -7579 -16579 -7545 -16132 2 VDD
port 41 nsew
rlabel locali s -7815 -16579 -7781 -16132 2 VDD
port 41 nsew
rlabel locali s -8051 -16579 -8017 -16132 2 VDD
port 41 nsew
rlabel locali s -8181 -16579 -8147 -16132 2 VDD
port 41 nsew
rlabel locali s -8417 -16579 -8383 -16132 2 VDD
port 41 nsew
rlabel locali s -8653 -16579 -8619 -16132 2 VDD
port 41 nsew
rlabel locali s -8889 -16579 -8855 -16132 2 VDD
port 41 nsew
rlabel locali s -9125 -16579 -9091 -16132 2 VDD
port 41 nsew
rlabel locali s -9255 -16579 -9221 -16132 2 VDD
port 41 nsew
rlabel locali s -9491 -16579 -9457 -16132 2 VDD
port 41 nsew
rlabel locali s -9727 -16579 -9693 -16132 2 VDD
port 41 nsew
rlabel locali s -9963 -16579 -9929 -16132 2 VDD
port 41 nsew
rlabel locali s -10199 -16579 -10165 -16132 2 VDD
port 41 nsew
rlabel locali s -10435 -16579 -10401 -16132 2 VDD
port 41 nsew
rlabel locali s -10671 -16579 -10637 -16132 2 VDD
port 41 nsew
rlabel locali s -10907 -16579 -10873 -16132 2 VDD
port 41 nsew
rlabel locali s -11143 -16579 -11109 -16132 2 VDD
port 41 nsew
rlabel locali s -11391 -16579 -11357 -16132 2 VDD
port 41 nsew
rlabel locali s -11627 -16579 -11593 -16132 2 VDD
port 41 nsew
rlabel locali s -11863 -16579 -11829 -16132 2 VDD
port 41 nsew
rlabel locali s -12099 -16579 -12065 -16132 2 VDD
port 41 nsew
rlabel locali s -12335 -16579 -12301 -16132 2 VDD
port 41 nsew
rlabel locali s -12571 -16579 -12537 -16132 2 VDD
port 41 nsew
rlabel locali s -12807 -16579 -12773 -16132 2 VDD
port 41 nsew
rlabel locali s -13043 -16579 -13009 -16132 2 VDD
port 41 nsew
rlabel locali s -13279 -16579 -13245 -16132 2 VDD
port 41 nsew
rlabel locali s -13515 -16579 -13481 -16132 2 VDD
port 41 nsew
rlabel locali s -13751 -16579 -13717 -16132 2 VDD
port 41 nsew
rlabel locali s -13987 -16579 -13953 -16132 2 VDD
port 41 nsew
rlabel locali s -14223 -16579 -14189 -16132 2 VDD
port 41 nsew
rlabel locali s -14459 -16579 -14425 -16132 2 VDD
port 41 nsew
rlabel locali s -14695 -16579 -14661 -16132 2 VDD
port 41 nsew
rlabel locali s -14931 -16579 -14897 -16132 2 VDD
port 41 nsew
rlabel locali s 81378 -16058 84526 -15816 8 VDD
port 41 nsew
rlabel locali s 81378 -15816 98798 -12668 8 VDD
port 41 nsew
rlabel locali s 95829 -12668 98798 -7667 8 VDD
port 41 nsew
rlabel locali s 95743 -7667 98798 -4698 8 VDD
port 41 nsew
rlabel locali s 95829 -4698 98798 1398 8 VDD
port 41 nsew
rlabel locali s 63602 -4326 64823 -4274 8 VDD
port 41 nsew
rlabel locali s 64771 -4274 64823 -2677 8 VDD
port 41 nsew
rlabel locali s 64166 -4274 64701 -4262 8 VDD
port 41 nsew
rlabel locali s 63602 -4274 63729 -4268 8 VDD
port 41 nsew
rlabel locali s 63234 -4268 63729 -4200 8 VDD
port 41 nsew
rlabel locali s 63635 -4200 63669 -3909 8 VDD
port 41 nsew
rlabel locali s 63439 -4200 63473 -3909 8 VDD
port 41 nsew
rlabel locali s 63243 -4200 63277 -3909 8 VDD
port 41 nsew
rlabel locali s 63635 -3042 63669 -2751 8 VDD
port 41 nsew
rlabel locali s 63439 -3042 63473 -2751 8 VDD
port 41 nsew
rlabel locali s 63243 -3042 63277 -2751 8 VDD
port 41 nsew
rlabel locali s 62785 -3042 62819 -2751 8 VDD
port 41 nsew
rlabel locali s 62589 -3042 62623 -2751 8 VDD
port 41 nsew
rlabel locali s 62393 -3042 62427 -2751 8 VDD
port 41 nsew
rlabel locali s 58045 -3328 58079 -2881 8 VDD
port 41 nsew
rlabel locali s 57809 -3328 57843 -2881 8 VDD
port 41 nsew
rlabel locali s 57573 -3328 57607 -2881 8 VDD
port 41 nsew
rlabel locali s 57337 -3328 57371 -2881 8 VDD
port 41 nsew
rlabel locali s 57101 -3328 57135 -2881 8 VDD
port 41 nsew
rlabel locali s 56865 -3328 56899 -2881 8 VDD
port 41 nsew
rlabel locali s 56629 -3328 56663 -2881 8 VDD
port 41 nsew
rlabel locali s 56393 -3328 56427 -2881 8 VDD
port 41 nsew
rlabel locali s 56157 -3328 56191 -2881 8 VDD
port 41 nsew
rlabel locali s 55921 -3328 55955 -2881 8 VDD
port 41 nsew
rlabel locali s 55685 -3328 55719 -2881 8 VDD
port 41 nsew
rlabel locali s 55449 -3328 55483 -2881 8 VDD
port 41 nsew
rlabel locali s 55213 -3328 55247 -2881 8 VDD
port 41 nsew
rlabel locali s 54977 -3328 55011 -2881 8 VDD
port 41 nsew
rlabel locali s 54741 -3328 54775 -2881 8 VDD
port 41 nsew
rlabel locali s 54505 -3328 54539 -2881 8 VDD
port 41 nsew
rlabel locali s 54257 -3328 54291 -2881 8 VDD
port 41 nsew
rlabel locali s 54021 -3328 54055 -2881 8 VDD
port 41 nsew
rlabel locali s 53785 -3328 53819 -2881 8 VDD
port 41 nsew
rlabel locali s 53549 -3328 53583 -2881 8 VDD
port 41 nsew
rlabel locali s 53313 -3328 53347 -2881 8 VDD
port 41 nsew
rlabel locali s 53077 -3328 53111 -2881 8 VDD
port 41 nsew
rlabel locali s 52841 -3328 52875 -2881 8 VDD
port 41 nsew
rlabel locali s 52605 -3328 52639 -2881 8 VDD
port 41 nsew
rlabel locali s 52369 -3328 52403 -2881 8 VDD
port 41 nsew
rlabel locali s 52239 -3328 52273 -2881 8 VDD
port 41 nsew
rlabel locali s 52003 -3328 52037 -2881 8 VDD
port 41 nsew
rlabel locali s 51767 -3328 51801 -2881 8 VDD
port 41 nsew
rlabel locali s 51531 -3328 51565 -2881 8 VDD
port 41 nsew
rlabel locali s 51295 -3328 51329 -2881 8 VDD
port 41 nsew
rlabel locali s 51165 -3328 51199 -2881 8 VDD
port 41 nsew
rlabel locali s 50929 -3328 50963 -2881 8 VDD
port 41 nsew
rlabel locali s 50693 -3328 50727 -2881 8 VDD
port 41 nsew
rlabel locali s 50693 -2881 58245 -2833 8 VDD
port 41 nsew
rlabel locali s 57088 -2833 57147 -2761 8 VDD
port 41 nsew
rlabel locali s 56611 -2833 56670 -2761 8 VDD
port 41 nsew
rlabel locali s 56380 -2833 56439 -2761 8 VDD
port 41 nsew
rlabel locali s 56144 -2833 56203 -2761 8 VDD
port 41 nsew
rlabel locali s 55906 -2833 55965 -2761 8 VDD
port 41 nsew
rlabel locali s 55666 -2833 55725 -2761 8 VDD
port 41 nsew
rlabel locali s 55436 -2833 55495 -2761 8 VDD
port 41 nsew
rlabel locali s 55199 -2833 55258 -2761 8 VDD
port 41 nsew
rlabel locali s 54965 -2833 55024 -2761 8 VDD
port 41 nsew
rlabel locali s 54731 -2833 54790 -2761 8 VDD
port 41 nsew
rlabel locali s 54006 -2833 54065 -2761 8 VDD
port 41 nsew
rlabel locali s 53775 -2833 53834 -2761 8 VDD
port 41 nsew
rlabel locali s 53539 -2833 53598 -2761 8 VDD
port 41 nsew
rlabel locali s 53304 -2833 53363 -2761 8 VDD
port 41 nsew
rlabel locali s 53065 -2833 53124 -2761 8 VDD
port 41 nsew
rlabel locali s 52836 -2833 52895 -2761 8 VDD
port 41 nsew
rlabel locali s 52230 -2833 52289 -2761 8 VDD
port 41 nsew
rlabel locali s 51998 -2833 52057 -2761 8 VDD
port 41 nsew
rlabel locali s 51757 -2833 51816 -2761 8 VDD
port 41 nsew
rlabel locali s 51486 -2833 51545 -2761 8 VDD
port 41 nsew
rlabel locali s 50898 -2833 50957 -2761 8 VDD
port 41 nsew
rlabel locali s 64166 -2689 64701 -2677 8 VDD
port 41 nsew
rlabel locali s 62384 -2751 63729 -2683 8 VDD
port 41 nsew
rlabel locali s 50697 -2761 58135 -2731 8 VDD
port 41 nsew
rlabel locali s 50697 -2731 58307 -2695 8 VDD
port 41 nsew
rlabel locali s 63602 -2683 63729 -2677 8 VDD
port 41 nsew
rlabel locali s 62867 -2683 63256 -2682 8 VDD
port 41 nsew
rlabel locali s 63602 -2677 64823 -2625 8 VDD
port 41 nsew
rlabel locali s 64082 -2625 64533 -1968 8 VDD
port 41 nsew
rlabel locali s 57856 -2695 58307 -1968 8 VDD
port 41 nsew
rlabel locali s 56669 -2695 57120 -1968 8 VDD
port 41 nsew
rlabel locali s 55332 -2695 55783 -1968 8 VDD
port 41 nsew
rlabel locali s 53892 -2695 54343 -1968 8 VDD
port 41 nsew
rlabel locali s 53892 -1968 64533 -1517 8 VDD
port 41 nsew
rlabel locali s 5739 -1965 6960 -1913 8 VDD
port 41 nsew
rlabel locali s 64082 -1517 64533 859 8 VDD
port 41 nsew
rlabel locali s 57856 -1517 58307 -1516 8 VDD
port 41 nsew
rlabel locali s 56669 -1517 57120 -1516 8 VDD
port 41 nsew
rlabel locali s 55332 -1517 55783 -1516 8 VDD
port 41 nsew
rlabel locali s 21175 -1460 22396 -1408 8 VDD
port 41 nsew
rlabel locali s 58045 -281 58079 166 8 VDD
port 41 nsew
rlabel locali s 57809 -281 57843 166 8 VDD
port 41 nsew
rlabel locali s 57573 -281 57607 166 8 VDD
port 41 nsew
rlabel locali s 57337 -281 57371 166 8 VDD
port 41 nsew
rlabel locali s 57101 -281 57135 166 8 VDD
port 41 nsew
rlabel locali s 56865 -281 56899 166 8 VDD
port 41 nsew
rlabel locali s 56629 -281 56663 166 8 VDD
port 41 nsew
rlabel locali s 56393 -281 56427 166 8 VDD
port 41 nsew
rlabel locali s 56157 -281 56191 166 8 VDD
port 41 nsew
rlabel locali s 55921 -281 55955 166 8 VDD
port 41 nsew
rlabel locali s 55685 -281 55719 166 8 VDD
port 41 nsew
rlabel locali s 55449 -281 55483 166 8 VDD
port 41 nsew
rlabel locali s 55213 -281 55247 166 8 VDD
port 41 nsew
rlabel locali s 54977 -281 55011 166 8 VDD
port 41 nsew
rlabel locali s 54741 -281 54775 166 8 VDD
port 41 nsew
rlabel locali s 54505 -281 54539 166 8 VDD
port 41 nsew
rlabel locali s 54257 -281 54291 166 8 VDD
port 41 nsew
rlabel locali s 54021 -281 54055 166 8 VDD
port 41 nsew
rlabel locali s 53785 -281 53819 166 8 VDD
port 41 nsew
rlabel locali s 53549 -281 53583 166 8 VDD
port 41 nsew
rlabel locali s 53313 -281 53347 166 8 VDD
port 41 nsew
rlabel locali s 53077 -281 53111 166 8 VDD
port 41 nsew
rlabel locali s 52841 -281 52875 166 8 VDD
port 41 nsew
rlabel locali s 52605 -281 52639 166 8 VDD
port 41 nsew
rlabel locali s 52369 -281 52403 166 8 VDD
port 41 nsew
rlabel locali s 52239 -281 52273 166 8 VDD
port 41 nsew
rlabel locali s 52003 -281 52037 166 8 VDD
port 41 nsew
rlabel locali s 51767 -281 51801 166 8 VDD
port 41 nsew
rlabel locali s 51531 -281 51565 166 8 VDD
port 41 nsew
rlabel locali s 51295 -281 51329 166 8 VDD
port 41 nsew
rlabel locali s 51165 -281 51199 166 8 VDD
port 41 nsew
rlabel locali s 50929 -281 50963 166 8 VDD
port 41 nsew
rlabel locali s 50693 -281 50727 166 8 VDD
port 41 nsew
rlabel locali s 32461 -152 32623 -140 8 VDD
port 41 nsew
rlabel locali s 26988 -166 27304 -149 8 VDD
port 41 nsew
rlabel locali s 32461 -140 32775 -72 8 VDD
port 41 nsew
rlabel locali s 27605 -149 27767 -133 8 VDD
port 41 nsew
rlabel locali s 32622 -72 32775 -66 8 VDD
port 41 nsew
rlabel locali s 27605 -133 27920 -69 8 VDD
port 41 nsew
rlabel locali s 26885 -149 27304 -69 8 VDD
port 41 nsew
rlabel locali s 27767 -69 27920 -59 8 VDD
port 41 nsew
rlabel locali s 26988 -69 27304 -38 8 VDD
port 41 nsew
rlabel locali s 50693 166 58245 214 6 VDD
port 41 nsew
rlabel locali s 22344 -1408 22396 189 8 VDD
port 41 nsew
rlabel locali s 21739 -1408 22274 -1396 8 VDD
port 41 nsew
rlabel locali s 21175 -1408 21302 -1402 8 VDD
port 41 nsew
rlabel locali s 20807 -1402 21302 -1334 8 VDD
port 41 nsew
rlabel locali s 21208 -1334 21242 -1043 8 VDD
port 41 nsew
rlabel locali s 21012 -1334 21046 -1043 8 VDD
port 41 nsew
rlabel locali s 20816 -1334 20850 -1043 8 VDD
port 41 nsew
rlabel locali s 14929 -903 14963 -456 8 VDD
port 41 nsew
rlabel locali s 14693 -903 14727 -456 8 VDD
port 41 nsew
rlabel locali s 14457 -903 14491 -456 8 VDD
port 41 nsew
rlabel locali s 14221 -903 14255 -456 8 VDD
port 41 nsew
rlabel locali s 13985 -903 14019 -456 8 VDD
port 41 nsew
rlabel locali s 13749 -903 13783 -456 8 VDD
port 41 nsew
rlabel locali s 13513 -903 13547 -456 8 VDD
port 41 nsew
rlabel locali s 13277 -903 13311 -456 8 VDD
port 41 nsew
rlabel locali s 13041 -903 13075 -456 8 VDD
port 41 nsew
rlabel locali s 12805 -903 12839 -456 8 VDD
port 41 nsew
rlabel locali s 12569 -903 12603 -456 8 VDD
port 41 nsew
rlabel locali s 12333 -903 12367 -456 8 VDD
port 41 nsew
rlabel locali s 12097 -903 12131 -456 8 VDD
port 41 nsew
rlabel locali s 11861 -903 11895 -456 8 VDD
port 41 nsew
rlabel locali s 11625 -903 11659 -456 8 VDD
port 41 nsew
rlabel locali s 11389 -903 11423 -456 8 VDD
port 41 nsew
rlabel locali s 11141 -903 11175 -456 8 VDD
port 41 nsew
rlabel locali s 10905 -903 10939 -456 8 VDD
port 41 nsew
rlabel locali s 10669 -903 10703 -456 8 VDD
port 41 nsew
rlabel locali s 10433 -903 10467 -456 8 VDD
port 41 nsew
rlabel locali s 10197 -903 10231 -456 8 VDD
port 41 nsew
rlabel locali s 9961 -903 9995 -456 8 VDD
port 41 nsew
rlabel locali s 9725 -903 9759 -456 8 VDD
port 41 nsew
rlabel locali s 9489 -903 9523 -456 8 VDD
port 41 nsew
rlabel locali s 9253 -903 9287 -456 8 VDD
port 41 nsew
rlabel locali s 9123 -903 9157 -456 8 VDD
port 41 nsew
rlabel locali s 8887 -903 8921 -456 8 VDD
port 41 nsew
rlabel locali s 8651 -903 8685 -456 8 VDD
port 41 nsew
rlabel locali s 8415 -903 8449 -456 8 VDD
port 41 nsew
rlabel locali s 8179 -903 8213 -456 8 VDD
port 41 nsew
rlabel locali s 8049 -903 8083 -456 8 VDD
port 41 nsew
rlabel locali s 7813 -903 7847 -456 8 VDD
port 41 nsew
rlabel locali s 7577 -903 7611 -456 8 VDD
port 41 nsew
rlabel locali s 7577 -456 15129 -408 8 VDD
port 41 nsew
rlabel locali s 13972 -408 14031 -336 8 VDD
port 41 nsew
rlabel locali s 13495 -408 13554 -336 8 VDD
port 41 nsew
rlabel locali s 13264 -408 13323 -336 8 VDD
port 41 nsew
rlabel locali s 13028 -408 13087 -336 8 VDD
port 41 nsew
rlabel locali s 12790 -408 12849 -336 8 VDD
port 41 nsew
rlabel locali s 12550 -408 12609 -336 8 VDD
port 41 nsew
rlabel locali s 12320 -408 12379 -336 8 VDD
port 41 nsew
rlabel locali s 12083 -408 12142 -336 8 VDD
port 41 nsew
rlabel locali s 11849 -408 11908 -336 8 VDD
port 41 nsew
rlabel locali s 11615 -408 11674 -336 8 VDD
port 41 nsew
rlabel locali s 10890 -408 10949 -336 8 VDD
port 41 nsew
rlabel locali s 10659 -408 10718 -336 8 VDD
port 41 nsew
rlabel locali s 10423 -408 10482 -336 8 VDD
port 41 nsew
rlabel locali s 10188 -408 10247 -336 8 VDD
port 41 nsew
rlabel locali s 9949 -408 10008 -336 8 VDD
port 41 nsew
rlabel locali s 9720 -408 9779 -336 8 VDD
port 41 nsew
rlabel locali s 9114 -408 9173 -336 8 VDD
port 41 nsew
rlabel locali s 8882 -408 8941 -336 8 VDD
port 41 nsew
rlabel locali s 8641 -408 8700 -336 8 VDD
port 41 nsew
rlabel locali s 8370 -408 8429 -336 8 VDD
port 41 nsew
rlabel locali s 7782 -408 7841 -336 8 VDD
port 41 nsew
rlabel locali s 7581 -336 15019 -270 8 VDD
port 41 nsew
rlabel locali s 6908 -1913 6960 -316 8 VDD
port 41 nsew
rlabel locali s 6303 -1913 6838 -1901 8 VDD
port 41 nsew
rlabel locali s 5739 -1913 5866 -1907 8 VDD
port 41 nsew
rlabel locali s 5371 -1907 5866 -1839 8 VDD
port 41 nsew
rlabel locali s 5772 -1839 5806 -1548 8 VDD
port 41 nsew
rlabel locali s 5576 -1839 5610 -1548 8 VDD
port 41 nsew
rlabel locali s 5380 -1839 5414 -1548 8 VDD
port 41 nsew
rlabel locali s -3843 -1823 -2622 -1771 2 VDD
port 41 nsew
rlabel locali s 5772 -681 5806 -390 8 VDD
port 41 nsew
rlabel locali s 5576 -681 5610 -390 8 VDD
port 41 nsew
rlabel locali s 5380 -681 5414 -390 8 VDD
port 41 nsew
rlabel locali s 4922 -681 4956 -390 8 VDD
port 41 nsew
rlabel locali s 4726 -681 4760 -390 8 VDD
port 41 nsew
rlabel locali s 4530 -681 4564 -390 8 VDD
port 41 nsew
rlabel locali s 6303 -328 6838 -316 8 VDD
port 41 nsew
rlabel locali s 4521 -390 5866 -322 8 VDD
port 41 nsew
rlabel locali s 5739 -322 5866 -316 8 VDD
port 41 nsew
rlabel locali s 5004 -322 5393 -321 8 VDD
port 41 nsew
rlabel locali s 15818 -209 16268 -176 8 VDD
port 41 nsew
rlabel locali s 13848 -270 14299 -176 8 VDD
port 41 nsew
rlabel locali s 12650 -270 13101 -176 8 VDD
port 41 nsew
rlabel locali s 11432 -270 11883 -176 8 VDD
port 41 nsew
rlabel locali s 9891 -270 10342 -176 8 VDD
port 41 nsew
rlabel locali s 8303 -270 8754 -176 8 VDD
port 41 nsew
rlabel locali s 5739 -316 6960 -264 8 VDD
port 41 nsew
rlabel locali s 5877 -264 6211 -176 8 VDD
port 41 nsew
rlabel locali s 21208 -176 21242 115 8 VDD
port 41 nsew
rlabel locali s 21012 -176 21046 115 8 VDD
port 41 nsew
rlabel locali s 20816 -176 20850 115 8 VDD
port 41 nsew
rlabel locali s 20358 -176 20392 115 8 VDD
port 41 nsew
rlabel locali s 20162 -176 20196 115 8 VDD
port 41 nsew
rlabel locali s 19966 -176 20000 115 8 VDD
port 41 nsew
rlabel locali s 21739 177 22274 189 6 VDD
port 41 nsew
rlabel locali s 19957 115 21302 183 6 VDD
port 41 nsew
rlabel locali s 21175 183 21302 189 6 VDD
port 41 nsew
rlabel locali s 20440 183 20829 184 6 VDD
port 41 nsew
rlabel locali s 57088 214 57147 286 6 VDD
port 41 nsew
rlabel locali s 56611 214 56670 286 6 VDD
port 41 nsew
rlabel locali s 56380 214 56439 286 6 VDD
port 41 nsew
rlabel locali s 56144 214 56203 286 6 VDD
port 41 nsew
rlabel locali s 55906 214 55965 286 6 VDD
port 41 nsew
rlabel locali s 55666 214 55725 286 6 VDD
port 41 nsew
rlabel locali s 55436 214 55495 286 6 VDD
port 41 nsew
rlabel locali s 55199 214 55258 286 6 VDD
port 41 nsew
rlabel locali s 54965 214 55024 286 6 VDD
port 41 nsew
rlabel locali s 54731 214 54790 286 6 VDD
port 41 nsew
rlabel locali s 54006 214 54065 286 6 VDD
port 41 nsew
rlabel locali s 53775 214 53834 286 6 VDD
port 41 nsew
rlabel locali s 53539 214 53598 286 6 VDD
port 41 nsew
rlabel locali s 53304 214 53363 286 6 VDD
port 41 nsew
rlabel locali s 53065 214 53124 286 6 VDD
port 41 nsew
rlabel locali s 52836 214 52895 286 6 VDD
port 41 nsew
rlabel locali s 52230 214 52289 286 6 VDD
port 41 nsew
rlabel locali s 51998 214 52057 286 6 VDD
port 41 nsew
rlabel locali s 51757 214 51816 286 6 VDD
port 41 nsew
rlabel locali s 51486 214 51545 286 6 VDD
port 41 nsew
rlabel locali s 50898 214 50957 286 6 VDD
port 41 nsew
rlabel locali s 21175 189 22396 241 6 VDD
port 41 nsew
rlabel locali s 50697 286 58135 352 6 VDD
port 41 nsew
rlabel locali s 57259 352 57897 859 6 VDD
port 41 nsew
rlabel locali s 56173 352 56811 859 6 VDD
port 41 nsew
rlabel locali s 54759 352 55397 859 6 VDD
port 41 nsew
rlabel locali s 53362 352 54000 859 6 VDD
port 41 nsew
rlabel locali s 53362 859 64533 1310 6 VDD
port 41 nsew
rlabel locali s 38050 502 38084 1060 6 VDD
port 41 nsew
rlabel locali s 37734 502 37768 1060 6 VDD
port 41 nsew
rlabel locali s 37418 502 37452 1060 6 VDD
port 41 nsew
rlabel locali s 37102 502 37136 1060 6 VDD
port 41 nsew
rlabel locali s 36786 502 36820 947 6 VDD
port 41 nsew
rlabel locali s 36329 459 36363 947 6 VDD
port 41 nsew
rlabel locali s 36329 947 36820 1011 6 VDD
port 41 nsew
rlabel locali s 36786 1011 36820 1060 6 VDD
port 41 nsew
rlabel locali s 36329 1011 36363 1017 6 VDD
port 41 nsew
rlabel locali s 36013 459 36047 1017 6 VDD
port 41 nsew
rlabel locali s 35697 459 35731 1017 6 VDD
port 41 nsew
rlabel locali s 35381 459 35415 1017 6 VDD
port 41 nsew
rlabel locali s 35065 459 35099 1017 6 VDD
port 41 nsew
rlabel locali s 31594 436 31628 994 6 VDD
port 41 nsew
rlabel locali s 31278 436 31312 994 6 VDD
port 41 nsew
rlabel locali s 30962 436 30996 994 6 VDD
port 41 nsew
rlabel locali s 30646 436 30680 994 6 VDD
port 41 nsew
rlabel locali s 30330 436 30364 994 6 VDD
port 41 nsew
rlabel locali s 36777 1060 38084 1242 6 VDD
port 41 nsew
rlabel locali s 36777 1242 40098 1262 6 VDD
port 41 nsew
rlabel locali s 36777 1262 45284 1265 6 VDD
port 41 nsew
rlabel locali s 35056 1017 36363 1124 6 VDD
port 41 nsew
rlabel locali s 30321 994 31628 1101 6 VDD
port 41 nsew
rlabel locali s 36329 1124 36363 1201 6 VDD
port 41 nsew
rlabel locali s 36013 1124 36047 1201 6 VDD
port 41 nsew
rlabel locali s 35697 1124 35731 1201 6 VDD
port 41 nsew
rlabel locali s 35381 1124 35415 1201 6 VDD
port 41 nsew
rlabel locali s 35065 1124 35099 1201 6 VDD
port 41 nsew
rlabel locali s 60670 1310 61121 1398 6 VDD
port 41 nsew
rlabel locali s 38049 1265 45284 1325 6 VDD
port 41 nsew
rlabel locali s 43711 1325 45284 1330 6 VDD
port 41 nsew
rlabel locali s 41011 1325 42813 1330 6 VDD
port 41 nsew
rlabel locali s 38049 1325 40098 1326 6 VDD
port 41 nsew
rlabel locali s 60670 1398 98798 4290 6 VDD
port 41 nsew
rlabel locali s 45570 1352 46065 1415 6 VDD
port 41 nsew
rlabel locali s 45195 1330 45284 1415 6 VDD
port 41 nsew
rlabel locali s 45195 1415 46065 1420 6 VDD
port 41 nsew
rlabel locali s 45971 1420 46005 1711 6 VDD
port 41 nsew
rlabel locali s 45775 1420 45809 1711 6 VDD
port 41 nsew
rlabel locali s 45195 1420 45613 1472 6 VDD
port 41 nsew
rlabel locali s 45579 1472 45613 1711 6 VDD
port 41 nsew
rlabel locali s 58248 2630 58282 3077 6 VDD
port 41 nsew
rlabel locali s 58012 2630 58046 3077 6 VDD
port 41 nsew
rlabel locali s 57776 2630 57810 3077 6 VDD
port 41 nsew
rlabel locali s 57540 2630 57574 3077 6 VDD
port 41 nsew
rlabel locali s 57304 2630 57338 3077 6 VDD
port 41 nsew
rlabel locali s 57068 2630 57102 3077 6 VDD
port 41 nsew
rlabel locali s 56832 2630 56866 3077 6 VDD
port 41 nsew
rlabel locali s 56596 2630 56630 3077 6 VDD
port 41 nsew
rlabel locali s 56360 2630 56394 3077 6 VDD
port 41 nsew
rlabel locali s 56124 2630 56158 3077 6 VDD
port 41 nsew
rlabel locali s 55888 2630 55922 3077 6 VDD
port 41 nsew
rlabel locali s 55652 2630 55686 3077 6 VDD
port 41 nsew
rlabel locali s 55416 2630 55450 3077 6 VDD
port 41 nsew
rlabel locali s 55180 2630 55214 3077 6 VDD
port 41 nsew
rlabel locali s 54944 2630 54978 3077 6 VDD
port 41 nsew
rlabel locali s 54708 2630 54742 3077 6 VDD
port 41 nsew
rlabel locali s 54460 2630 54494 3077 6 VDD
port 41 nsew
rlabel locali s 54224 2630 54258 3077 6 VDD
port 41 nsew
rlabel locali s 53988 2630 54022 3077 6 VDD
port 41 nsew
rlabel locali s 53752 2630 53786 3077 6 VDD
port 41 nsew
rlabel locali s 53516 2630 53550 3077 6 VDD
port 41 nsew
rlabel locali s 53280 2630 53314 3077 6 VDD
port 41 nsew
rlabel locali s 53044 2630 53078 3077 6 VDD
port 41 nsew
rlabel locali s 52808 2630 52842 3077 6 VDD
port 41 nsew
rlabel locali s 52572 2630 52606 3077 6 VDD
port 41 nsew
rlabel locali s 52442 2630 52476 3077 6 VDD
port 41 nsew
rlabel locali s 52206 2630 52240 3077 6 VDD
port 41 nsew
rlabel locali s 51970 2630 52004 3077 6 VDD
port 41 nsew
rlabel locali s 51734 2630 51768 3077 6 VDD
port 41 nsew
rlabel locali s 51498 2630 51532 3077 6 VDD
port 41 nsew
rlabel locali s 51368 2630 51402 3077 6 VDD
port 41 nsew
rlabel locali s 51132 2630 51166 3077 6 VDD
port 41 nsew
rlabel locali s 50896 2630 50930 3077 6 VDD
port 41 nsew
rlabel locali s 50896 3077 58448 3125 6 VDD
port 41 nsew
rlabel locali s 45195 1472 45284 3025 6 VDD
port 41 nsew
rlabel locali s 45001 1330 45035 1621 6 VDD
port 41 nsew
rlabel locali s 44805 1330 44839 1621 6 VDD
port 41 nsew
rlabel locali s 44609 1330 44643 1621 6 VDD
port 41 nsew
rlabel locali s 44164 1330 44198 1621 6 VDD
port 41 nsew
rlabel locali s 43968 1330 44002 1621 6 VDD
port 41 nsew
rlabel locali s 43772 1330 43806 1621 6 VDD
port 41 nsew
rlabel locali s 42301 1330 42335 1621 6 VDD
port 41 nsew
rlabel locali s 42105 1330 42139 1621 6 VDD
port 41 nsew
rlabel locali s 41909 1330 41943 1621 6 VDD
port 41 nsew
rlabel locali s 41464 1330 41498 1621 6 VDD
port 41 nsew
rlabel locali s 41268 1330 41302 1621 6 VDD
port 41 nsew
rlabel locali s 41072 1330 41106 1621 6 VDD
port 41 nsew
rlabel locali s 38050 1326 38084 1823 6 VDD
port 41 nsew
rlabel locali s 37734 1265 37768 1823 6 VDD
port 41 nsew
rlabel locali s 37418 1265 37452 1823 6 VDD
port 41 nsew
rlabel locali s 37102 1265 37136 1823 6 VDD
port 41 nsew
rlabel locali s 36786 1265 36820 1299 6 VDD
port 41 nsew
rlabel locali s 35056 1201 36363 1299 6 VDD
port 41 nsew
rlabel locali s 35056 1299 36820 1308 6 VDD
port 41 nsew
rlabel locali s 30321 1179 31628 1286 6 VDD
port 41 nsew
rlabel locali s 36329 1308 36820 1363 6 VDD
port 41 nsew
rlabel locali s 36786 1363 36820 1823 6 VDD
port 41 nsew
rlabel locali s 36329 1363 36363 1866 6 VDD
port 41 nsew
rlabel locali s 36013 1308 36047 1866 6 VDD
port 41 nsew
rlabel locali s 35697 1308 35731 1866 6 VDD
port 41 nsew
rlabel locali s 35381 1308 35415 1866 6 VDD
port 41 nsew
rlabel locali s 35065 1308 35099 1866 6 VDD
port 41 nsew
rlabel locali s 34330 1456 34364 1664 6 VDD
port 41 nsew
rlabel locali s 34172 1456 34206 1664 6 VDD
port 41 nsew
rlabel locali s 33884 1457 33918 1665 6 VDD
port 41 nsew
rlabel locali s 33438 1457 33472 1665 6 VDD
port 41 nsew
rlabel locali s 33122 1457 33156 1665 6 VDD
port 41 nsew
rlabel locali s 34326 1851 34360 2116 6 VDD
port 41 nsew
rlabel locali s 34168 1851 34202 2059 6 VDD
port 41 nsew
rlabel locali s 34214 2116 34360 2189 6 VDD
port 41 nsew
rlabel locali s 33884 1851 33918 2142 6 VDD
port 41 nsew
rlabel locali s 33438 1846 33472 2142 6 VDD
port 41 nsew
rlabel locali s 33122 1846 33156 2142 6 VDD
port 41 nsew
rlabel locali s 32734 1457 32768 2030 6 VDD
port 41 nsew
rlabel locali s 32576 1457 32610 2030 6 VDD
port 41 nsew
rlabel locali s 31594 1286 31628 1844 6 VDD
port 41 nsew
rlabel locali s 31278 1286 31312 1844 6 VDD
port 41 nsew
rlabel locali s 30962 1286 30996 1844 6 VDD
port 41 nsew
rlabel locali s 30646 1286 30680 1844 6 VDD
port 41 nsew
rlabel locali s 30330 1286 30364 1844 6 VDD
port 41 nsew
rlabel locali s 29475 1463 29509 1671 6 VDD
port 41 nsew
rlabel locali s 29317 1463 29351 1671 6 VDD
port 41 nsew
rlabel locali s 29029 1464 29063 1672 6 VDD
port 41 nsew
rlabel locali s 28583 1464 28617 1672 6 VDD
port 41 nsew
rlabel locali s 28267 1464 28301 1672 6 VDD
port 41 nsew
rlabel locali s 32576 2030 32769 2099 6 VDD
port 41 nsew
rlabel locali s 33122 2142 33918 2176 6 VDD
port 41 nsew
rlabel locali s 34326 2189 34360 2268 6 VDD
port 41 nsew
rlabel locali s 33587 2176 33628 2255 6 VDD
port 41 nsew
rlabel locali s 33191 2176 33232 2255 6 VDD
port 41 nsew
rlabel locali s 32987 2255 33988 2268 6 VDD
port 41 nsew
rlabel locali s 32987 2268 34360 2273 6 VDD
port 41 nsew
rlabel locali s 32576 2099 32610 2273 6 VDD
port 41 nsew
rlabel locali s 32576 2273 34360 2302 6 VDD
port 41 nsew
rlabel locali s 32576 2302 33988 2307 6 VDD
port 41 nsew
rlabel locali s 29471 1858 29505 2123 6 VDD
port 41 nsew
rlabel locali s 29313 1858 29347 2066 6 VDD
port 41 nsew
rlabel locali s 29359 2123 29505 2196 6 VDD
port 41 nsew
rlabel locali s 29029 1858 29063 2149 6 VDD
port 41 nsew
rlabel locali s 28583 1853 28617 2149 6 VDD
port 41 nsew
rlabel locali s 28267 1853 28301 2149 6 VDD
port 41 nsew
rlabel locali s 27879 1464 27913 2037 6 VDD
port 41 nsew
rlabel locali s 27721 1464 27755 2037 6 VDD
port 41 nsew
rlabel locali s 21915 241 22067 1890 6 VDD
port 41 nsew
rlabel locali s 21288 241 21541 1890 6 VDD
port 41 nsew
rlabel locali s 5857 -176 16268 275 6 VDD
port 41 nsew
rlabel locali s -2674 -1771 -2622 -174 2 VDD
port 41 nsew
rlabel locali s -3279 -1771 -2744 -1759 2 VDD
port 41 nsew
rlabel locali s -3843 -1771 -3716 -1765 2 VDD
port 41 nsew
rlabel locali s -4211 -1765 -3716 -1697 2 VDD
port 41 nsew
rlabel locali s -3810 -1697 -3776 -1406 2 VDD
port 41 nsew
rlabel locali s -4006 -1697 -3972 -1406 2 VDD
port 41 nsew
rlabel locali s -4202 -1697 -4168 -1406 2 VDD
port 41 nsew
rlabel locali s -3810 -539 -3776 -248 2 VDD
port 41 nsew
rlabel locali s -4006 -539 -3972 -248 2 VDD
port 41 nsew
rlabel locali s -4202 -539 -4168 -248 2 VDD
port 41 nsew
rlabel locali s -4660 -539 -4626 -248 2 VDD
port 41 nsew
rlabel locali s -4856 -539 -4822 -248 2 VDD
port 41 nsew
rlabel locali s -5052 -539 -5018 -248 2 VDD
port 41 nsew
rlabel locali s -3279 -186 -2744 -174 2 VDD
port 41 nsew
rlabel locali s -5061 -248 -3716 -180 2 VDD
port 41 nsew
rlabel locali s -3843 -180 -3716 -174 2 VDD
port 41 nsew
rlabel locali s -4578 -180 -4189 -179 2 VDD
port 41 nsew
rlabel locali s -3843 -174 -2622 -122 2 VDD
port 41 nsew
rlabel locali s -3192 -122 -2863 35 2 VDD
port 41 nsew
rlabel locali s 15818 275 16268 345 6 VDD
port 41 nsew
rlabel locali s -3192 35 -2075 364 4 VDD
port 41 nsew
rlabel locali s -2404 364 -2075 549 4 VDD
port 41 nsew
rlabel locali s -2404 549 -1154 601 4 VDD
port 41 nsew
rlabel locali s 5730 686 6208 725 6 VDD
port 41 nsew
rlabel locali s 5724 725 6945 777 6 VDD
port 41 nsew
rlabel locali s 27721 2037 27914 2106 6 VDD
port 41 nsew
rlabel locali s 28267 2149 29063 2183 6 VDD
port 41 nsew
rlabel locali s 29471 2196 29505 2275 6 VDD
port 41 nsew
rlabel locali s 28732 2183 28773 2262 6 VDD
port 41 nsew
rlabel locali s 28336 2183 28377 2262 6 VDD
port 41 nsew
rlabel locali s 28132 2262 29133 2275 6 VDD
port 41 nsew
rlabel locali s 28132 2275 29505 2280 6 VDD
port 41 nsew
rlabel locali s 27721 2106 27755 2280 6 VDD
port 41 nsew
rlabel locali s 32987 2307 33988 2320 6 VDD
port 41 nsew
rlabel locali s 27721 2280 29505 2309 6 VDD
port 41 nsew
rlabel locali s 27721 2309 29133 2314 6 VDD
port 41 nsew
rlabel locali s 21003 1890 22224 1942 6 VDD
port 41 nsew
rlabel locali s 28132 2314 29133 2327 6 VDD
port 41 nsew
rlabel locali s 27825 2314 28014 2669 6 VDD
port 41 nsew
rlabel locali s 26688 2653 26963 2669 6 VDD
port 41 nsew
rlabel locali s 44903 2731 44937 3022 6 VDD
port 41 nsew
rlabel locali s 44707 2731 44741 3022 6 VDD
port 41 nsew
rlabel locali s 44511 2731 44545 3022 6 VDD
port 41 nsew
rlabel locali s 43160 2731 43194 3022 6 VDD
port 41 nsew
rlabel locali s 42964 2731 42998 3022 6 VDD
port 41 nsew
rlabel locali s 42768 2731 42802 3022 6 VDD
port 41 nsew
rlabel locali s 42203 2731 42237 3022 6 VDD
port 41 nsew
rlabel locali s 42007 2731 42041 3022 6 VDD
port 41 nsew
rlabel locali s 41811 2731 41845 3022 6 VDD
port 41 nsew
rlabel locali s 40460 2731 40494 3022 6 VDD
port 41 nsew
rlabel locali s 40264 2731 40298 3022 6 VDD
port 41 nsew
rlabel locali s 40068 2731 40102 3022 6 VDD
port 41 nsew
rlabel locali s 39578 2731 39612 3022 6 VDD
port 41 nsew
rlabel locali s 39382 2731 39416 3022 6 VDD
port 41 nsew
rlabel locali s 39186 2731 39220 3022 6 VDD
port 41 nsew
rlabel locali s 26688 2669 28014 2858 6 VDD
port 41 nsew
rlabel locali s 26688 2858 26963 2876 6 VDD
port 41 nsew
rlabel locali s 44502 3022 44997 3025 6 VDD
port 41 nsew
rlabel locali s 41802 3022 43255 3023 6 VDD
port 41 nsew
rlabel locali s 44180 3025 45284 3027 6 VDD
port 41 nsew
rlabel locali s 41489 3023 43255 3027 6 VDD
port 41 nsew
rlabel locali s 39177 3022 40555 3027 6 VDD
port 41 nsew
rlabel locali s 39177 3027 45284 3090 6 VDD
port 41 nsew
rlabel locali s 41489 3090 45284 3091 6 VDD
port 41 nsew
rlabel locali s 41815 3091 45284 3093 6 VDD
port 41 nsew
rlabel locali s 57291 3125 57350 3197 6 VDD
port 41 nsew
rlabel locali s 56814 3125 56873 3197 6 VDD
port 41 nsew
rlabel locali s 56583 3125 56642 3197 6 VDD
port 41 nsew
rlabel locali s 56347 3125 56406 3197 6 VDD
port 41 nsew
rlabel locali s 56109 3125 56168 3197 6 VDD
port 41 nsew
rlabel locali s 55869 3125 55928 3197 6 VDD
port 41 nsew
rlabel locali s 55639 3125 55698 3197 6 VDD
port 41 nsew
rlabel locali s 55402 3125 55461 3197 6 VDD
port 41 nsew
rlabel locali s 55168 3125 55227 3197 6 VDD
port 41 nsew
rlabel locali s 54934 3125 54993 3197 6 VDD
port 41 nsew
rlabel locali s 54209 3125 54268 3197 6 VDD
port 41 nsew
rlabel locali s 53978 3125 54037 3197 6 VDD
port 41 nsew
rlabel locali s 53742 3125 53801 3197 6 VDD
port 41 nsew
rlabel locali s 53507 3125 53566 3197 6 VDD
port 41 nsew
rlabel locali s 53268 3125 53327 3197 6 VDD
port 41 nsew
rlabel locali s 53039 3125 53098 3197 6 VDD
port 41 nsew
rlabel locali s 52433 3125 52492 3197 6 VDD
port 41 nsew
rlabel locali s 52201 3125 52260 3197 6 VDD
port 41 nsew
rlabel locali s 51960 3125 52019 3197 6 VDD
port 41 nsew
rlabel locali s 51689 3125 51748 3197 6 VDD
port 41 nsew
rlabel locali s 51101 3125 51160 3197 6 VDD
port 41 nsew
rlabel locali s 50900 3197 58338 3263 6 VDD
port 41 nsew
rlabel locali s 41815 3093 44205 3238 6 VDD
port 41 nsew
rlabel locali s 57618 3263 58213 4290 6 VDD
port 41 nsew
rlabel locali s 55261 3263 55856 4290 6 VDD
port 41 nsew
rlabel locali s 53312 3263 53907 4290 6 VDD
port 41 nsew
rlabel locali s 51135 3263 51730 4290 6 VDD
port 41 nsew
rlabel locali s 22172 1942 22224 3539 6 VDD
port 41 nsew
rlabel locali s 21567 1942 22102 1954 6 VDD
port 41 nsew
rlabel locali s 21003 1942 21130 1948 6 VDD
port 41 nsew
rlabel locali s 20635 1948 21130 2016 6 VDD
port 41 nsew
rlabel locali s 21036 2016 21070 2307 6 VDD
port 41 nsew
rlabel locali s 20840 2016 20874 2307 6 VDD
port 41 nsew
rlabel locali s 20644 2016 20678 2307 6 VDD
port 41 nsew
rlabel locali s 14970 1853 15004 2300 6 VDD
port 41 nsew
rlabel locali s 14734 1853 14768 2300 6 VDD
port 41 nsew
rlabel locali s 14498 1853 14532 2300 6 VDD
port 41 nsew
rlabel locali s 14262 1853 14296 2300 6 VDD
port 41 nsew
rlabel locali s 14026 1853 14060 2300 6 VDD
port 41 nsew
rlabel locali s 13790 1853 13824 2300 6 VDD
port 41 nsew
rlabel locali s 13554 1853 13588 2300 6 VDD
port 41 nsew
rlabel locali s 13318 1853 13352 2300 6 VDD
port 41 nsew
rlabel locali s 13082 1853 13116 2300 6 VDD
port 41 nsew
rlabel locali s 12846 1853 12880 2300 6 VDD
port 41 nsew
rlabel locali s 12610 1853 12644 2300 6 VDD
port 41 nsew
rlabel locali s 12374 1853 12408 2300 6 VDD
port 41 nsew
rlabel locali s 12138 1853 12172 2300 6 VDD
port 41 nsew
rlabel locali s 11902 1853 11936 2300 6 VDD
port 41 nsew
rlabel locali s 11666 1853 11700 2300 6 VDD
port 41 nsew
rlabel locali s 11430 1853 11464 2300 6 VDD
port 41 nsew
rlabel locali s 11182 1853 11216 2300 6 VDD
port 41 nsew
rlabel locali s 10946 1853 10980 2300 6 VDD
port 41 nsew
rlabel locali s 10710 1853 10744 2300 6 VDD
port 41 nsew
rlabel locali s 10474 1853 10508 2300 6 VDD
port 41 nsew
rlabel locali s 10238 1853 10272 2300 6 VDD
port 41 nsew
rlabel locali s 10002 1853 10036 2300 6 VDD
port 41 nsew
rlabel locali s 9766 1853 9800 2300 6 VDD
port 41 nsew
rlabel locali s 9530 1853 9564 2300 6 VDD
port 41 nsew
rlabel locali s 9294 1853 9328 2300 6 VDD
port 41 nsew
rlabel locali s 9164 1853 9198 2300 6 VDD
port 41 nsew
rlabel locali s 8928 1853 8962 2300 6 VDD
port 41 nsew
rlabel locali s 8692 1853 8726 2300 6 VDD
port 41 nsew
rlabel locali s 8456 1853 8490 2300 6 VDD
port 41 nsew
rlabel locali s 8220 1853 8254 2300 6 VDD
port 41 nsew
rlabel locali s 8090 1853 8124 2300 6 VDD
port 41 nsew
rlabel locali s 7854 1853 7888 2300 6 VDD
port 41 nsew
rlabel locali s 7618 1853 7652 2300 6 VDD
port 41 nsew
rlabel locali s 7618 2300 15170 2348 6 VDD
port 41 nsew
rlabel locali s 14013 2348 14072 2420 6 VDD
port 41 nsew
rlabel locali s 13536 2348 13595 2420 6 VDD
port 41 nsew
rlabel locali s 13305 2348 13364 2420 6 VDD
port 41 nsew
rlabel locali s 13069 2348 13128 2420 6 VDD
port 41 nsew
rlabel locali s 12831 2348 12890 2420 6 VDD
port 41 nsew
rlabel locali s 12591 2348 12650 2420 6 VDD
port 41 nsew
rlabel locali s 12361 2348 12420 2420 6 VDD
port 41 nsew
rlabel locali s 12124 2348 12183 2420 6 VDD
port 41 nsew
rlabel locali s 11890 2348 11949 2420 6 VDD
port 41 nsew
rlabel locali s 11656 2348 11715 2420 6 VDD
port 41 nsew
rlabel locali s 10931 2348 10990 2420 6 VDD
port 41 nsew
rlabel locali s 10700 2348 10759 2420 6 VDD
port 41 nsew
rlabel locali s 10464 2348 10523 2420 6 VDD
port 41 nsew
rlabel locali s 10229 2348 10288 2420 6 VDD
port 41 nsew
rlabel locali s 9990 2348 10049 2420 6 VDD
port 41 nsew
rlabel locali s 9761 2348 9820 2420 6 VDD
port 41 nsew
rlabel locali s 9155 2348 9214 2420 6 VDD
port 41 nsew
rlabel locali s 8923 2348 8982 2420 6 VDD
port 41 nsew
rlabel locali s 8682 2348 8741 2420 6 VDD
port 41 nsew
rlabel locali s 8411 2348 8470 2420 6 VDD
port 41 nsew
rlabel locali s 7823 2348 7882 2420 6 VDD
port 41 nsew
rlabel locali s 6893 777 6945 2374 6 VDD
port 41 nsew
rlabel locali s 6288 777 6823 789 6 VDD
port 41 nsew
rlabel locali s 5724 777 5851 783 6 VDD
port 41 nsew
rlabel locali s 5356 783 5851 851 6 VDD
port 41 nsew
rlabel locali s 5757 851 5791 1142 6 VDD
port 41 nsew
rlabel locali s 5561 851 5595 1142 6 VDD
port 41 nsew
rlabel locali s 5365 851 5399 1142 6 VDD
port 41 nsew
rlabel locali s 2809 1037 2843 1271 6 VDD
port 41 nsew
rlabel locali s 2500 1037 2534 1271 6 VDD
port 41 nsew
rlabel locali s 3500 1279 3875 1319 6 VDD
port 41 nsew
rlabel locali s 2452 1271 2979 1286 6 VDD
port 41 nsew
rlabel locali s 1836 1039 1870 1286 6 VDD
port 41 nsew
rlabel locali s 1690 1039 1724 1286 6 VDD
port 41 nsew
rlabel locali s 1401 1039 1435 1286 6 VDD
port 41 nsew
rlabel locali s 1401 1286 2979 1319 6 VDD
port 41 nsew
rlabel locali s 1401 1319 3875 1323 6 VDD
port 41 nsew
rlabel locali s 1225 1039 1259 1323 6 VDD
port 41 nsew
rlabel locali s 1049 1039 1083 1286 6 VDD
port 41 nsew
rlabel locali s 713 1037 747 1271 6 VDD
port 41 nsew
rlabel locali s 577 1271 795 1286 6 VDD
port 41 nsew
rlabel locali s 577 1286 1083 1323 6 VDD
port 41 nsew
rlabel locali s 577 1323 3875 1539 6 VDD
port 41 nsew
rlabel locali s 1401 1539 3875 1574 6 VDD
port 41 nsew
rlabel locali s 3500 1574 3875 1654 6 VDD
port 41 nsew
rlabel locali s 1401 1574 2979 1576 6 VDD
port 41 nsew
rlabel locali s 2452 1576 2979 1591 6 VDD
port 41 nsew
rlabel locali s 2809 1591 2843 1825 6 VDD
port 41 nsew
rlabel locali s 2500 1591 2534 1825 6 VDD
port 41 nsew
rlabel locali s 1836 1576 1870 1823 6 VDD
port 41 nsew
rlabel locali s 1690 1576 1724 1823 6 VDD
port 41 nsew
rlabel locali s 1401 1576 1435 1823 6 VDD
port 41 nsew
rlabel locali s 1225 1539 1259 1823 6 VDD
port 41 nsew
rlabel locali s 577 1539 1083 1576 6 VDD
port 41 nsew
rlabel locali s 1049 1576 1083 1823 6 VDD
port 41 nsew
rlabel locali s 577 1576 795 1591 6 VDD
port 41 nsew
rlabel locali s 713 1591 747 1825 6 VDD
port 41 nsew
rlabel locali s 5757 2009 5791 2300 6 VDD
port 41 nsew
rlabel locali s 5561 2009 5595 2300 6 VDD
port 41 nsew
rlabel locali s 5365 2009 5399 2300 6 VDD
port 41 nsew
rlabel locali s 4907 2009 4941 2300 6 VDD
port 41 nsew
rlabel locali s 4711 2009 4745 2300 6 VDD
port 41 nsew
rlabel locali s 4515 2009 4549 2300 6 VDD
port 41 nsew
rlabel locali s -1206 601 -1154 2198 4 VDD
port 41 nsew
rlabel locali s -1811 601 -1276 613 4 VDD
port 41 nsew
rlabel locali s -2404 601 -2248 607 4 VDD
port 41 nsew
rlabel locali s -2743 607 -2248 675 4 VDD
port 41 nsew
rlabel locali s -2342 675 -2308 966 4 VDD
port 41 nsew
rlabel locali s -2538 675 -2504 966 4 VDD
port 41 nsew
rlabel locali s -2734 675 -2700 966 4 VDD
port 41 nsew
rlabel locali s -2342 1833 -2308 2124 4 VDD
port 41 nsew
rlabel locali s -2538 1833 -2504 2124 4 VDD
port 41 nsew
rlabel locali s -2734 1833 -2700 2124 4 VDD
port 41 nsew
rlabel locali s -3192 1833 -3158 2124 4 VDD
port 41 nsew
rlabel locali s -3388 1833 -3354 2124 4 VDD
port 41 nsew
rlabel locali s -3584 1833 -3550 2124 4 VDD
port 41 nsew
rlabel locali s -5939 1571 -5905 2018 4 VDD
port 41 nsew
rlabel locali s -6175 1571 -6141 2018 4 VDD
port 41 nsew
rlabel locali s -6411 1571 -6377 2018 4 VDD
port 41 nsew
rlabel locali s -6541 1571 -6507 2018 4 VDD
port 41 nsew
rlabel locali s -6777 1571 -6743 2018 4 VDD
port 41 nsew
rlabel locali s -7013 1571 -6979 2018 4 VDD
port 41 nsew
rlabel locali s -7249 1571 -7215 2018 4 VDD
port 41 nsew
rlabel locali s -7485 1571 -7451 2018 4 VDD
port 41 nsew
rlabel locali s -7615 1571 -7581 2018 4 VDD
port 41 nsew
rlabel locali s -7851 1571 -7817 2018 4 VDD
port 41 nsew
rlabel locali s -8087 1571 -8053 2018 4 VDD
port 41 nsew
rlabel locali s -8323 1571 -8289 2018 4 VDD
port 41 nsew
rlabel locali s -8559 1571 -8525 2018 4 VDD
port 41 nsew
rlabel locali s -8795 1571 -8761 2018 4 VDD
port 41 nsew
rlabel locali s -9031 1571 -8997 2018 4 VDD
port 41 nsew
rlabel locali s -9267 1571 -9233 2018 4 VDD
port 41 nsew
rlabel locali s -9503 1571 -9469 2018 4 VDD
port 41 nsew
rlabel locali s -9751 1571 -9717 2018 4 VDD
port 41 nsew
rlabel locali s -9987 1571 -9953 2018 4 VDD
port 41 nsew
rlabel locali s -10223 1571 -10189 2018 4 VDD
port 41 nsew
rlabel locali s -10459 1571 -10425 2018 4 VDD
port 41 nsew
rlabel locali s -10695 1571 -10661 2018 4 VDD
port 41 nsew
rlabel locali s -10931 1571 -10897 2018 4 VDD
port 41 nsew
rlabel locali s -11167 1571 -11133 2018 4 VDD
port 41 nsew
rlabel locali s -11403 1571 -11369 2018 4 VDD
port 41 nsew
rlabel locali s -11639 1571 -11605 2018 4 VDD
port 41 nsew
rlabel locali s -11875 1571 -11841 2018 4 VDD
port 41 nsew
rlabel locali s -12111 1571 -12077 2018 4 VDD
port 41 nsew
rlabel locali s -12347 1571 -12313 2018 4 VDD
port 41 nsew
rlabel locali s -12583 1571 -12549 2018 4 VDD
port 41 nsew
rlabel locali s -12819 1571 -12785 2018 4 VDD
port 41 nsew
rlabel locali s -13055 1571 -13021 2018 4 VDD
port 41 nsew
rlabel locali s -13291 1571 -13257 2018 4 VDD
port 41 nsew
rlabel locali s -13457 2018 -5905 2066 4 VDD
port 41 nsew
rlabel locali s -1811 2186 -1276 2198 4 VDD
port 41 nsew
rlabel locali s -3593 2124 -2248 2192 4 VDD
port 41 nsew
rlabel locali s -6169 2066 -6110 2138 4 VDD
port 41 nsew
rlabel locali s -6757 2066 -6698 2138 4 VDD
port 41 nsew
rlabel locali s -7028 2066 -6969 2138 4 VDD
port 41 nsew
rlabel locali s -7269 2066 -7210 2138 4 VDD
port 41 nsew
rlabel locali s -7501 2066 -7442 2138 4 VDD
port 41 nsew
rlabel locali s -8107 2066 -8048 2138 4 VDD
port 41 nsew
rlabel locali s -8336 2066 -8277 2138 4 VDD
port 41 nsew
rlabel locali s -8575 2066 -8516 2138 4 VDD
port 41 nsew
rlabel locali s -8810 2066 -8751 2138 4 VDD
port 41 nsew
rlabel locali s -9046 2066 -8987 2138 4 VDD
port 41 nsew
rlabel locali s -9277 2066 -9218 2138 4 VDD
port 41 nsew
rlabel locali s -10002 2066 -9943 2138 4 VDD
port 41 nsew
rlabel locali s -10236 2066 -10177 2138 4 VDD
port 41 nsew
rlabel locali s -10470 2066 -10411 2138 4 VDD
port 41 nsew
rlabel locali s -10707 2066 -10648 2138 4 VDD
port 41 nsew
rlabel locali s -10937 2066 -10878 2138 4 VDD
port 41 nsew
rlabel locali s -11177 2066 -11118 2138 4 VDD
port 41 nsew
rlabel locali s -11415 2066 -11356 2138 4 VDD
port 41 nsew
rlabel locali s -11651 2066 -11592 2138 4 VDD
port 41 nsew
rlabel locali s -11882 2066 -11823 2138 4 VDD
port 41 nsew
rlabel locali s -12359 2066 -12300 2138 4 VDD
port 41 nsew
rlabel locali s -2375 2192 -2248 2198 4 VDD
port 41 nsew
rlabel locali s -3110 2192 -2721 2193 4 VDD
port 41 nsew
rlabel locali s -2375 2198 -1154 2250 4 VDD
port 41 nsew
rlabel locali s -13347 2138 -5909 2204 4 VDD
port 41 nsew
rlabel locali s 6288 2362 6823 2374 6 VDD
port 41 nsew
rlabel locali s 4506 2300 5851 2368 6 VDD
port 41 nsew
rlabel locali s 5724 2368 5851 2374 6 VDD
port 41 nsew
rlabel locali s 4989 2368 5378 2369 6 VDD
port 41 nsew
rlabel locali s 7622 2420 15060 2486 6 VDD
port 41 nsew
rlabel locali s 5724 2374 6945 2426 6 VDD
port 41 nsew
rlabel locali s 21036 3174 21070 3465 6 VDD
port 41 nsew
rlabel locali s 20840 3174 20874 3465 6 VDD
port 41 nsew
rlabel locali s 20644 3174 20678 3465 6 VDD
port 41 nsew
rlabel locali s 20186 3174 20220 3465 6 VDD
port 41 nsew
rlabel locali s 19990 3174 20024 3465 6 VDD
port 41 nsew
rlabel locali s 19794 3174 19828 3465 6 VDD
port 41 nsew
rlabel locali s 11748 2486 12550 3241 6 VDD
port 41 nsew
rlabel locali s 6011 2426 6354 3241 6 VDD
port 41 nsew
rlabel locali s -2198 2250 -1747 3241 4 VDD
port 41 nsew
rlabel locali s -13326 2204 -9322 2305 4 VDD
port 41 nsew
rlabel locali s 21567 3527 22102 3539 6 VDD
port 41 nsew
rlabel locali s 19785 3465 21130 3533 6 VDD
port 41 nsew
rlabel locali s 21003 3533 21130 3539 6 VDD
port 41 nsew
rlabel locali s 20268 3533 20657 3534 6 VDD
port 41 nsew
rlabel locali s 21003 3539 22224 3591 6 VDD
port 41 nsew
rlabel locali s 21388 3591 21612 3717 6 VDD
port 41 nsew
rlabel locali s -13207 3241 15270 3692 6 VDD
port 41 nsew
rlabel locali s 14819 3692 15270 3717 6 VDD
port 41 nsew
rlabel locali s 14819 3717 24380 4168 6 VDD
port 41 nsew
rlabel locali s 23929 4168 24380 4290 6 VDD
port 41 nsew
rlabel locali s 15817 4168 16331 4171 6 VDD
port 41 nsew
rlabel locali s 23929 4290 98798 4367 6 VDD
port 41 nsew
rlabel locali s 23929 4367 61121 4741 6 VDD
port 41 nsew
rlabel locali s -12975 5372 -11404 5558 4 VDD
port 41 nsew
rlabel locali s 12622 6692 12656 7658 6 VDD
port 41 nsew
rlabel locali s 11576 6692 11740 7658 6 VDD
port 41 nsew
rlabel locali s 9860 6692 9894 7658 6 VDD
port 41 nsew
rlabel locali s 8144 6692 8178 7658 6 VDD
port 41 nsew
rlabel locali s -12975 5558 -2388 6803 4 VDD
port 41 nsew
rlabel locali s -12975 6803 -11404 6943 4 VDD
port 41 nsew
rlabel locali s 8144 7658 12714 7659 6 VDD
port 41 nsew
rlabel locali s 3375 7565 4103 7659 6 VDD
port 41 nsew
rlabel locali s 3375 7659 12714 7840 6 VDD
port 41 nsew
rlabel locali s 3375 7840 8854 7918 6 VDD
port 41 nsew
rlabel locali s 3375 7918 4103 8200 6 VDD
port 41 nsew
rlabel locali s 15722 8972 15890 9006 6 VDD
port 41 nsew
rlabel locali s 15833 9006 15867 9101 6 VDD
port 41 nsew
rlabel locali s 15584 9101 15867 9135 6 VDD
port 41 nsew
rlabel locali s 15833 9135 15867 9617 6 VDD
port 41 nsew
rlabel locali s 14469 9053 14662 9172 6 VDD
port 41 nsew
rlabel locali s 3428 8200 4063 9172 6 VDD
port 41 nsew
rlabel locali s 3428 9172 14662 9359 6 VDD
port 41 nsew
rlabel locali s 3428 9359 14989 9393 6 VDD
port 41 nsew
rlabel locali s 15584 9617 15867 9651 6 VDD
port 41 nsew
rlabel locali s 15833 9651 15867 10133 6 VDD
port 41 nsew
rlabel locali s 3428 9393 14662 9807 6 VDD
port 41 nsew
rlabel locali s -7534 8962 -5338 9234 4 VDD
port 41 nsew
rlabel locali s 14469 9807 14662 9875 6 VDD
port 41 nsew
rlabel locali s 14469 9875 14989 9909 6 VDD
port 41 nsew
rlabel locali s 15584 10133 15867 10167 6 VDD
port 41 nsew
rlabel locali s 15833 10167 15867 10257 6 VDD
port 41 nsew
rlabel locali s 14469 9909 14662 10215 6 VDD
port 41 nsew
rlabel locali s 14597 10215 14631 10257 6 VDD
port 41 nsew
rlabel locali s 14597 10257 15867 10291 6 VDD
port 41 nsew
rlabel locali s -5561 9234 -5338 10575 4 VDD
port 41 nsew
rlabel locali s -5857 10575 -5338 10609 4 VDD
port 41 nsew
rlabel locali s -5561 10609 -5338 10771 4 VDD
port 41 nsew
rlabel locali s -7534 9234 -7302 10622 4 VDD
port 41 nsew
rlabel locali s -14051 10350 -13984 10360 4 VDD
port 41 nsew
rlabel locali s -7571 10622 -7302 10632 4 VDD
port 41 nsew
rlabel locali s -7988 10632 -7302 10666 4 VDD
port 41 nsew
rlabel locali s -5857 10771 -5338 10805 4 VDD
port 41 nsew
rlabel locali s -5561 10805 -5338 10967 4 VDD
port 41 nsew
rlabel locali s -7571 10666 -7302 10828 4 VDD
port 41 nsew
rlabel locali s -10498 10378 -10331 10748 4 VDD
port 41 nsew
rlabel locali s -14051 10360 -13692 10394 4 VDD
port 41 nsew
rlabel locali s -14051 10394 -13984 10538 4 VDD
port 41 nsew
rlabel locali s -14060 10538 -13968 10556 4 VDD
port 41 nsew
rlabel locali s -14060 10556 -13692 10590 4 VDD
port 41 nsew
rlabel locali s -10882 10688 -10637 10697 4 VDD
port 41 nsew
rlabel locali s -11482 10697 -10637 10731 4 VDD
port 41 nsew
rlabel locali s -10882 10731 -10637 10741 4 VDD
port 41 nsew
rlabel locali s -10770 10741 -10637 10748 4 VDD
port 41 nsew
rlabel locali s -7988 10828 -7302 10862 4 VDD
port 41 nsew
rlabel locali s -5857 10967 -5338 11001 4 VDD
port 41 nsew
rlabel locali s -5561 11001 -5338 11163 4 VDD
port 41 nsew
rlabel locali s -7571 10862 -7302 11024 4 VDD
port 41 nsew
rlabel locali s -10770 10748 -10331 10884 4 VDD
port 41 nsew
rlabel locali s -10898 10884 -10331 10893 4 VDD
port 41 nsew
rlabel locali s -11482 10893 -10331 10927 4 VDD
port 41 nsew
rlabel locali s -10898 10927 -10331 10937 4 VDD
port 41 nsew
rlabel locali s -7988 11024 -7302 11058 4 VDD
port 41 nsew
rlabel locali s -5857 11163 -5338 11197 4 VDD
port 41 nsew
rlabel locali s -5551 11197 -5338 11700 4 VDD
port 41 nsew
rlabel locali s -7621 11058 -7302 11241 4 VDD
port 41 nsew
rlabel locali s -7787 11241 -7302 11275 4 VDD
port 41 nsew
rlabel locali s -7621 11275 -7302 11437 4 VDD
port 41 nsew
rlabel locali s -7787 11437 -7302 11471 4 VDD
port 41 nsew
rlabel locali s -7621 11471 -7302 11633 4 VDD
port 41 nsew
rlabel locali s -10770 10937 -10331 11530 4 VDD
port 41 nsew
rlabel locali s -14060 10590 -13968 11098 4 VDD
port 41 nsew
rlabel locali s -14060 11098 -13692 11132 4 VDD
port 41 nsew
rlabel locali s -14060 11132 -13968 11294 4 VDD
port 41 nsew
rlabel locali s -14060 11294 -13692 11328 4 VDD
port 41 nsew
rlabel locali s -14060 11328 -13968 11490 4 VDD
port 41 nsew
rlabel locali s -14060 11490 -13692 11524 4 VDD
port 41 nsew
rlabel locali s -7787 11633 -7302 11667 4 VDD
port 41 nsew
rlabel locali s -5565 11700 -5338 11705 4 VDD
port 41 nsew
rlabel locali s -5857 11705 -5338 11739 4 VDD
port 41 nsew
rlabel locali s -5565 11739 -5338 11901 4 VDD
port 41 nsew
rlabel locali s -7621 11667 -7302 11829 4 VDD
port 41 nsew
rlabel locali s -7787 11829 -7302 11863 4 VDD
port 41 nsew
rlabel locali s -5857 11901 -5338 11935 4 VDD
port 41 nsew
rlabel locali s -7621 11863 -7302 11911 4 VDD
port 41 nsew
rlabel locali s -10498 11530 -10331 11906 4 VDD
port 41 nsew
rlabel locali s -10770 11530 -10637 11556 4 VDD
port 41 nsew
rlabel locali s -14060 11524 -13968 11686 4 VDD
port 41 nsew
rlabel locali s -14060 11686 -13692 11720 4 VDD
port 41 nsew
rlabel locali s -10693 11891 -10624 11896 4 VDD
port 41 nsew
rlabel locali s -10820 11896 -10624 11903 4 VDD
port 41 nsew
rlabel locali s -11211 11903 -10624 11906 4 VDD
port 41 nsew
rlabel locali s -5565 11935 -5338 11945 4 VDD
port 41 nsew
rlabel locali s -5551 11945 -5338 12522 4 VDD
port 41 nsew
rlabel locali s -7534 11911 -7302 12405 4 VDD
port 41 nsew
rlabel locali s -11211 11906 -10331 11937 4 VDD
port 41 nsew
rlabel locali s -10820 11937 -10331 11944 4 VDD
port 41 nsew
rlabel locali s -10693 11944 -10331 12093 4 VDD
port 41 nsew
rlabel locali s -10826 12093 -10331 12099 4 VDD
port 41 nsew
rlabel locali s -11211 12099 -10331 12133 4 VDD
port 41 nsew
rlabel locali s -10826 12133 -10331 12141 4 VDD
port 41 nsew
rlabel locali s -7793 12405 -7302 12439 4 VDD
port 41 nsew
rlabel locali s -10693 12141 -10331 12424 4 VDD
port 41 nsew
rlabel locali s -5668 12522 -5338 12574 4 VDD
port 41 nsew
rlabel locali s -6079 12574 -5338 12608 4 VDD
port 41 nsew
rlabel locali s -7534 12439 -7302 12601 4 VDD
port 41 nsew
rlabel locali s -5668 12608 -5338 12770 4 VDD
port 41 nsew
rlabel locali s -7793 12601 -7302 12635 4 VDD
port 41 nsew
rlabel locali s -6079 12770 -5338 12804 4 VDD
port 41 nsew
rlabel locali s -7534 12635 -7302 12797 4 VDD
port 41 nsew
rlabel locali s -10498 12424 -10331 12795 4 VDD
port 41 nsew
rlabel locali s -10693 12424 -10624 12445 4 VDD
port 41 nsew
rlabel locali s -10666 12795 -10331 12796 4 VDD
port 41 nsew
rlabel locali s -5668 12804 -5338 12966 4 VDD
port 41 nsew
rlabel locali s -7793 12797 -7302 12831 4 VDD
port 41 nsew
rlabel locali s -10694 12796 -10331 12801 4 VDD
port 41 nsew
rlabel locali s -10821 12801 -10331 12808 4 VDD
port 41 nsew
rlabel locali s -6079 12966 -5338 13000 4 VDD
port 41 nsew
rlabel locali s -7534 12831 -7302 12993 4 VDD
port 41 nsew
rlabel locali s -11212 12808 -10331 12842 4 VDD
port 41 nsew
rlabel locali s -10821 12842 -10331 12849 4 VDD
port 41 nsew
rlabel locali s -5712 13000 -5338 13183 4 VDD
port 41 nsew
rlabel locali s -7793 12993 -7302 13027 4 VDD
port 41 nsew
rlabel locali s -10694 12849 -10331 12998 4 VDD
port 41 nsew
rlabel locali s -13516 12964 -13429 12966 4 VDD
port 41 nsew
rlabel locali s -10827 12998 -10331 13004 4 VDD
port 41 nsew
rlabel locali s -5878 13183 -5338 13217 4 VDD
port 41 nsew
rlabel locali s -5712 13217 -5338 13379 4 VDD
port 41 nsew
rlabel locali s -5878 13379 -5338 13413 4 VDD
port 41 nsew
rlabel locali s -5712 13413 -5338 13575 4 VDD
port 41 nsew
rlabel locali s -7534 13027 -7302 13535 4 VDD
port 41 nsew
rlabel locali s -11212 13004 -10331 13038 4 VDD
port 41 nsew
rlabel locali s -10827 13038 -10331 13046 4 VDD
port 41 nsew
rlabel locali s -10694 13046 -10331 13348 4 VDD
port 41 nsew
rlabel locali s -7793 13535 -7302 13569 4 VDD
port 41 nsew
rlabel locali s -5878 13575 -5338 13609 4 VDD
port 41 nsew
rlabel locali s -5712 13609 -5338 13771 4 VDD
port 41 nsew
rlabel locali s -7534 13569 -7302 13731 4 VDD
port 41 nsew
rlabel locali s -7793 13731 -7302 13765 4 VDD
port 41 nsew
rlabel locali s -5878 13771 -5338 13805 4 VDD
port 41 nsew
rlabel locali s -7501 13765 -7302 13775 4 VDD
port 41 nsew
rlabel locali s -5712 13805 -5338 13849 4 VDD
port 41 nsew
rlabel locali s -5551 13849 -5338 17925 4 VDD
port 41 nsew
rlabel locali s -5712 13849 -5613 13853 4 VDD
port 41 nsew
rlabel locali s -7415 13775 -7302 14200 4 VDD
port 41 nsew
rlabel locali s -7214 14200 -7150 14210 4 VDD
port 41 nsew
rlabel locali s -7214 14210 -6733 14244 4 VDD
port 41 nsew
rlabel locali s -7214 14244 -7150 14406 4 VDD
port 41 nsew
rlabel locali s -7214 14406 -6733 14440 4 VDD
port 41 nsew
rlabel locali s -7214 14440 -7150 14602 4 VDD
port 41 nsew
rlabel locali s -7415 14200 -7262 14370 4 VDD
port 41 nsew
rlabel locali s -7704 14188 -7605 14236 4 VDD
port 41 nsew
rlabel locali s -7970 14236 -7605 14270 4 VDD
port 41 nsew
rlabel locali s -7704 14270 -7605 14370 4 VDD
port 41 nsew
rlabel locali s -7704 14370 -7262 14432 4 VDD
port 41 nsew
rlabel locali s -7970 14432 -7262 14466 4 VDD
port 41 nsew
rlabel locali s -7704 14466 -7262 14542 4 VDD
port 41 nsew
rlabel locali s -7415 14542 -7262 14602 4 VDD
port 41 nsew
rlabel locali s -7214 14602 -6733 14636 4 VDD
port 41 nsew
rlabel locali s -7214 14636 -7100 14642 4 VDD
port 41 nsew
rlabel locali s -7415 14602 -7255 14639 4 VDD
port 41 nsew
rlabel locali s -7199 14642 -7100 14819 4 VDD
port 41 nsew
rlabel locali s -7199 14819 -6934 14853 4 VDD
port 41 nsew
rlabel locali s -7415 14639 -7248 14828 4 VDD
port 41 nsew
rlabel locali s -7199 14853 -7100 15015 4 VDD
port 41 nsew
rlabel locali s -7199 15015 -6934 15049 4 VDD
port 41 nsew
rlabel locali s -7199 15049 -7100 15211 4 VDD
port 41 nsew
rlabel locali s -7199 15211 -6934 15245 4 VDD
port 41 nsew
rlabel locali s -7199 15245 -7100 15407 4 VDD
port 41 nsew
rlabel locali s -7199 15407 -6934 15441 4 VDD
port 41 nsew
rlabel locali s -7199 15441 -7100 15489 4 VDD
port 41 nsew
rlabel locali s -7415 14828 -7262 15198 4 VDD
port 41 nsew
rlabel locali s -7704 14542 -7605 14628 4 VDD
port 41 nsew
rlabel locali s -7970 14628 -7605 14662 4 VDD
port 41 nsew
rlabel locali s -7704 14662 -7605 14824 4 VDD
port 41 nsew
rlabel locali s -7970 14824 -7605 14858 4 VDD
port 41 nsew
rlabel locali s -7704 14858 -7605 14906 4 VDD
port 41 nsew
rlabel locali s -7461 15198 -7262 15199 4 VDD
port 41 nsew
rlabel locali s -7524 15199 -7262 15209 4 VDD
port 41 nsew
rlabel locali s -7941 15209 -7262 15243 4 VDD
port 41 nsew
rlabel locali s -7524 15243 -7262 15405 4 VDD
port 41 nsew
rlabel locali s -7941 15405 -7262 15439 4 VDD
port 41 nsew
rlabel locali s -7524 15439 -7262 15601 4 VDD
port 41 nsew
rlabel locali s -7941 15601 -7262 15635 4 VDD
port 41 nsew
rlabel locali s -7574 15635 -7262 15641 4 VDD
port 41 nsew
rlabel locali s -7432 15641 -7262 15646 4 VDD
port 41 nsew
rlabel locali s -7432 15646 -7238 15652 4 VDD
port 41 nsew
rlabel locali s -7432 15652 -7112 15657 4 VDD
port 41 nsew
rlabel locali s -7432 15657 -6522 15691 4 VDD
port 41 nsew
rlabel locali s -7432 15691 -7112 15697 4 VDD
port 41 nsew
rlabel locali s -7432 15697 -7238 15816 4 VDD
port 41 nsew
rlabel locali s -7415 15816 -7238 15847 4 VDD
port 41 nsew
rlabel locali s -7415 15847 -7115 15853 4 VDD
port 41 nsew
rlabel locali s -7415 15853 -6522 15887 4 VDD
port 41 nsew
rlabel locali s -7415 15887 -7115 15892 4 VDD
port 41 nsew
rlabel locali s -7415 15892 -7238 16269 4 VDD
port 41 nsew
rlabel locali s -7415 16269 -7114 16276 4 VDD
port 41 nsew
rlabel locali s -7415 16276 -6522 16310 4 VDD
port 41 nsew
rlabel locali s -7415 16310 -7114 16311 4 VDD
port 41 nsew
rlabel locali s -7574 15641 -7475 15818 4 VDD
port 41 nsew
rlabel locali s -7740 15818 -7475 15852 4 VDD
port 41 nsew
rlabel locali s -7574 15852 -7475 16014 4 VDD
port 41 nsew
rlabel locali s -7740 16014 -7475 16048 4 VDD
port 41 nsew
rlabel locali s -7574 16048 -7475 16210 4 VDD
port 41 nsew
rlabel locali s -7740 16210 -7475 16244 4 VDD
port 41 nsew
rlabel locali s -7304 16311 -7114 16314 4 VDD
port 41 nsew
rlabel locali s -7304 16314 -7238 16415 4 VDD
port 41 nsew
rlabel locali s -7574 16244 -7475 16406 4 VDD
port 41 nsew
rlabel locali s -7740 16406 -7475 16440 4 VDD
port 41 nsew
rlabel locali s -7574 16440 -7475 16488 4 VDD
port 41 nsew
rlabel locali s -10498 13348 -10331 17925 4 VDD
port 41 nsew
rlabel locali s -10694 13348 -10625 13350 4 VDD
port 41 nsew
rlabel locali s -13516 12966 -12262 13138 4 VDD
port 41 nsew
rlabel locali s -12214 14200 -12150 14210 4 VDD
port 41 nsew
rlabel locali s -12214 14210 -11733 14244 4 VDD
port 41 nsew
rlabel locali s -12214 14244 -12150 14406 4 VDD
port 41 nsew
rlabel locali s -12214 14406 -11733 14440 4 VDD
port 41 nsew
rlabel locali s -12214 14440 -12150 14602 4 VDD
port 41 nsew
rlabel locali s -12434 13138 -12262 14370 4 VDD
port 41 nsew
rlabel locali s -13516 13138 -13429 13140 4 VDD
port 41 nsew
rlabel locali s -14060 11720 -13968 13140 4 VDD
port 41 nsew
rlabel locali s -12704 14188 -12605 14236 4 VDD
port 41 nsew
rlabel locali s -12970 14236 -12605 14270 4 VDD
port 41 nsew
rlabel locali s -12704 14270 -12605 14370 4 VDD
port 41 nsew
rlabel locali s -12704 14370 -12262 14432 4 VDD
port 41 nsew
rlabel locali s -12970 14432 -12262 14466 4 VDD
port 41 nsew
rlabel locali s -12704 14466 -12262 14542 4 VDD
port 41 nsew
rlabel locali s -12415 14542 -12262 14602 4 VDD
port 41 nsew
rlabel locali s -12214 14602 -11733 14636 4 VDD
port 41 nsew
rlabel locali s -12214 14636 -12100 14642 4 VDD
port 41 nsew
rlabel locali s -12415 14602 -12255 14639 4 VDD
port 41 nsew
rlabel locali s -12199 14642 -12100 14819 4 VDD
port 41 nsew
rlabel locali s -12199 14819 -11934 14853 4 VDD
port 41 nsew
rlabel locali s -12415 14639 -12248 14828 4 VDD
port 41 nsew
rlabel locali s -12199 14853 -12100 15015 4 VDD
port 41 nsew
rlabel locali s -12199 15015 -11934 15049 4 VDD
port 41 nsew
rlabel locali s -12199 15049 -12100 15211 4 VDD
port 41 nsew
rlabel locali s -12199 15211 -11934 15245 4 VDD
port 41 nsew
rlabel locali s -12199 15245 -12100 15407 4 VDD
port 41 nsew
rlabel locali s -12199 15407 -11934 15441 4 VDD
port 41 nsew
rlabel locali s -12199 15441 -12100 15489 4 VDD
port 41 nsew
rlabel locali s -12415 14828 -12262 15198 4 VDD
port 41 nsew
rlabel locali s -12704 14542 -12605 14628 4 VDD
port 41 nsew
rlabel locali s -12970 14628 -12605 14662 4 VDD
port 41 nsew
rlabel locali s -12704 14662 -12605 14824 4 VDD
port 41 nsew
rlabel locali s -12970 14824 -12605 14858 4 VDD
port 41 nsew
rlabel locali s -12704 14858 -12605 14906 4 VDD
port 41 nsew
rlabel locali s -12461 15198 -12262 15199 4 VDD
port 41 nsew
rlabel locali s -12524 15199 -12262 15209 4 VDD
port 41 nsew
rlabel locali s -12941 15209 -12262 15243 4 VDD
port 41 nsew
rlabel locali s -12524 15243 -12262 15405 4 VDD
port 41 nsew
rlabel locali s -12941 15405 -12262 15439 4 VDD
port 41 nsew
rlabel locali s -12524 15439 -12262 15601 4 VDD
port 41 nsew
rlabel locali s -12941 15601 -12262 15635 4 VDD
port 41 nsew
rlabel locali s -12574 15635 -12262 15641 4 VDD
port 41 nsew
rlabel locali s -12432 15641 -12262 15646 4 VDD
port 41 nsew
rlabel locali s -12432 15646 -12238 15652 4 VDD
port 41 nsew
rlabel locali s -12432 15652 -12112 15657 4 VDD
port 41 nsew
rlabel locali s -12432 15657 -11522 15691 4 VDD
port 41 nsew
rlabel locali s -12432 15691 -12112 15697 4 VDD
port 41 nsew
rlabel locali s -12432 15697 -12238 15816 4 VDD
port 41 nsew
rlabel locali s -12415 15816 -12238 15847 4 VDD
port 41 nsew
rlabel locali s -12415 15847 -12115 15853 4 VDD
port 41 nsew
rlabel locali s -12415 15853 -11522 15887 4 VDD
port 41 nsew
rlabel locali s -12415 15887 -12115 15892 4 VDD
port 41 nsew
rlabel locali s -12415 15892 -12238 16269 4 VDD
port 41 nsew
rlabel locali s -12415 16269 -12114 16276 4 VDD
port 41 nsew
rlabel locali s -12415 16276 -11522 16310 4 VDD
port 41 nsew
rlabel locali s -12415 16310 -12114 16311 4 VDD
port 41 nsew
rlabel locali s -12574 15641 -12475 15818 4 VDD
port 41 nsew
rlabel locali s -12740 15818 -12475 15852 4 VDD
port 41 nsew
rlabel locali s -12574 15852 -12475 16014 4 VDD
port 41 nsew
rlabel locali s -12740 16014 -12475 16048 4 VDD
port 41 nsew
rlabel locali s -12574 16048 -12475 16210 4 VDD
port 41 nsew
rlabel locali s -12740 16210 -12475 16244 4 VDD
port 41 nsew
rlabel locali s -12304 16311 -12114 16314 4 VDD
port 41 nsew
rlabel locali s -12304 16314 -12238 16415 4 VDD
port 41 nsew
rlabel locali s -12574 16244 -12475 16406 4 VDD
port 41 nsew
rlabel locali s -12740 16406 -12475 16440 4 VDD
port 41 nsew
rlabel locali s -12574 16440 -12475 16488 4 VDD
port 41 nsew
rlabel locali s -6542 17925 -4711 18014 4 VDD
port 41 nsew
rlabel locali s -4779 18014 -4711 18174 4 VDD
port 41 nsew
rlabel locali s -5070 18174 -4711 18208 4 VDD
port 41 nsew
rlabel locali s -4779 18208 -4711 18370 4 VDD
port 41 nsew
rlabel locali s -6542 18014 -6474 18212 4 VDD
port 41 nsew
rlabel locali s -6542 18212 -6471 18272 4 VDD
port 41 nsew
rlabel locali s -6542 18272 -6180 18306 4 VDD
port 41 nsew
rlabel locali s -5070 18370 -4711 18404 4 VDD
port 41 nsew
rlabel locali s -6542 18306 -6471 18387 4 VDD
port 41 nsew
rlabel locali s -11469 17925 -9638 18014 4 VDD
port 41 nsew
rlabel locali s -9706 18014 -9638 18174 4 VDD
port 41 nsew
rlabel locali s -10498 18014 -10331 18015 4 VDD
port 41 nsew
rlabel locali s -9997 18174 -9638 18208 4 VDD
port 41 nsew
rlabel locali s -9706 18208 -9638 18370 4 VDD
port 41 nsew
rlabel locali s -11469 18014 -11401 18212 4 VDD
port 41 nsew
rlabel locali s -11469 18212 -11398 18272 4 VDD
port 41 nsew
rlabel locali s -11469 18272 -11107 18306 4 VDD
port 41 nsew
rlabel locali s -9997 18370 -9638 18387 4 VDD
port 41 nsew
rlabel locali s -9997 18387 -6471 18404 4 VDD
port 41 nsew
rlabel locali s -4779 18404 -4711 18566 4 VDD
port 41 nsew
rlabel locali s -9706 18404 -6471 18468 4 VDD
port 41 nsew
rlabel locali s -11469 18306 -11398 18468 4 VDD
port 41 nsew
rlabel locali s -9706 18468 -6180 18502 4 VDD
port 41 nsew
rlabel locali s -11469 18468 -11107 18502 4 VDD
port 41 nsew
rlabel locali s -9706 18502 -6471 18540 4 VDD
port 41 nsew
rlabel locali s -5070 18566 -4711 18600 4 VDD
port 41 nsew
rlabel locali s -4779 18600 -4711 19011 4 VDD
port 41 nsew
rlabel locali s -6542 18540 -6471 18664 4 VDD
port 41 nsew
rlabel locali s -6542 18664 -6180 18698 4 VDD
port 41 nsew
rlabel locali s -6542 18698 -6471 18707 4 VDD
port 41 nsew
rlabel locali s -5070 19011 -4711 19045 4 VDD
port 41 nsew
rlabel locali s -6542 18707 -6474 19029 4 VDD
port 41 nsew
rlabel locali s -4779 19045 -4711 19207 4 VDD
port 41 nsew
rlabel locali s -5070 19207 -4711 19241 4 VDD
port 41 nsew
rlabel locali s -4779 19241 -4711 19403 4 VDD
port 41 nsew
rlabel locali s -5070 19403 -4711 19437 4 VDD
port 41 nsew
rlabel locali s -4779 19437 -4711 19498 4 VDD
port 41 nsew
rlabel locali s -4774 19498 -4711 20396 4 VDD
port 41 nsew
rlabel locali s -6539 19029 -6476 19954 4 VDD
port 41 nsew
rlabel locali s -8190 19189 -8126 19199 4 VDD
port 41 nsew
rlabel locali s -8190 19199 -7709 19233 4 VDD
port 41 nsew
rlabel locali s -8190 19233 -8126 19395 4 VDD
port 41 nsew
rlabel locali s -8190 19395 -7709 19429 4 VDD
port 41 nsew
rlabel locali s -8190 19429 -8126 19591 4 VDD
port 41 nsew
rlabel locali s -8391 18540 -8238 19359 4 VDD
port 41 nsew
rlabel locali s -9706 18540 -9638 18566 4 VDD
port 41 nsew
rlabel locali s -9997 18566 -9638 18600 4 VDD
port 41 nsew
rlabel locali s -9706 18600 -9638 19011 4 VDD
port 41 nsew
rlabel locali s -11469 18502 -11398 18664 4 VDD
port 41 nsew
rlabel locali s -11469 18664 -11107 18698 4 VDD
port 41 nsew
rlabel locali s -11469 18698 -11398 18707 4 VDD
port 41 nsew
rlabel locali s -9997 19011 -9638 19045 4 VDD
port 41 nsew
rlabel locali s -11469 18707 -11401 19029 4 VDD
port 41 nsew
rlabel locali s -8680 19177 -8581 19225 4 VDD
port 41 nsew
rlabel locali s -9706 19045 -9638 19207 4 VDD
port 41 nsew
rlabel locali s -8946 19225 -8581 19259 4 VDD
port 41 nsew
rlabel locali s -9997 19207 -9638 19241 4 VDD
port 41 nsew
rlabel locali s -8680 19259 -8581 19359 4 VDD
port 41 nsew
rlabel locali s -8680 19359 -8238 19421 4 VDD
port 41 nsew
rlabel locali s -9706 19241 -9638 19403 4 VDD
port 41 nsew
rlabel locali s -8946 19421 -8238 19455 4 VDD
port 41 nsew
rlabel locali s -9997 19403 -9638 19437 4 VDD
port 41 nsew
rlabel locali s -8680 19455 -8238 19531 4 VDD
port 41 nsew
rlabel locali s -8391 19531 -8238 19591 4 VDD
port 41 nsew
rlabel locali s -8190 19591 -7709 19625 4 VDD
port 41 nsew
rlabel locali s -8190 19625 -8076 19631 4 VDD
port 41 nsew
rlabel locali s -8391 19591 -8231 19628 4 VDD
port 41 nsew
rlabel locali s -8175 19631 -8076 19808 4 VDD
port 41 nsew
rlabel locali s -8175 19808 -7910 19842 4 VDD
port 41 nsew
rlabel locali s -8391 19628 -8224 19817 4 VDD
port 41 nsew
rlabel locali s -6539 19954 -6471 20015 4 VDD
port 41 nsew
rlabel locali s -8175 19842 -8076 20004 4 VDD
port 41 nsew
rlabel locali s -6539 20015 -6180 20049 4 VDD
port 41 nsew
rlabel locali s -8175 20004 -7910 20038 4 VDD
port 41 nsew
rlabel locali s -6539 20049 -6471 20211 4 VDD
port 41 nsew
rlabel locali s -8175 20038 -8076 20200 4 VDD
port 41 nsew
rlabel locali s -6539 20211 -6180 20245 4 VDD
port 41 nsew
rlabel locali s -8175 20200 -7910 20234 4 VDD
port 41 nsew
rlabel locali s -4779 20396 -4711 20874 4 VDD
port 41 nsew
rlabel locali s -6539 20245 -6471 20407 4 VDD
port 41 nsew
rlabel locali s -8175 20234 -8076 20396 4 VDD
port 41 nsew
rlabel locali s -6539 20407 -6180 20441 4 VDD
port 41 nsew
rlabel locali s -8175 20396 -7910 20430 4 VDD
port 41 nsew
rlabel locali s -5070 20874 -4711 20908 4 VDD
port 41 nsew
rlabel locali s -4779 20908 -4711 21070 4 VDD
port 41 nsew
rlabel locali s -6539 20441 -6471 20972 4 VDD
port 41 nsew
rlabel locali s -8175 20430 -8076 20478 4 VDD
port 41 nsew
rlabel locali s -8391 19817 -8238 20187 4 VDD
port 41 nsew
rlabel locali s -8680 19531 -8581 19617 4 VDD
port 41 nsew
rlabel locali s -9706 19437 -9638 19498 4 VDD
port 41 nsew
rlabel locali s -8946 19617 -8581 19651 4 VDD
port 41 nsew
rlabel locali s -8680 19651 -8581 19813 4 VDD
port 41 nsew
rlabel locali s -8946 19813 -8581 19847 4 VDD
port 41 nsew
rlabel locali s -8680 19847 -8581 19895 4 VDD
port 41 nsew
rlabel locali s -8437 20187 -8238 20188 4 VDD
port 41 nsew
rlabel locali s -8500 20188 -8238 20198 4 VDD
port 41 nsew
rlabel locali s -8917 20198 -8238 20232 4 VDD
port 41 nsew
rlabel locali s -8500 20232 -8238 20394 4 VDD
port 41 nsew
rlabel locali s -8917 20394 -8238 20428 4 VDD
port 41 nsew
rlabel locali s -9701 19498 -9638 20396 4 VDD
port 41 nsew
rlabel locali s -11466 19029 -11403 19954 4 VDD
port 41 nsew
rlabel locali s -11466 19954 -11398 20015 4 VDD
port 41 nsew
rlabel locali s -11466 20015 -11107 20049 4 VDD
port 41 nsew
rlabel locali s -11466 20049 -11398 20211 4 VDD
port 41 nsew
rlabel locali s -11466 20211 -11107 20245 4 VDD
port 41 nsew
rlabel locali s -8500 20428 -8238 20590 4 VDD
port 41 nsew
rlabel locali s -8917 20590 -8238 20624 4 VDD
port 41 nsew
rlabel locali s -8550 20624 -8238 20630 4 VDD
port 41 nsew
rlabel locali s -8408 20630 -8238 20635 4 VDD
port 41 nsew
rlabel locali s -8408 20635 -8214 20641 4 VDD
port 41 nsew
rlabel locali s -8408 20641 -8088 20646 4 VDD
port 41 nsew
rlabel locali s -8408 20646 -7498 20680 4 VDD
port 41 nsew
rlabel locali s -8408 20680 -8088 20686 4 VDD
port 41 nsew
rlabel locali s -8408 20686 -8214 20805 4 VDD
port 41 nsew
rlabel locali s -8391 20805 -8214 20836 4 VDD
port 41 nsew
rlabel locali s -8391 20836 -8091 20842 4 VDD
port 41 nsew
rlabel locali s -8391 20842 -7498 20876 4 VDD
port 41 nsew
rlabel locali s -8391 20876 -8091 20881 4 VDD
port 41 nsew
rlabel locali s -6539 20972 -6180 21006 4 VDD
port 41 nsew
rlabel locali s -5070 21070 -4711 21104 4 VDD
port 41 nsew
rlabel locali s -4779 21104 -4711 21266 4 VDD
port 41 nsew
rlabel locali s -6539 21006 -6471 21168 4 VDD
port 41 nsew
rlabel locali s -6539 21168 -6180 21202 4 VDD
port 41 nsew
rlabel locali s -6539 21202 -6471 21247 4 VDD
port 41 nsew
rlabel locali s -5070 21266 -4711 21300 4 VDD
port 41 nsew
rlabel locali s -4779 21300 -4711 21711 4 VDD
port 41 nsew
rlabel locali s -6540 21247 -6471 21364 4 VDD
port 41 nsew
rlabel locali s -8391 20881 -8214 21258 4 VDD
port 41 nsew
rlabel locali s -8391 21258 -8090 21265 4 VDD
port 41 nsew
rlabel locali s -8391 21265 -7498 21299 4 VDD
port 41 nsew
rlabel locali s -8391 21299 -8090 21300 4 VDD
port 41 nsew
rlabel locali s -8550 20630 -8451 20807 4 VDD
port 41 nsew
rlabel locali s -8716 20807 -8451 20841 4 VDD
port 41 nsew
rlabel locali s -8550 20841 -8451 21003 4 VDD
port 41 nsew
rlabel locali s -9706 20396 -9638 20874 4 VDD
port 41 nsew
rlabel locali s -11466 20245 -11398 20407 4 VDD
port 41 nsew
rlabel locali s -11466 20407 -11107 20441 4 VDD
port 41 nsew
rlabel locali s -9997 20874 -9638 20908 4 VDD
port 41 nsew
rlabel locali s -8716 21003 -8451 21037 4 VDD
port 41 nsew
rlabel locali s -8550 21037 -8451 21199 4 VDD
port 41 nsew
rlabel locali s -9706 20908 -9638 21070 4 VDD
port 41 nsew
rlabel locali s -11466 20441 -11398 20972 4 VDD
port 41 nsew
rlabel locali s -11466 20972 -11107 21006 4 VDD
port 41 nsew
rlabel locali s -9997 21070 -9638 21104 4 VDD
port 41 nsew
rlabel locali s -8716 21199 -8451 21233 4 VDD
port 41 nsew
rlabel locali s -8280 21300 -8090 21303 4 VDD
port 41 nsew
rlabel locali s -6540 21364 -6180 21398 4 VDD
port 41 nsew
rlabel locali s -6540 21398 -6471 21407 4 VDD
port 41 nsew
rlabel locali s -8280 21303 -8214 21404 4 VDD
port 41 nsew
rlabel locali s -8550 21233 -8451 21395 4 VDD
port 41 nsew
rlabel locali s -9706 21104 -9638 21266 4 VDD
port 41 nsew
rlabel locali s -11466 21006 -11398 21168 4 VDD
port 41 nsew
rlabel locali s -11466 21168 -11107 21202 4 VDD
port 41 nsew
rlabel locali s -11466 21202 -11398 21247 4 VDD
port 41 nsew
rlabel locali s -9997 21266 -9638 21300 4 VDD
port 41 nsew
rlabel locali s -5070 21711 -4711 21745 4 VDD
port 41 nsew
rlabel locali s -6540 21407 -6472 21720 4 VDD
port 41 nsew
rlabel locali s -8716 21395 -8451 21429 4 VDD
port 41 nsew
rlabel locali s -8550 21429 -8451 21477 4 VDD
port 41 nsew
rlabel locali s -9706 21300 -9638 21711 4 VDD
port 41 nsew
rlabel locali s -11467 21247 -11398 21364 4 VDD
port 41 nsew
rlabel locali s -11467 21364 -11107 21398 4 VDD
port 41 nsew
rlabel locali s -11467 21398 -11398 21407 4 VDD
port 41 nsew
rlabel locali s -4779 21745 -4711 21907 4 VDD
port 41 nsew
rlabel locali s -5070 21907 -4711 21941 4 VDD
port 41 nsew
rlabel locali s -4779 21941 -4711 22103 4 VDD
port 41 nsew
rlabel locali s -5070 22103 -4711 22137 4 VDD
port 41 nsew
rlabel locali s -4779 22137 -4711 22198 4 VDD
port 41 nsew
rlabel locali s -4774 22198 -4711 22950 4 VDD
port 41 nsew
rlabel locali s -6539 21720 -6476 22654 4 VDD
port 41 nsew
rlabel locali s -9997 21711 -9638 21745 4 VDD
port 41 nsew
rlabel locali s -11467 21407 -11399 21720 4 VDD
port 41 nsew
rlabel locali s -9706 21745 -9638 21907 4 VDD
port 41 nsew
rlabel locali s -9997 21907 -9638 21941 4 VDD
port 41 nsew
rlabel locali s -9706 21941 -9638 22003 4 VDD
port 41 nsew
rlabel locali s -6539 22654 -6471 22715 4 VDD
port 41 nsew
rlabel locali s -6539 22715 -6180 22749 4 VDD
port 41 nsew
rlabel locali s -6539 22749 -6471 22911 4 VDD
port 41 nsew
rlabel locali s -6539 22911 -6180 22945 4 VDD
port 41 nsew
rlabel locali s -4774 22950 -4675 23150 4 VDD
port 41 nsew
rlabel locali s -6539 22945 -6471 23107 4 VDD
port 41 nsew
rlabel locali s -6539 23107 -6180 23141 4 VDD
port 41 nsew
rlabel locali s -4764 23150 -4675 24532 4 VDD
port 41 nsew
rlabel locali s -6539 23141 -6471 23597 4 VDD
port 41 nsew
rlabel locali s -6539 23597 -6180 23631 4 VDD
port 41 nsew
rlabel locali s -6539 23631 -6471 23793 4 VDD
port 41 nsew
rlabel locali s -6539 23793 -6180 23827 4 VDD
port 41 nsew
rlabel locali s -6539 23827 -6471 23989 4 VDD
port 41 nsew
rlabel locali s -6539 23989 -6180 24023 4 VDD
port 41 nsew
rlabel locali s -6539 24023 -6471 24032 4 VDD
port 41 nsew
rlabel locali s -9706 22003 -9616 22103 4 VDD
port 41 nsew
rlabel locali s -9997 22103 -9616 22137 4 VDD
port 41 nsew
rlabel locali s -9706 22137 -9616 22198 4 VDD
port 41 nsew
rlabel locali s -4888 24532 -4675 24536 4 VDD
port 41 nsew
rlabel locali s -5480 24536 -4675 24570 4 VDD
port 41 nsew
rlabel locali s -9701 22198 -9616 24559 4 VDD
port 41 nsew
rlabel locali s -11466 21720 -11403 22654 4 VDD
port 41 nsew
rlabel locali s -11466 22654 -11398 22715 4 VDD
port 41 nsew
rlabel locali s -11466 22715 -11107 22749 4 VDD
port 41 nsew
rlabel locali s -11466 22749 -11398 22911 4 VDD
port 41 nsew
rlabel locali s -11466 22911 -11107 22945 4 VDD
port 41 nsew
rlabel locali s -11466 22945 -11398 23107 4 VDD
port 41 nsew
rlabel locali s -11466 23107 -11107 23141 4 VDD
port 41 nsew
rlabel locali s -11466 23141 -11398 23597 4 VDD
port 41 nsew
rlabel locali s -11466 23597 -11107 23631 4 VDD
port 41 nsew
rlabel locali s -11466 23631 -11398 23793 4 VDD
port 41 nsew
rlabel locali s -11466 23793 -11107 23827 4 VDD
port 41 nsew
rlabel locali s -11466 23827 -11398 23989 4 VDD
port 41 nsew
rlabel locali s -11466 23989 -11107 24023 4 VDD
port 41 nsew
rlabel locali s -11466 24023 -11398 24032 4 VDD
port 41 nsew
rlabel locali s -9822 24559 -9616 24563 4 VDD
port 41 nsew
rlabel locali s -4888 24570 -4675 24577 4 VDD
port 41 nsew
rlabel locali s -4764 24577 -4675 24954 4 VDD
port 41 nsew
rlabel locali s -10414 24563 -9616 24597 4 VDD
port 41 nsew
rlabel locali s -9822 24597 -9616 24604 4 VDD
port 41 nsew
rlabel locali s -4887 24954 -4675 24959 4 VDD
port 41 nsew
rlabel locali s -5480 24959 -4675 24993 4 VDD
port 41 nsew
rlabel locali s -9701 24604 -9616 24981 4 VDD
port 41 nsew
rlabel locali s -9821 24981 -9616 24986 4 VDD
port 41 nsew
rlabel locali s -4887 24993 -4675 24999 4 VDD
port 41 nsew
rlabel locali s -4764 24999 -4675 25149 4 VDD
port 41 nsew
rlabel locali s -10414 24986 -9616 25020 4 VDD
port 41 nsew
rlabel locali s -9821 25020 -9616 25026 4 VDD
port 41 nsew
rlabel locali s -4890 25149 -4675 25155 4 VDD
port 41 nsew
rlabel locali s -5480 25155 -4675 25189 4 VDD
port 41 nsew
rlabel locali s -9701 25026 -9616 25176 4 VDD
port 41 nsew
rlabel locali s -9824 25176 -9616 25182 4 VDD
port 41 nsew
rlabel locali s -4890 25189 -4675 25194 4 VDD
port 41 nsew
rlabel locali s -4764 25194 -4675 25279 4 VDD
port 41 nsew
rlabel locali s -10414 25182 -9616 25216 4 VDD
port 41 nsew
rlabel locali s -9824 25216 -9616 25221 4 VDD
port 41 nsew
rlabel locali s -4857 25279 -4675 25281 4 VDD
port 41 nsew
rlabel locali s -4857 25281 -4664 26644 4 VDD
port 41 nsew
rlabel locali s -9701 25221 -9616 25799 4 VDD
port 41 nsew
rlabel locali s -11736 25799 -7146 25888 4 VDD
port 41 nsew
rlabel locali s -7214 25888 -7146 26086 4 VDD
port 41 nsew
rlabel locali s -8977 25888 -8909 26048 4 VDD
port 41 nsew
rlabel locali s -9973 25888 -9816 25889 4 VDD
port 41 nsew
rlabel locali s -8977 26048 -8618 26082 4 VDD
port 41 nsew
rlabel locali s -7217 26086 -7146 26146 4 VDD
port 41 nsew
rlabel locali s -8977 26082 -8909 26087 4 VDD
port 41 nsew
rlabel locali s -9973 25889 -9905 26048 4 VDD
port 41 nsew
rlabel locali s -10264 26048 -9905 26082 4 VDD
port 41 nsew
rlabel locali s -9973 26082 -9905 26087 4 VDD
port 41 nsew
rlabel locali s -11736 25888 -11668 26086 4 VDD
port 41 nsew
rlabel locali s -7508 26146 -7146 26180 4 VDD
port 41 nsew
rlabel locali s -6756 26296 -6688 26305 4 VDD
port 41 nsew
rlabel locali s -6756 26305 -6397 26312 4 VDD
port 41 nsew
rlabel locali s -7217 26180 -7146 26312 4 VDD
port 41 nsew
rlabel locali s -9973 26087 -8909 26244 4 VDD
port 41 nsew
rlabel locali s -11736 26086 -11665 26146 4 VDD
port 41 nsew
rlabel locali s -11736 26146 -11374 26180 4 VDD
port 41 nsew
rlabel locali s -10264 26244 -8618 26278 4 VDD
port 41 nsew
rlabel locali s -7217 26312 -6397 26339 4 VDD
port 41 nsew
rlabel locali s -7217 26339 -6688 26342 4 VDD
port 41 nsew
rlabel locali s -7508 26342 -6688 26376 4 VDD
port 41 nsew
rlabel locali s -9973 26278 -8909 26356 4 VDD
port 41 nsew
rlabel locali s -11736 26180 -11665 26342 4 VDD
port 41 nsew
rlabel locali s -7217 26376 -6688 26400 4 VDD
port 41 nsew
rlabel locali s -6756 26400 -6688 26495 4 VDD
port 41 nsew
rlabel locali s -7217 26400 -7146 26495 4 VDD
port 41 nsew
rlabel locali s -8977 26356 -8909 26440 4 VDD
port 41 nsew
rlabel locali s -8977 26440 -8618 26474 4 VDD
port 41 nsew
rlabel locali s -7217 26495 -6688 26501 4 VDD
port 41 nsew
rlabel locali s -7217 26501 -6397 26535 4 VDD
port 41 nsew
rlabel locali s -7217 26535 -6688 26538 4 VDD
port 41 nsew
rlabel locali s -7508 26538 -6688 26572 4 VDD
port 41 nsew
rlabel locali s -7217 26572 -6688 26581 4 VDD
port 41 nsew
rlabel locali s -7214 26581 -6688 26583 4 VDD
port 41 nsew
rlabel locali s -5276 26644 -4664 26678 4 VDD
port 41 nsew
rlabel locali s -6756 26583 -6688 26677 4 VDD
port 41 nsew
rlabel locali s -7214 26583 -7146 26677 4 VDD
port 41 nsew
rlabel locali s -5093 26678 -4664 26684 4 VDD
port 41 nsew
rlabel locali s -4964 26684 -4664 26833 4 VDD
port 41 nsew
rlabel locali s -7214 26677 -6688 26697 4 VDD
port 41 nsew
rlabel locali s -7214 26697 -6397 26731 4 VDD
port 41 nsew
rlabel locali s -7214 26731 -6688 26765 4 VDD
port 41 nsew
rlabel locali s -6756 26765 -6688 26791 4 VDD
port 41 nsew
rlabel locali s -5093 26833 -4664 26840 4 VDD
port 41 nsew
rlabel locali s -5276 26840 -4664 26874 4 VDD
port 41 nsew
rlabel locali s -5093 26874 -4664 26879 4 VDD
port 41 nsew
rlabel locali s -4964 26879 -4664 27031 4 VDD
port 41 nsew
rlabel locali s -7214 26765 -7146 26903 4 VDD
port 41 nsew
rlabel locali s -8977 26474 -8909 26633 4 VDD
port 41 nsew
rlabel locali s -9973 26356 -9905 26440 4 VDD
port 41 nsew
rlabel locali s -11736 26342 -11374 26376 4 VDD
port 41 nsew
rlabel locali s -10264 26440 -9905 26474 4 VDD
port 41 nsew
rlabel locali s -9973 26474 -9905 26633 4 VDD
port 41 nsew
rlabel locali s -11736 26376 -11665 26538 4 VDD
port 41 nsew
rlabel locali s -11736 26538 -11374 26572 4 VDD
port 41 nsew
rlabel locali s -11736 26572 -11665 26581 4 VDD
port 41 nsew
rlabel locali s -9973 26633 -8909 26885 4 VDD
port 41 nsew
rlabel locali s -10264 26885 -8618 26902 4 VDD
port 41 nsew
rlabel locali s -5089 27031 -4664 27036 4 VDD
port 41 nsew
rlabel locali s -5276 27036 -4664 27070 4 VDD
port 41 nsew
rlabel locali s -5089 27070 -4664 27077 4 VDD
port 41 nsew
rlabel locali s -4964 27077 -4664 27144 4 VDD
port 41 nsew
rlabel locali s -5093 27144 -4664 27150 4 VDD
port 41 nsew
rlabel locali s -5276 27150 -4664 27184 4 VDD
port 41 nsew
rlabel locali s -5093 27184 -4664 27190 4 VDD
port 41 nsew
rlabel locali s -4964 27190 -4664 27340 4 VDD
port 41 nsew
rlabel locali s -5088 27340 -4664 27346 4 VDD
port 41 nsew
rlabel locali s -5276 27346 -4664 27380 4 VDD
port 41 nsew
rlabel locali s -5088 27380 -4664 27386 4 VDD
port 41 nsew
rlabel locali s -4964 27386 -4664 27453 4 VDD
port 41 nsew
rlabel locali s -5098 27453 -4664 27459 4 VDD
port 41 nsew
rlabel locali s -5276 27459 -4664 27493 4 VDD
port 41 nsew
rlabel locali s -5098 27493 -4664 27499 4 VDD
port 41 nsew
rlabel locali s -4964 27499 -4664 27650 4 VDD
port 41 nsew
rlabel locali s -5086 27650 -4664 27655 4 VDD
port 41 nsew
rlabel locali s -5276 27655 -4664 27689 4 VDD
port 41 nsew
rlabel locali s -5086 27689 -4664 27696 4 VDD
port 41 nsew
rlabel locali s -4857 27696 -4664 27971 4 VDD
port 41 nsew
rlabel locali s -7212 26903 -7149 27828 4 VDD
port 41 nsew
rlabel locali s -8977 26902 -8618 26919 4 VDD
port 41 nsew
rlabel locali s -8977 26919 -8909 27081 4 VDD
port 41 nsew
rlabel locali s -8977 27081 -8618 27115 4 VDD
port 41 nsew
rlabel locali s -8977 27115 -8909 27277 4 VDD
port 41 nsew
rlabel locali s -8977 27277 -8618 27311 4 VDD
port 41 nsew
rlabel locali s -8977 27311 -8909 27372 4 VDD
port 41 nsew
rlabel locali s -8977 27372 -8914 27510 4 VDD
port 41 nsew
rlabel locali s -10264 26902 -9905 26919 4 VDD
port 41 nsew
rlabel locali s -11736 26581 -11668 26903 4 VDD
port 41 nsew
rlabel locali s -14218 25779 -14025 26644 4 VDD
port 41 nsew
rlabel locali s -14218 26644 -13606 26678 4 VDD
port 41 nsew
rlabel locali s -14218 26678 -13789 26684 4 VDD
port 41 nsew
rlabel locali s -14218 26684 -13918 26833 4 VDD
port 41 nsew
rlabel locali s -14218 26833 -13789 26840 4 VDD
port 41 nsew
rlabel locali s -14218 26840 -13606 26874 4 VDD
port 41 nsew
rlabel locali s -14218 26874 -13789 26879 4 VDD
port 41 nsew
rlabel locali s -9973 26919 -9905 27081 4 VDD
port 41 nsew
rlabel locali s -10264 27081 -9905 27115 4 VDD
port 41 nsew
rlabel locali s -9973 27115 -9905 27277 4 VDD
port 41 nsew
rlabel locali s -10264 27277 -9905 27311 4 VDD
port 41 nsew
rlabel locali s -9973 27311 -9905 27372 4 VDD
port 41 nsew
rlabel locali s -9968 27372 -9905 27510 4 VDD
port 41 nsew
rlabel locali s -9968 27510 -8914 27779 4 VDD
port 41 nsew
rlabel locali s -7217 27828 -7149 27889 4 VDD
port 41 nsew
rlabel locali s -7508 27889 -7149 27923 4 VDD
port 41 nsew
rlabel locali s -5830 27966 -5694 27971 4 VDD
port 41 nsew
rlabel locali s -5830 27971 -4664 28086 4 VDD
port 41 nsew
rlabel locali s -4857 28086 -4664 29458 4 VDD
port 41 nsew
rlabel locali s -5830 28086 -5694 28089 4 VDD
port 41 nsew
rlabel locali s -6597 27965 -6461 27970 4 VDD
port 41 nsew
rlabel locali s -7217 27923 -7149 27970 4 VDD
port 41 nsew
rlabel locali s -7217 27970 -6461 28085 4 VDD
port 41 nsew
rlabel locali s -6597 28085 -6461 28088 4 VDD
port 41 nsew
rlabel locali s -7508 28085 -7149 28119 4 VDD
port 41 nsew
rlabel locali s -7217 28119 -7149 28281 4 VDD
port 41 nsew
rlabel locali s -8977 27779 -8914 28270 4 VDD
port 41 nsew
rlabel locali s -7508 28281 -7149 28315 4 VDD
port 41 nsew
rlabel locali s -7217 28315 -7149 28846 4 VDD
port 41 nsew
rlabel locali s -8977 28270 -8909 28372 4 VDD
port 41 nsew
rlabel locali s -9968 27779 -9905 28270 4 VDD
port 41 nsew
rlabel locali s -11733 26903 -11670 27828 4 VDD
port 41 nsew
rlabel locali s -14218 26879 -13918 27031 4 VDD
port 41 nsew
rlabel locali s -14218 27031 -13793 27036 4 VDD
port 41 nsew
rlabel locali s -14218 27036 -13606 27070 4 VDD
port 41 nsew
rlabel locali s -14218 27070 -13793 27077 4 VDD
port 41 nsew
rlabel locali s -14218 27077 -13918 27144 4 VDD
port 41 nsew
rlabel locali s -14218 27144 -13789 27150 4 VDD
port 41 nsew
rlabel locali s -14218 27150 -13606 27184 4 VDD
port 41 nsew
rlabel locali s -14218 27184 -13789 27190 4 VDD
port 41 nsew
rlabel locali s -14218 27190 -13918 27340 4 VDD
port 41 nsew
rlabel locali s -14218 27340 -13794 27346 4 VDD
port 41 nsew
rlabel locali s -14218 27346 -13606 27380 4 VDD
port 41 nsew
rlabel locali s -14218 27380 -13794 27386 4 VDD
port 41 nsew
rlabel locali s -14218 27386 -13918 27453 4 VDD
port 41 nsew
rlabel locali s -14218 27453 -13784 27459 4 VDD
port 41 nsew
rlabel locali s -14218 27459 -13606 27493 4 VDD
port 41 nsew
rlabel locali s -14218 27493 -13784 27499 4 VDD
port 41 nsew
rlabel locali s -14218 27499 -13918 27650 4 VDD
port 41 nsew
rlabel locali s -14218 27650 -13796 27655 4 VDD
port 41 nsew
rlabel locali s -14218 27655 -13606 27689 4 VDD
port 41 nsew
rlabel locali s -14218 27689 -13796 27696 4 VDD
port 41 nsew
rlabel locali s -11733 27828 -11665 27889 4 VDD
port 41 nsew
rlabel locali s -11733 27889 -11374 27923 4 VDD
port 41 nsew
rlabel locali s -11733 27923 -11665 27970 4 VDD
port 41 nsew
rlabel locali s -12421 27965 -12285 27970 4 VDD
port 41 nsew
rlabel locali s -12421 27970 -11665 28085 4 VDD
port 41 nsew
rlabel locali s -11733 28085 -11374 28119 4 VDD
port 41 nsew
rlabel locali s -12421 28085 -12285 28088 4 VDD
port 41 nsew
rlabel locali s -13188 27966 -13052 27971 4 VDD
port 41 nsew
rlabel locali s -14218 27696 -14025 27971 4 VDD
port 41 nsew
rlabel locali s -14218 27971 -13052 28086 4 VDD
port 41 nsew
rlabel locali s -13188 28086 -13052 28089 4 VDD
port 41 nsew
rlabel locali s -9973 28270 -9905 28372 4 VDD
port 41 nsew
rlabel locali s -11733 28119 -11665 28281 4 VDD
port 41 nsew
rlabel locali s -11733 28281 -11374 28315 4 VDD
port 41 nsew
rlabel locali s -9973 28372 -8909 28641 4 VDD
port 41 nsew
rlabel locali s -8977 28641 -8909 28748 4 VDD
port 41 nsew
rlabel locali s -8977 28748 -8618 28782 4 VDD
port 41 nsew
rlabel locali s -7508 28846 -7149 28880 4 VDD
port 41 nsew
rlabel locali s -7217 28880 -7149 29042 4 VDD
port 41 nsew
rlabel locali s -8977 28782 -8909 28944 4 VDD
port 41 nsew
rlabel locali s -8977 28944 -8618 28978 4 VDD
port 41 nsew
rlabel locali s -7508 29042 -7149 29076 4 VDD
port 41 nsew
rlabel locali s -7217 29076 -7149 29121 4 VDD
port 41 nsew
rlabel locali s -5276 29144 -4895 29178 4 VDD
port 41 nsew
rlabel locali s -5093 29178 -4895 29184 4 VDD
port 41 nsew
rlabel locali s -4964 29184 -4895 29333 4 VDD
port 41 nsew
rlabel locali s -7217 29121 -7148 29238 4 VDD
port 41 nsew
rlabel locali s -8977 28978 -8909 29140 4 VDD
port 41 nsew
rlabel locali s -8977 29140 -8618 29174 4 VDD
port 41 nsew
rlabel locali s -7508 29238 -7148 29272 4 VDD
port 41 nsew
rlabel locali s -7217 29272 -7148 29281 4 VDD
port 41 nsew
rlabel locali s -8977 29174 -8909 29275 4 VDD
port 41 nsew
rlabel locali s -9973 28641 -9905 28748 4 VDD
port 41 nsew
rlabel locali s -10264 28748 -9905 28782 4 VDD
port 41 nsew
rlabel locali s -9973 28782 -9905 28944 4 VDD
port 41 nsew
rlabel locali s -11733 28315 -11665 28846 4 VDD
port 41 nsew
rlabel locali s -11733 28846 -11374 28880 4 VDD
port 41 nsew
rlabel locali s -10264 28944 -9905 28978 4 VDD
port 41 nsew
rlabel locali s -9973 28978 -9905 29140 4 VDD
port 41 nsew
rlabel locali s -11733 28880 -11665 29042 4 VDD
port 41 nsew
rlabel locali s -11733 29042 -11374 29076 4 VDD
port 41 nsew
rlabel locali s -11733 29076 -11665 29121 4 VDD
port 41 nsew
rlabel locali s -10264 29140 -9905 29174 4 VDD
port 41 nsew
rlabel locali s -9973 29174 -9905 29275 4 VDD
port 41 nsew
rlabel locali s -11734 29121 -11665 29238 4 VDD
port 41 nsew
rlabel locali s -13987 29144 -13606 29178 4 VDD
port 41 nsew
rlabel locali s -13987 29178 -13789 29184 4 VDD
port 41 nsew
rlabel locali s -11734 29238 -11374 29272 4 VDD
port 41 nsew
rlabel locali s -5093 29333 -4895 29340 4 VDD
port 41 nsew
rlabel locali s -5276 29340 -4895 29374 4 VDD
port 41 nsew
rlabel locali s -5093 29374 -4895 29379 4 VDD
port 41 nsew
rlabel locali s -4964 29379 -4895 29458 4 VDD
port 41 nsew
rlabel locali s -4964 29458 -4664 29531 4 VDD
port 41 nsew
rlabel locali s -5089 29531 -4664 29536 4 VDD
port 41 nsew
rlabel locali s -5276 29536 -4664 29570 4 VDD
port 41 nsew
rlabel locali s -5089 29570 -4664 29577 4 VDD
port 41 nsew
rlabel locali s -4964 29577 -4664 29644 4 VDD
port 41 nsew
rlabel locali s -7216 29281 -7148 29594 4 VDD
port 41 nsew
rlabel locali s -9973 29275 -8909 29544 4 VDD
port 41 nsew
rlabel locali s -11734 29272 -11665 29281 4 VDD
port 41 nsew
rlabel locali s -8977 29544 -8909 29585 4 VDD
port 41 nsew
rlabel locali s -5093 29644 -4664 29650 4 VDD
port 41 nsew
rlabel locali s -5276 29650 -4664 29684 4 VDD
port 41 nsew
rlabel locali s -5093 29684 -4664 29690 4 VDD
port 41 nsew
rlabel locali s -4964 29690 -4664 29840 4 VDD
port 41 nsew
rlabel locali s -5088 29840 -4664 29846 4 VDD
port 41 nsew
rlabel locali s -5276 29846 -4664 29880 4 VDD
port 41 nsew
rlabel locali s -5088 29880 -4664 29886 4 VDD
port 41 nsew
rlabel locali s -4964 29886 -4664 29953 4 VDD
port 41 nsew
rlabel locali s -5098 29953 -4664 29959 4 VDD
port 41 nsew
rlabel locali s -5276 29959 -4664 29993 4 VDD
port 41 nsew
rlabel locali s -5098 29993 -4664 29999 4 VDD
port 41 nsew
rlabel locali s -4964 29999 -4664 30051 4 VDD
port 41 nsew
rlabel locali s -4857 30051 -4664 30539 4 VDD
port 41 nsew
rlabel locali s -4964 30051 -4895 30150 4 VDD
port 41 nsew
rlabel locali s -5086 30150 -4895 30155 4 VDD
port 41 nsew
rlabel locali s -5276 30155 -4895 30189 4 VDD
port 41 nsew
rlabel locali s -5086 30189 -4895 30196 4 VDD
port 41 nsew
rlabel locali s -7212 29594 -7149 30528 4 VDD
port 41 nsew
rlabel locali s -8977 29585 -8618 29619 4 VDD
port 41 nsew
rlabel locali s -8977 29619 -8909 29781 4 VDD
port 41 nsew
rlabel locali s -8977 29781 -8618 29815 4 VDD
port 41 nsew
rlabel locali s -8977 29815 -8909 29977 4 VDD
port 41 nsew
rlabel locali s -8977 29977 -8618 30011 4 VDD
port 41 nsew
rlabel locali s -8977 30011 -8909 30072 4 VDD
port 41 nsew
rlabel locali s -8977 30072 -8914 30306 4 VDD
port 41 nsew
rlabel locali s -9973 29544 -9905 29585 4 VDD
port 41 nsew
rlabel locali s -10264 29585 -9905 29619 4 VDD
port 41 nsew
rlabel locali s -11734 29281 -11666 29594 4 VDD
port 41 nsew
rlabel locali s -13987 29184 -13918 29333 4 VDD
port 41 nsew
rlabel locali s -13987 29333 -13789 29340 4 VDD
port 41 nsew
rlabel locali s -13987 29340 -13606 29374 4 VDD
port 41 nsew
rlabel locali s -13987 29374 -13789 29379 4 VDD
port 41 nsew
rlabel locali s -13987 29379 -13918 29458 4 VDD
port 41 nsew
rlabel locali s -14218 28086 -14025 29458 4 VDD
port 41 nsew
rlabel locali s -14218 29458 -13918 29531 4 VDD
port 41 nsew
rlabel locali s -14218 29531 -13793 29536 4 VDD
port 41 nsew
rlabel locali s -14218 29536 -13606 29570 4 VDD
port 41 nsew
rlabel locali s -14218 29570 -13793 29577 4 VDD
port 41 nsew
rlabel locali s -9973 29619 -9905 29781 4 VDD
port 41 nsew
rlabel locali s -10264 29781 -9905 29815 4 VDD
port 41 nsew
rlabel locali s -9973 29815 -9905 29977 4 VDD
port 41 nsew
rlabel locali s -10264 29977 -9905 30011 4 VDD
port 41 nsew
rlabel locali s -9973 30011 -9905 30072 4 VDD
port 41 nsew
rlabel locali s -9968 30072 -9905 30306 4 VDD
port 41 nsew
rlabel locali s -5865 30533 -5729 30539 4 VDD
port 41 nsew
rlabel locali s -5865 30539 -4664 30653 4 VDD
port 41 nsew
rlabel locali s -4857 30653 -4664 31974 4 VDD
port 41 nsew
rlabel locali s -5865 30653 -5729 30656 4 VDD
port 41 nsew
rlabel locali s -6453 30532 -6317 30536 4 VDD
port 41 nsew
rlabel locali s -7217 30528 -7149 30536 4 VDD
port 41 nsew
rlabel locali s -7217 30536 -6317 30589 4 VDD
port 41 nsew
rlabel locali s -9968 30306 -8914 30575 4 VDD
port 41 nsew
rlabel locali s -11733 29594 -11670 30528 4 VDD
port 41 nsew
rlabel locali s -14218 29577 -13918 29644 4 VDD
port 41 nsew
rlabel locali s -14218 29644 -13789 29650 4 VDD
port 41 nsew
rlabel locali s -14218 29650 -13606 29684 4 VDD
port 41 nsew
rlabel locali s -14218 29684 -13789 29690 4 VDD
port 41 nsew
rlabel locali s -14218 29690 -13918 29840 4 VDD
port 41 nsew
rlabel locali s -14218 29840 -13794 29846 4 VDD
port 41 nsew
rlabel locali s -14218 29846 -13606 29880 4 VDD
port 41 nsew
rlabel locali s -14218 29880 -13794 29886 4 VDD
port 41 nsew
rlabel locali s -14218 29886 -13918 29953 4 VDD
port 41 nsew
rlabel locali s -14218 29953 -13784 29959 4 VDD
port 41 nsew
rlabel locali s -14218 29959 -13606 29993 4 VDD
port 41 nsew
rlabel locali s -14218 29993 -13784 29999 4 VDD
port 41 nsew
rlabel locali s -14218 29999 -13918 30051 4 VDD
port 41 nsew
rlabel locali s -13987 30051 -13918 30150 4 VDD
port 41 nsew
rlabel locali s -13987 30150 -13796 30155 4 VDD
port 41 nsew
rlabel locali s -13987 30155 -13606 30189 4 VDD
port 41 nsew
rlabel locali s -13987 30189 -13796 30196 4 VDD
port 41 nsew
rlabel locali s -7508 30589 -6317 30623 4 VDD
port 41 nsew
rlabel locali s -7217 30623 -6317 30651 4 VDD
port 41 nsew
rlabel locali s -6453 30651 -6317 30655 4 VDD
port 41 nsew
rlabel locali s -7217 30651 -7149 30785 4 VDD
port 41 nsew
rlabel locali s -7508 30785 -7149 30819 4 VDD
port 41 nsew
rlabel locali s -7217 30819 -7149 30981 4 VDD
port 41 nsew
rlabel locali s -7508 30981 -7149 31015 4 VDD
port 41 nsew
rlabel locali s -7217 31015 -7149 31471 4 VDD
port 41 nsew
rlabel locali s -8977 30575 -8914 31024 4 VDD
port 41 nsew
rlabel locali s -9968 30575 -9905 31024 4 VDD
port 41 nsew
rlabel locali s -11733 30528 -11665 30536 4 VDD
port 41 nsew
rlabel locali s -12565 30532 -12429 30536 4 VDD
port 41 nsew
rlabel locali s -12565 30536 -11665 30589 4 VDD
port 41 nsew
rlabel locali s -12565 30589 -11374 30623 4 VDD
port 41 nsew
rlabel locali s -12565 30623 -11665 30651 4 VDD
port 41 nsew
rlabel locali s -11733 30651 -11665 30785 4 VDD
port 41 nsew
rlabel locali s -12565 30651 -12429 30655 4 VDD
port 41 nsew
rlabel locali s -13153 30533 -13017 30539 4 VDD
port 41 nsew
rlabel locali s -14218 30051 -14025 30539 4 VDD
port 41 nsew
rlabel locali s -14218 30539 -13017 30653 4 VDD
port 41 nsew
rlabel locali s -13153 30653 -13017 30656 4 VDD
port 41 nsew
rlabel locali s -11733 30785 -11374 30819 4 VDD
port 41 nsew
rlabel locali s -11733 30819 -11665 30981 4 VDD
port 41 nsew
rlabel locali s -11733 30981 -11374 31015 4 VDD
port 41 nsew
rlabel locali s -11733 31015 -11665 31471 4 VDD
port 41 nsew
rlabel locali s -7508 31471 -7149 31505 4 VDD
port 41 nsew
rlabel locali s -11733 31471 -11374 31505 4 VDD
port 41 nsew
rlabel locali s -5276 31644 -4895 31678 4 VDD
port 41 nsew
rlabel locali s -7217 31505 -7149 31667 4 VDD
port 41 nsew
rlabel locali s -11733 31505 -11665 31667 4 VDD
port 41 nsew
rlabel locali s -5093 31678 -4895 31684 4 VDD
port 41 nsew
rlabel locali s -4964 31684 -4895 31833 4 VDD
port 41 nsew
rlabel locali s -7508 31667 -7149 31701 4 VDD
port 41 nsew
rlabel locali s -11733 31667 -11374 31701 4 VDD
port 41 nsew
rlabel locali s -13987 31644 -13606 31678 4 VDD
port 41 nsew
rlabel locali s -13987 31678 -13789 31684 4 VDD
port 41 nsew
rlabel locali s -7217 31701 -7149 31791 4 VDD
port 41 nsew
rlabel locali s -11733 31701 -11665 31791 4 VDD
port 41 nsew
rlabel locali s -5093 31833 -4895 31840 4 VDD
port 41 nsew
rlabel locali s -5276 31840 -4895 31874 4 VDD
port 41 nsew
rlabel locali s -7263 31791 -7127 31863 4 VDD
port 41 nsew
rlabel locali s -11755 31791 -11619 31863 4 VDD
port 41 nsew
rlabel locali s -13987 31684 -13918 31833 4 VDD
port 41 nsew
rlabel locali s -13987 31833 -13789 31840 4 VDD
port 41 nsew
rlabel locali s -5093 31874 -4895 31879 4 VDD
port 41 nsew
rlabel locali s -4964 31879 -4895 31974 4 VDD
port 41 nsew
rlabel locali s -7508 31863 -7127 31897 4 VDD
port 41 nsew
rlabel locali s -11755 31863 -11374 31897 4 VDD
port 41 nsew
rlabel locali s -13987 31840 -13606 31874 4 VDD
port 41 nsew
rlabel locali s -13987 31874 -13789 31879 4 VDD
port 41 nsew
rlabel locali s -7263 31897 -7127 31914 4 VDD
port 41 nsew
rlabel locali s -11755 31897 -11619 31914 4 VDD
port 41 nsew
rlabel locali s -4964 31974 -4664 32031 4 VDD
port 41 nsew
rlabel locali s -13987 31879 -13918 31974 4 VDD
port 41 nsew
rlabel locali s -14218 30653 -14025 31974 4 VDD
port 41 nsew
rlabel locali s -14218 31974 -13918 32031 4 VDD
port 41 nsew
rlabel locali s -5089 32031 -4664 32036 4 VDD
port 41 nsew
rlabel locali s -14218 32031 -13793 32036 4 VDD
port 41 nsew
rlabel locali s -5276 32036 -4664 32070 4 VDD
port 41 nsew
rlabel locali s -14218 32036 -13606 32070 4 VDD
port 41 nsew
rlabel locali s -5089 32070 -4664 32077 4 VDD
port 41 nsew
rlabel locali s -14218 32070 -13793 32077 4 VDD
port 41 nsew
rlabel locali s -4964 32077 -4664 32144 4 VDD
port 41 nsew
rlabel locali s -5093 32144 -4664 32150 4 VDD
port 41 nsew
rlabel locali s -5276 32150 -4664 32184 4 VDD
port 41 nsew
rlabel locali s -5093 32184 -4664 32190 4 VDD
port 41 nsew
rlabel locali s -4964 32190 -4664 32340 4 VDD
port 41 nsew
rlabel locali s -7262 32085 -7126 32205 4 VDD
port 41 nsew
rlabel locali s -11756 32085 -11620 32205 4 VDD
port 41 nsew
rlabel locali s -14218 32077 -13918 32144 4 VDD
port 41 nsew
rlabel locali s -14218 32144 -13789 32150 4 VDD
port 41 nsew
rlabel locali s -14218 32150 -13606 32184 4 VDD
port 41 nsew
rlabel locali s -14218 32184 -13789 32190 4 VDD
port 41 nsew
rlabel locali s -7525 32205 -7126 32208 4 VDD
port 41 nsew
rlabel locali s -7525 32208 -7153 32239 4 VDD
port 41 nsew
rlabel locali s -11756 32205 -11357 32208 4 VDD
port 41 nsew
rlabel locali s -11729 32208 -11357 32239 4 VDD
port 41 nsew
rlabel locali s -5088 32340 -4664 32346 4 VDD
port 41 nsew
rlabel locali s -5276 32346 -4664 32380 4 VDD
port 41 nsew
rlabel locali s -5088 32380 -4664 32386 4 VDD
port 41 nsew
rlabel locali s -4964 32386 -4664 32453 4 VDD
port 41 nsew
rlabel locali s -7233 32239 -7153 32401 4 VDD
port 41 nsew
rlabel locali s -11729 32239 -11649 32401 4 VDD
port 41 nsew
rlabel locali s -14218 32190 -13918 32340 4 VDD
port 41 nsew
rlabel locali s -14218 32340 -13794 32346 4 VDD
port 41 nsew
rlabel locali s -14218 32346 -13606 32380 4 VDD
port 41 nsew
rlabel locali s -14218 32380 -13794 32386 4 VDD
port 41 nsew
rlabel locali s -7525 32401 -7153 32435 4 VDD
port 41 nsew
rlabel locali s -11729 32401 -11357 32435 4 VDD
port 41 nsew
rlabel locali s -7233 32435 -7153 32440 4 VDD
port 41 nsew
rlabel locali s -11729 32435 -11649 32440 4 VDD
port 41 nsew
rlabel locali s -5098 32453 -4664 32459 4 VDD
port 41 nsew
rlabel locali s -5276 32459 -4664 32493 4 VDD
port 41 nsew
rlabel locali s -5098 32493 -4664 32499 4 VDD
port 41 nsew
rlabel locali s -4964 32499 -4664 32567 4 VDD
port 41 nsew
rlabel locali s -4857 32567 -4664 33021 4 VDD
port 41 nsew
rlabel locali s -4964 32567 -4895 32650 4 VDD
port 41 nsew
rlabel locali s -5086 32650 -4895 32655 4 VDD
port 41 nsew
rlabel locali s -5276 32655 -4895 32689 4 VDD
port 41 nsew
rlabel locali s -5086 32689 -4895 32696 4 VDD
port 41 nsew
rlabel locali s -7232 32440 -7153 32943 4 VDD
port 41 nsew
rlabel locali s -11729 32440 -11650 32943 4 VDD
port 41 nsew
rlabel locali s -14218 32386 -13918 32453 4 VDD
port 41 nsew
rlabel locali s -14218 32453 -13784 32459 4 VDD
port 41 nsew
rlabel locali s -14218 32459 -13606 32493 4 VDD
port 41 nsew
rlabel locali s -14218 32493 -13784 32499 4 VDD
port 41 nsew
rlabel locali s -14218 32499 -13918 32567 4 VDD
port 41 nsew
rlabel locali s -13987 32567 -13918 32650 4 VDD
port 41 nsew
rlabel locali s -13987 32650 -13796 32655 4 VDD
port 41 nsew
rlabel locali s -13987 32655 -13606 32689 4 VDD
port 41 nsew
rlabel locali s -13987 32689 -13796 32696 4 VDD
port 41 nsew
rlabel locali s -7525 32943 -7153 32977 4 VDD
port 41 nsew
rlabel locali s -11729 32943 -11357 32977 4 VDD
port 41 nsew
rlabel locali s -5865 33016 -5729 33021 4 VDD
port 41 nsew
rlabel locali s -5865 33021 -4664 33136 4 VDD
port 41 nsew
rlabel locali s -4857 33136 -4664 34508 4 VDD
port 41 nsew
rlabel locali s -5865 33136 -5729 33139 4 VDD
port 41 nsew
rlabel locali s -6345 33015 -6282 33020 4 VDD
port 41 nsew
rlabel locali s -7232 32977 -7153 33020 4 VDD
port 41 nsew
rlabel locali s -7232 33020 -6282 33135 4 VDD
port 41 nsew
rlabel locali s -6345 33135 -6282 33138 4 VDD
port 41 nsew
rlabel locali s -6345 33138 -6283 33321 4 VDD
port 41 nsew
rlabel locali s -7232 33135 -7153 33139 4 VDD
port 41 nsew
rlabel locali s -11729 32977 -11650 33020 4 VDD
port 41 nsew
rlabel locali s -12600 33015 -12537 33020 4 VDD
port 41 nsew
rlabel locali s -12600 33020 -11650 33135 4 VDD
port 41 nsew
rlabel locali s -11729 33135 -11650 33139 4 VDD
port 41 nsew
rlabel locali s -7525 33139 -7153 33173 4 VDD
port 41 nsew
rlabel locali s -11729 33139 -11357 33173 4 VDD
port 41 nsew
rlabel locali s -7232 33173 -7153 33335 4 VDD
port 41 nsew
rlabel locali s -11729 33173 -11650 33335 4 VDD
port 41 nsew
rlabel locali s -12600 33135 -12537 33138 4 VDD
port 41 nsew
rlabel locali s -13153 33016 -13017 33021 4 VDD
port 41 nsew
rlabel locali s -14218 32567 -14025 33021 4 VDD
port 41 nsew
rlabel locali s -14218 33021 -13017 33136 4 VDD
port 41 nsew
rlabel locali s -12599 33138 -12537 33321 4 VDD
port 41 nsew
rlabel locali s -13153 33136 -13017 33139 4 VDD
port 41 nsew
rlabel locali s -7525 33335 -7153 33369 4 VDD
port 41 nsew
rlabel locali s -11729 33335 -11357 33369 4 VDD
port 41 nsew
rlabel locali s -7232 33369 -7153 33531 4 VDD
port 41 nsew
rlabel locali s -11729 33369 -11650 33531 4 VDD
port 41 nsew
rlabel locali s -7525 33531 -7153 33565 4 VDD
port 41 nsew
rlabel locali s -11729 33531 -11357 33565 4 VDD
port 41 nsew
rlabel locali s -7232 33565 -7153 33890 4 VDD
port 41 nsew
rlabel locali s -11729 33565 -11650 33890 4 VDD
port 41 nsew
rlabel locali s -7272 33890 -7153 33938 4 VDD
port 41 nsew
rlabel locali s -11729 33890 -11610 33938 4 VDD
port 41 nsew
rlabel locali s -7438 33938 -7153 33972 4 VDD
port 41 nsew
rlabel locali s -11729 33938 -11444 33972 4 VDD
port 41 nsew
rlabel locali s -7272 33972 -7153 34134 4 VDD
port 41 nsew
rlabel locali s -11729 33972 -11610 34134 4 VDD
port 41 nsew
rlabel locali s -5276 34144 -4895 34178 4 VDD
port 41 nsew
rlabel locali s -7438 34134 -7153 34168 4 VDD
port 41 nsew
rlabel locali s -11729 34134 -11444 34168 4 VDD
port 41 nsew
rlabel locali s -5093 34178 -4895 34184 4 VDD
port 41 nsew
rlabel locali s -4964 34184 -4895 34333 4 VDD
port 41 nsew
rlabel locali s -7272 34168 -7153 34330 4 VDD
port 41 nsew
rlabel locali s -11729 34168 -11610 34330 4 VDD
port 41 nsew
rlabel locali s -13987 34144 -13606 34178 4 VDD
port 41 nsew
rlabel locali s -13987 34178 -13789 34184 4 VDD
port 41 nsew
rlabel locali s -5093 34333 -4895 34340 4 VDD
port 41 nsew
rlabel locali s -5276 34340 -4895 34374 4 VDD
port 41 nsew
rlabel locali s -7438 34330 -7153 34364 4 VDD
port 41 nsew
rlabel locali s -11729 34330 -11444 34364 4 VDD
port 41 nsew
rlabel locali s -13987 34184 -13918 34333 4 VDD
port 41 nsew
rlabel locali s -13987 34333 -13789 34340 4 VDD
port 41 nsew
rlabel locali s -5093 34374 -4895 34379 4 VDD
port 41 nsew
rlabel locali s -4964 34379 -4895 34508 4 VDD
port 41 nsew
rlabel locali s -4964 34508 -4664 34531 4 VDD
port 41 nsew
rlabel locali s -7272 34364 -7153 34526 4 VDD
port 41 nsew
rlabel locali s -11729 34364 -11610 34526 4 VDD
port 41 nsew
rlabel locali s -13987 34340 -13606 34374 4 VDD
port 41 nsew
rlabel locali s -13987 34374 -13789 34379 4 VDD
port 41 nsew
rlabel locali s -5089 34531 -4664 34536 4 VDD
port 41 nsew
rlabel locali s -5276 34536 -4664 34570 4 VDD
port 41 nsew
rlabel locali s -7438 34526 -7153 34560 4 VDD
port 41 nsew
rlabel locali s -11729 34526 -11444 34560 4 VDD
port 41 nsew
rlabel locali s -13987 34379 -13918 34508 4 VDD
port 41 nsew
rlabel locali s -14218 33136 -14025 34508 4 VDD
port 41 nsew
rlabel locali s -14218 34508 -13918 34531 4 VDD
port 41 nsew
rlabel locali s -14218 34531 -13793 34536 4 VDD
port 41 nsew
rlabel locali s -5089 34570 -4664 34577 4 VDD
port 41 nsew
rlabel locali s -4964 34577 -4664 34644 4 VDD
port 41 nsew
rlabel locali s -5093 34644 -4664 34650 4 VDD
port 41 nsew
rlabel locali s -5276 34650 -4664 34684 4 VDD
port 41 nsew
rlabel locali s -5093 34684 -4664 34690 4 VDD
port 41 nsew
rlabel locali s -4964 34690 -4664 34840 4 VDD
port 41 nsew
rlabel locali s -7272 34560 -7153 34743 4 VDD
port 41 nsew
rlabel locali s -11729 34560 -11610 34743 4 VDD
port 41 nsew
rlabel locali s -14218 34536 -13606 34570 4 VDD
port 41 nsew
rlabel locali s -14218 34570 -13793 34577 4 VDD
port 41 nsew
rlabel locali s -14218 34577 -13918 34644 4 VDD
port 41 nsew
rlabel locali s -14218 34644 -13789 34650 4 VDD
port 41 nsew
rlabel locali s -14218 34650 -13606 34684 4 VDD
port 41 nsew
rlabel locali s -14218 34684 -13789 34690 4 VDD
port 41 nsew
rlabel locali s -7639 34743 -7153 34777 4 VDD
port 41 nsew
rlabel locali s -11729 34743 -11243 34777 4 VDD
port 41 nsew
rlabel locali s -5088 34840 -4664 34846 4 VDD
port 41 nsew
rlabel locali s -5276 34846 -4664 34880 4 VDD
port 41 nsew
rlabel locali s -5088 34880 -4664 34886 4 VDD
port 41 nsew
rlabel locali s -4964 34886 -4664 34953 4 VDD
port 41 nsew
rlabel locali s -7232 34777 -7153 34939 4 VDD
port 41 nsew
rlabel locali s -11729 34777 -11650 34939 4 VDD
port 41 nsew
rlabel locali s -14218 34690 -13918 34840 4 VDD
port 41 nsew
rlabel locali s -14218 34840 -13794 34846 4 VDD
port 41 nsew
rlabel locali s -14218 34846 -13606 34880 4 VDD
port 41 nsew
rlabel locali s -14218 34880 -13794 34886 4 VDD
port 41 nsew
rlabel locali s -5098 34953 -4664 34959 4 VDD
port 41 nsew
rlabel locali s -5276 34959 -4664 34993 4 VDD
port 41 nsew
rlabel locali s -7639 34939 -7153 34973 4 VDD
port 41 nsew
rlabel locali s -11729 34939 -11243 34973 4 VDD
port 41 nsew
rlabel locali s -14218 34886 -13918 34953 4 VDD
port 41 nsew
rlabel locali s -14218 34953 -13784 34959 4 VDD
port 41 nsew
rlabel locali s -5098 34993 -4664 34999 4 VDD
port 41 nsew
rlabel locali s -4964 34999 -4664 35101 4 VDD
port 41 nsew
rlabel locali s -7232 34973 -7153 35063 4 VDD
port 41 nsew
rlabel locali s -11729 34973 -11650 35063 4 VDD
port 41 nsew
rlabel locali s -14218 34959 -13606 34993 4 VDD
port 41 nsew
rlabel locali s -14218 34993 -13784 34999 4 VDD
port 41 nsew
rlabel locali s -4857 35101 -4664 36921 4 VDD
port 41 nsew
rlabel locali s -4964 35101 -4895 35150 4 VDD
port 41 nsew
rlabel locali s -7275 35063 -7139 35135 4 VDD
port 41 nsew
rlabel locali s -11743 35063 -11607 35135 4 VDD
port 41 nsew
rlabel locali s -5086 35150 -4895 35155 4 VDD
port 41 nsew
rlabel locali s -5276 35155 -4895 35189 4 VDD
port 41 nsew
rlabel locali s -7639 35135 -7139 35169 4 VDD
port 41 nsew
rlabel locali s -11743 35135 -11243 35169 4 VDD
port 41 nsew
rlabel locali s -14218 34999 -13918 35101 4 VDD
port 41 nsew
rlabel locali s -13987 35101 -13918 35150 4 VDD
port 41 nsew
rlabel locali s -13987 35150 -13796 35155 4 VDD
port 41 nsew
rlabel locali s -7275 35169 -7139 35186 4 VDD
port 41 nsew
rlabel locali s -11743 35169 -11607 35186 4 VDD
port 41 nsew
rlabel locali s -13987 35155 -13606 35189 4 VDD
port 41 nsew
rlabel locali s -5086 35189 -4895 35196 4 VDD
port 41 nsew
rlabel locali s -13987 35189 -13796 35196 4 VDD
port 41 nsew
rlabel locali s -7274 35452 -7138 35543 4 VDD
port 41 nsew
rlabel locali s -11744 35452 -11608 35543 4 VDD
port 41 nsew
rlabel locali s -7440 35543 -7138 35575 4 VDD
port 41 nsew
rlabel locali s -7440 35575 -7175 35577 4 VDD
port 41 nsew
rlabel locali s -11744 35543 -11442 35575 4 VDD
port 41 nsew
rlabel locali s -11707 35575 -11442 35577 4 VDD
port 41 nsew
rlabel locali s -7274 35577 -7175 35739 4 VDD
port 41 nsew
rlabel locali s -11707 35577 -11608 35739 4 VDD
port 41 nsew
rlabel locali s -7440 35739 -7175 35773 4 VDD
port 41 nsew
rlabel locali s -11707 35739 -11442 35773 4 VDD
port 41 nsew
rlabel locali s -7274 35773 -7175 35935 4 VDD
port 41 nsew
rlabel locali s -11707 35773 -11608 35935 4 VDD
port 41 nsew
rlabel locali s -7440 35935 -7175 35969 4 VDD
port 41 nsew
rlabel locali s -11707 35935 -11442 35969 4 VDD
port 41 nsew
rlabel locali s -7274 35969 -7175 36131 4 VDD
port 41 nsew
rlabel locali s -11707 35969 -11608 36131 4 VDD
port 41 nsew
rlabel locali s -7440 36131 -7175 36165 4 VDD
port 41 nsew
rlabel locali s -11707 36131 -11442 36165 4 VDD
port 41 nsew
rlabel locali s -7274 36165 -7175 36342 4 VDD
port 41 nsew
rlabel locali s -7274 36342 -7160 36348 4 VDD
port 41 nsew
rlabel locali s -11707 36165 -11608 36342 4 VDD
port 41 nsew
rlabel locali s -11722 36342 -11608 36348 4 VDD
port 41 nsew
rlabel locali s -7641 36348 -7160 36382 4 VDD
port 41 nsew
rlabel locali s -11722 36348 -11241 36382 4 VDD
port 41 nsew
rlabel locali s -7224 36382 -7160 36544 4 VDD
port 41 nsew
rlabel locali s -11722 36382 -11658 36544 4 VDD
port 41 nsew
rlabel locali s -7641 36544 -7160 36578 4 VDD
port 41 nsew
rlabel locali s -11722 36544 -11241 36578 4 VDD
port 41 nsew
rlabel locali s -5276 36644 -4895 36678 4 VDD
port 41 nsew
rlabel locali s -5093 36678 -4895 36684 4 VDD
port 41 nsew
rlabel locali s -7224 36578 -7160 36680 4 VDD
port 41 nsew
rlabel locali s -11722 36578 -11658 36680 4 VDD
port 41 nsew
rlabel locali s -13987 36644 -13606 36678 4 VDD
port 41 nsew
rlabel locali s -4964 36684 -4895 36833 4 VDD
port 41 nsew
rlabel locali s -7251 36680 -7115 36740 4 VDD
port 41 nsew
rlabel locali s -11767 36680 -11631 36740 4 VDD
port 41 nsew
rlabel locali s -13987 36678 -13789 36684 4 VDD
port 41 nsew
rlabel locali s -7641 36740 -7115 36774 4 VDD
port 41 nsew
rlabel locali s -11767 36740 -11241 36774 4 VDD
port 41 nsew
rlabel locali s -7251 36774 -7115 36803 4 VDD
port 41 nsew
rlabel locali s -11767 36774 -11631 36803 4 VDD
port 41 nsew
rlabel locali s -13987 36684 -13918 36833 4 VDD
port 41 nsew
rlabel locali s -5093 36833 -4895 36840 4 VDD
port 41 nsew
rlabel locali s -13987 36833 -13789 36840 4 VDD
port 41 nsew
rlabel locali s -5276 36840 -4895 36874 4 VDD
port 41 nsew
rlabel locali s -13987 36840 -13606 36874 4 VDD
port 41 nsew
rlabel locali s -5093 36874 -4895 36879 4 VDD
port 41 nsew
rlabel locali s -13987 36874 -13789 36879 4 VDD
port 41 nsew
rlabel locali s -4964 36879 -4895 36921 4 VDD
port 41 nsew
rlabel locali s -4964 36921 -4664 37031 4 VDD
port 41 nsew
rlabel locali s -13987 36879 -13918 36921 4 VDD
port 41 nsew
rlabel locali s -14218 35101 -14025 36921 4 VDD
port 41 nsew
rlabel locali s -14218 36921 -13918 37031 4 VDD
port 41 nsew
rlabel locali s -5089 37031 -4664 37036 4 VDD
port 41 nsew
rlabel locali s -14218 37031 -13793 37036 4 VDD
port 41 nsew
rlabel locali s -5276 37036 -4664 37070 4 VDD
port 41 nsew
rlabel locali s -14218 37036 -13606 37070 4 VDD
port 41 nsew
rlabel locali s -5089 37070 -4664 37077 4 VDD
port 41 nsew
rlabel locali s -14218 37070 -13793 37077 4 VDD
port 41 nsew
rlabel locali s -4964 37077 -4664 37144 4 VDD
port 41 nsew
rlabel locali s -5093 37144 -4664 37150 4 VDD
port 41 nsew
rlabel locali s -5276 37150 -4664 37184 4 VDD
port 41 nsew
rlabel locali s -7249 37081 -7113 37167 4 VDD
port 41 nsew
rlabel locali s -11769 37081 -11633 37167 4 VDD
port 41 nsew
rlabel locali s -14218 37077 -13918 37144 4 VDD
port 41 nsew
rlabel locali s -14218 37144 -13789 37150 4 VDD
port 41 nsew
rlabel locali s -5093 37184 -4664 37190 4 VDD
port 41 nsew
rlabel locali s -4964 37190 -4664 37340 4 VDD
port 41 nsew
rlabel locali s -7516 37167 -7113 37201 4 VDD
port 41 nsew
rlabel locali s -11769 37167 -11366 37201 4 VDD
port 41 nsew
rlabel locali s -14218 37150 -13606 37184 4 VDD
port 41 nsew
rlabel locali s -14218 37184 -13789 37190 4 VDD
port 41 nsew
rlabel locali s -7249 37201 -7113 37204 4 VDD
port 41 nsew
rlabel locali s -11769 37201 -11633 37204 4 VDD
port 41 nsew
rlabel locali s -5088 37340 -4664 37346 4 VDD
port 41 nsew
rlabel locali s -5276 37346 -4664 37380 4 VDD
port 41 nsew
rlabel locali s -7224 37204 -7146 37363 4 VDD
port 41 nsew
rlabel locali s -11736 37204 -11658 37363 4 VDD
port 41 nsew
rlabel locali s -14218 37190 -13918 37340 4 VDD
port 41 nsew
rlabel locali s -14218 37340 -13794 37346 4 VDD
port 41 nsew
rlabel locali s -5088 37380 -4664 37386 4 VDD
port 41 nsew
rlabel locali s -4964 37386 -4664 37453 4 VDD
port 41 nsew
rlabel locali s -7516 37363 -7146 37397 4 VDD
port 41 nsew
rlabel locali s -11736 37363 -11366 37397 4 VDD
port 41 nsew
rlabel locali s -14218 37346 -13606 37380 4 VDD
port 41 nsew
rlabel locali s -14218 37380 -13794 37386 4 VDD
port 41 nsew
rlabel locali s -7224 37397 -7146 37402 4 VDD
port 41 nsew
rlabel locali s -11736 37397 -11658 37402 4 VDD
port 41 nsew
rlabel locali s -5098 37453 -4664 37459 4 VDD
port 41 nsew
rlabel locali s -5276 37459 -4664 37493 4 VDD
port 41 nsew
rlabel locali s -5098 37493 -4664 37499 4 VDD
port 41 nsew
rlabel locali s -4964 37499 -4664 37514 4 VDD
port 41 nsew
rlabel locali s -3742 39356 -2527 39510 4 VDD
port 41 nsew
rlabel locali s -4857 37514 -4664 39510 4 VDD
port 41 nsew
rlabel locali s -4964 37514 -4895 37650 4 VDD
port 41 nsew
rlabel locali s -5086 37650 -4895 37655 4 VDD
port 41 nsew
rlabel locali s -5276 37655 -4895 37689 4 VDD
port 41 nsew
rlabel locali s -5086 37689 -4895 37696 4 VDD
port 41 nsew
rlabel locali s -7219 37402 -7146 37905 4 VDD
port 41 nsew
rlabel locali s -11736 37402 -11663 37905 4 VDD
port 41 nsew
rlabel locali s -14218 37386 -13918 37453 4 VDD
port 41 nsew
rlabel locali s -14218 37453 -13784 37459 4 VDD
port 41 nsew
rlabel locali s -14218 37459 -13606 37493 4 VDD
port 41 nsew
rlabel locali s -14218 37493 -13784 37499 4 VDD
port 41 nsew
rlabel locali s -14218 37499 -13918 37514 4 VDD
port 41 nsew
rlabel locali s -13987 37514 -13918 37650 4 VDD
port 41 nsew
rlabel locali s -13987 37650 -13796 37655 4 VDD
port 41 nsew
rlabel locali s -13987 37655 -13606 37689 4 VDD
port 41 nsew
rlabel locali s -13987 37689 -13796 37696 4 VDD
port 41 nsew
rlabel locali s -7516 37905 -7146 37939 4 VDD
port 41 nsew
rlabel locali s -11736 37905 -11366 37939 4 VDD
port 41 nsew
rlabel locali s -7220 37939 -7146 37977 4 VDD
port 41 nsew
rlabel locali s -7220 37977 -7151 38101 4 VDD
port 41 nsew
rlabel locali s -11736 37939 -11662 37977 4 VDD
port 41 nsew
rlabel locali s -11731 37977 -11662 38101 4 VDD
port 41 nsew
rlabel locali s -7516 38101 -7151 38135 4 VDD
port 41 nsew
rlabel locali s -11731 38101 -11366 38135 4 VDD
port 41 nsew
rlabel locali s -7220 38135 -7151 38297 4 VDD
port 41 nsew
rlabel locali s -11731 38135 -11662 38297 4 VDD
port 41 nsew
rlabel locali s -7516 38297 -7151 38331 4 VDD
port 41 nsew
rlabel locali s -11731 38297 -11366 38331 4 VDD
port 41 nsew
rlabel locali s -7220 38331 -7151 38437 4 VDD
port 41 nsew
rlabel locali s -11731 38331 -11662 38437 4 VDD
port 41 nsew
rlabel locali s -7254 38437 -7118 38493 4 VDD
port 41 nsew
rlabel locali s -11764 38437 -11628 38493 4 VDD
port 41 nsew
rlabel locali s -7516 38493 -7118 38527 4 VDD
port 41 nsew
rlabel locali s -11764 38493 -11366 38527 4 VDD
port 41 nsew
rlabel locali s -7254 38527 -7118 38560 4 VDD
port 41 nsew
rlabel locali s -11764 38527 -11628 38560 4 VDD
port 41 nsew
rlabel locali s -4857 39510 -2527 39644 4 VDD
port 41 nsew
rlabel locali s -14218 37514 -14025 39644 4 VDD
port 41 nsew
rlabel locali s -5276 39644 -2527 39678 4 VDD
port 41 nsew
rlabel locali s -7255 39653 -7119 39654 4 VDD
port 41 nsew
rlabel locali s -11763 39653 -11627 39654 4 VDD
port 41 nsew
rlabel locali s -5093 39678 -2527 39684 4 VDD
port 41 nsew
rlabel locali s -4964 39684 -2527 39833 4 VDD
port 41 nsew
rlabel locali s -7527 39654 -7119 39688 4 VDD
port 41 nsew
rlabel locali s -11763 39654 -11355 39688 4 VDD
port 41 nsew
rlabel locali s -14218 39644 -13606 39678 4 VDD
port 41 nsew
rlabel locali s -14218 39678 -13789 39684 4 VDD
port 41 nsew
rlabel locali s -7344 39688 -7119 39694 4 VDD
port 41 nsew
rlabel locali s -11763 39688 -11538 39694 4 VDD
port 41 nsew
rlabel locali s -7255 39694 -7119 39776 4 VDD
port 41 nsew
rlabel locali s -11763 39694 -11627 39776 4 VDD
port 41 nsew
rlabel locali s -5093 39833 -2527 39840 4 VDD
port 41 nsew
rlabel locali s -5276 39840 -2527 39874 4 VDD
port 41 nsew
rlabel locali s -7215 39776 -7146 39843 4 VDD
port 41 nsew
rlabel locali s -11736 39776 -11667 39843 4 VDD
port 41 nsew
rlabel locali s -14218 39684 -13918 39833 4 VDD
port 41 nsew
rlabel locali s -14218 39833 -13789 39840 4 VDD
port 41 nsew
rlabel locali s -7344 39843 -7146 39850 4 VDD
port 41 nsew
rlabel locali s -11736 39843 -11538 39850 4 VDD
port 41 nsew
rlabel locali s -5093 39874 -2527 39879 4 VDD
port 41 nsew
rlabel locali s -4964 39879 -2527 40031 4 VDD
port 41 nsew
rlabel locali s -7527 39850 -7146 39884 4 VDD
port 41 nsew
rlabel locali s -11736 39850 -11355 39884 4 VDD
port 41 nsew
rlabel locali s -14218 39840 -13606 39874 4 VDD
port 41 nsew
rlabel locali s -14218 39874 -13789 39879 4 VDD
port 41 nsew
rlabel locali s -7344 39884 -7146 39889 4 VDD
port 41 nsew
rlabel locali s -11736 39884 -11538 39889 4 VDD
port 41 nsew
rlabel locali s -5089 40031 -2527 40036 4 VDD
port 41 nsew
rlabel locali s -5276 40036 -2527 40070 4 VDD
port 41 nsew
rlabel locali s -7215 39889 -7146 40041 4 VDD
port 41 nsew
rlabel locali s -11736 39889 -11667 40041 4 VDD
port 41 nsew
rlabel locali s -14218 39879 -13918 40031 4 VDD
port 41 nsew
rlabel locali s -14218 40031 -13793 40036 4 VDD
port 41 nsew
rlabel locali s -7340 40041 -7146 40046 4 VDD
port 41 nsew
rlabel locali s -11736 40041 -11542 40046 4 VDD
port 41 nsew
rlabel locali s -5089 40070 -2527 40077 4 VDD
port 41 nsew
rlabel locali s -4964 40077 -2527 40144 4 VDD
port 41 nsew
rlabel locali s -7527 40046 -7146 40080 4 VDD
port 41 nsew
rlabel locali s -11736 40046 -11355 40080 4 VDD
port 41 nsew
rlabel locali s -14218 40036 -13606 40070 4 VDD
port 41 nsew
rlabel locali s -14218 40070 -13793 40077 4 VDD
port 41 nsew
rlabel locali s -7340 40080 -7146 40087 4 VDD
port 41 nsew
rlabel locali s -11736 40080 -11542 40087 4 VDD
port 41 nsew
rlabel locali s -5093 40144 -2527 40150 4 VDD
port 41 nsew
rlabel locali s -5276 40150 -2527 40184 4 VDD
port 41 nsew
rlabel locali s -7215 40087 -7146 40154 4 VDD
port 41 nsew
rlabel locali s -11736 40087 -11667 40154 4 VDD
port 41 nsew
rlabel locali s -14218 40077 -13918 40144 4 VDD
port 41 nsew
rlabel locali s -14218 40144 -13789 40150 4 VDD
port 41 nsew
rlabel locali s -7344 40154 -7146 40160 4 VDD
port 41 nsew
rlabel locali s -11736 40154 -11538 40160 4 VDD
port 41 nsew
rlabel locali s -5093 40184 -2527 40190 4 VDD
port 41 nsew
rlabel locali s -4964 40190 -2527 40272 4 VDD
port 41 nsew
rlabel locali s -3742 40272 -2527 40571 4 VDD
port 41 nsew
rlabel locali s -4964 40272 -4664 40340 4 VDD
port 41 nsew
rlabel locali s -7527 40160 -7146 40194 4 VDD
port 41 nsew
rlabel locali s -11736 40160 -11355 40194 4 VDD
port 41 nsew
rlabel locali s -14218 40150 -13606 40184 4 VDD
port 41 nsew
rlabel locali s -14218 40184 -13789 40190 4 VDD
port 41 nsew
rlabel locali s -7344 40194 -7146 40200 4 VDD
port 41 nsew
rlabel locali s -11736 40194 -11538 40200 4 VDD
port 41 nsew
rlabel locali s -5088 40340 -4664 40346 4 VDD
port 41 nsew
rlabel locali s -5276 40346 -4664 40380 4 VDD
port 41 nsew
rlabel locali s -7215 40200 -7146 40350 4 VDD
port 41 nsew
rlabel locali s -11736 40200 -11667 40350 4 VDD
port 41 nsew
rlabel locali s -14218 40190 -13918 40340 4 VDD
port 41 nsew
rlabel locali s -14218 40340 -13794 40346 4 VDD
port 41 nsew
rlabel locali s -7339 40350 -7146 40356 4 VDD
port 41 nsew
rlabel locali s -11736 40350 -11543 40356 4 VDD
port 41 nsew
rlabel locali s -5088 40380 -4664 40386 4 VDD
port 41 nsew
rlabel locali s -4964 40386 -4664 40453 4 VDD
port 41 nsew
rlabel locali s -7527 40356 -7146 40390 4 VDD
port 41 nsew
rlabel locali s -11736 40356 -11355 40390 4 VDD
port 41 nsew
rlabel locali s -14218 40346 -13606 40380 4 VDD
port 41 nsew
rlabel locali s -14218 40380 -13794 40386 4 VDD
port 41 nsew
rlabel locali s -7339 40390 -7146 40396 4 VDD
port 41 nsew
rlabel locali s -11736 40390 -11543 40396 4 VDD
port 41 nsew
rlabel locali s -5098 40453 -4664 40459 4 VDD
port 41 nsew
rlabel locali s -5276 40459 -4664 40493 4 VDD
port 41 nsew
rlabel locali s -7215 40396 -7146 40463 4 VDD
port 41 nsew
rlabel locali s -11736 40396 -11667 40463 4 VDD
port 41 nsew
rlabel locali s -14218 40386 -13918 40453 4 VDD
port 41 nsew
rlabel locali s -14218 40453 -13784 40459 4 VDD
port 41 nsew
rlabel locali s -7349 40463 -7146 40469 4 VDD
port 41 nsew
rlabel locali s -11736 40463 -11533 40469 4 VDD
port 41 nsew
rlabel locali s -5098 40493 -4664 40499 4 VDD
port 41 nsew
rlabel locali s -3510 40571 -2748 58538 4 VDD
port 41 nsew
rlabel locali s -4964 40499 -4664 40650 4 VDD
port 41 nsew
rlabel locali s -7527 40469 -7146 40503 4 VDD
port 41 nsew
rlabel locali s -11736 40469 -11355 40503 4 VDD
port 41 nsew
rlabel locali s -14218 40459 -13606 40493 4 VDD
port 41 nsew
rlabel locali s -14218 40493 -13784 40499 4 VDD
port 41 nsew
rlabel locali s -7349 40503 -7146 40509 4 VDD
port 41 nsew
rlabel locali s -11736 40503 -11533 40509 4 VDD
port 41 nsew
rlabel locali s -5086 40650 -4664 40655 4 VDD
port 41 nsew
rlabel locali s -5276 40655 -4664 40689 4 VDD
port 41 nsew
rlabel locali s -7215 40509 -7146 40660 4 VDD
port 41 nsew
rlabel locali s -11736 40509 -11667 40660 4 VDD
port 41 nsew
rlabel locali s -14218 40499 -13918 40650 4 VDD
port 41 nsew
rlabel locali s -14218 40650 -13796 40655 4 VDD
port 41 nsew
rlabel locali s -7337 40660 -7146 40665 4 VDD
port 41 nsew
rlabel locali s -11736 40660 -11545 40665 4 VDD
port 41 nsew
rlabel locali s -5086 40689 -4664 40696 4 VDD
port 41 nsew
rlabel locali s -4857 40696 -4664 40741 4 VDD
port 41 nsew
rlabel locali s -7527 40665 -7146 40699 4 VDD
port 41 nsew
rlabel locali s -11736 40665 -11355 40699 4 VDD
port 41 nsew
rlabel locali s -14218 40655 -13606 40689 4 VDD
port 41 nsew
rlabel locali s -14218 40689 -13796 40696 4 VDD
port 41 nsew
rlabel locali s -7337 40699 -7146 40706 4 VDD
port 41 nsew
rlabel locali s -11736 40699 -11545 40706 4 VDD
port 41 nsew
rlabel locali s -14218 40696 -14025 40741 4 VDD
port 41 nsew
rlabel locali s -12042 43876 -11974 43885 4 VDD
port 41 nsew
rlabel locali s -12333 43885 -11974 43919 4 VDD
port 41 nsew
rlabel locali s -12042 43919 -11974 44081 4 VDD
port 41 nsew
rlabel locali s -12333 44081 -11974 44115 4 VDD
port 41 nsew
rlabel locali s -12042 44115 -11974 44277 4 VDD
port 41 nsew
rlabel locali s -12333 44277 -11974 44311 4 VDD
port 41 nsew
rlabel locali s -12042 44311 -11974 44767 4 VDD
port 41 nsew
rlabel locali s -12333 44767 -11974 44801 4 VDD
port 41 nsew
rlabel locali s -12042 44801 -11974 44963 4 VDD
port 41 nsew
rlabel locali s -12333 44963 -11974 44997 4 VDD
port 41 nsew
rlabel locali s -12042 44997 -11974 45159 4 VDD
port 41 nsew
rlabel locali s -12333 45159 -11974 45193 4 VDD
port 41 nsew
rlabel locali s -12042 45193 -11974 45254 4 VDD
port 41 nsew
rlabel locali s -12037 45254 -11974 46188 4 VDD
port 41 nsew
rlabel locali s -13802 44758 -13739 45710 4 VDD
port 41 nsew
rlabel locali s -13802 45710 -13734 45771 4 VDD
port 41 nsew
rlabel locali s -13802 45771 -13443 45805 4 VDD
port 41 nsew
rlabel locali s -13802 45805 -13734 45967 4 VDD
port 41 nsew
rlabel locali s -13802 45967 -13443 46001 4 VDD
port 41 nsew
rlabel locali s -13802 46001 -13734 46163 4 VDD
port 41 nsew
rlabel locali s -12041 46188 -11973 46501 4 VDD
port 41 nsew
rlabel locali s -13802 46163 -13443 46197 4 VDD
port 41 nsew
rlabel locali s -12042 46501 -11973 46510 4 VDD
port 41 nsew
rlabel locali s -12333 46510 -11973 46544 4 VDD
port 41 nsew
rlabel locali s -12042 46544 -11973 46661 4 VDD
port 41 nsew
rlabel locali s -13802 46197 -13734 46608 4 VDD
port 41 nsew
rlabel locali s -13802 46608 -13443 46642 4 VDD
port 41 nsew
rlabel locali s -12042 46661 -11974 46706 4 VDD
port 41 nsew
rlabel locali s -12333 46706 -11974 46740 4 VDD
port 41 nsew
rlabel locali s -12042 46740 -11974 46902 4 VDD
port 41 nsew
rlabel locali s -13802 46642 -13734 46804 4 VDD
port 41 nsew
rlabel locali s -13802 46804 -13443 46838 4 VDD
port 41 nsew
rlabel locali s -12333 46902 -11974 46936 4 VDD
port 41 nsew
rlabel locali s -12042 46936 -11974 47467 4 VDD
port 41 nsew
rlabel locali s -13802 46838 -13734 47000 4 VDD
port 41 nsew
rlabel locali s -13802 47000 -13443 47034 4 VDD
port 41 nsew
rlabel locali s -12333 47467 -11974 47501 4 VDD
port 41 nsew
rlabel locali s -12042 47501 -11974 47663 4 VDD
port 41 nsew
rlabel locali s -13802 47034 -13734 47512 4 VDD
port 41 nsew
rlabel locali s -12333 47663 -11974 47697 4 VDD
port 41 nsew
rlabel locali s -12042 47697 -11974 47859 4 VDD
port 41 nsew
rlabel locali s -12333 47859 -11974 47893 4 VDD
port 41 nsew
rlabel locali s -12042 47893 -11974 47954 4 VDD
port 41 nsew
rlabel locali s -12037 47954 -11974 48879 4 VDD
port 41 nsew
rlabel locali s -13802 47512 -13739 48410 4 VDD
port 41 nsew
rlabel locali s -13802 48410 -13734 48471 4 VDD
port 41 nsew
rlabel locali s -13802 48471 -13443 48505 4 VDD
port 41 nsew
rlabel locali s -13802 48505 -13734 48667 4 VDD
port 41 nsew
rlabel locali s -13802 48667 -13443 48701 4 VDD
port 41 nsew
rlabel locali s -13802 48701 -13734 48863 4 VDD
port 41 nsew
rlabel locali s -12039 48879 -11971 49201 4 VDD
port 41 nsew
rlabel locali s -13802 48863 -13443 48897 4 VDD
port 41 nsew
rlabel locali s -12042 49201 -11971 49210 4 VDD
port 41 nsew
rlabel locali s -12333 49210 -11971 49244 4 VDD
port 41 nsew
rlabel locali s -12042 49244 -11971 49406 4 VDD
port 41 nsew
rlabel locali s -13802 48897 -13734 49308 4 VDD
port 41 nsew
rlabel locali s -13802 49308 -13443 49342 4 VDD
port 41 nsew
rlabel locali s -12333 49406 -11971 49440 4 VDD
port 41 nsew
rlabel locali s -12042 49440 -11971 49602 4 VDD
port 41 nsew
rlabel locali s -13802 49342 -13734 49504 4 VDD
port 41 nsew
rlabel locali s -13802 49504 -13443 49538 4 VDD
port 41 nsew
rlabel locali s -12333 49602 -11971 49636 4 VDD
port 41 nsew
rlabel locali s -12042 49636 -11971 49696 4 VDD
port 41 nsew
rlabel locali s -12039 49696 -11971 49857 4 VDD
port 41 nsew
rlabel locali s -13802 49538 -13734 49700 4 VDD
port 41 nsew
rlabel locali s -13802 49700 -13443 49734 4 VDD
port 41 nsew
rlabel locali s -12039 49857 -11431 49894 4 VDD
port 41 nsew
rlabel locali s -13802 49734 -13734 49894 4 VDD
port 41 nsew
rlabel locali s -13802 49894 -11431 49983 4 VDD
port 41 nsew
rlabel locali s -11500 49983 -11431 50680 4 VDD
port 41 nsew
rlabel locali s -9212 50683 -8967 50692 4 VDD
port 41 nsew
rlabel locali s -11500 50680 -11304 50687 4 VDD
port 41 nsew
rlabel locali s -9212 50692 -8367 50726 4 VDD
port 41 nsew
rlabel locali s -11500 50687 -10913 50721 4 VDD
port 41 nsew
rlabel locali s -9212 50726 -8967 50736 4 VDD
port 41 nsew
rlabel locali s -11500 50721 -11304 50728 4 VDD
port 41 nsew
rlabel locali s -9212 50736 -9079 50879 4 VDD
port 41 nsew
rlabel locali s -11500 50728 -11431 50877 4 VDD
port 41 nsew
rlabel locali s -9212 50879 -8951 50888 4 VDD
port 41 nsew
rlabel locali s -11500 50877 -11298 50883 4 VDD
port 41 nsew
rlabel locali s -9212 50888 -8367 50922 4 VDD
port 41 nsew
rlabel locali s -11500 50883 -10913 50917 4 VDD
port 41 nsew
rlabel locali s -9212 50922 -8951 50932 4 VDD
port 41 nsew
rlabel locali s -11500 50917 -11298 50925 4 VDD
port 41 nsew
rlabel locali s -9212 50932 -9079 51551 4 VDD
port 41 nsew
rlabel locali s -11500 50925 -11431 51626 4 VDD
port 41 nsew
rlabel locali s -11500 51626 -11304 51633 4 VDD
port 41 nsew
rlabel locali s -11500 51633 -10913 51667 4 VDD
port 41 nsew
rlabel locali s -11500 51667 -11304 51674 4 VDD
port 41 nsew
rlabel locali s -11500 51674 -11431 51823 4 VDD
port 41 nsew
rlabel locali s -11500 51823 -11298 51829 4 VDD
port 41 nsew
rlabel locali s -11500 51829 -10913 51863 4 VDD
port 41 nsew
rlabel locali s -11500 51863 -11298 51871 4 VDD
port 41 nsew
rlabel locali s -9246 52004 -9178 52013 4 VDD
port 41 nsew
rlabel locali s -9246 52013 -8887 52047 4 VDD
port 41 nsew
rlabel locali s -9246 52047 -9178 52209 4 VDD
port 41 nsew
rlabel locali s -9246 52209 -8887 52243 4 VDD
port 41 nsew
rlabel locali s -9246 52243 -9178 52405 4 VDD
port 41 nsew
rlabel locali s -11500 51871 -11431 52304 4 VDD
port 41 nsew
rlabel locali s -11516 52304 -11423 52390 4 VDD
port 41 nsew
rlabel locali s -9246 52405 -8887 52439 4 VDD
port 41 nsew
rlabel locali s -7481 52886 -7418 53838 4 VDD
port 41 nsew
rlabel locali s -9246 52439 -9178 52895 4 VDD
port 41 nsew
rlabel locali s -11512 52390 -11443 52549 4 VDD
port 41 nsew
rlabel locali s -11512 52549 -11147 52583 4 VDD
port 41 nsew
rlabel locali s -11512 52583 -11443 52745 4 VDD
port 41 nsew
rlabel locali s -11512 52745 -11147 52779 4 VDD
port 41 nsew
rlabel locali s -9246 52895 -8887 52929 4 VDD
port 41 nsew
rlabel locali s -9246 52929 -9178 53091 4 VDD
port 41 nsew
rlabel locali s -11512 52779 -11443 52941 4 VDD
port 41 nsew
rlabel locali s -11512 52941 -11147 52975 4 VDD
port 41 nsew
rlabel locali s -9246 53091 -8887 53125 4 VDD
port 41 nsew
rlabel locali s -9246 53125 -9178 53287 4 VDD
port 41 nsew
rlabel locali s -11512 52975 -11443 53137 4 VDD
port 41 nsew
rlabel locali s -11512 53137 -11147 53171 4 VDD
port 41 nsew
rlabel locali s -9246 53287 -8887 53321 4 VDD
port 41 nsew
rlabel locali s -9246 53321 -9178 53382 4 VDD
port 41 nsew
rlabel locali s -7486 53838 -7418 53899 4 VDD
port 41 nsew
rlabel locali s -7777 53899 -7418 53933 4 VDD
port 41 nsew
rlabel locali s -7486 53933 -7418 54095 4 VDD
port 41 nsew
rlabel locali s -7777 54095 -7418 54129 4 VDD
port 41 nsew
rlabel locali s -7486 54129 -7418 54291 4 VDD
port 41 nsew
rlabel locali s -7777 54291 -7418 54325 4 VDD
port 41 nsew
rlabel locali s -9246 53382 -9183 54316 4 VDD
port 41 nsew
rlabel locali s -11512 53171 -11443 53424 4 VDD
port 41 nsew
rlabel locali s -11523 53424 -11425 53487 4 VDD
port 41 nsew
rlabel locali s -11506 53487 -11439 53679 4 VDD
port 41 nsew
rlabel locali s -11506 53679 -11147 53713 4 VDD
port 41 nsew
rlabel locali s -11506 53713 -11439 53875 4 VDD
port 41 nsew
rlabel locali s -11506 53875 -11147 53909 4 VDD
port 41 nsew
rlabel locali s -11506 53909 -11439 54105 4 VDD
port 41 nsew
rlabel locali s -11512 54105 -11425 54179 4 VDD
port 41 nsew
rlabel locali s -7486 54325 -7418 54736 4 VDD
port 41 nsew
rlabel locali s -9247 54316 -9179 54506 4 VDD
port 41 nsew
rlabel locali s -11499 54179 -11431 54408 4 VDD
port 41 nsew
rlabel locali s -11499 54408 -11140 54442 4 VDD
port 41 nsew
rlabel locali s -9530 54448 -9466 54458 4 VDD
port 41 nsew
rlabel locali s -10047 54458 -9466 54492 4 VDD
port 41 nsew
rlabel locali s -9530 54492 -9466 54506 4 VDD
port 41 nsew
rlabel locali s -9530 54506 -9179 54629 4 VDD
port 41 nsew
rlabel locali s -11499 54442 -11431 54604 4 VDD
port 41 nsew
rlabel locali s -9530 54629 -9178 54638 4 VDD
port 41 nsew
rlabel locali s -11499 54604 -11140 54638 4 VDD
port 41 nsew
rlabel locali s -9530 54638 -8887 54654 4 VDD
port 41 nsew
rlabel locali s -10047 54654 -8887 54672 4 VDD
port 41 nsew
rlabel locali s -10047 54672 -9178 54688 4 VDD
port 41 nsew
rlabel locali s -7777 54736 -7418 54770 4 VDD
port 41 nsew
rlabel locali s -9530 54688 -9178 54738 4 VDD
port 41 nsew
rlabel locali s -7486 54770 -7418 54932 4 VDD
port 41 nsew
rlabel locali s -9247 54738 -9178 54789 4 VDD
port 41 nsew
rlabel locali s -9246 54789 -9178 54834 4 VDD
port 41 nsew
rlabel locali s -9246 54834 -8887 54868 4 VDD
port 41 nsew
rlabel locali s -7777 54932 -7418 54966 4 VDD
port 41 nsew
rlabel locali s -7486 54966 -7418 55128 4 VDD
port 41 nsew
rlabel locali s -9246 54868 -9178 55030 4 VDD
port 41 nsew
rlabel locali s -9530 54738 -9466 54850 4 VDD
port 41 nsew
rlabel locali s -11499 54638 -11431 54800 4 VDD
port 41 nsew
rlabel locali s -11499 54800 -11140 54822 4 VDD
port 41 nsew
rlabel locali s -11507 54822 -11140 54834 4 VDD
port 41 nsew
rlabel locali s -10047 54850 -9466 54884 4 VDD
port 41 nsew
rlabel locali s -9530 54884 -9466 54890 4 VDD
port 41 nsew
rlabel locali s -9246 55030 -8887 55064 4 VDD
port 41 nsew
rlabel locali s -7777 55128 -7418 55162 4 VDD
port 41 nsew
rlabel locali s -7486 55162 -7418 55640 4 VDD
port 41 nsew
rlabel locali s -9246 55064 -9178 55595 4 VDD
port 41 nsew
rlabel locali s -11507 54834 -11404 55288 4 VDD
port 41 nsew
rlabel locali s -11507 55288 -10569 55322 4 VDD
port 41 nsew
rlabel locali s -11507 55322 -11404 55484 4 VDD
port 41 nsew
rlabel locali s -11507 55484 -10569 55518 4 VDD
port 41 nsew
rlabel locali s -9246 55595 -8887 55629 4 VDD
port 41 nsew
rlabel locali s -7481 55640 -7418 56538 4 VDD
port 41 nsew
rlabel locali s -9246 55629 -9178 55791 4 VDD
port 41 nsew
rlabel locali s -11507 55518 -11404 55688 4 VDD
port 41 nsew
rlabel locali s -11507 55688 -10569 55722 4 VDD
port 41 nsew
rlabel locali s -9246 55791 -8887 55825 4 VDD
port 41 nsew
rlabel locali s -9246 55825 -9178 55987 4 VDD
port 41 nsew
rlabel locali s -11507 55722 -11404 55884 4 VDD
port 41 nsew
rlabel locali s -11507 55884 -10569 55918 4 VDD
port 41 nsew
rlabel locali s -9246 55987 -8887 56021 4 VDD
port 41 nsew
rlabel locali s -9246 56021 -9178 56082 4 VDD
port 41 nsew
rlabel locali s -7486 56538 -7418 56599 4 VDD
port 41 nsew
rlabel locali s -7777 56599 -7418 56633 4 VDD
port 41 nsew
rlabel locali s -7486 56633 -7418 56795 4 VDD
port 41 nsew
rlabel locali s -7777 56795 -7418 56829 4 VDD
port 41 nsew
rlabel locali s -7486 56829 -7418 56991 4 VDD
port 41 nsew
rlabel locali s -7777 56991 -7418 57025 4 VDD
port 41 nsew
rlabel locali s -9246 56082 -9183 57007 4 VDD
port 41 nsew
rlabel locali s -11507 55918 -11404 56288 4 VDD
port 41 nsew
rlabel locali s -11507 56288 -10569 56322 4 VDD
port 41 nsew
rlabel locali s -11507 56322 -11404 56484 4 VDD
port 41 nsew
rlabel locali s -11507 56484 -10569 56518 4 VDD
port 41 nsew
rlabel locali s -11507 56518 -11404 56688 4 VDD
port 41 nsew
rlabel locali s -11507 56688 -10569 56722 4 VDD
port 41 nsew
rlabel locali s -11507 56722 -11404 56884 4 VDD
port 41 nsew
rlabel locali s -11507 56884 -10569 56918 4 VDD
port 41 nsew
rlabel locali s -7486 57025 -7418 57436 4 VDD
port 41 nsew
rlabel locali s -9249 57007 -9181 57329 4 VDD
port 41 nsew
rlabel locali s -11507 56918 -11404 57288 4 VDD
port 41 nsew
rlabel locali s -11507 57288 -10569 57322 4 VDD
port 41 nsew
rlabel locali s -9249 57329 -9178 57338 4 VDD
port 41 nsew
rlabel locali s -9249 57338 -8887 57372 4 VDD
port 41 nsew
rlabel locali s -7777 57436 -7418 57470 4 VDD
port 41 nsew
rlabel locali s -7486 57470 -7418 57632 4 VDD
port 41 nsew
rlabel locali s -9249 57372 -9178 57534 4 VDD
port 41 nsew
rlabel locali s -11507 57322 -11404 57484 4 VDD
port 41 nsew
rlabel locali s -11507 57484 -10569 57518 4 VDD
port 41 nsew
rlabel locali s -9249 57534 -8887 57568 4 VDD
port 41 nsew
rlabel locali s -7777 57632 -7418 57666 4 VDD
port 41 nsew
rlabel locali s -7486 57666 -7418 57828 4 VDD
port 41 nsew
rlabel locali s -9249 57568 -9178 57730 4 VDD
port 41 nsew
rlabel locali s -11507 57518 -11404 57688 4 VDD
port 41 nsew
rlabel locali s -11507 57688 -10569 57722 4 VDD
port 41 nsew
rlabel locali s -9249 57730 -8887 57764 4 VDD
port 41 nsew
rlabel locali s -9249 57764 -9178 57824 4 VDD
port 41 nsew
rlabel locali s -7777 57828 -7418 57862 4 VDD
port 41 nsew
rlabel locali s -7486 57862 -7418 58022 4 VDD
port 41 nsew
rlabel locali s -9249 57824 -9181 58022 4 VDD
port 41 nsew
rlabel locali s -11507 57722 -11404 57884 4 VDD
port 41 nsew
rlabel locali s -11507 57884 -10569 57918 4 VDD
port 41 nsew
rlabel locali s -11507 57918 -11404 58022 4 VDD
port 41 nsew
rlabel locali s -11507 58022 -7418 58111 4 VDD
port 41 nsew
rlabel locali s -5019 58538 -2527 59641 4 VDD
port 41 nsew
rlabel locali s -3630 59641 -2527 119211 4 VDD
port 41 nsew
rlabel locali s -7840 58111 -7546 60223 4 VDD
port 41 nsew
rlabel locali s -7840 60223 -7482 60235 4 VDD
port 41 nsew
rlabel locali s -7924 60235 -7482 60271 4 VDD
port 41 nsew
rlabel locali s -7924 60271 -7216 60305 4 VDD
port 41 nsew
rlabel locali s -7924 60305 -7482 60467 4 VDD
port 41 nsew
rlabel locali s -7924 60467 -7216 60501 4 VDD
port 41 nsew
rlabel locali s -7924 60501 -7482 60577 4 VDD
port 41 nsew
rlabel locali s -7581 60577 -7482 60663 4 VDD
port 41 nsew
rlabel locali s -7581 60663 -7216 60697 4 VDD
port 41 nsew
rlabel locali s -7581 60697 -7482 60859 4 VDD
port 41 nsew
rlabel locali s -7581 60859 -7216 60893 4 VDD
port 41 nsew
rlabel locali s -7581 60893 -7482 60941 4 VDD
port 41 nsew
rlabel locali s -7924 60577 -7771 60637 4 VDD
port 41 nsew
rlabel locali s -8036 60235 -7972 60245 4 VDD
port 41 nsew
rlabel locali s -8453 60245 -7972 60279 4 VDD
port 41 nsew
rlabel locali s -11034 60215 -10935 60263 4 VDD
port 41 nsew
rlabel locali s -8036 60279 -7972 60441 4 VDD
port 41 nsew
rlabel locali s -11034 60263 -10669 60297 4 VDD
port 41 nsew
rlabel locali s -11034 60297 -10935 60397 4 VDD
port 41 nsew
rlabel locali s -11377 60227 -11224 60397 4 VDD
port 41 nsew
rlabel locali s -8453 60441 -7972 60475 4 VDD
port 41 nsew
rlabel locali s -11377 60397 -10935 60459 4 VDD
port 41 nsew
rlabel locali s -8036 60475 -7972 60637 4 VDD
port 41 nsew
rlabel locali s -11377 60459 -10669 60493 4 VDD
port 41 nsew
rlabel locali s -11377 60493 -10935 60569 4 VDD
port 41 nsew
rlabel locali s -7931 60637 -7771 60674 4 VDD
port 41 nsew
rlabel locali s -8453 60637 -7972 60671 4 VDD
port 41 nsew
rlabel locali s -11034 60569 -10935 60655 4 VDD
port 41 nsew
rlabel locali s -7938 60674 -7771 60863 4 VDD
port 41 nsew
rlabel locali s -8086 60671 -7972 60677 4 VDD
port 41 nsew
rlabel locali s -8086 60677 -7987 60854 4 VDD
port 41 nsew
rlabel locali s -11034 60655 -10669 60689 4 VDD
port 41 nsew
rlabel locali s -11034 60689 -10935 60851 4 VDD
port 41 nsew
rlabel locali s -7924 60863 -7771 61233 4 VDD
port 41 nsew
rlabel locali s -7924 61233 -7725 61234 4 VDD
port 41 nsew
rlabel locali s -7924 61234 -7662 61244 4 VDD
port 41 nsew
rlabel locali s -7924 61244 -7245 61278 4 VDD
port 41 nsew
rlabel locali s -7924 61278 -7662 61440 4 VDD
port 41 nsew
rlabel locali s -7924 61440 -7245 61474 4 VDD
port 41 nsew
rlabel locali s -7924 61474 -7662 61636 4 VDD
port 41 nsew
rlabel locali s -8252 60854 -7987 60888 4 VDD
port 41 nsew
rlabel locali s -11034 60851 -10669 60885 4 VDD
port 41 nsew
rlabel locali s -8086 60888 -7987 61050 4 VDD
port 41 nsew
rlabel locali s -11034 60885 -10935 60933 4 VDD
port 41 nsew
rlabel locali s -11377 60569 -11224 60629 4 VDD
port 41 nsew
rlabel locali s -11489 60227 -11425 60237 4 VDD
port 41 nsew
rlabel locali s -11906 60237 -11425 60271 4 VDD
port 41 nsew
rlabel locali s -11489 60271 -11425 60433 4 VDD
port 41 nsew
rlabel locali s -11906 60433 -11425 60467 4 VDD
port 41 nsew
rlabel locali s -11489 60467 -11425 60629 4 VDD
port 41 nsew
rlabel locali s -11384 60629 -11224 60666 4 VDD
port 41 nsew
rlabel locali s -11906 60629 -11425 60663 4 VDD
port 41 nsew
rlabel locali s -11391 60666 -11224 60855 4 VDD
port 41 nsew
rlabel locali s -11539 60663 -11425 60669 4 VDD
port 41 nsew
rlabel locali s -11539 60669 -11440 60846 4 VDD
port 41 nsew
rlabel locali s -8252 61050 -7987 61084 4 VDD
port 41 nsew
rlabel locali s -8086 61084 -7987 61246 4 VDD
port 41 nsew
rlabel locali s -11377 60855 -11224 61225 4 VDD
port 41 nsew
rlabel locali s -11377 61225 -11178 61226 4 VDD
port 41 nsew
rlabel locali s -11377 61226 -11115 61236 4 VDD
port 41 nsew
rlabel locali s -8252 61246 -7987 61280 4 VDD
port 41 nsew
rlabel locali s -11377 61236 -10698 61270 4 VDD
port 41 nsew
rlabel locali s -8086 61280 -7987 61442 4 VDD
port 41 nsew
rlabel locali s -11377 61270 -11115 61432 4 VDD
port 41 nsew
rlabel locali s -8252 61442 -7987 61476 4 VDD
port 41 nsew
rlabel locali s -11377 61432 -10698 61466 4 VDD
port 41 nsew
rlabel locali s -8086 61476 -7987 61524 4 VDD
port 41 nsew
rlabel locali s -11377 61466 -11115 61628 4 VDD
port 41 nsew
rlabel locali s -11705 60846 -11440 60880 4 VDD
port 41 nsew
rlabel locali s -11539 60880 -11440 61042 4 VDD
port 41 nsew
rlabel locali s -11705 61042 -11440 61076 4 VDD
port 41 nsew
rlabel locali s -11539 61076 -11440 61238 4 VDD
port 41 nsew
rlabel locali s -11705 61238 -11440 61272 4 VDD
port 41 nsew
rlabel locali s -11539 61272 -11440 61434 4 VDD
port 41 nsew
rlabel locali s -11705 61434 -11440 61468 4 VDD
port 41 nsew
rlabel locali s -11539 61468 -11440 61516 4 VDD
port 41 nsew
rlabel locali s -7924 61636 -7245 61670 4 VDD
port 41 nsew
rlabel locali s -11377 61628 -10698 61662 4 VDD
port 41 nsew
rlabel locali s -7924 61670 -7612 61676 4 VDD
port 41 nsew
rlabel locali s -7711 61676 -7612 61853 4 VDD
port 41 nsew
rlabel locali s -7924 61676 -7754 61681 4 VDD
port 41 nsew
rlabel locali s -11377 61662 -11065 61668 4 VDD
port 41 nsew
rlabel locali s -7948 61681 -7754 61687 4 VDD
port 41 nsew
rlabel locali s -8074 61687 -7754 61692 4 VDD
port 41 nsew
rlabel locali s -8664 61692 -7754 61726 4 VDD
port 41 nsew
rlabel locali s -8074 61726 -7754 61732 4 VDD
port 41 nsew
rlabel locali s -7948 61732 -7754 61851 4 VDD
port 41 nsew
rlabel locali s -11164 61668 -11065 61845 4 VDD
port 41 nsew
rlabel locali s -11377 61668 -11207 61673 4 VDD
port 41 nsew
rlabel locali s -11401 61673 -11207 61679 4 VDD
port 41 nsew
rlabel locali s -11527 61679 -11207 61684 4 VDD
port 41 nsew
rlabel locali s -12117 61684 -11207 61718 4 VDD
port 41 nsew
rlabel locali s -11527 61718 -11207 61724 4 VDD
port 41 nsew
rlabel locali s -11401 61724 -11207 61843 4 VDD
port 41 nsew
rlabel locali s -7711 61853 -7446 61887 4 VDD
port 41 nsew
rlabel locali s -7711 61887 -7612 62049 4 VDD
port 41 nsew
rlabel locali s -7711 62049 -7446 62083 4 VDD
port 41 nsew
rlabel locali s -7711 62083 -7612 62245 4 VDD
port 41 nsew
rlabel locali s -7711 62245 -7446 62279 4 VDD
port 41 nsew
rlabel locali s -7711 62279 -7612 62441 4 VDD
port 41 nsew
rlabel locali s -7948 61851 -7771 61882 4 VDD
port 41 nsew
rlabel locali s -11164 61845 -10899 61879 4 VDD
port 41 nsew
rlabel locali s -8071 61882 -7771 61888 4 VDD
port 41 nsew
rlabel locali s -8664 61888 -7771 61922 4 VDD
port 41 nsew
rlabel locali s -8071 61922 -7771 61927 4 VDD
port 41 nsew
rlabel locali s -7948 61927 -7771 62304 4 VDD
port 41 nsew
rlabel locali s -11164 61879 -11065 62041 4 VDD
port 41 nsew
rlabel locali s -11164 62041 -10899 62075 4 VDD
port 41 nsew
rlabel locali s -11164 62075 -11065 62237 4 VDD
port 41 nsew
rlabel locali s -11164 62237 -10899 62271 4 VDD
port 41 nsew
rlabel locali s -8072 62304 -7771 62311 4 VDD
port 41 nsew
rlabel locali s -8664 62311 -7771 62345 4 VDD
port 41 nsew
rlabel locali s -8072 62345 -7771 62346 4 VDD
port 41 nsew
rlabel locali s -7711 62441 -7446 62475 4 VDD
port 41 nsew
rlabel locali s -8072 62346 -7882 62349 4 VDD
port 41 nsew
rlabel locali s -7948 62349 -7882 62450 4 VDD
port 41 nsew
rlabel locali s -11164 62271 -11065 62433 4 VDD
port 41 nsew
rlabel locali s -11401 61843 -11224 61874 4 VDD
port 41 nsew
rlabel locali s -11524 61874 -11224 61880 4 VDD
port 41 nsew
rlabel locali s -12117 61880 -11224 61914 4 VDD
port 41 nsew
rlabel locali s -11524 61914 -11224 61919 4 VDD
port 41 nsew
rlabel locali s -11401 61919 -11224 62296 4 VDD
port 41 nsew
rlabel locali s -11525 62296 -11224 62303 4 VDD
port 41 nsew
rlabel locali s -12117 62303 -11224 62337 4 VDD
port 41 nsew
rlabel locali s -11525 62337 -11224 62338 4 VDD
port 41 nsew
rlabel locali s -7711 62475 -7612 62523 4 VDD
port 41 nsew
rlabel locali s -7941 62450 -7889 62523 4 VDD
port 41 nsew
rlabel locali s -11164 62433 -10899 62467 4 VDD
port 41 nsew
rlabel locali s -11525 62338 -11335 62341 4 VDD
port 41 nsew
rlabel locali s -11401 62341 -11335 62442 4 VDD
port 41 nsew
rlabel locali s -11164 62467 -11065 62515 4 VDD
port 41 nsew
rlabel locali s -7955 62523 -7861 62585 4 VDD
port 41 nsew
rlabel locali s -7967 62751 -7841 62849 4 VDD
port 41 nsew
rlabel locali s -11373 62741 -11260 62758 4 VDD
port 41 nsew
rlabel locali s -11373 62758 -9893 62824 4 VDD
port 41 nsew
rlabel locali s -7961 62849 -7844 63314 4 VDD
port 41 nsew
rlabel locali s -9959 62824 -9893 63094 4 VDD
port 41 nsew
rlabel locali s -11373 62824 -11260 62825 4 VDD
port 41 nsew
rlabel locali s -11355 63094 -9893 63160 4 VDD
port 41 nsew
rlabel locali s -7961 63314 -7717 63431 4 VDD
port 41 nsew
rlabel locali s -7834 63431 -7717 63681 4 VDD
port 41 nsew
rlabel locali s -7929 63681 -7647 63684 4 VDD
port 41 nsew
rlabel locali s -8422 63684 -7647 63718 4 VDD
port 41 nsew
rlabel locali s -7929 63718 -7647 63719 4 VDD
port 41 nsew
rlabel locali s -7770 63719 -7647 63878 4 VDD
port 41 nsew
rlabel locali s -7927 63878 -7647 63880 4 VDD
port 41 nsew
rlabel locali s -8422 63880 -7647 63914 4 VDD
port 41 nsew
rlabel locali s -7927 63914 -7647 63916 4 VDD
port 41 nsew
rlabel locali s -7770 63916 -7647 64470 4 VDD
port 41 nsew
rlabel locali s -11065 63883 -10966 63931 4 VDD
port 41 nsew
rlabel locali s -11355 63160 -11289 63895 4 VDD
port 41 nsew
rlabel locali s -11065 63931 -10700 63965 4 VDD
port 41 nsew
rlabel locali s -11065 63965 -10966 64065 4 VDD
port 41 nsew
rlabel locali s -11408 63895 -11255 64065 4 VDD
port 41 nsew
rlabel locali s -11408 64065 -10966 64127 4 VDD
port 41 nsew
rlabel locali s -11408 64127 -10700 64161 4 VDD
port 41 nsew
rlabel locali s -11408 64161 -10966 64237 4 VDD
port 41 nsew
rlabel locali s -11065 64237 -10966 64323 4 VDD
port 41 nsew
rlabel locali s -11065 64323 -10700 64357 4 VDD
port 41 nsew
rlabel locali s -7950 64470 -7647 64475 4 VDD
port 41 nsew
rlabel locali s -8422 64475 -7647 64509 4 VDD
port 41 nsew
rlabel locali s -7950 64509 -7647 64520 4 VDD
port 41 nsew
rlabel locali s -11065 64357 -10966 64519 4 VDD
port 41 nsew
rlabel locali s -7770 64520 -7647 64596 4 VDD
port 41 nsew
rlabel locali s -11065 64519 -10700 64553 4 VDD
port 41 nsew
rlabel locali s -7947 64596 -7647 64605 4 VDD
port 41 nsew
rlabel locali s -11065 64553 -10966 64601 4 VDD
port 41 nsew
rlabel locali s -11408 64237 -11255 64297 4 VDD
port 41 nsew
rlabel locali s -11520 63895 -11456 63905 4 VDD
port 41 nsew
rlabel locali s -11937 63905 -11456 63939 4 VDD
port 41 nsew
rlabel locali s -11520 63939 -11456 64101 4 VDD
port 41 nsew
rlabel locali s -11937 64101 -11456 64135 4 VDD
port 41 nsew
rlabel locali s -11520 64135 -11456 64297 4 VDD
port 41 nsew
rlabel locali s -11415 64297 -11255 64334 4 VDD
port 41 nsew
rlabel locali s -11937 64297 -11456 64331 4 VDD
port 41 nsew
rlabel locali s -11422 64334 -11255 64523 4 VDD
port 41 nsew
rlabel locali s -11570 64331 -11456 64337 4 VDD
port 41 nsew
rlabel locali s -11570 64337 -11471 64514 4 VDD
port 41 nsew
rlabel locali s -8422 64605 -7647 64639 4 VDD
port 41 nsew
rlabel locali s -7947 64639 -7647 64646 4 VDD
port 41 nsew
rlabel locali s -7770 64646 -7647 64827 4 VDD
port 41 nsew
rlabel locali s -7932 64827 -7647 64833 4 VDD
port 41 nsew
rlabel locali s -8222 64833 -7647 64867 4 VDD
port 41 nsew
rlabel locali s -7932 64867 -7647 64870 4 VDD
port 41 nsew
rlabel locali s -7770 64870 -7647 65024 4 VDD
port 41 nsew
rlabel locali s -11408 64523 -11255 64893 4 VDD
port 41 nsew
rlabel locali s -11408 64893 -11209 64894 4 VDD
port 41 nsew
rlabel locali s -11408 64894 -11146 64904 4 VDD
port 41 nsew
rlabel locali s -11408 64904 -10729 64938 4 VDD
port 41 nsew
rlabel locali s -7930 65024 -7647 65029 4 VDD
port 41 nsew
rlabel locali s -8222 65029 -7647 65063 4 VDD
port 41 nsew
rlabel locali s -7930 65063 -7647 65067 4 VDD
port 41 nsew
rlabel locali s -7769 65067 -7647 65991 4 VDD
port 41 nsew
rlabel locali s -11408 64938 -11146 65100 4 VDD
port 41 nsew
rlabel locali s -11408 65100 -10729 65134 4 VDD
port 41 nsew
rlabel locali s -11408 65134 -11146 65296 4 VDD
port 41 nsew
rlabel locali s -11736 64514 -11471 64548 4 VDD
port 41 nsew
rlabel locali s -11570 64548 -11471 64710 4 VDD
port 41 nsew
rlabel locali s -11736 64710 -11471 64744 4 VDD
port 41 nsew
rlabel locali s -11570 64744 -11471 64906 4 VDD
port 41 nsew
rlabel locali s -11736 64906 -11471 64940 4 VDD
port 41 nsew
rlabel locali s -11570 64940 -11471 65102 4 VDD
port 41 nsew
rlabel locali s -11736 65102 -11471 65136 4 VDD
port 41 nsew
rlabel locali s -11570 65136 -11471 65184 4 VDD
port 41 nsew
rlabel locali s -11408 65296 -10729 65330 4 VDD
port 41 nsew
rlabel locali s -11408 65330 -11096 65336 4 VDD
port 41 nsew
rlabel locali s -11195 65336 -11096 65513 4 VDD
port 41 nsew
rlabel locali s -11408 65336 -11238 65341 4 VDD
port 41 nsew
rlabel locali s -11432 65341 -11238 65347 4 VDD
port 41 nsew
rlabel locali s -11558 65347 -11238 65352 4 VDD
port 41 nsew
rlabel locali s -12148 65352 -11238 65386 4 VDD
port 41 nsew
rlabel locali s -11558 65386 -11238 65392 4 VDD
port 41 nsew
rlabel locali s -11432 65392 -11238 65511 4 VDD
port 41 nsew
rlabel locali s -11195 65513 -10930 65547 4 VDD
port 41 nsew
rlabel locali s -11195 65547 -11096 65709 4 VDD
port 41 nsew
rlabel locali s -11195 65709 -10930 65743 4 VDD
port 41 nsew
rlabel locali s -11195 65743 -11096 65905 4 VDD
port 41 nsew
rlabel locali s -11195 65905 -10930 65939 4 VDD
port 41 nsew
rlabel locali s -10288 65991 -7647 66113 4 VDD
port 41 nsew
rlabel locali s -11195 65939 -11096 66101 4 VDD
port 41 nsew
rlabel locali s -11432 65511 -11255 65542 4 VDD
port 41 nsew
rlabel locali s -11555 65542 -11255 65548 4 VDD
port 41 nsew
rlabel locali s -12148 65548 -11255 65582 4 VDD
port 41 nsew
rlabel locali s -11555 65582 -11255 65587 4 VDD
port 41 nsew
rlabel locali s -11432 65587 -11255 65964 4 VDD
port 41 nsew
rlabel locali s -11556 65964 -11255 65971 4 VDD
port 41 nsew
rlabel locali s -12148 65971 -11255 66005 4 VDD
port 41 nsew
rlabel locali s -11556 66005 -11255 66006 4 VDD
port 41 nsew
rlabel locali s -11556 66006 -11366 66009 4 VDD
port 41 nsew
rlabel locali s -11432 66009 -11366 66061 4 VDD
port 41 nsew
rlabel locali s -7592 68663 -7493 68711 4 VDD
port 41 nsew
rlabel locali s -7592 68711 -7227 68745 4 VDD
port 41 nsew
rlabel locali s -7592 68745 -7493 68845 4 VDD
port 41 nsew
rlabel locali s -7935 66113 -7782 68845 4 VDD
port 41 nsew
rlabel locali s -10288 66113 -10166 66501 4 VDD
port 41 nsew
rlabel locali s -11195 66101 -10930 66135 4 VDD
port 41 nsew
rlabel locali s -11195 66135 -11096 66183 4 VDD
port 41 nsew
rlabel locali s -11432 66061 -11330 66110 4 VDD
port 41 nsew
rlabel locali s -11413 66110 -11330 66161 4 VDD
port 41 nsew
rlabel locali s -11438 66161 -11299 66240 4 VDD
port 41 nsew
rlabel locali s -11451 66411 -11284 66501 4 VDD
port 41 nsew
rlabel locali s -11451 66501 -10166 66550 4 VDD
port 41 nsew
rlabel locali s -11423 66550 -10166 66623 4 VDD
port 41 nsew
rlabel locali s -7935 68845 -7493 68907 4 VDD
port 41 nsew
rlabel locali s -7935 68907 -7227 68941 4 VDD
port 41 nsew
rlabel locali s -7935 68941 -7493 69017 4 VDD
port 41 nsew
rlabel locali s -7592 69017 -7493 69103 4 VDD
port 41 nsew
rlabel locali s -7592 69103 -7227 69137 4 VDD
port 41 nsew
rlabel locali s -7592 69137 -7493 69299 4 VDD
port 41 nsew
rlabel locali s -7592 69299 -7227 69333 4 VDD
port 41 nsew
rlabel locali s -7592 69333 -7493 69381 4 VDD
port 41 nsew
rlabel locali s -7935 69017 -7782 69077 4 VDD
port 41 nsew
rlabel locali s -8047 68675 -7983 68685 4 VDD
port 41 nsew
rlabel locali s -8464 68685 -7983 68719 4 VDD
port 41 nsew
rlabel locali s -11045 68655 -10946 68703 4 VDD
port 41 nsew
rlabel locali s -8047 68719 -7983 68881 4 VDD
port 41 nsew
rlabel locali s -11045 68703 -10680 68737 4 VDD
port 41 nsew
rlabel locali s -11045 68737 -10946 68837 4 VDD
port 41 nsew
rlabel locali s -11388 68667 -11235 68837 4 VDD
port 41 nsew
rlabel locali s -8464 68881 -7983 68915 4 VDD
port 41 nsew
rlabel locali s -11388 68837 -10946 68899 4 VDD
port 41 nsew
rlabel locali s -8047 68915 -7983 69077 4 VDD
port 41 nsew
rlabel locali s -11388 68899 -10680 68933 4 VDD
port 41 nsew
rlabel locali s -11388 68933 -10946 69009 4 VDD
port 41 nsew
rlabel locali s -7942 69077 -7782 69114 4 VDD
port 41 nsew
rlabel locali s -8464 69077 -7983 69111 4 VDD
port 41 nsew
rlabel locali s -11045 69009 -10946 69095 4 VDD
port 41 nsew
rlabel locali s -7949 69114 -7782 69303 4 VDD
port 41 nsew
rlabel locali s -8097 69111 -7983 69117 4 VDD
port 41 nsew
rlabel locali s -8097 69117 -7998 69294 4 VDD
port 41 nsew
rlabel locali s -11045 69095 -10680 69129 4 VDD
port 41 nsew
rlabel locali s -11045 69129 -10946 69291 4 VDD
port 41 nsew
rlabel locali s -7935 69303 -7782 69673 4 VDD
port 41 nsew
rlabel locali s -7935 69673 -7736 69674 4 VDD
port 41 nsew
rlabel locali s -7935 69674 -7673 69684 4 VDD
port 41 nsew
rlabel locali s -7935 69684 -7256 69718 4 VDD
port 41 nsew
rlabel locali s -7935 69718 -7673 69880 4 VDD
port 41 nsew
rlabel locali s -7935 69880 -7256 69914 4 VDD
port 41 nsew
rlabel locali s -7935 69914 -7673 70076 4 VDD
port 41 nsew
rlabel locali s -8263 69294 -7998 69328 4 VDD
port 41 nsew
rlabel locali s -11045 69291 -10680 69325 4 VDD
port 41 nsew
rlabel locali s -8097 69328 -7998 69490 4 VDD
port 41 nsew
rlabel locali s -11045 69325 -10946 69373 4 VDD
port 41 nsew
rlabel locali s -11388 69009 -11235 69069 4 VDD
port 41 nsew
rlabel locali s -11500 68667 -11436 68677 4 VDD
port 41 nsew
rlabel locali s -11917 68677 -11436 68711 4 VDD
port 41 nsew
rlabel locali s -11500 68711 -11436 68873 4 VDD
port 41 nsew
rlabel locali s -11917 68873 -11436 68907 4 VDD
port 41 nsew
rlabel locali s -11500 68907 -11436 69069 4 VDD
port 41 nsew
rlabel locali s -11395 69069 -11235 69106 4 VDD
port 41 nsew
rlabel locali s -11917 69069 -11436 69103 4 VDD
port 41 nsew
rlabel locali s -11402 69106 -11235 69295 4 VDD
port 41 nsew
rlabel locali s -11550 69103 -11436 69109 4 VDD
port 41 nsew
rlabel locali s -11550 69109 -11451 69286 4 VDD
port 41 nsew
rlabel locali s -8263 69490 -7998 69524 4 VDD
port 41 nsew
rlabel locali s -8097 69524 -7998 69686 4 VDD
port 41 nsew
rlabel locali s -11388 69295 -11235 69665 4 VDD
port 41 nsew
rlabel locali s -11388 69665 -11189 69666 4 VDD
port 41 nsew
rlabel locali s -11388 69666 -11126 69676 4 VDD
port 41 nsew
rlabel locali s -8263 69686 -7998 69720 4 VDD
port 41 nsew
rlabel locali s -11388 69676 -10709 69710 4 VDD
port 41 nsew
rlabel locali s -8097 69720 -7998 69882 4 VDD
port 41 nsew
rlabel locali s -11388 69710 -11126 69872 4 VDD
port 41 nsew
rlabel locali s -8263 69882 -7998 69916 4 VDD
port 41 nsew
rlabel locali s -11388 69872 -10709 69906 4 VDD
port 41 nsew
rlabel locali s -8097 69916 -7998 69964 4 VDD
port 41 nsew
rlabel locali s -11388 69906 -11126 70068 4 VDD
port 41 nsew
rlabel locali s -11716 69286 -11451 69320 4 VDD
port 41 nsew
rlabel locali s -11550 69320 -11451 69482 4 VDD
port 41 nsew
rlabel locali s -11716 69482 -11451 69516 4 VDD
port 41 nsew
rlabel locali s -11550 69516 -11451 69678 4 VDD
port 41 nsew
rlabel locali s -11716 69678 -11451 69712 4 VDD
port 41 nsew
rlabel locali s -11550 69712 -11451 69874 4 VDD
port 41 nsew
rlabel locali s -11716 69874 -11451 69908 4 VDD
port 41 nsew
rlabel locali s -11550 69908 -11451 69956 4 VDD
port 41 nsew
rlabel locali s -7935 70076 -7256 70110 4 VDD
port 41 nsew
rlabel locali s -11388 70068 -10709 70102 4 VDD
port 41 nsew
rlabel locali s -7935 70110 -7623 70116 4 VDD
port 41 nsew
rlabel locali s -7722 70116 -7623 70293 4 VDD
port 41 nsew
rlabel locali s -7935 70116 -7765 70121 4 VDD
port 41 nsew
rlabel locali s -11388 70102 -11076 70108 4 VDD
port 41 nsew
rlabel locali s -7959 70121 -7765 70127 4 VDD
port 41 nsew
rlabel locali s -8085 70127 -7765 70132 4 VDD
port 41 nsew
rlabel locali s -8675 70132 -7765 70166 4 VDD
port 41 nsew
rlabel locali s -8085 70166 -7765 70172 4 VDD
port 41 nsew
rlabel locali s -7959 70172 -7765 70291 4 VDD
port 41 nsew
rlabel locali s -11175 70108 -11076 70285 4 VDD
port 41 nsew
rlabel locali s -11388 70108 -11218 70113 4 VDD
port 41 nsew
rlabel locali s -11412 70113 -11218 70119 4 VDD
port 41 nsew
rlabel locali s -11538 70119 -11218 70124 4 VDD
port 41 nsew
rlabel locali s -12128 70124 -11218 70158 4 VDD
port 41 nsew
rlabel locali s -11538 70158 -11218 70164 4 VDD
port 41 nsew
rlabel locali s -11412 70164 -11218 70283 4 VDD
port 41 nsew
rlabel locali s -7722 70293 -7457 70327 4 VDD
port 41 nsew
rlabel locali s -7722 70327 -7623 70489 4 VDD
port 41 nsew
rlabel locali s -7722 70489 -7457 70523 4 VDD
port 41 nsew
rlabel locali s -7722 70523 -7623 70685 4 VDD
port 41 nsew
rlabel locali s -7722 70685 -7457 70719 4 VDD
port 41 nsew
rlabel locali s -7722 70719 -7623 70881 4 VDD
port 41 nsew
rlabel locali s -7959 70291 -7782 70322 4 VDD
port 41 nsew
rlabel locali s -11175 70285 -10910 70319 4 VDD
port 41 nsew
rlabel locali s -8082 70322 -7782 70328 4 VDD
port 41 nsew
rlabel locali s -8675 70328 -7782 70362 4 VDD
port 41 nsew
rlabel locali s -8082 70362 -7782 70367 4 VDD
port 41 nsew
rlabel locali s -7959 70367 -7782 70744 4 VDD
port 41 nsew
rlabel locali s -11175 70319 -11076 70481 4 VDD
port 41 nsew
rlabel locali s -11175 70481 -10910 70515 4 VDD
port 41 nsew
rlabel locali s -11175 70515 -11076 70677 4 VDD
port 41 nsew
rlabel locali s -11175 70677 -10910 70711 4 VDD
port 41 nsew
rlabel locali s -8083 70744 -7782 70751 4 VDD
port 41 nsew
rlabel locali s -8675 70751 -7782 70785 4 VDD
port 41 nsew
rlabel locali s -8083 70785 -7782 70786 4 VDD
port 41 nsew
rlabel locali s -7722 70881 -7457 70915 4 VDD
port 41 nsew
rlabel locali s -8083 70786 -7893 70789 4 VDD
port 41 nsew
rlabel locali s -7959 70789 -7893 70890 4 VDD
port 41 nsew
rlabel locali s -11175 70711 -11076 70873 4 VDD
port 41 nsew
rlabel locali s -11412 70283 -11235 70314 4 VDD
port 41 nsew
rlabel locali s -11535 70314 -11235 70320 4 VDD
port 41 nsew
rlabel locali s -12128 70320 -11235 70354 4 VDD
port 41 nsew
rlabel locali s -11535 70354 -11235 70359 4 VDD
port 41 nsew
rlabel locali s -11412 70359 -11235 70736 4 VDD
port 41 nsew
rlabel locali s -11536 70736 -11235 70743 4 VDD
port 41 nsew
rlabel locali s -12128 70743 -11235 70777 4 VDD
port 41 nsew
rlabel locali s -11536 70777 -11235 70778 4 VDD
port 41 nsew
rlabel locali s -7722 70915 -7623 70963 4 VDD
port 41 nsew
rlabel locali s -7952 70890 -7900 70963 4 VDD
port 41 nsew
rlabel locali s -11175 70873 -10910 70907 4 VDD
port 41 nsew
rlabel locali s -11536 70778 -11346 70781 4 VDD
port 41 nsew
rlabel locali s -11412 70781 -11346 70882 4 VDD
port 41 nsew
rlabel locali s -11175 70907 -11076 70955 4 VDD
port 41 nsew
rlabel locali s -7966 70963 -7872 71025 4 VDD
port 41 nsew
rlabel locali s -7978 71191 -7852 71289 4 VDD
port 41 nsew
rlabel locali s -11384 71181 -11271 71198 4 VDD
port 41 nsew
rlabel locali s -11384 71198 -9904 71264 4 VDD
port 41 nsew
rlabel locali s -7972 71289 -7855 71754 4 VDD
port 41 nsew
rlabel locali s -9970 71264 -9904 71534 4 VDD
port 41 nsew
rlabel locali s -11384 71264 -11271 71265 4 VDD
port 41 nsew
rlabel locali s -11366 71534 -9904 71600 4 VDD
port 41 nsew
rlabel locali s -7972 71754 -7728 71871 4 VDD
port 41 nsew
rlabel locali s -7845 71871 -7728 72121 4 VDD
port 41 nsew
rlabel locali s -7940 72121 -7658 72124 4 VDD
port 41 nsew
rlabel locali s -8433 72124 -7658 72158 4 VDD
port 41 nsew
rlabel locali s -7940 72158 -7658 72159 4 VDD
port 41 nsew
rlabel locali s -7781 72159 -7658 72318 4 VDD
port 41 nsew
rlabel locali s -7938 72318 -7658 72320 4 VDD
port 41 nsew
rlabel locali s -8433 72320 -7658 72354 4 VDD
port 41 nsew
rlabel locali s -7938 72354 -7658 72356 4 VDD
port 41 nsew
rlabel locali s -7781 72356 -7658 72910 4 VDD
port 41 nsew
rlabel locali s -11076 72323 -10977 72371 4 VDD
port 41 nsew
rlabel locali s -11366 71600 -11300 72335 4 VDD
port 41 nsew
rlabel locali s -11076 72371 -10711 72405 4 VDD
port 41 nsew
rlabel locali s -11076 72405 -10977 72505 4 VDD
port 41 nsew
rlabel locali s -11419 72335 -11266 72505 4 VDD
port 41 nsew
rlabel locali s -11419 72505 -10977 72567 4 VDD
port 41 nsew
rlabel locali s -11419 72567 -10711 72601 4 VDD
port 41 nsew
rlabel locali s -11419 72601 -10977 72677 4 VDD
port 41 nsew
rlabel locali s -11076 72677 -10977 72763 4 VDD
port 41 nsew
rlabel locali s -11076 72763 -10711 72797 4 VDD
port 41 nsew
rlabel locali s -7961 72910 -7658 72915 4 VDD
port 41 nsew
rlabel locali s -8433 72915 -7658 72949 4 VDD
port 41 nsew
rlabel locali s -7961 72949 -7658 72960 4 VDD
port 41 nsew
rlabel locali s -11076 72797 -10977 72959 4 VDD
port 41 nsew
rlabel locali s -7781 72960 -7658 73036 4 VDD
port 41 nsew
rlabel locali s -11076 72959 -10711 72993 4 VDD
port 41 nsew
rlabel locali s -7958 73036 -7658 73045 4 VDD
port 41 nsew
rlabel locali s -11076 72993 -10977 73041 4 VDD
port 41 nsew
rlabel locali s -11419 72677 -11266 72737 4 VDD
port 41 nsew
rlabel locali s -11531 72335 -11467 72345 4 VDD
port 41 nsew
rlabel locali s -11948 72345 -11467 72379 4 VDD
port 41 nsew
rlabel locali s -11531 72379 -11467 72541 4 VDD
port 41 nsew
rlabel locali s -11948 72541 -11467 72575 4 VDD
port 41 nsew
rlabel locali s -11531 72575 -11467 72737 4 VDD
port 41 nsew
rlabel locali s -11426 72737 -11266 72774 4 VDD
port 41 nsew
rlabel locali s -11948 72737 -11467 72771 4 VDD
port 41 nsew
rlabel locali s -11433 72774 -11266 72963 4 VDD
port 41 nsew
rlabel locali s -11581 72771 -11467 72777 4 VDD
port 41 nsew
rlabel locali s -11581 72777 -11482 72954 4 VDD
port 41 nsew
rlabel locali s -8433 73045 -7658 73079 4 VDD
port 41 nsew
rlabel locali s -7958 73079 -7658 73086 4 VDD
port 41 nsew
rlabel locali s -7781 73086 -7658 73267 4 VDD
port 41 nsew
rlabel locali s -7943 73267 -7658 73273 4 VDD
port 41 nsew
rlabel locali s -8233 73273 -7658 73307 4 VDD
port 41 nsew
rlabel locali s -7943 73307 -7658 73310 4 VDD
port 41 nsew
rlabel locali s -7781 73310 -7658 73464 4 VDD
port 41 nsew
rlabel locali s -11419 72963 -11266 73333 4 VDD
port 41 nsew
rlabel locali s -11419 73333 -11220 73334 4 VDD
port 41 nsew
rlabel locali s -11419 73334 -11157 73344 4 VDD
port 41 nsew
rlabel locali s -11419 73344 -10740 73378 4 VDD
port 41 nsew
rlabel locali s -7941 73464 -7658 73469 4 VDD
port 41 nsew
rlabel locali s -8233 73469 -7658 73493 4 VDD
port 41 nsew
rlabel locali s -8233 73493 -7616 73503 4 VDD
port 41 nsew
rlabel locali s -7941 73503 -7616 73507 4 VDD
port 41 nsew
rlabel locali s -7870 73507 -7616 74431 4 VDD
port 41 nsew
rlabel locali s -11419 73378 -11157 73540 4 VDD
port 41 nsew
rlabel locali s -11419 73540 -10740 73574 4 VDD
port 41 nsew
rlabel locali s -11419 73574 -11157 73736 4 VDD
port 41 nsew
rlabel locali s -11747 72954 -11482 72988 4 VDD
port 41 nsew
rlabel locali s -11581 72988 -11482 73150 4 VDD
port 41 nsew
rlabel locali s -11747 73150 -11482 73184 4 VDD
port 41 nsew
rlabel locali s -11581 73184 -11482 73346 4 VDD
port 41 nsew
rlabel locali s -11747 73346 -11482 73380 4 VDD
port 41 nsew
rlabel locali s -11581 73380 -11482 73542 4 VDD
port 41 nsew
rlabel locali s -11747 73542 -11482 73576 4 VDD
port 41 nsew
rlabel locali s -11581 73576 -11482 73624 4 VDD
port 41 nsew
rlabel locali s -11419 73736 -10740 73770 4 VDD
port 41 nsew
rlabel locali s -11419 73770 -11107 73776 4 VDD
port 41 nsew
rlabel locali s -11206 73776 -11107 73953 4 VDD
port 41 nsew
rlabel locali s -11419 73776 -11249 73781 4 VDD
port 41 nsew
rlabel locali s -11443 73781 -11249 73787 4 VDD
port 41 nsew
rlabel locali s -11569 73787 -11249 73792 4 VDD
port 41 nsew
rlabel locali s -12159 73792 -11249 73826 4 VDD
port 41 nsew
rlabel locali s -11569 73826 -11249 73832 4 VDD
port 41 nsew
rlabel locali s -11443 73832 -11249 73951 4 VDD
port 41 nsew
rlabel locali s -11206 73953 -10941 73987 4 VDD
port 41 nsew
rlabel locali s -11206 73987 -11107 74149 4 VDD
port 41 nsew
rlabel locali s -11206 74149 -10941 74183 4 VDD
port 41 nsew
rlabel locali s -11206 74183 -11107 74345 4 VDD
port 41 nsew
rlabel locali s -11206 74345 -10941 74379 4 VDD
port 41 nsew
rlabel locali s -10299 74431 -7616 74553 4 VDD
port 41 nsew
rlabel locali s -11206 74379 -11107 74541 4 VDD
port 41 nsew
rlabel locali s -11443 73951 -11266 73982 4 VDD
port 41 nsew
rlabel locali s -11566 73982 -11266 73988 4 VDD
port 41 nsew
rlabel locali s -12159 73988 -11266 74022 4 VDD
port 41 nsew
rlabel locali s -11566 74022 -11266 74027 4 VDD
port 41 nsew
rlabel locali s -11443 74027 -11266 74404 4 VDD
port 41 nsew
rlabel locali s -11567 74404 -11266 74411 4 VDD
port 41 nsew
rlabel locali s -12159 74411 -11266 74445 4 VDD
port 41 nsew
rlabel locali s -11567 74445 -11266 74446 4 VDD
port 41 nsew
rlabel locali s -11567 74446 -11377 74449 4 VDD
port 41 nsew
rlabel locali s -11443 74449 -11377 74501 4 VDD
port 41 nsew
rlabel locali s -7870 74553 -7616 77526 4 VDD
port 41 nsew
rlabel locali s -10299 74553 -10177 74941 4 VDD
port 41 nsew
rlabel locali s -11206 74541 -10941 74575 4 VDD
port 41 nsew
rlabel locali s -11206 74575 -11107 74623 4 VDD
port 41 nsew
rlabel locali s -11443 74501 -11341 74550 4 VDD
port 41 nsew
rlabel locali s -11424 74550 -11341 74601 4 VDD
port 41 nsew
rlabel locali s -11449 74601 -11310 74680 4 VDD
port 41 nsew
rlabel locali s -11462 74851 -11295 74941 4 VDD
port 41 nsew
rlabel locali s -11462 74941 -10177 74990 4 VDD
port 41 nsew
rlabel locali s -11434 74990 -10177 75063 4 VDD
port 41 nsew
rlabel locali s -7870 77526 -7532 77538 4 VDD
port 41 nsew
rlabel locali s -7974 77538 -7532 77574 4 VDD
port 41 nsew
rlabel locali s -7974 77574 -7266 77608 4 VDD
port 41 nsew
rlabel locali s -7974 77608 -7532 77770 4 VDD
port 41 nsew
rlabel locali s -7974 77770 -7266 77804 4 VDD
port 41 nsew
rlabel locali s -7974 77804 -7532 77880 4 VDD
port 41 nsew
rlabel locali s -7631 77880 -7532 77966 4 VDD
port 41 nsew
rlabel locali s -7631 77966 -7266 78000 4 VDD
port 41 nsew
rlabel locali s -7631 78000 -7532 78162 4 VDD
port 41 nsew
rlabel locali s -7631 78162 -7266 78196 4 VDD
port 41 nsew
rlabel locali s -7631 78196 -7532 78244 4 VDD
port 41 nsew
rlabel locali s -7974 77880 -7821 77940 4 VDD
port 41 nsew
rlabel locali s -8086 77538 -8022 77548 4 VDD
port 41 nsew
rlabel locali s -8503 77548 -8022 77582 4 VDD
port 41 nsew
rlabel locali s -11084 77518 -10985 77566 4 VDD
port 41 nsew
rlabel locali s -8086 77582 -8022 77744 4 VDD
port 41 nsew
rlabel locali s -11084 77566 -10719 77600 4 VDD
port 41 nsew
rlabel locali s -11084 77600 -10985 77700 4 VDD
port 41 nsew
rlabel locali s -11427 77530 -11274 77700 4 VDD
port 41 nsew
rlabel locali s -8503 77744 -8022 77778 4 VDD
port 41 nsew
rlabel locali s -11427 77700 -10985 77762 4 VDD
port 41 nsew
rlabel locali s -8086 77778 -8022 77940 4 VDD
port 41 nsew
rlabel locali s -11427 77762 -10719 77796 4 VDD
port 41 nsew
rlabel locali s -11427 77796 -10985 77872 4 VDD
port 41 nsew
rlabel locali s -7981 77940 -7821 77977 4 VDD
port 41 nsew
rlabel locali s -8503 77940 -8022 77974 4 VDD
port 41 nsew
rlabel locali s -11084 77872 -10985 77958 4 VDD
port 41 nsew
rlabel locali s -7988 77977 -7821 78166 4 VDD
port 41 nsew
rlabel locali s -8136 77974 -8022 77980 4 VDD
port 41 nsew
rlabel locali s -8136 77980 -8037 78157 4 VDD
port 41 nsew
rlabel locali s -11084 77958 -10719 77992 4 VDD
port 41 nsew
rlabel locali s -11084 77992 -10985 78154 4 VDD
port 41 nsew
rlabel locali s -7974 78166 -7821 78536 4 VDD
port 41 nsew
rlabel locali s -7974 78536 -7775 78537 4 VDD
port 41 nsew
rlabel locali s -7974 78537 -7712 78547 4 VDD
port 41 nsew
rlabel locali s -7974 78547 -7295 78581 4 VDD
port 41 nsew
rlabel locali s -7974 78581 -7712 78743 4 VDD
port 41 nsew
rlabel locali s -7974 78743 -7295 78777 4 VDD
port 41 nsew
rlabel locali s -7974 78777 -7712 78939 4 VDD
port 41 nsew
rlabel locali s -8302 78157 -8037 78191 4 VDD
port 41 nsew
rlabel locali s -11084 78154 -10719 78188 4 VDD
port 41 nsew
rlabel locali s -8136 78191 -8037 78353 4 VDD
port 41 nsew
rlabel locali s -11084 78188 -10985 78236 4 VDD
port 41 nsew
rlabel locali s -11427 77872 -11274 77932 4 VDD
port 41 nsew
rlabel locali s -11539 77530 -11475 77540 4 VDD
port 41 nsew
rlabel locali s -11956 77540 -11475 77574 4 VDD
port 41 nsew
rlabel locali s -11539 77574 -11475 77736 4 VDD
port 41 nsew
rlabel locali s -11956 77736 -11475 77770 4 VDD
port 41 nsew
rlabel locali s -11539 77770 -11475 77932 4 VDD
port 41 nsew
rlabel locali s -11434 77932 -11274 77969 4 VDD
port 41 nsew
rlabel locali s -11956 77932 -11475 77966 4 VDD
port 41 nsew
rlabel locali s -11441 77969 -11274 78158 4 VDD
port 41 nsew
rlabel locali s -11589 77966 -11475 77972 4 VDD
port 41 nsew
rlabel locali s -11589 77972 -11490 78149 4 VDD
port 41 nsew
rlabel locali s -8302 78353 -8037 78387 4 VDD
port 41 nsew
rlabel locali s -8136 78387 -8037 78549 4 VDD
port 41 nsew
rlabel locali s -11427 78158 -11274 78528 4 VDD
port 41 nsew
rlabel locali s -11427 78528 -11228 78529 4 VDD
port 41 nsew
rlabel locali s -11427 78529 -11165 78539 4 VDD
port 41 nsew
rlabel locali s -8302 78549 -8037 78583 4 VDD
port 41 nsew
rlabel locali s -11427 78539 -10748 78573 4 VDD
port 41 nsew
rlabel locali s -8136 78583 -8037 78745 4 VDD
port 41 nsew
rlabel locali s -11427 78573 -11165 78735 4 VDD
port 41 nsew
rlabel locali s -8302 78745 -8037 78779 4 VDD
port 41 nsew
rlabel locali s -11427 78735 -10748 78769 4 VDD
port 41 nsew
rlabel locali s -8136 78779 -8037 78827 4 VDD
port 41 nsew
rlabel locali s -11427 78769 -11165 78931 4 VDD
port 41 nsew
rlabel locali s -11755 78149 -11490 78183 4 VDD
port 41 nsew
rlabel locali s -11589 78183 -11490 78345 4 VDD
port 41 nsew
rlabel locali s -11755 78345 -11490 78379 4 VDD
port 41 nsew
rlabel locali s -11589 78379 -11490 78541 4 VDD
port 41 nsew
rlabel locali s -11755 78541 -11490 78575 4 VDD
port 41 nsew
rlabel locali s -11589 78575 -11490 78737 4 VDD
port 41 nsew
rlabel locali s -11755 78737 -11490 78771 4 VDD
port 41 nsew
rlabel locali s -11589 78771 -11490 78819 4 VDD
port 41 nsew
rlabel locali s -7974 78939 -7295 78973 4 VDD
port 41 nsew
rlabel locali s -11427 78931 -10748 78965 4 VDD
port 41 nsew
rlabel locali s -7974 78973 -7662 78979 4 VDD
port 41 nsew
rlabel locali s -7761 78979 -7662 79156 4 VDD
port 41 nsew
rlabel locali s -7974 78979 -7804 78984 4 VDD
port 41 nsew
rlabel locali s -11427 78965 -11115 78971 4 VDD
port 41 nsew
rlabel locali s -7998 78984 -7804 78990 4 VDD
port 41 nsew
rlabel locali s -8124 78990 -7804 78995 4 VDD
port 41 nsew
rlabel locali s -8714 78995 -7804 79029 4 VDD
port 41 nsew
rlabel locali s -8124 79029 -7804 79035 4 VDD
port 41 nsew
rlabel locali s -7998 79035 -7804 79154 4 VDD
port 41 nsew
rlabel locali s -11214 78971 -11115 79148 4 VDD
port 41 nsew
rlabel locali s -11427 78971 -11257 78976 4 VDD
port 41 nsew
rlabel locali s -11451 78976 -11257 78982 4 VDD
port 41 nsew
rlabel locali s -11577 78982 -11257 78987 4 VDD
port 41 nsew
rlabel locali s -12167 78987 -11257 79021 4 VDD
port 41 nsew
rlabel locali s -11577 79021 -11257 79027 4 VDD
port 41 nsew
rlabel locali s -11451 79027 -11257 79146 4 VDD
port 41 nsew
rlabel locali s -7761 79156 -7496 79190 4 VDD
port 41 nsew
rlabel locali s -7761 79190 -7662 79352 4 VDD
port 41 nsew
rlabel locali s -7761 79352 -7496 79386 4 VDD
port 41 nsew
rlabel locali s -7761 79386 -7662 79548 4 VDD
port 41 nsew
rlabel locali s -7761 79548 -7496 79582 4 VDD
port 41 nsew
rlabel locali s -7761 79582 -7662 79744 4 VDD
port 41 nsew
rlabel locali s -7998 79154 -7821 79185 4 VDD
port 41 nsew
rlabel locali s -11214 79148 -10949 79182 4 VDD
port 41 nsew
rlabel locali s -8121 79185 -7821 79191 4 VDD
port 41 nsew
rlabel locali s -8714 79191 -7821 79225 4 VDD
port 41 nsew
rlabel locali s -8121 79225 -7821 79230 4 VDD
port 41 nsew
rlabel locali s -7998 79230 -7821 79607 4 VDD
port 41 nsew
rlabel locali s -11214 79182 -11115 79344 4 VDD
port 41 nsew
rlabel locali s -11214 79344 -10949 79378 4 VDD
port 41 nsew
rlabel locali s -11214 79378 -11115 79540 4 VDD
port 41 nsew
rlabel locali s -11214 79540 -10949 79574 4 VDD
port 41 nsew
rlabel locali s -8122 79607 -7821 79614 4 VDD
port 41 nsew
rlabel locali s -8714 79614 -7821 79648 4 VDD
port 41 nsew
rlabel locali s -8122 79648 -7821 79649 4 VDD
port 41 nsew
rlabel locali s -7761 79744 -7496 79778 4 VDD
port 41 nsew
rlabel locali s -8122 79649 -7932 79652 4 VDD
port 41 nsew
rlabel locali s -7998 79652 -7932 79753 4 VDD
port 41 nsew
rlabel locali s -11214 79574 -11115 79736 4 VDD
port 41 nsew
rlabel locali s -11451 79146 -11274 79177 4 VDD
port 41 nsew
rlabel locali s -11574 79177 -11274 79183 4 VDD
port 41 nsew
rlabel locali s -12167 79183 -11274 79217 4 VDD
port 41 nsew
rlabel locali s -11574 79217 -11274 79222 4 VDD
port 41 nsew
rlabel locali s -11451 79222 -11274 79599 4 VDD
port 41 nsew
rlabel locali s -11575 79599 -11274 79606 4 VDD
port 41 nsew
rlabel locali s -12167 79606 -11274 79640 4 VDD
port 41 nsew
rlabel locali s -11575 79640 -11274 79641 4 VDD
port 41 nsew
rlabel locali s -7761 79778 -7662 79826 4 VDD
port 41 nsew
rlabel locali s -7991 79753 -7939 79826 4 VDD
port 41 nsew
rlabel locali s -11214 79736 -10949 79770 4 VDD
port 41 nsew
rlabel locali s -11575 79641 -11385 79644 4 VDD
port 41 nsew
rlabel locali s -11451 79644 -11385 79745 4 VDD
port 41 nsew
rlabel locali s -11214 79770 -11115 79818 4 VDD
port 41 nsew
rlabel locali s -8005 79826 -7911 79888 4 VDD
port 41 nsew
rlabel locali s -8017 80054 -7891 80152 4 VDD
port 41 nsew
rlabel locali s -11423 80044 -11310 80061 4 VDD
port 41 nsew
rlabel locali s -11423 80061 -9943 80127 4 VDD
port 41 nsew
rlabel locali s -8011 80152 -7894 80617 4 VDD
port 41 nsew
rlabel locali s -10009 80127 -9943 80397 4 VDD
port 41 nsew
rlabel locali s -11423 80127 -11310 80128 4 VDD
port 41 nsew
rlabel locali s -11405 80397 -9943 80463 4 VDD
port 41 nsew
rlabel locali s -8011 80617 -7767 80734 4 VDD
port 41 nsew
rlabel locali s -7884 80734 -7767 80984 4 VDD
port 41 nsew
rlabel locali s -7979 80984 -7697 80987 4 VDD
port 41 nsew
rlabel locali s -8472 80987 -7697 81021 4 VDD
port 41 nsew
rlabel locali s -7979 81021 -7697 81022 4 VDD
port 41 nsew
rlabel locali s -7820 81022 -7697 81181 4 VDD
port 41 nsew
rlabel locali s -7977 81181 -7697 81183 4 VDD
port 41 nsew
rlabel locali s -8472 81183 -7697 81217 4 VDD
port 41 nsew
rlabel locali s -7977 81217 -7697 81219 4 VDD
port 41 nsew
rlabel locali s -7820 81219 -7697 81773 4 VDD
port 41 nsew
rlabel locali s -11115 81186 -11016 81234 4 VDD
port 41 nsew
rlabel locali s -11405 80463 -11339 81198 4 VDD
port 41 nsew
rlabel locali s -11115 81234 -10750 81268 4 VDD
port 41 nsew
rlabel locali s -11115 81268 -11016 81368 4 VDD
port 41 nsew
rlabel locali s -11458 81198 -11305 81368 4 VDD
port 41 nsew
rlabel locali s -11458 81368 -11016 81430 4 VDD
port 41 nsew
rlabel locali s -11458 81430 -10750 81464 4 VDD
port 41 nsew
rlabel locali s -11458 81464 -11016 81540 4 VDD
port 41 nsew
rlabel locali s -11115 81540 -11016 81626 4 VDD
port 41 nsew
rlabel locali s -11115 81626 -10750 81660 4 VDD
port 41 nsew
rlabel locali s -8000 81773 -7697 81778 4 VDD
port 41 nsew
rlabel locali s -8472 81778 -7697 81812 4 VDD
port 41 nsew
rlabel locali s -8000 81812 -7697 81823 4 VDD
port 41 nsew
rlabel locali s -11115 81660 -11016 81822 4 VDD
port 41 nsew
rlabel locali s -7820 81823 -7697 81899 4 VDD
port 41 nsew
rlabel locali s -11115 81822 -10750 81856 4 VDD
port 41 nsew
rlabel locali s -7997 81899 -7697 81908 4 VDD
port 41 nsew
rlabel locali s -11115 81856 -11016 81904 4 VDD
port 41 nsew
rlabel locali s -11458 81540 -11305 81600 4 VDD
port 41 nsew
rlabel locali s -11570 81198 -11506 81208 4 VDD
port 41 nsew
rlabel locali s -11987 81208 -11506 81242 4 VDD
port 41 nsew
rlabel locali s -11570 81242 -11506 81404 4 VDD
port 41 nsew
rlabel locali s -11987 81404 -11506 81438 4 VDD
port 41 nsew
rlabel locali s -11570 81438 -11506 81600 4 VDD
port 41 nsew
rlabel locali s -11465 81600 -11305 81637 4 VDD
port 41 nsew
rlabel locali s -11987 81600 -11506 81634 4 VDD
port 41 nsew
rlabel locali s -11472 81637 -11305 81826 4 VDD
port 41 nsew
rlabel locali s -11620 81634 -11506 81640 4 VDD
port 41 nsew
rlabel locali s -11620 81640 -11521 81817 4 VDD
port 41 nsew
rlabel locali s -8472 81908 -7697 81942 4 VDD
port 41 nsew
rlabel locali s -7997 81942 -7697 81949 4 VDD
port 41 nsew
rlabel locali s -7820 81949 -7697 82130 4 VDD
port 41 nsew
rlabel locali s -7982 82130 -7697 82136 4 VDD
port 41 nsew
rlabel locali s -8272 82136 -7697 82170 4 VDD
port 41 nsew
rlabel locali s -7982 82170 -7697 82173 4 VDD
port 41 nsew
rlabel locali s -7820 82173 -7697 82327 4 VDD
port 41 nsew
rlabel locali s -11458 81826 -11305 82196 4 VDD
port 41 nsew
rlabel locali s -11458 82196 -11259 82197 4 VDD
port 41 nsew
rlabel locali s -11458 82197 -11196 82207 4 VDD
port 41 nsew
rlabel locali s -11458 82207 -10779 82241 4 VDD
port 41 nsew
rlabel locali s -7980 82327 -7697 82332 4 VDD
port 41 nsew
rlabel locali s -8272 82332 -7697 82344 4 VDD
port 41 nsew
rlabel locali s -8272 82344 -7566 82366 4 VDD
port 41 nsew
rlabel locali s -7980 82366 -7566 82370 4 VDD
port 41 nsew
rlabel locali s -7880 82370 -7566 83294 4 VDD
port 41 nsew
rlabel locali s -11458 82241 -11196 82403 4 VDD
port 41 nsew
rlabel locali s -11458 82403 -10779 82437 4 VDD
port 41 nsew
rlabel locali s -11458 82437 -11196 82599 4 VDD
port 41 nsew
rlabel locali s -11786 81817 -11521 81851 4 VDD
port 41 nsew
rlabel locali s -11620 81851 -11521 82013 4 VDD
port 41 nsew
rlabel locali s -11786 82013 -11521 82047 4 VDD
port 41 nsew
rlabel locali s -11620 82047 -11521 82209 4 VDD
port 41 nsew
rlabel locali s -11786 82209 -11521 82243 4 VDD
port 41 nsew
rlabel locali s -11620 82243 -11521 82405 4 VDD
port 41 nsew
rlabel locali s -11786 82405 -11521 82439 4 VDD
port 41 nsew
rlabel locali s -11620 82439 -11521 82487 4 VDD
port 41 nsew
rlabel locali s -11458 82599 -10779 82633 4 VDD
port 41 nsew
rlabel locali s -11458 82633 -11146 82639 4 VDD
port 41 nsew
rlabel locali s -11245 82639 -11146 82816 4 VDD
port 41 nsew
rlabel locali s -11458 82639 -11288 82644 4 VDD
port 41 nsew
rlabel locali s -11482 82644 -11288 82650 4 VDD
port 41 nsew
rlabel locali s -11608 82650 -11288 82655 4 VDD
port 41 nsew
rlabel locali s -12198 82655 -11288 82689 4 VDD
port 41 nsew
rlabel locali s -11608 82689 -11288 82695 4 VDD
port 41 nsew
rlabel locali s -11482 82695 -11288 82814 4 VDD
port 41 nsew
rlabel locali s -11245 82816 -10980 82850 4 VDD
port 41 nsew
rlabel locali s -11245 82850 -11146 83012 4 VDD
port 41 nsew
rlabel locali s -11245 83012 -10980 83046 4 VDD
port 41 nsew
rlabel locali s -11245 83046 -11146 83208 4 VDD
port 41 nsew
rlabel locali s -11245 83208 -10980 83242 4 VDD
port 41 nsew
rlabel locali s -10338 83294 -7566 83416 4 VDD
port 41 nsew
rlabel locali s -11245 83242 -11146 83404 4 VDD
port 41 nsew
rlabel locali s -11482 82814 -11305 82845 4 VDD
port 41 nsew
rlabel locali s -11605 82845 -11305 82851 4 VDD
port 41 nsew
rlabel locali s -12198 82851 -11305 82885 4 VDD
port 41 nsew
rlabel locali s -11605 82885 -11305 82890 4 VDD
port 41 nsew
rlabel locali s -11482 82890 -11305 83267 4 VDD
port 41 nsew
rlabel locali s -11606 83267 -11305 83274 4 VDD
port 41 nsew
rlabel locali s -12198 83274 -11305 83308 4 VDD
port 41 nsew
rlabel locali s -11606 83308 -11305 83309 4 VDD
port 41 nsew
rlabel locali s -11606 83309 -11416 83312 4 VDD
port 41 nsew
rlabel locali s -11482 83312 -11416 83364 4 VDD
port 41 nsew
rlabel locali s -7880 83416 -7566 86724 4 VDD
port 41 nsew
rlabel locali s -10338 83416 -10216 83804 4 VDD
port 41 nsew
rlabel locali s -11245 83404 -10980 83438 4 VDD
port 41 nsew
rlabel locali s -11245 83438 -11146 83486 4 VDD
port 41 nsew
rlabel locali s -11482 83364 -11380 83413 4 VDD
port 41 nsew
rlabel locali s -11463 83413 -11380 83464 4 VDD
port 41 nsew
rlabel locali s -11488 83464 -11349 83543 4 VDD
port 41 nsew
rlabel locali s -11501 83714 -11334 83804 4 VDD
port 41 nsew
rlabel locali s -11501 83804 -10216 83853 4 VDD
port 41 nsew
rlabel locali s -11473 83853 -10216 83926 4 VDD
port 41 nsew
rlabel locali s -7880 86724 -7498 86736 4 VDD
port 41 nsew
rlabel locali s -7940 86736 -7498 86772 4 VDD
port 41 nsew
rlabel locali s -7940 86772 -7232 86806 4 VDD
port 41 nsew
rlabel locali s -7940 86806 -7498 86968 4 VDD
port 41 nsew
rlabel locali s -7940 86968 -7232 87002 4 VDD
port 41 nsew
rlabel locali s -7940 87002 -7498 87078 4 VDD
port 41 nsew
rlabel locali s -7597 87078 -7498 87164 4 VDD
port 41 nsew
rlabel locali s -7597 87164 -7232 87198 4 VDD
port 41 nsew
rlabel locali s -7597 87198 -7498 87360 4 VDD
port 41 nsew
rlabel locali s -7597 87360 -7232 87394 4 VDD
port 41 nsew
rlabel locali s -7597 87394 -7498 87442 4 VDD
port 41 nsew
rlabel locali s -7940 87078 -7787 87138 4 VDD
port 41 nsew
rlabel locali s -8052 86736 -7988 86746 4 VDD
port 41 nsew
rlabel locali s -8469 86746 -7988 86780 4 VDD
port 41 nsew
rlabel locali s -11050 86716 -10951 86764 4 VDD
port 41 nsew
rlabel locali s -8052 86780 -7988 86942 4 VDD
port 41 nsew
rlabel locali s -11050 86764 -10685 86798 4 VDD
port 41 nsew
rlabel locali s -11050 86798 -10951 86898 4 VDD
port 41 nsew
rlabel locali s -11393 86728 -11240 86898 4 VDD
port 41 nsew
rlabel locali s -8469 86942 -7988 86976 4 VDD
port 41 nsew
rlabel locali s -11393 86898 -10951 86960 4 VDD
port 41 nsew
rlabel locali s -8052 86976 -7988 87138 4 VDD
port 41 nsew
rlabel locali s -11393 86960 -10685 86994 4 VDD
port 41 nsew
rlabel locali s -11393 86994 -10951 87070 4 VDD
port 41 nsew
rlabel locali s -7947 87138 -7787 87175 4 VDD
port 41 nsew
rlabel locali s -8469 87138 -7988 87172 4 VDD
port 41 nsew
rlabel locali s -11050 87070 -10951 87156 4 VDD
port 41 nsew
rlabel locali s -7954 87175 -7787 87364 4 VDD
port 41 nsew
rlabel locali s -8102 87172 -7988 87178 4 VDD
port 41 nsew
rlabel locali s -8102 87178 -8003 87355 4 VDD
port 41 nsew
rlabel locali s -11050 87156 -10685 87190 4 VDD
port 41 nsew
rlabel locali s -11050 87190 -10951 87352 4 VDD
port 41 nsew
rlabel locali s -7940 87364 -7787 87734 4 VDD
port 41 nsew
rlabel locali s -7940 87734 -7741 87735 4 VDD
port 41 nsew
rlabel locali s -7940 87735 -7678 87745 4 VDD
port 41 nsew
rlabel locali s -7940 87745 -7261 87779 4 VDD
port 41 nsew
rlabel locali s -7940 87779 -7678 87941 4 VDD
port 41 nsew
rlabel locali s -7940 87941 -7261 87975 4 VDD
port 41 nsew
rlabel locali s -7940 87975 -7678 88137 4 VDD
port 41 nsew
rlabel locali s -8268 87355 -8003 87389 4 VDD
port 41 nsew
rlabel locali s -11050 87352 -10685 87386 4 VDD
port 41 nsew
rlabel locali s -8102 87389 -8003 87551 4 VDD
port 41 nsew
rlabel locali s -11050 87386 -10951 87434 4 VDD
port 41 nsew
rlabel locali s -11393 87070 -11240 87130 4 VDD
port 41 nsew
rlabel locali s -11505 86728 -11441 86738 4 VDD
port 41 nsew
rlabel locali s -11922 86738 -11441 86772 4 VDD
port 41 nsew
rlabel locali s -11505 86772 -11441 86934 4 VDD
port 41 nsew
rlabel locali s -11922 86934 -11441 86968 4 VDD
port 41 nsew
rlabel locali s -11505 86968 -11441 87130 4 VDD
port 41 nsew
rlabel locali s -11400 87130 -11240 87167 4 VDD
port 41 nsew
rlabel locali s -11922 87130 -11441 87164 4 VDD
port 41 nsew
rlabel locali s -11407 87167 -11240 87356 4 VDD
port 41 nsew
rlabel locali s -11555 87164 -11441 87170 4 VDD
port 41 nsew
rlabel locali s -11555 87170 -11456 87347 4 VDD
port 41 nsew
rlabel locali s -8268 87551 -8003 87585 4 VDD
port 41 nsew
rlabel locali s -8102 87585 -8003 87747 4 VDD
port 41 nsew
rlabel locali s -11393 87356 -11240 87726 4 VDD
port 41 nsew
rlabel locali s -11393 87726 -11194 87727 4 VDD
port 41 nsew
rlabel locali s -11393 87727 -11131 87737 4 VDD
port 41 nsew
rlabel locali s -8268 87747 -8003 87781 4 VDD
port 41 nsew
rlabel locali s -11393 87737 -10714 87771 4 VDD
port 41 nsew
rlabel locali s -8102 87781 -8003 87943 4 VDD
port 41 nsew
rlabel locali s -11393 87771 -11131 87933 4 VDD
port 41 nsew
rlabel locali s -8268 87943 -8003 87977 4 VDD
port 41 nsew
rlabel locali s -11393 87933 -10714 87967 4 VDD
port 41 nsew
rlabel locali s -8102 87977 -8003 88025 4 VDD
port 41 nsew
rlabel locali s -11393 87967 -11131 88129 4 VDD
port 41 nsew
rlabel locali s -11721 87347 -11456 87381 4 VDD
port 41 nsew
rlabel locali s -11555 87381 -11456 87543 4 VDD
port 41 nsew
rlabel locali s -11721 87543 -11456 87577 4 VDD
port 41 nsew
rlabel locali s -11555 87577 -11456 87739 4 VDD
port 41 nsew
rlabel locali s -11721 87739 -11456 87773 4 VDD
port 41 nsew
rlabel locali s -11555 87773 -11456 87935 4 VDD
port 41 nsew
rlabel locali s -11721 87935 -11456 87969 4 VDD
port 41 nsew
rlabel locali s -11555 87969 -11456 88017 4 VDD
port 41 nsew
rlabel locali s -7940 88137 -7261 88171 4 VDD
port 41 nsew
rlabel locali s -11393 88129 -10714 88163 4 VDD
port 41 nsew
rlabel locali s -7940 88171 -7628 88177 4 VDD
port 41 nsew
rlabel locali s -7727 88177 -7628 88354 4 VDD
port 41 nsew
rlabel locali s -7940 88177 -7770 88182 4 VDD
port 41 nsew
rlabel locali s -11393 88163 -11081 88169 4 VDD
port 41 nsew
rlabel locali s -7964 88182 -7770 88188 4 VDD
port 41 nsew
rlabel locali s -8090 88188 -7770 88193 4 VDD
port 41 nsew
rlabel locali s -8680 88193 -7770 88227 4 VDD
port 41 nsew
rlabel locali s -8090 88227 -7770 88233 4 VDD
port 41 nsew
rlabel locali s -7964 88233 -7770 88352 4 VDD
port 41 nsew
rlabel locali s -11180 88169 -11081 88346 4 VDD
port 41 nsew
rlabel locali s -11393 88169 -11223 88174 4 VDD
port 41 nsew
rlabel locali s -11417 88174 -11223 88180 4 VDD
port 41 nsew
rlabel locali s -11543 88180 -11223 88185 4 VDD
port 41 nsew
rlabel locali s -12133 88185 -11223 88219 4 VDD
port 41 nsew
rlabel locali s -11543 88219 -11223 88225 4 VDD
port 41 nsew
rlabel locali s -11417 88225 -11223 88344 4 VDD
port 41 nsew
rlabel locali s -7727 88354 -7462 88388 4 VDD
port 41 nsew
rlabel locali s -7727 88388 -7628 88550 4 VDD
port 41 nsew
rlabel locali s -7727 88550 -7462 88584 4 VDD
port 41 nsew
rlabel locali s -7727 88584 -7628 88746 4 VDD
port 41 nsew
rlabel locali s -7727 88746 -7462 88780 4 VDD
port 41 nsew
rlabel locali s -7727 88780 -7628 88942 4 VDD
port 41 nsew
rlabel locali s -7964 88352 -7787 88383 4 VDD
port 41 nsew
rlabel locali s -11180 88346 -10915 88380 4 VDD
port 41 nsew
rlabel locali s -8087 88383 -7787 88389 4 VDD
port 41 nsew
rlabel locali s -8680 88389 -7787 88423 4 VDD
port 41 nsew
rlabel locali s -8087 88423 -7787 88428 4 VDD
port 41 nsew
rlabel locali s -7964 88428 -7787 88805 4 VDD
port 41 nsew
rlabel locali s -11180 88380 -11081 88542 4 VDD
port 41 nsew
rlabel locali s -11180 88542 -10915 88576 4 VDD
port 41 nsew
rlabel locali s -11180 88576 -11081 88738 4 VDD
port 41 nsew
rlabel locali s -11180 88738 -10915 88772 4 VDD
port 41 nsew
rlabel locali s -8088 88805 -7787 88812 4 VDD
port 41 nsew
rlabel locali s -8680 88812 -7787 88846 4 VDD
port 41 nsew
rlabel locali s -8088 88846 -7787 88847 4 VDD
port 41 nsew
rlabel locali s -7727 88942 -7462 88976 4 VDD
port 41 nsew
rlabel locali s -8088 88847 -7898 88850 4 VDD
port 41 nsew
rlabel locali s -7964 88850 -7898 88951 4 VDD
port 41 nsew
rlabel locali s -11180 88772 -11081 88934 4 VDD
port 41 nsew
rlabel locali s -11417 88344 -11240 88375 4 VDD
port 41 nsew
rlabel locali s -11540 88375 -11240 88381 4 VDD
port 41 nsew
rlabel locali s -12133 88381 -11240 88415 4 VDD
port 41 nsew
rlabel locali s -11540 88415 -11240 88420 4 VDD
port 41 nsew
rlabel locali s -11417 88420 -11240 88797 4 VDD
port 41 nsew
rlabel locali s -11541 88797 -11240 88804 4 VDD
port 41 nsew
rlabel locali s -12133 88804 -11240 88838 4 VDD
port 41 nsew
rlabel locali s -11541 88838 -11240 88839 4 VDD
port 41 nsew
rlabel locali s -7727 88976 -7628 89024 4 VDD
port 41 nsew
rlabel locali s -7957 88951 -7905 89024 4 VDD
port 41 nsew
rlabel locali s -11180 88934 -10915 88968 4 VDD
port 41 nsew
rlabel locali s -11541 88839 -11351 88842 4 VDD
port 41 nsew
rlabel locali s -11417 88842 -11351 88943 4 VDD
port 41 nsew
rlabel locali s -11180 88968 -11081 89016 4 VDD
port 41 nsew
rlabel locali s -7971 89024 -7877 89086 4 VDD
port 41 nsew
rlabel locali s -7983 89252 -7857 89350 4 VDD
port 41 nsew
rlabel locali s -11389 89242 -11276 89259 4 VDD
port 41 nsew
rlabel locali s -11389 89259 -9909 89325 4 VDD
port 41 nsew
rlabel locali s -7977 89350 -7860 89815 4 VDD
port 41 nsew
rlabel locali s -9975 89325 -9909 89595 4 VDD
port 41 nsew
rlabel locali s -11389 89325 -11276 89326 4 VDD
port 41 nsew
rlabel locali s -11371 89595 -9909 89661 4 VDD
port 41 nsew
rlabel locali s -7977 89815 -7733 89932 4 VDD
port 41 nsew
rlabel locali s -7850 89932 -7733 90182 4 VDD
port 41 nsew
rlabel locali s -7945 90182 -7663 90185 4 VDD
port 41 nsew
rlabel locali s -8438 90185 -7663 90219 4 VDD
port 41 nsew
rlabel locali s -7945 90219 -7663 90220 4 VDD
port 41 nsew
rlabel locali s -7786 90220 -7663 90379 4 VDD
port 41 nsew
rlabel locali s -7943 90379 -7663 90381 4 VDD
port 41 nsew
rlabel locali s -8438 90381 -7663 90415 4 VDD
port 41 nsew
rlabel locali s -7943 90415 -7663 90417 4 VDD
port 41 nsew
rlabel locali s -7786 90417 -7663 90971 4 VDD
port 41 nsew
rlabel locali s -11081 90384 -10982 90432 4 VDD
port 41 nsew
rlabel locali s -11371 89661 -11305 90396 4 VDD
port 41 nsew
rlabel locali s -11081 90432 -10716 90466 4 VDD
port 41 nsew
rlabel locali s -11081 90466 -10982 90566 4 VDD
port 41 nsew
rlabel locali s -11424 90396 -11271 90566 4 VDD
port 41 nsew
rlabel locali s -11424 90566 -10982 90628 4 VDD
port 41 nsew
rlabel locali s -11424 90628 -10716 90662 4 VDD
port 41 nsew
rlabel locali s -11424 90662 -10982 90738 4 VDD
port 41 nsew
rlabel locali s -11081 90738 -10982 90824 4 VDD
port 41 nsew
rlabel locali s -11081 90824 -10716 90858 4 VDD
port 41 nsew
rlabel locali s -7966 90971 -7663 90976 4 VDD
port 41 nsew
rlabel locali s -8438 90976 -7663 91010 4 VDD
port 41 nsew
rlabel locali s -7966 91010 -7663 91021 4 VDD
port 41 nsew
rlabel locali s -11081 90858 -10982 91020 4 VDD
port 41 nsew
rlabel locali s -7786 91021 -7663 91097 4 VDD
port 41 nsew
rlabel locali s -11081 91020 -10716 91054 4 VDD
port 41 nsew
rlabel locali s -7963 91097 -7663 91106 4 VDD
port 41 nsew
rlabel locali s -11081 91054 -10982 91102 4 VDD
port 41 nsew
rlabel locali s -11424 90738 -11271 90798 4 VDD
port 41 nsew
rlabel locali s -11536 90396 -11472 90406 4 VDD
port 41 nsew
rlabel locali s -11953 90406 -11472 90440 4 VDD
port 41 nsew
rlabel locali s -11536 90440 -11472 90602 4 VDD
port 41 nsew
rlabel locali s -11953 90602 -11472 90636 4 VDD
port 41 nsew
rlabel locali s -11536 90636 -11472 90798 4 VDD
port 41 nsew
rlabel locali s -11431 90798 -11271 90835 4 VDD
port 41 nsew
rlabel locali s -11953 90798 -11472 90832 4 VDD
port 41 nsew
rlabel locali s -11438 90835 -11271 91024 4 VDD
port 41 nsew
rlabel locali s -11586 90832 -11472 90838 4 VDD
port 41 nsew
rlabel locali s -11586 90838 -11487 91015 4 VDD
port 41 nsew
rlabel locali s -8438 91106 -7663 91140 4 VDD
port 41 nsew
rlabel locali s -7963 91140 -7663 91147 4 VDD
port 41 nsew
rlabel locali s -7786 91147 -7663 91328 4 VDD
port 41 nsew
rlabel locali s -7948 91328 -7663 91334 4 VDD
port 41 nsew
rlabel locali s -8238 91334 -7663 91368 4 VDD
port 41 nsew
rlabel locali s -7948 91368 -7663 91371 4 VDD
port 41 nsew
rlabel locali s -7786 91371 -7663 91525 4 VDD
port 41 nsew
rlabel locali s -11424 91024 -11271 91394 4 VDD
port 41 nsew
rlabel locali s -11424 91394 -11225 91395 4 VDD
port 41 nsew
rlabel locali s -11424 91395 -11162 91405 4 VDD
port 41 nsew
rlabel locali s -11424 91405 -10745 91439 4 VDD
port 41 nsew
rlabel locali s -7946 91525 -7663 91527 4 VDD
port 41 nsew
rlabel locali s -7946 91527 -7469 91530 4 VDD
port 41 nsew
rlabel locali s -8238 91530 -7469 91564 4 VDD
port 41 nsew
rlabel locali s -7946 91564 -7469 91568 4 VDD
port 41 nsew
rlabel locali s -7848 91568 -7469 92492 4 VDD
port 41 nsew
rlabel locali s -11424 91439 -11162 91601 4 VDD
port 41 nsew
rlabel locali s -11424 91601 -10745 91635 4 VDD
port 41 nsew
rlabel locali s -11424 91635 -11162 91797 4 VDD
port 41 nsew
rlabel locali s -11752 91015 -11487 91049 4 VDD
port 41 nsew
rlabel locali s -11586 91049 -11487 91211 4 VDD
port 41 nsew
rlabel locali s -11752 91211 -11487 91245 4 VDD
port 41 nsew
rlabel locali s -11586 91245 -11487 91407 4 VDD
port 41 nsew
rlabel locali s -11752 91407 -11487 91441 4 VDD
port 41 nsew
rlabel locali s -11586 91441 -11487 91603 4 VDD
port 41 nsew
rlabel locali s -11752 91603 -11487 91637 4 VDD
port 41 nsew
rlabel locali s -11586 91637 -11487 91685 4 VDD
port 41 nsew
rlabel locali s -11424 91797 -10745 91831 4 VDD
port 41 nsew
rlabel locali s -11424 91831 -11112 91837 4 VDD
port 41 nsew
rlabel locali s -11211 91837 -11112 92014 4 VDD
port 41 nsew
rlabel locali s -11424 91837 -11254 91842 4 VDD
port 41 nsew
rlabel locali s -11448 91842 -11254 91848 4 VDD
port 41 nsew
rlabel locali s -11574 91848 -11254 91853 4 VDD
port 41 nsew
rlabel locali s -12164 91853 -11254 91887 4 VDD
port 41 nsew
rlabel locali s -11574 91887 -11254 91893 4 VDD
port 41 nsew
rlabel locali s -11448 91893 -11254 92012 4 VDD
port 41 nsew
rlabel locali s -11211 92014 -10946 92048 4 VDD
port 41 nsew
rlabel locali s -11211 92048 -11112 92210 4 VDD
port 41 nsew
rlabel locali s -11211 92210 -10946 92244 4 VDD
port 41 nsew
rlabel locali s -11211 92244 -11112 92406 4 VDD
port 41 nsew
rlabel locali s -11211 92406 -10946 92440 4 VDD
port 41 nsew
rlabel locali s -10304 92492 -7469 92614 4 VDD
port 41 nsew
rlabel locali s -11211 92440 -11112 92602 4 VDD
port 41 nsew
rlabel locali s -11448 92012 -11271 92043 4 VDD
port 41 nsew
rlabel locali s -11571 92043 -11271 92049 4 VDD
port 41 nsew
rlabel locali s -12164 92049 -11271 92083 4 VDD
port 41 nsew
rlabel locali s -11571 92083 -11271 92088 4 VDD
port 41 nsew
rlabel locali s -11448 92088 -11271 92465 4 VDD
port 41 nsew
rlabel locali s -11572 92465 -11271 92472 4 VDD
port 41 nsew
rlabel locali s -12164 92472 -11271 92506 4 VDD
port 41 nsew
rlabel locali s -11572 92506 -11271 92507 4 VDD
port 41 nsew
rlabel locali s -11572 92507 -11382 92510 4 VDD
port 41 nsew
rlabel locali s -11448 92510 -11382 92562 4 VDD
port 41 nsew
rlabel locali s -7848 92614 -7469 95478 4 VDD
port 41 nsew
rlabel locali s -10304 92614 -10182 93002 4 VDD
port 41 nsew
rlabel locali s -11211 92602 -10946 92636 4 VDD
port 41 nsew
rlabel locali s -11211 92636 -11112 92684 4 VDD
port 41 nsew
rlabel locali s -11448 92562 -11346 92611 4 VDD
port 41 nsew
rlabel locali s -11429 92611 -11346 92662 4 VDD
port 41 nsew
rlabel locali s -11454 92662 -11315 92741 4 VDD
port 41 nsew
rlabel locali s -11467 92912 -11300 93002 4 VDD
port 41 nsew
rlabel locali s -11467 93002 -10182 93051 4 VDD
port 41 nsew
rlabel locali s -11439 93051 -10182 93124 4 VDD
port 41 nsew
rlabel locali s -7848 95478 -7432 95490 4 VDD
port 41 nsew
rlabel locali s -7874 95490 -7432 95526 4 VDD
port 41 nsew
rlabel locali s -7874 95526 -7166 95560 4 VDD
port 41 nsew
rlabel locali s -7874 95560 -7432 95722 4 VDD
port 41 nsew
rlabel locali s -7874 95722 -7166 95756 4 VDD
port 41 nsew
rlabel locali s -7874 95756 -7432 95832 4 VDD
port 41 nsew
rlabel locali s -7531 95832 -7432 95918 4 VDD
port 41 nsew
rlabel locali s -7531 95918 -7166 95952 4 VDD
port 41 nsew
rlabel locali s -7531 95952 -7432 96114 4 VDD
port 41 nsew
rlabel locali s -7531 96114 -7166 96148 4 VDD
port 41 nsew
rlabel locali s -7531 96148 -7432 96196 4 VDD
port 41 nsew
rlabel locali s -7874 95832 -7721 95892 4 VDD
port 41 nsew
rlabel locali s -7986 95490 -7922 95500 4 VDD
port 41 nsew
rlabel locali s -8403 95500 -7922 95534 4 VDD
port 41 nsew
rlabel locali s -10984 95470 -10885 95518 4 VDD
port 41 nsew
rlabel locali s -7986 95534 -7922 95696 4 VDD
port 41 nsew
rlabel locali s -10984 95518 -10619 95552 4 VDD
port 41 nsew
rlabel locali s -10984 95552 -10885 95652 4 VDD
port 41 nsew
rlabel locali s -11327 95482 -11174 95652 4 VDD
port 41 nsew
rlabel locali s -8403 95696 -7922 95730 4 VDD
port 41 nsew
rlabel locali s -11327 95652 -10885 95714 4 VDD
port 41 nsew
rlabel locali s -7986 95730 -7922 95892 4 VDD
port 41 nsew
rlabel locali s -11327 95714 -10619 95748 4 VDD
port 41 nsew
rlabel locali s -11327 95748 -10885 95824 4 VDD
port 41 nsew
rlabel locali s -7881 95892 -7721 95929 4 VDD
port 41 nsew
rlabel locali s -8403 95892 -7922 95926 4 VDD
port 41 nsew
rlabel locali s -10984 95824 -10885 95910 4 VDD
port 41 nsew
rlabel locali s -7888 95929 -7721 96118 4 VDD
port 41 nsew
rlabel locali s -8036 95926 -7922 95932 4 VDD
port 41 nsew
rlabel locali s -8036 95932 -7937 96109 4 VDD
port 41 nsew
rlabel locali s -10984 95910 -10619 95944 4 VDD
port 41 nsew
rlabel locali s -10984 95944 -10885 96106 4 VDD
port 41 nsew
rlabel locali s -7874 96118 -7721 96488 4 VDD
port 41 nsew
rlabel locali s -7874 96488 -7675 96489 4 VDD
port 41 nsew
rlabel locali s -7874 96489 -7612 96499 4 VDD
port 41 nsew
rlabel locali s -7874 96499 -7195 96533 4 VDD
port 41 nsew
rlabel locali s -7874 96533 -7612 96695 4 VDD
port 41 nsew
rlabel locali s -7874 96695 -7195 96729 4 VDD
port 41 nsew
rlabel locali s -7874 96729 -7612 96891 4 VDD
port 41 nsew
rlabel locali s -8202 96109 -7937 96143 4 VDD
port 41 nsew
rlabel locali s -10984 96106 -10619 96140 4 VDD
port 41 nsew
rlabel locali s -8036 96143 -7937 96305 4 VDD
port 41 nsew
rlabel locali s -10984 96140 -10885 96188 4 VDD
port 41 nsew
rlabel locali s -11327 95824 -11174 95884 4 VDD
port 41 nsew
rlabel locali s -11439 95482 -11375 95492 4 VDD
port 41 nsew
rlabel locali s -11856 95492 -11375 95526 4 VDD
port 41 nsew
rlabel locali s -11439 95526 -11375 95688 4 VDD
port 41 nsew
rlabel locali s -11856 95688 -11375 95722 4 VDD
port 41 nsew
rlabel locali s -11439 95722 -11375 95884 4 VDD
port 41 nsew
rlabel locali s -11334 95884 -11174 95921 4 VDD
port 41 nsew
rlabel locali s -11856 95884 -11375 95918 4 VDD
port 41 nsew
rlabel locali s -11341 95921 -11174 96110 4 VDD
port 41 nsew
rlabel locali s -11489 95918 -11375 95924 4 VDD
port 41 nsew
rlabel locali s -11489 95924 -11390 96101 4 VDD
port 41 nsew
rlabel locali s -8202 96305 -7937 96339 4 VDD
port 41 nsew
rlabel locali s -8036 96339 -7937 96501 4 VDD
port 41 nsew
rlabel locali s -11327 96110 -11174 96480 4 VDD
port 41 nsew
rlabel locali s -11327 96480 -11128 96481 4 VDD
port 41 nsew
rlabel locali s -11327 96481 -11065 96491 4 VDD
port 41 nsew
rlabel locali s -8202 96501 -7937 96535 4 VDD
port 41 nsew
rlabel locali s -11327 96491 -10648 96525 4 VDD
port 41 nsew
rlabel locali s -8036 96535 -7937 96697 4 VDD
port 41 nsew
rlabel locali s -11327 96525 -11065 96687 4 VDD
port 41 nsew
rlabel locali s -8202 96697 -7937 96731 4 VDD
port 41 nsew
rlabel locali s -11327 96687 -10648 96721 4 VDD
port 41 nsew
rlabel locali s -8036 96731 -7937 96779 4 VDD
port 41 nsew
rlabel locali s -11327 96721 -11065 96883 4 VDD
port 41 nsew
rlabel locali s -11655 96101 -11390 96135 4 VDD
port 41 nsew
rlabel locali s -11489 96135 -11390 96297 4 VDD
port 41 nsew
rlabel locali s -11655 96297 -11390 96331 4 VDD
port 41 nsew
rlabel locali s -11489 96331 -11390 96493 4 VDD
port 41 nsew
rlabel locali s -11655 96493 -11390 96527 4 VDD
port 41 nsew
rlabel locali s -11489 96527 -11390 96689 4 VDD
port 41 nsew
rlabel locali s -11655 96689 -11390 96723 4 VDD
port 41 nsew
rlabel locali s -11489 96723 -11390 96771 4 VDD
port 41 nsew
rlabel locali s -7874 96891 -7195 96925 4 VDD
port 41 nsew
rlabel locali s -11327 96883 -10648 96917 4 VDD
port 41 nsew
rlabel locali s -7874 96925 -7562 96931 4 VDD
port 41 nsew
rlabel locali s -7661 96931 -7562 97108 4 VDD
port 41 nsew
rlabel locali s -7874 96931 -7704 96936 4 VDD
port 41 nsew
rlabel locali s -11327 96917 -11015 96923 4 VDD
port 41 nsew
rlabel locali s -7898 96936 -7704 96942 4 VDD
port 41 nsew
rlabel locali s -8024 96942 -7704 96947 4 VDD
port 41 nsew
rlabel locali s -8614 96947 -7704 96981 4 VDD
port 41 nsew
rlabel locali s -8024 96981 -7704 96987 4 VDD
port 41 nsew
rlabel locali s -7898 96987 -7704 97106 4 VDD
port 41 nsew
rlabel locali s -11114 96923 -11015 97100 4 VDD
port 41 nsew
rlabel locali s -11327 96923 -11157 96928 4 VDD
port 41 nsew
rlabel locali s -11351 96928 -11157 96934 4 VDD
port 41 nsew
rlabel locali s -11477 96934 -11157 96939 4 VDD
port 41 nsew
rlabel locali s -12067 96939 -11157 96973 4 VDD
port 41 nsew
rlabel locali s -11477 96973 -11157 96979 4 VDD
port 41 nsew
rlabel locali s -11351 96979 -11157 97098 4 VDD
port 41 nsew
rlabel locali s -7661 97108 -7396 97142 4 VDD
port 41 nsew
rlabel locali s -7661 97142 -7562 97304 4 VDD
port 41 nsew
rlabel locali s -7661 97304 -7396 97338 4 VDD
port 41 nsew
rlabel locali s -7661 97338 -7562 97500 4 VDD
port 41 nsew
rlabel locali s -7661 97500 -7396 97534 4 VDD
port 41 nsew
rlabel locali s -7661 97534 -7562 97696 4 VDD
port 41 nsew
rlabel locali s -7898 97106 -7721 97137 4 VDD
port 41 nsew
rlabel locali s -11114 97100 -10849 97134 4 VDD
port 41 nsew
rlabel locali s -8021 97137 -7721 97143 4 VDD
port 41 nsew
rlabel locali s -8614 97143 -7721 97177 4 VDD
port 41 nsew
rlabel locali s -8021 97177 -7721 97182 4 VDD
port 41 nsew
rlabel locali s -7898 97182 -7721 97559 4 VDD
port 41 nsew
rlabel locali s -11114 97134 -11015 97296 4 VDD
port 41 nsew
rlabel locali s -11114 97296 -10849 97330 4 VDD
port 41 nsew
rlabel locali s -11114 97330 -11015 97492 4 VDD
port 41 nsew
rlabel locali s -11114 97492 -10849 97526 4 VDD
port 41 nsew
rlabel locali s -8022 97559 -7721 97566 4 VDD
port 41 nsew
rlabel locali s -8614 97566 -7721 97600 4 VDD
port 41 nsew
rlabel locali s -8022 97600 -7721 97601 4 VDD
port 41 nsew
rlabel locali s -7661 97696 -7396 97730 4 VDD
port 41 nsew
rlabel locali s -8022 97601 -7832 97604 4 VDD
port 41 nsew
rlabel locali s -7898 97604 -7832 97705 4 VDD
port 41 nsew
rlabel locali s -11114 97526 -11015 97688 4 VDD
port 41 nsew
rlabel locali s -11351 97098 -11174 97129 4 VDD
port 41 nsew
rlabel locali s -11474 97129 -11174 97135 4 VDD
port 41 nsew
rlabel locali s -12067 97135 -11174 97169 4 VDD
port 41 nsew
rlabel locali s -11474 97169 -11174 97174 4 VDD
port 41 nsew
rlabel locali s -11351 97174 -11174 97551 4 VDD
port 41 nsew
rlabel locali s -11475 97551 -11174 97558 4 VDD
port 41 nsew
rlabel locali s -12067 97558 -11174 97592 4 VDD
port 41 nsew
rlabel locali s -11475 97592 -11174 97593 4 VDD
port 41 nsew
rlabel locali s -7661 97730 -7562 97778 4 VDD
port 41 nsew
rlabel locali s -7891 97705 -7839 97778 4 VDD
port 41 nsew
rlabel locali s -11114 97688 -10849 97722 4 VDD
port 41 nsew
rlabel locali s -11475 97593 -11285 97596 4 VDD
port 41 nsew
rlabel locali s -11351 97596 -11285 97697 4 VDD
port 41 nsew
rlabel locali s -11114 97722 -11015 97770 4 VDD
port 41 nsew
rlabel locali s -7905 97778 -7811 97840 4 VDD
port 41 nsew
rlabel locali s -7917 98006 -7791 98104 4 VDD
port 41 nsew
rlabel locali s -11323 97996 -11210 98013 4 VDD
port 41 nsew
rlabel locali s -11323 98013 -9843 98079 4 VDD
port 41 nsew
rlabel locali s -7911 98104 -7794 98569 4 VDD
port 41 nsew
rlabel locali s -9909 98079 -9843 98349 4 VDD
port 41 nsew
rlabel locali s -11323 98079 -11210 98080 4 VDD
port 41 nsew
rlabel locali s -11305 98349 -9843 98415 4 VDD
port 41 nsew
rlabel locali s -7911 98569 -7667 98686 4 VDD
port 41 nsew
rlabel locali s -7784 98686 -7667 98936 4 VDD
port 41 nsew
rlabel locali s -7879 98936 -7597 98939 4 VDD
port 41 nsew
rlabel locali s -8372 98939 -7597 98973 4 VDD
port 41 nsew
rlabel locali s -7879 98973 -7597 98974 4 VDD
port 41 nsew
rlabel locali s -7720 98974 -7597 99133 4 VDD
port 41 nsew
rlabel locali s -7877 99133 -7597 99135 4 VDD
port 41 nsew
rlabel locali s -8372 99135 -7597 99169 4 VDD
port 41 nsew
rlabel locali s -7877 99169 -7597 99171 4 VDD
port 41 nsew
rlabel locali s -7720 99171 -7597 99725 4 VDD
port 41 nsew
rlabel locali s -11015 99138 -10916 99186 4 VDD
port 41 nsew
rlabel locali s -11305 98415 -11239 99150 4 VDD
port 41 nsew
rlabel locali s -11015 99186 -10650 99220 4 VDD
port 41 nsew
rlabel locali s -11015 99220 -10916 99320 4 VDD
port 41 nsew
rlabel locali s -11358 99150 -11205 99320 4 VDD
port 41 nsew
rlabel locali s -11358 99320 -10916 99382 4 VDD
port 41 nsew
rlabel locali s -11358 99382 -10650 99416 4 VDD
port 41 nsew
rlabel locali s -11358 99416 -10916 99492 4 VDD
port 41 nsew
rlabel locali s -11015 99492 -10916 99578 4 VDD
port 41 nsew
rlabel locali s -11015 99578 -10650 99612 4 VDD
port 41 nsew
rlabel locali s -7900 99725 -7597 99730 4 VDD
port 41 nsew
rlabel locali s -8372 99730 -7597 99764 4 VDD
port 41 nsew
rlabel locali s -7900 99764 -7597 99775 4 VDD
port 41 nsew
rlabel locali s -11015 99612 -10916 99774 4 VDD
port 41 nsew
rlabel locali s -7720 99775 -7597 99851 4 VDD
port 41 nsew
rlabel locali s -11015 99774 -10650 99808 4 VDD
port 41 nsew
rlabel locali s -7897 99851 -7597 99860 4 VDD
port 41 nsew
rlabel locali s -11015 99808 -10916 99856 4 VDD
port 41 nsew
rlabel locali s -11358 99492 -11205 99552 4 VDD
port 41 nsew
rlabel locali s -11470 99150 -11406 99160 4 VDD
port 41 nsew
rlabel locali s -11887 99160 -11406 99194 4 VDD
port 41 nsew
rlabel locali s -11470 99194 -11406 99356 4 VDD
port 41 nsew
rlabel locali s -11887 99356 -11406 99390 4 VDD
port 41 nsew
rlabel locali s -11470 99390 -11406 99552 4 VDD
port 41 nsew
rlabel locali s -11365 99552 -11205 99589 4 VDD
port 41 nsew
rlabel locali s -11887 99552 -11406 99586 4 VDD
port 41 nsew
rlabel locali s -11372 99589 -11205 99778 4 VDD
port 41 nsew
rlabel locali s -11520 99586 -11406 99592 4 VDD
port 41 nsew
rlabel locali s -11520 99592 -11421 99769 4 VDD
port 41 nsew
rlabel locali s -8372 99860 -7597 99894 4 VDD
port 41 nsew
rlabel locali s -7897 99894 -7597 99901 4 VDD
port 41 nsew
rlabel locali s -7720 99901 -7597 100082 4 VDD
port 41 nsew
rlabel locali s -7882 100082 -7597 100088 4 VDD
port 41 nsew
rlabel locali s -8172 100088 -7597 100122 4 VDD
port 41 nsew
rlabel locali s -7882 100122 -7597 100125 4 VDD
port 41 nsew
rlabel locali s -7720 100125 -7597 100274 4 VDD
port 41 nsew
rlabel locali s -11358 99778 -11205 100148 4 VDD
port 41 nsew
rlabel locali s -11358 100148 -11159 100149 4 VDD
port 41 nsew
rlabel locali s -11358 100149 -11096 100159 4 VDD
port 41 nsew
rlabel locali s -11358 100159 -10679 100193 4 VDD
port 41 nsew
rlabel locali s -7754 100274 -7490 100279 4 VDD
port 41 nsew
rlabel locali s -7880 100279 -7490 100284 4 VDD
port 41 nsew
rlabel locali s -8172 100284 -7490 100318 4 VDD
port 41 nsew
rlabel locali s -7880 100318 -7490 100322 4 VDD
port 41 nsew
rlabel locali s -7754 100322 -7490 101246 4 VDD
port 41 nsew
rlabel locali s -11358 100193 -11096 100355 4 VDD
port 41 nsew
rlabel locali s -11358 100355 -10679 100389 4 VDD
port 41 nsew
rlabel locali s -11358 100389 -11096 100551 4 VDD
port 41 nsew
rlabel locali s -11686 99769 -11421 99803 4 VDD
port 41 nsew
rlabel locali s -11520 99803 -11421 99965 4 VDD
port 41 nsew
rlabel locali s -11686 99965 -11421 99999 4 VDD
port 41 nsew
rlabel locali s -11520 99999 -11421 100161 4 VDD
port 41 nsew
rlabel locali s -11686 100161 -11421 100195 4 VDD
port 41 nsew
rlabel locali s -11520 100195 -11421 100357 4 VDD
port 41 nsew
rlabel locali s -11686 100357 -11421 100391 4 VDD
port 41 nsew
rlabel locali s -11520 100391 -11421 100439 4 VDD
port 41 nsew
rlabel locali s -11358 100551 -10679 100585 4 VDD
port 41 nsew
rlabel locali s -11358 100585 -11046 100591 4 VDD
port 41 nsew
rlabel locali s -11145 100591 -11046 100768 4 VDD
port 41 nsew
rlabel locali s -11358 100591 -11188 100596 4 VDD
port 41 nsew
rlabel locali s -11382 100596 -11188 100602 4 VDD
port 41 nsew
rlabel locali s -11508 100602 -11188 100607 4 VDD
port 41 nsew
rlabel locali s -12098 100607 -11188 100641 4 VDD
port 41 nsew
rlabel locali s -11508 100641 -11188 100647 4 VDD
port 41 nsew
rlabel locali s -11382 100647 -11188 100766 4 VDD
port 41 nsew
rlabel locali s -11145 100768 -10880 100802 4 VDD
port 41 nsew
rlabel locali s -11145 100802 -11046 100964 4 VDD
port 41 nsew
rlabel locali s -11145 100964 -10880 100998 4 VDD
port 41 nsew
rlabel locali s -11145 100998 -11046 101160 4 VDD
port 41 nsew
rlabel locali s -11145 101160 -10880 101194 4 VDD
port 41 nsew
rlabel locali s -10238 101246 -7490 101368 4 VDD
port 41 nsew
rlabel locali s -11145 101194 -11046 101356 4 VDD
port 41 nsew
rlabel locali s -11382 100766 -11205 100797 4 VDD
port 41 nsew
rlabel locali s -11505 100797 -11205 100803 4 VDD
port 41 nsew
rlabel locali s -12098 100803 -11205 100837 4 VDD
port 41 nsew
rlabel locali s -11505 100837 -11205 100842 4 VDD
port 41 nsew
rlabel locali s -11382 100842 -11205 101219 4 VDD
port 41 nsew
rlabel locali s -11506 101219 -11205 101226 4 VDD
port 41 nsew
rlabel locali s -12098 101226 -11205 101260 4 VDD
port 41 nsew
rlabel locali s -11506 101260 -11205 101261 4 VDD
port 41 nsew
rlabel locali s -11506 101261 -11316 101264 4 VDD
port 41 nsew
rlabel locali s -11382 101264 -11316 101316 4 VDD
port 41 nsew
rlabel locali s -7754 101368 -7490 104631 4 VDD
port 41 nsew
rlabel locali s -10238 101368 -10116 101756 4 VDD
port 41 nsew
rlabel locali s -11145 101356 -10880 101390 4 VDD
port 41 nsew
rlabel locali s -11145 101390 -11046 101438 4 VDD
port 41 nsew
rlabel locali s -11382 101316 -11280 101365 4 VDD
port 41 nsew
rlabel locali s -11363 101365 -11280 101416 4 VDD
port 41 nsew
rlabel locali s -11388 101416 -11249 101495 4 VDD
port 41 nsew
rlabel locali s -11401 101666 -11234 101756 4 VDD
port 41 nsew
rlabel locali s -11401 101756 -10116 101805 4 VDD
port 41 nsew
rlabel locali s -11373 101805 -10116 101878 4 VDD
port 41 nsew
rlabel locali s -7754 104631 -7415 104643 4 VDD
port 41 nsew
rlabel locali s -7857 104643 -7415 104679 4 VDD
port 41 nsew
rlabel locali s -7857 104679 -7149 104713 4 VDD
port 41 nsew
rlabel locali s -7857 104713 -7415 104875 4 VDD
port 41 nsew
rlabel locali s -7857 104875 -7149 104909 4 VDD
port 41 nsew
rlabel locali s -7857 104909 -7415 104985 4 VDD
port 41 nsew
rlabel locali s -7514 104985 -7415 105071 4 VDD
port 41 nsew
rlabel locali s -7514 105071 -7149 105105 4 VDD
port 41 nsew
rlabel locali s -7514 105105 -7415 105267 4 VDD
port 41 nsew
rlabel locali s -7514 105267 -7149 105301 4 VDD
port 41 nsew
rlabel locali s -7514 105301 -7415 105349 4 VDD
port 41 nsew
rlabel locali s -7857 104985 -7704 105045 4 VDD
port 41 nsew
rlabel locali s -7969 104643 -7905 104653 4 VDD
port 41 nsew
rlabel locali s -8386 104653 -7905 104687 4 VDD
port 41 nsew
rlabel locali s -10967 104623 -10868 104671 4 VDD
port 41 nsew
rlabel locali s -7969 104687 -7905 104849 4 VDD
port 41 nsew
rlabel locali s -10967 104671 -10602 104705 4 VDD
port 41 nsew
rlabel locali s -10967 104705 -10868 104805 4 VDD
port 41 nsew
rlabel locali s -11310 104635 -11157 104805 4 VDD
port 41 nsew
rlabel locali s -8386 104849 -7905 104883 4 VDD
port 41 nsew
rlabel locali s -11310 104805 -10868 104867 4 VDD
port 41 nsew
rlabel locali s -7969 104883 -7905 105045 4 VDD
port 41 nsew
rlabel locali s -11310 104867 -10602 104901 4 VDD
port 41 nsew
rlabel locali s -11310 104901 -10868 104977 4 VDD
port 41 nsew
rlabel locali s -7864 105045 -7704 105082 4 VDD
port 41 nsew
rlabel locali s -8386 105045 -7905 105079 4 VDD
port 41 nsew
rlabel locali s -10967 104977 -10868 105063 4 VDD
port 41 nsew
rlabel locali s -7871 105082 -7704 105271 4 VDD
port 41 nsew
rlabel locali s -8019 105079 -7905 105085 4 VDD
port 41 nsew
rlabel locali s -8019 105085 -7920 105262 4 VDD
port 41 nsew
rlabel locali s -10967 105063 -10602 105097 4 VDD
port 41 nsew
rlabel locali s -10967 105097 -10868 105259 4 VDD
port 41 nsew
rlabel locali s -7857 105271 -7704 105641 4 VDD
port 41 nsew
rlabel locali s -7857 105641 -7658 105642 4 VDD
port 41 nsew
rlabel locali s -7857 105642 -7595 105652 4 VDD
port 41 nsew
rlabel locali s -7857 105652 -7178 105686 4 VDD
port 41 nsew
rlabel locali s -7857 105686 -7595 105848 4 VDD
port 41 nsew
rlabel locali s -7857 105848 -7178 105882 4 VDD
port 41 nsew
rlabel locali s -7857 105882 -7595 106044 4 VDD
port 41 nsew
rlabel locali s -8185 105262 -7920 105296 4 VDD
port 41 nsew
rlabel locali s -10967 105259 -10602 105293 4 VDD
port 41 nsew
rlabel locali s -8019 105296 -7920 105458 4 VDD
port 41 nsew
rlabel locali s -10967 105293 -10868 105341 4 VDD
port 41 nsew
rlabel locali s -11310 104977 -11157 105037 4 VDD
port 41 nsew
rlabel locali s -11422 104635 -11358 104645 4 VDD
port 41 nsew
rlabel locali s -11839 104645 -11358 104679 4 VDD
port 41 nsew
rlabel locali s -11422 104679 -11358 104841 4 VDD
port 41 nsew
rlabel locali s -11839 104841 -11358 104875 4 VDD
port 41 nsew
rlabel locali s -11422 104875 -11358 105037 4 VDD
port 41 nsew
rlabel locali s -11317 105037 -11157 105074 4 VDD
port 41 nsew
rlabel locali s -11839 105037 -11358 105071 4 VDD
port 41 nsew
rlabel locali s -11324 105074 -11157 105263 4 VDD
port 41 nsew
rlabel locali s -11472 105071 -11358 105077 4 VDD
port 41 nsew
rlabel locali s -11472 105077 -11373 105254 4 VDD
port 41 nsew
rlabel locali s -8185 105458 -7920 105492 4 VDD
port 41 nsew
rlabel locali s -8019 105492 -7920 105654 4 VDD
port 41 nsew
rlabel locali s -11310 105263 -11157 105633 4 VDD
port 41 nsew
rlabel locali s -11310 105633 -11111 105634 4 VDD
port 41 nsew
rlabel locali s -11310 105634 -11048 105644 4 VDD
port 41 nsew
rlabel locali s -8185 105654 -7920 105688 4 VDD
port 41 nsew
rlabel locali s -11310 105644 -10631 105678 4 VDD
port 41 nsew
rlabel locali s -8019 105688 -7920 105850 4 VDD
port 41 nsew
rlabel locali s -11310 105678 -11048 105840 4 VDD
port 41 nsew
rlabel locali s -8185 105850 -7920 105884 4 VDD
port 41 nsew
rlabel locali s -11310 105840 -10631 105874 4 VDD
port 41 nsew
rlabel locali s -8019 105884 -7920 105932 4 VDD
port 41 nsew
rlabel locali s -11310 105874 -11048 106036 4 VDD
port 41 nsew
rlabel locali s -11638 105254 -11373 105288 4 VDD
port 41 nsew
rlabel locali s -11472 105288 -11373 105450 4 VDD
port 41 nsew
rlabel locali s -11638 105450 -11373 105484 4 VDD
port 41 nsew
rlabel locali s -11472 105484 -11373 105646 4 VDD
port 41 nsew
rlabel locali s -11638 105646 -11373 105680 4 VDD
port 41 nsew
rlabel locali s -11472 105680 -11373 105842 4 VDD
port 41 nsew
rlabel locali s -11638 105842 -11373 105876 4 VDD
port 41 nsew
rlabel locali s -11472 105876 -11373 105924 4 VDD
port 41 nsew
rlabel locali s -7857 106044 -7178 106078 4 VDD
port 41 nsew
rlabel locali s -11310 106036 -10631 106070 4 VDD
port 41 nsew
rlabel locali s -7857 106078 -7545 106084 4 VDD
port 41 nsew
rlabel locali s -7644 106084 -7545 106261 4 VDD
port 41 nsew
rlabel locali s -7857 106084 -7687 106089 4 VDD
port 41 nsew
rlabel locali s -11310 106070 -10998 106076 4 VDD
port 41 nsew
rlabel locali s -7881 106089 -7687 106095 4 VDD
port 41 nsew
rlabel locali s -8007 106095 -7687 106100 4 VDD
port 41 nsew
rlabel locali s -8597 106100 -7687 106134 4 VDD
port 41 nsew
rlabel locali s -8007 106134 -7687 106140 4 VDD
port 41 nsew
rlabel locali s -7881 106140 -7687 106259 4 VDD
port 41 nsew
rlabel locali s -11097 106076 -10998 106253 4 VDD
port 41 nsew
rlabel locali s -11310 106076 -11140 106081 4 VDD
port 41 nsew
rlabel locali s -11334 106081 -11140 106087 4 VDD
port 41 nsew
rlabel locali s -11460 106087 -11140 106092 4 VDD
port 41 nsew
rlabel locali s -12050 106092 -11140 106126 4 VDD
port 41 nsew
rlabel locali s -11460 106126 -11140 106132 4 VDD
port 41 nsew
rlabel locali s -11334 106132 -11140 106251 4 VDD
port 41 nsew
rlabel locali s -7644 106261 -7379 106295 4 VDD
port 41 nsew
rlabel locali s -7644 106295 -7545 106457 4 VDD
port 41 nsew
rlabel locali s -7644 106457 -7379 106491 4 VDD
port 41 nsew
rlabel locali s -7644 106491 -7545 106653 4 VDD
port 41 nsew
rlabel locali s -7644 106653 -7379 106687 4 VDD
port 41 nsew
rlabel locali s -7644 106687 -7545 106849 4 VDD
port 41 nsew
rlabel locali s -7881 106259 -7704 106290 4 VDD
port 41 nsew
rlabel locali s -11097 106253 -10832 106287 4 VDD
port 41 nsew
rlabel locali s -8004 106290 -7704 106296 4 VDD
port 41 nsew
rlabel locali s -8597 106296 -7704 106330 4 VDD
port 41 nsew
rlabel locali s -8004 106330 -7704 106335 4 VDD
port 41 nsew
rlabel locali s -7881 106335 -7704 106712 4 VDD
port 41 nsew
rlabel locali s -11097 106287 -10998 106449 4 VDD
port 41 nsew
rlabel locali s -11097 106449 -10832 106483 4 VDD
port 41 nsew
rlabel locali s -11097 106483 -10998 106645 4 VDD
port 41 nsew
rlabel locali s -11097 106645 -10832 106679 4 VDD
port 41 nsew
rlabel locali s -8005 106712 -7704 106719 4 VDD
port 41 nsew
rlabel locali s -8597 106719 -7704 106753 4 VDD
port 41 nsew
rlabel locali s -8005 106753 -7704 106754 4 VDD
port 41 nsew
rlabel locali s -7644 106849 -7379 106883 4 VDD
port 41 nsew
rlabel locali s -8005 106754 -7815 106757 4 VDD
port 41 nsew
rlabel locali s -7881 106757 -7815 106858 4 VDD
port 41 nsew
rlabel locali s -11097 106679 -10998 106841 4 VDD
port 41 nsew
rlabel locali s -11334 106251 -11157 106282 4 VDD
port 41 nsew
rlabel locali s -11457 106282 -11157 106288 4 VDD
port 41 nsew
rlabel locali s -12050 106288 -11157 106322 4 VDD
port 41 nsew
rlabel locali s -11457 106322 -11157 106327 4 VDD
port 41 nsew
rlabel locali s -11334 106327 -11157 106704 4 VDD
port 41 nsew
rlabel locali s -11458 106704 -11157 106711 4 VDD
port 41 nsew
rlabel locali s -12050 106711 -11157 106745 4 VDD
port 41 nsew
rlabel locali s -11458 106745 -11157 106746 4 VDD
port 41 nsew
rlabel locali s -7644 106883 -7545 106931 4 VDD
port 41 nsew
rlabel locali s -7874 106858 -7822 106931 4 VDD
port 41 nsew
rlabel locali s -11097 106841 -10832 106875 4 VDD
port 41 nsew
rlabel locali s -11458 106746 -11268 106749 4 VDD
port 41 nsew
rlabel locali s -11334 106749 -11268 106850 4 VDD
port 41 nsew
rlabel locali s -11097 106875 -10998 106923 4 VDD
port 41 nsew
rlabel locali s -7888 106931 -7794 106993 4 VDD
port 41 nsew
rlabel locali s -7900 107159 -7774 107257 4 VDD
port 41 nsew
rlabel locali s -11306 107149 -11193 107166 4 VDD
port 41 nsew
rlabel locali s -11306 107166 -9826 107232 4 VDD
port 41 nsew
rlabel locali s -7894 107257 -7777 107722 4 VDD
port 41 nsew
rlabel locali s -9892 107232 -9826 107502 4 VDD
port 41 nsew
rlabel locali s -11306 107232 -11193 107233 4 VDD
port 41 nsew
rlabel locali s -11288 107502 -9826 107568 4 VDD
port 41 nsew
rlabel locali s -7894 107722 -7650 107839 4 VDD
port 41 nsew
rlabel locali s -7767 107839 -7650 108089 4 VDD
port 41 nsew
rlabel locali s -7862 108089 -7580 108092 4 VDD
port 41 nsew
rlabel locali s -8355 108092 -7580 108126 4 VDD
port 41 nsew
rlabel locali s -7862 108126 -7580 108127 4 VDD
port 41 nsew
rlabel locali s -7703 108127 -7580 108286 4 VDD
port 41 nsew
rlabel locali s -7860 108286 -7580 108288 4 VDD
port 41 nsew
rlabel locali s -8355 108288 -7580 108322 4 VDD
port 41 nsew
rlabel locali s -7860 108322 -7580 108324 4 VDD
port 41 nsew
rlabel locali s -7703 108324 -7580 108878 4 VDD
port 41 nsew
rlabel locali s -10998 108291 -10899 108339 4 VDD
port 41 nsew
rlabel locali s -11288 107568 -11222 108303 4 VDD
port 41 nsew
rlabel locali s -10998 108339 -10633 108373 4 VDD
port 41 nsew
rlabel locali s -10998 108373 -10899 108473 4 VDD
port 41 nsew
rlabel locali s -11341 108303 -11188 108473 4 VDD
port 41 nsew
rlabel locali s -11341 108473 -10899 108535 4 VDD
port 41 nsew
rlabel locali s -11341 108535 -10633 108569 4 VDD
port 41 nsew
rlabel locali s -11341 108569 -10899 108645 4 VDD
port 41 nsew
rlabel locali s -10998 108645 -10899 108731 4 VDD
port 41 nsew
rlabel locali s -10998 108731 -10633 108765 4 VDD
port 41 nsew
rlabel locali s -7883 108878 -7580 108883 4 VDD
port 41 nsew
rlabel locali s -8355 108883 -7580 108917 4 VDD
port 41 nsew
rlabel locali s -7883 108917 -7580 108928 4 VDD
port 41 nsew
rlabel locali s -10998 108765 -10899 108927 4 VDD
port 41 nsew
rlabel locali s -7703 108928 -7580 109004 4 VDD
port 41 nsew
rlabel locali s -10998 108927 -10633 108961 4 VDD
port 41 nsew
rlabel locali s -7880 109004 -7580 109013 4 VDD
port 41 nsew
rlabel locali s -10998 108961 -10899 109009 4 VDD
port 41 nsew
rlabel locali s -11341 108645 -11188 108705 4 VDD
port 41 nsew
rlabel locali s -11453 108303 -11389 108313 4 VDD
port 41 nsew
rlabel locali s -11870 108313 -11389 108347 4 VDD
port 41 nsew
rlabel locali s -11453 108347 -11389 108509 4 VDD
port 41 nsew
rlabel locali s -11870 108509 -11389 108543 4 VDD
port 41 nsew
rlabel locali s -11453 108543 -11389 108705 4 VDD
port 41 nsew
rlabel locali s -11348 108705 -11188 108742 4 VDD
port 41 nsew
rlabel locali s -11870 108705 -11389 108739 4 VDD
port 41 nsew
rlabel locali s -11355 108742 -11188 108931 4 VDD
port 41 nsew
rlabel locali s -11503 108739 -11389 108745 4 VDD
port 41 nsew
rlabel locali s -11503 108745 -11404 108922 4 VDD
port 41 nsew
rlabel locali s -8355 109013 -7580 109047 4 VDD
port 41 nsew
rlabel locali s -7880 109047 -7580 109054 4 VDD
port 41 nsew
rlabel locali s -7703 109054 -7580 109235 4 VDD
port 41 nsew
rlabel locali s -7865 109235 -7580 109241 4 VDD
port 41 nsew
rlabel locali s -8155 109241 -7580 109275 4 VDD
port 41 nsew
rlabel locali s -7865 109275 -7580 109278 4 VDD
port 41 nsew
rlabel locali s -7703 109278 -7580 109432 4 VDD
port 41 nsew
rlabel locali s -11341 108931 -11188 109301 4 VDD
port 41 nsew
rlabel locali s -11341 109301 -11142 109302 4 VDD
port 41 nsew
rlabel locali s -11341 109302 -11079 109312 4 VDD
port 41 nsew
rlabel locali s -11341 109312 -10662 109346 4 VDD
port 41 nsew
rlabel locali s -7863 109432 -7580 109436 4 VDD
port 41 nsew
rlabel locali s -7863 109436 -7421 109437 4 VDD
port 41 nsew
rlabel locali s -8155 109437 -7421 109471 4 VDD
port 41 nsew
rlabel locali s -7863 109471 -7421 109475 4 VDD
port 41 nsew
rlabel locali s -7763 109475 -7421 110399 4 VDD
port 41 nsew
rlabel locali s -11341 109346 -11079 109508 4 VDD
port 41 nsew
rlabel locali s -11341 109508 -10662 109542 4 VDD
port 41 nsew
rlabel locali s -11341 109542 -11079 109704 4 VDD
port 41 nsew
rlabel locali s -11669 108922 -11404 108956 4 VDD
port 41 nsew
rlabel locali s -11503 108956 -11404 109118 4 VDD
port 41 nsew
rlabel locali s -11669 109118 -11404 109152 4 VDD
port 41 nsew
rlabel locali s -11503 109152 -11404 109314 4 VDD
port 41 nsew
rlabel locali s -11669 109314 -11404 109348 4 VDD
port 41 nsew
rlabel locali s -11503 109348 -11404 109510 4 VDD
port 41 nsew
rlabel locali s -11669 109510 -11404 109544 4 VDD
port 41 nsew
rlabel locali s -11503 109544 -11404 109592 4 VDD
port 41 nsew
rlabel locali s -11341 109704 -10662 109738 4 VDD
port 41 nsew
rlabel locali s -11341 109738 -11029 109744 4 VDD
port 41 nsew
rlabel locali s -11128 109744 -11029 109921 4 VDD
port 41 nsew
rlabel locali s -11341 109744 -11171 109749 4 VDD
port 41 nsew
rlabel locali s -11365 109749 -11171 109755 4 VDD
port 41 nsew
rlabel locali s -11491 109755 -11171 109760 4 VDD
port 41 nsew
rlabel locali s -12081 109760 -11171 109794 4 VDD
port 41 nsew
rlabel locali s -11491 109794 -11171 109800 4 VDD
port 41 nsew
rlabel locali s -11365 109800 -11171 109919 4 VDD
port 41 nsew
rlabel locali s -11128 109921 -10863 109955 4 VDD
port 41 nsew
rlabel locali s -11128 109955 -11029 110117 4 VDD
port 41 nsew
rlabel locali s -11128 110117 -10863 110151 4 VDD
port 41 nsew
rlabel locali s -11128 110151 -11029 110313 4 VDD
port 41 nsew
rlabel locali s -11128 110313 -10863 110347 4 VDD
port 41 nsew
rlabel locali s -10221 110399 -7421 110521 4 VDD
port 41 nsew
rlabel locali s -11128 110347 -11029 110509 4 VDD
port 41 nsew
rlabel locali s -11365 109919 -11188 109950 4 VDD
port 41 nsew
rlabel locali s -11488 109950 -11188 109956 4 VDD
port 41 nsew
rlabel locali s -12081 109956 -11188 109990 4 VDD
port 41 nsew
rlabel locali s -11488 109990 -11188 109995 4 VDD
port 41 nsew
rlabel locali s -11365 109995 -11188 110372 4 VDD
port 41 nsew
rlabel locali s -11489 110372 -11188 110379 4 VDD
port 41 nsew
rlabel locali s -12081 110379 -11188 110413 4 VDD
port 41 nsew
rlabel locali s -11489 110413 -11188 110414 4 VDD
port 41 nsew
rlabel locali s -11489 110414 -11299 110417 4 VDD
port 41 nsew
rlabel locali s -11365 110417 -11299 110469 4 VDD
port 41 nsew
rlabel locali s -7763 110521 -7421 113995 4 VDD
port 41 nsew
rlabel locali s -10221 110521 -10099 110909 4 VDD
port 41 nsew
rlabel locali s -11128 110509 -10863 110543 4 VDD
port 41 nsew
rlabel locali s -11128 110543 -11029 110591 4 VDD
port 41 nsew
rlabel locali s -11365 110469 -11263 110518 4 VDD
port 41 nsew
rlabel locali s -11346 110518 -11263 110569 4 VDD
port 41 nsew
rlabel locali s -11371 110569 -11232 110648 4 VDD
port 41 nsew
rlabel locali s -11384 110819 -11217 110909 4 VDD
port 41 nsew
rlabel locali s -11384 110909 -10099 110958 4 VDD
port 41 nsew
rlabel locali s -11356 110958 -10099 111031 4 VDD
port 41 nsew
rlabel locali s -7763 113995 -7377 114007 4 VDD
port 41 nsew
rlabel locali s -7819 114007 -7377 114043 4 VDD
port 41 nsew
rlabel locali s -7819 114043 -7111 114077 4 VDD
port 41 nsew
rlabel locali s -7819 114077 -7377 114239 4 VDD
port 41 nsew
rlabel locali s -7819 114239 -7111 114273 4 VDD
port 41 nsew
rlabel locali s -7819 114273 -7377 114349 4 VDD
port 41 nsew
rlabel locali s -7476 114349 -7377 114435 4 VDD
port 41 nsew
rlabel locali s -7476 114435 -7111 114469 4 VDD
port 41 nsew
rlabel locali s -7476 114469 -7377 114631 4 VDD
port 41 nsew
rlabel locali s -7476 114631 -7111 114665 4 VDD
port 41 nsew
rlabel locali s -7476 114665 -7377 114713 4 VDD
port 41 nsew
rlabel locali s -7819 114349 -7666 114409 4 VDD
port 41 nsew
rlabel locali s -7931 114007 -7867 114017 4 VDD
port 41 nsew
rlabel locali s -8348 114017 -7867 114051 4 VDD
port 41 nsew
rlabel locali s -10929 113987 -10830 114035 4 VDD
port 41 nsew
rlabel locali s -7931 114051 -7867 114213 4 VDD
port 41 nsew
rlabel locali s -10929 114035 -10564 114069 4 VDD
port 41 nsew
rlabel locali s -10929 114069 -10830 114169 4 VDD
port 41 nsew
rlabel locali s -11272 113999 -11119 114169 4 VDD
port 41 nsew
rlabel locali s -8348 114213 -7867 114247 4 VDD
port 41 nsew
rlabel locali s -11272 114169 -10830 114231 4 VDD
port 41 nsew
rlabel locali s -7931 114247 -7867 114409 4 VDD
port 41 nsew
rlabel locali s -11272 114231 -10564 114265 4 VDD
port 41 nsew
rlabel locali s -11272 114265 -10830 114341 4 VDD
port 41 nsew
rlabel locali s -7826 114409 -7666 114446 4 VDD
port 41 nsew
rlabel locali s -8348 114409 -7867 114443 4 VDD
port 41 nsew
rlabel locali s -10929 114341 -10830 114427 4 VDD
port 41 nsew
rlabel locali s -7833 114446 -7666 114635 4 VDD
port 41 nsew
rlabel locali s -7981 114443 -7867 114449 4 VDD
port 41 nsew
rlabel locali s -7981 114449 -7882 114626 4 VDD
port 41 nsew
rlabel locali s -10929 114427 -10564 114461 4 VDD
port 41 nsew
rlabel locali s -10929 114461 -10830 114623 4 VDD
port 41 nsew
rlabel locali s -7819 114635 -7666 115005 4 VDD
port 41 nsew
rlabel locali s -7819 115005 -7620 115006 4 VDD
port 41 nsew
rlabel locali s -7819 115006 -7557 115016 4 VDD
port 41 nsew
rlabel locali s -7819 115016 -7140 115050 4 VDD
port 41 nsew
rlabel locali s -7819 115050 -7557 115212 4 VDD
port 41 nsew
rlabel locali s -7819 115212 -7140 115246 4 VDD
port 41 nsew
rlabel locali s -7819 115246 -7557 115408 4 VDD
port 41 nsew
rlabel locali s -8147 114626 -7882 114660 4 VDD
port 41 nsew
rlabel locali s -10929 114623 -10564 114657 4 VDD
port 41 nsew
rlabel locali s -7981 114660 -7882 114822 4 VDD
port 41 nsew
rlabel locali s -10929 114657 -10830 114705 4 VDD
port 41 nsew
rlabel locali s -11272 114341 -11119 114401 4 VDD
port 41 nsew
rlabel locali s -11384 113999 -11320 114009 4 VDD
port 41 nsew
rlabel locali s -11801 114009 -11320 114043 4 VDD
port 41 nsew
rlabel locali s -11384 114043 -11320 114205 4 VDD
port 41 nsew
rlabel locali s -11801 114205 -11320 114239 4 VDD
port 41 nsew
rlabel locali s -11384 114239 -11320 114401 4 VDD
port 41 nsew
rlabel locali s -11279 114401 -11119 114438 4 VDD
port 41 nsew
rlabel locali s -11801 114401 -11320 114435 4 VDD
port 41 nsew
rlabel locali s -11286 114438 -11119 114627 4 VDD
port 41 nsew
rlabel locali s -11434 114435 -11320 114441 4 VDD
port 41 nsew
rlabel locali s -11434 114441 -11335 114618 4 VDD
port 41 nsew
rlabel locali s -8147 114822 -7882 114856 4 VDD
port 41 nsew
rlabel locali s -7981 114856 -7882 115018 4 VDD
port 41 nsew
rlabel locali s -11272 114627 -11119 114997 4 VDD
port 41 nsew
rlabel locali s -11272 114997 -11073 114998 4 VDD
port 41 nsew
rlabel locali s -11272 114998 -11010 115008 4 VDD
port 41 nsew
rlabel locali s -8147 115018 -7882 115052 4 VDD
port 41 nsew
rlabel locali s -11272 115008 -10593 115042 4 VDD
port 41 nsew
rlabel locali s -7981 115052 -7882 115214 4 VDD
port 41 nsew
rlabel locali s -11272 115042 -11010 115204 4 VDD
port 41 nsew
rlabel locali s -8147 115214 -7882 115248 4 VDD
port 41 nsew
rlabel locali s -11272 115204 -10593 115238 4 VDD
port 41 nsew
rlabel locali s -7981 115248 -7882 115296 4 VDD
port 41 nsew
rlabel locali s -11272 115238 -11010 115400 4 VDD
port 41 nsew
rlabel locali s -11600 114618 -11335 114652 4 VDD
port 41 nsew
rlabel locali s -11434 114652 -11335 114814 4 VDD
port 41 nsew
rlabel locali s -11600 114814 -11335 114848 4 VDD
port 41 nsew
rlabel locali s -11434 114848 -11335 115010 4 VDD
port 41 nsew
rlabel locali s -11600 115010 -11335 115044 4 VDD
port 41 nsew
rlabel locali s -11434 115044 -11335 115206 4 VDD
port 41 nsew
rlabel locali s -11600 115206 -11335 115240 4 VDD
port 41 nsew
rlabel locali s -11434 115240 -11335 115288 4 VDD
port 41 nsew
rlabel locali s -7819 115408 -7140 115442 4 VDD
port 41 nsew
rlabel locali s -11272 115400 -10593 115434 4 VDD
port 41 nsew
rlabel locali s -7819 115442 -7507 115448 4 VDD
port 41 nsew
rlabel locali s -7606 115448 -7507 115625 4 VDD
port 41 nsew
rlabel locali s -7819 115448 -7649 115453 4 VDD
port 41 nsew
rlabel locali s -11272 115434 -10960 115440 4 VDD
port 41 nsew
rlabel locali s -7843 115453 -7649 115459 4 VDD
port 41 nsew
rlabel locali s -7969 115459 -7649 115464 4 VDD
port 41 nsew
rlabel locali s -8559 115464 -7649 115498 4 VDD
port 41 nsew
rlabel locali s -7969 115498 -7649 115504 4 VDD
port 41 nsew
rlabel locali s -7843 115504 -7649 115623 4 VDD
port 41 nsew
rlabel locali s -11059 115440 -10960 115617 4 VDD
port 41 nsew
rlabel locali s -11272 115440 -11102 115445 4 VDD
port 41 nsew
rlabel locali s -11296 115445 -11102 115451 4 VDD
port 41 nsew
rlabel locali s -11422 115451 -11102 115456 4 VDD
port 41 nsew
rlabel locali s -12012 115456 -11102 115490 4 VDD
port 41 nsew
rlabel locali s -11422 115490 -11102 115496 4 VDD
port 41 nsew
rlabel locali s -11296 115496 -11102 115615 4 VDD
port 41 nsew
rlabel locali s -7606 115625 -7341 115659 4 VDD
port 41 nsew
rlabel locali s -7606 115659 -7507 115821 4 VDD
port 41 nsew
rlabel locali s -7606 115821 -7341 115855 4 VDD
port 41 nsew
rlabel locali s -7606 115855 -7507 116017 4 VDD
port 41 nsew
rlabel locali s -7606 116017 -7341 116051 4 VDD
port 41 nsew
rlabel locali s -7606 116051 -7507 116213 4 VDD
port 41 nsew
rlabel locali s -7843 115623 -7666 115654 4 VDD
port 41 nsew
rlabel locali s -11059 115617 -10794 115651 4 VDD
port 41 nsew
rlabel locali s -7966 115654 -7666 115660 4 VDD
port 41 nsew
rlabel locali s -8559 115660 -7666 115694 4 VDD
port 41 nsew
rlabel locali s -7966 115694 -7666 115699 4 VDD
port 41 nsew
rlabel locali s -7843 115699 -7666 116076 4 VDD
port 41 nsew
rlabel locali s -11059 115651 -10960 115813 4 VDD
port 41 nsew
rlabel locali s -11059 115813 -10794 115847 4 VDD
port 41 nsew
rlabel locali s -11059 115847 -10960 116009 4 VDD
port 41 nsew
rlabel locali s -11059 116009 -10794 116043 4 VDD
port 41 nsew
rlabel locali s -7967 116076 -7666 116083 4 VDD
port 41 nsew
rlabel locali s -8559 116083 -7666 116117 4 VDD
port 41 nsew
rlabel locali s -7967 116117 -7666 116118 4 VDD
port 41 nsew
rlabel locali s -7606 116213 -7341 116247 4 VDD
port 41 nsew
rlabel locali s -7967 116118 -7777 116121 4 VDD
port 41 nsew
rlabel locali s -7843 116121 -7777 116222 4 VDD
port 41 nsew
rlabel locali s -11059 116043 -10960 116205 4 VDD
port 41 nsew
rlabel locali s -11296 115615 -11119 115646 4 VDD
port 41 nsew
rlabel locali s -11419 115646 -11119 115652 4 VDD
port 41 nsew
rlabel locali s -12012 115652 -11119 115686 4 VDD
port 41 nsew
rlabel locali s -11419 115686 -11119 115691 4 VDD
port 41 nsew
rlabel locali s -11296 115691 -11119 116068 4 VDD
port 41 nsew
rlabel locali s -11420 116068 -11119 116075 4 VDD
port 41 nsew
rlabel locali s -12012 116075 -11119 116109 4 VDD
port 41 nsew
rlabel locali s -11420 116109 -11119 116110 4 VDD
port 41 nsew
rlabel locali s -7606 116247 -7507 116295 4 VDD
port 41 nsew
rlabel locali s -7836 116222 -7784 116295 4 VDD
port 41 nsew
rlabel locali s -11059 116205 -10794 116239 4 VDD
port 41 nsew
rlabel locali s -11420 116110 -11230 116113 4 VDD
port 41 nsew
rlabel locali s -11296 116113 -11230 116214 4 VDD
port 41 nsew
rlabel locali s -11059 116239 -10960 116287 4 VDD
port 41 nsew
rlabel locali s -7850 116295 -7756 116357 4 VDD
port 41 nsew
rlabel locali s -7862 116523 -7736 116621 4 VDD
port 41 nsew
rlabel locali s -11268 116513 -11155 116530 4 VDD
port 41 nsew
rlabel locali s -11268 116530 -9788 116596 4 VDD
port 41 nsew
rlabel locali s -7856 116621 -7739 117086 4 VDD
port 41 nsew
rlabel locali s -9854 116596 -9788 116866 4 VDD
port 41 nsew
rlabel locali s -11268 116596 -11155 116597 4 VDD
port 41 nsew
rlabel locali s -11250 116866 -9788 116932 4 VDD
port 41 nsew
rlabel locali s -7856 117086 -7612 117203 4 VDD
port 41 nsew
rlabel locali s -7729 117203 -7612 117453 4 VDD
port 41 nsew
rlabel locali s -7824 117453 -7542 117456 4 VDD
port 41 nsew
rlabel locali s -8317 117456 -7542 117490 4 VDD
port 41 nsew
rlabel locali s -7824 117490 -7542 117491 4 VDD
port 41 nsew
rlabel locali s -7665 117491 -7542 117650 4 VDD
port 41 nsew
rlabel locali s -7822 117650 -7542 117652 4 VDD
port 41 nsew
rlabel locali s -8317 117652 -7542 117686 4 VDD
port 41 nsew
rlabel locali s -7822 117686 -7542 117688 4 VDD
port 41 nsew
rlabel locali s -7665 117688 -7542 118242 4 VDD
port 41 nsew
rlabel locali s -10960 117655 -10861 117703 4 VDD
port 41 nsew
rlabel locali s -11250 116932 -11184 117667 4 VDD
port 41 nsew
rlabel locali s -10960 117703 -10595 117737 4 VDD
port 41 nsew
rlabel locali s -10960 117737 -10861 117837 4 VDD
port 41 nsew
rlabel locali s -11303 117667 -11150 117837 4 VDD
port 41 nsew
rlabel locali s -11303 117837 -10861 117899 4 VDD
port 41 nsew
rlabel locali s -11303 117899 -10595 117933 4 VDD
port 41 nsew
rlabel locali s -11303 117933 -10861 118009 4 VDD
port 41 nsew
rlabel locali s -10960 118009 -10861 118095 4 VDD
port 41 nsew
rlabel locali s -10960 118095 -10595 118129 4 VDD
port 41 nsew
rlabel locali s -7845 118242 -7542 118247 4 VDD
port 41 nsew
rlabel locali s -8317 118247 -7542 118281 4 VDD
port 41 nsew
rlabel locali s -7845 118281 -7542 118292 4 VDD
port 41 nsew
rlabel locali s -10960 118129 -10861 118291 4 VDD
port 41 nsew
rlabel locali s -7665 118292 -7542 118368 4 VDD
port 41 nsew
rlabel locali s -10960 118291 -10595 118325 4 VDD
port 41 nsew
rlabel locali s -7842 118368 -7542 118377 4 VDD
port 41 nsew
rlabel locali s -10960 118325 -10861 118373 4 VDD
port 41 nsew
rlabel locali s -11303 118009 -11150 118069 4 VDD
port 41 nsew
rlabel locali s -11415 117667 -11351 117677 4 VDD
port 41 nsew
rlabel locali s -11832 117677 -11351 117711 4 VDD
port 41 nsew
rlabel locali s -11415 117711 -11351 117873 4 VDD
port 41 nsew
rlabel locali s -11832 117873 -11351 117907 4 VDD
port 41 nsew
rlabel locali s -11415 117907 -11351 118069 4 VDD
port 41 nsew
rlabel locali s -11310 118069 -11150 118106 4 VDD
port 41 nsew
rlabel locali s -11832 118069 -11351 118103 4 VDD
port 41 nsew
rlabel locali s -11317 118106 -11150 118295 4 VDD
port 41 nsew
rlabel locali s -11465 118103 -11351 118109 4 VDD
port 41 nsew
rlabel locali s -11465 118109 -11366 118286 4 VDD
port 41 nsew
rlabel locali s -8317 118377 -7542 118411 4 VDD
port 41 nsew
rlabel locali s -7842 118411 -7542 118418 4 VDD
port 41 nsew
rlabel locali s -7665 118418 -7542 118599 4 VDD
port 41 nsew
rlabel locali s -7827 118599 -7542 118605 4 VDD
port 41 nsew
rlabel locali s -8117 118605 -7542 118639 4 VDD
port 41 nsew
rlabel locali s -7827 118639 -7542 118642 4 VDD
port 41 nsew
rlabel locali s -7665 118642 -7542 118796 4 VDD
port 41 nsew
rlabel locali s -11303 118295 -11150 118665 4 VDD
port 41 nsew
rlabel locali s -11303 118665 -11104 118666 4 VDD
port 41 nsew
rlabel locali s -11303 118666 -11041 118676 4 VDD
port 41 nsew
rlabel locali s -11303 118676 -10624 118710 4 VDD
port 41 nsew
rlabel locali s -7825 118796 -7542 118801 4 VDD
port 41 nsew
rlabel locali s -8117 118801 -7542 118835 4 VDD
port 41 nsew
rlabel locali s -7825 118835 -7542 118839 4 VDD
port 41 nsew
rlabel locali s -7664 118839 -7542 119211 4 VDD
port 41 nsew
rlabel locali s -11303 118710 -11041 118872 4 VDD
port 41 nsew
rlabel locali s -11303 118872 -10624 118906 4 VDD
port 41 nsew
rlabel locali s -11303 118906 -11041 119068 4 VDD
port 41 nsew
rlabel locali s -11631 118286 -11366 118320 4 VDD
port 41 nsew
rlabel locali s -11465 118320 -11366 118482 4 VDD
port 41 nsew
rlabel locali s -11631 118482 -11366 118516 4 VDD
port 41 nsew
rlabel locali s -11465 118516 -11366 118678 4 VDD
port 41 nsew
rlabel locali s -11631 118678 -11366 118712 4 VDD
port 41 nsew
rlabel locali s -11465 118712 -11366 118874 4 VDD
port 41 nsew
rlabel locali s -11631 118874 -11366 118908 4 VDD
port 41 nsew
rlabel locali s -11465 118908 -11366 118956 4 VDD
port 41 nsew
rlabel locali s -11303 119068 -10624 119102 4 VDD
port 41 nsew
rlabel locali s -7664 119211 -2527 119686 4 VDD
port 41 nsew
rlabel locali s -11303 119102 -10991 119108 4 VDD
port 41 nsew
rlabel locali s -11090 119108 -10991 119285 4 VDD
port 41 nsew
rlabel locali s -11303 119108 -11133 119113 4 VDD
port 41 nsew
rlabel locali s -11327 119113 -11133 119119 4 VDD
port 41 nsew
rlabel locali s -11453 119119 -11133 119124 4 VDD
port 41 nsew
rlabel locali s -12043 119124 -11133 119158 4 VDD
port 41 nsew
rlabel locali s -11453 119158 -11133 119164 4 VDD
port 41 nsew
rlabel locali s -11327 119164 -11133 119283 4 VDD
port 41 nsew
rlabel locali s -11090 119285 -10825 119319 4 VDD
port 41 nsew
rlabel locali s -11090 119319 -10991 119481 4 VDD
port 41 nsew
rlabel locali s -11090 119481 -10825 119515 4 VDD
port 41 nsew
rlabel locali s -11090 119515 -10991 119677 4 VDD
port 41 nsew
rlabel locali s -7664 119686 -7542 119763 4 VDD
port 41 nsew
rlabel locali s -11090 119677 -10825 119711 4 VDD
port 41 nsew
rlabel locali s -10183 119763 -7542 119885 4 VDD
port 41 nsew
rlabel locali s -11090 119711 -10991 119873 4 VDD
port 41 nsew
rlabel locali s -11327 119283 -11150 119314 4 VDD
port 41 nsew
rlabel locali s -11450 119314 -11150 119320 4 VDD
port 41 nsew
rlabel locali s -12043 119320 -11150 119354 4 VDD
port 41 nsew
rlabel locali s -11450 119354 -11150 119359 4 VDD
port 41 nsew
rlabel locali s -11327 119359 -11150 119736 4 VDD
port 41 nsew
rlabel locali s -11451 119736 -11150 119743 4 VDD
port 41 nsew
rlabel locali s -12043 119743 -11150 119777 4 VDD
port 41 nsew
rlabel locali s -11451 119777 -11150 119778 4 VDD
port 41 nsew
rlabel locali s -11451 119778 -11261 119781 4 VDD
port 41 nsew
rlabel locali s -11327 119781 -11261 119833 4 VDD
port 41 nsew
rlabel locali s -10183 119885 -10061 120273 4 VDD
port 41 nsew
rlabel locali s -11090 119873 -10825 119907 4 VDD
port 41 nsew
rlabel locali s -11090 119907 -10991 119955 4 VDD
port 41 nsew
rlabel locali s -11327 119833 -11225 119882 4 VDD
port 41 nsew
rlabel locali s -11308 119882 -11225 119933 4 VDD
port 41 nsew
rlabel locali s -11333 119933 -11194 120012 4 VDD
port 41 nsew
rlabel locali s -11346 120183 -11179 120273 4 VDD
port 41 nsew
rlabel locali s -11346 120273 -10061 120322 4 VDD
port 41 nsew
rlabel locali s -11318 120322 -10061 120395 4 VDD
port 41 nsew
rlabel nwell s -21569 -62326 -20144 -62325 2 VDD
port 41 nsew
rlabel nwell s 15134 -62072 17870 -62071 8 VDD
port 41 nsew
rlabel nwell s 12808 -62071 17870 -61618 8 VDD
port 41 nsew
rlabel nwell s 6907 -62256 8825 -61854 8 VDD
port 41 nsew
rlabel nwell s 3907 -62256 5825 -61854 8 VDD
port 41 nsew
rlabel nwell s 1407 -62256 3325 -61854 8 VDD
port 41 nsew
rlabel nwell s -1093 -62256 825 -61854 2 VDD
port 41 nsew
rlabel nwell s -3593 -62256 -1675 -61854 2 VDD
port 41 nsew
rlabel nwell s -6093 -62256 -4175 -61854 2 VDD
port 41 nsew
rlabel nwell s -21600 -62325 -20144 -61867 2 VDD
port 41 nsew
rlabel nwell s 6908 -61854 8825 -61781 8 VDD
port 41 nsew
rlabel nwell s 3908 -61854 5825 -61781 8 VDD
port 41 nsew
rlabel nwell s 1408 -61854 3325 -61781 8 VDD
port 41 nsew
rlabel nwell s -1092 -61854 825 -61781 2 VDD
port 41 nsew
rlabel nwell s -3592 -61854 -1675 -61781 2 VDD
port 41 nsew
rlabel nwell s -6092 -61854 -4175 -61781 2 VDD
port 41 nsew
rlabel nwell s 14328 -61618 15169 -61612 8 VDD
port 41 nsew
rlabel nwell s -16751 -61232 -16229 -61217 2 VDD
port 41 nsew
rlabel nwell s -17724 -61261 -17006 -61217 2 VDD
port 41 nsew
rlabel nwell s -17724 -61217 -16229 -61038 2 VDD
port 41 nsew
rlabel nwell s -17724 -61038 -16142 -61031 2 VDD
port 41 nsew
rlabel nwell s -17724 -61031 -15424 -60851 2 VDD
port 41 nsew
rlabel nwell s -17750 -60851 -15424 -60657 2 VDD
port 41 nsew
rlabel nwell s 12529 -60635 12870 -60624 8 VDD
port 41 nsew
rlabel nwell s 87164 -60334 88011 -59929 8 VDD
port 41 nsew
rlabel nwell s 85717 -60123 86239 -59929 8 VDD
port 41 nsew
rlabel nwell s 86946 -59929 88011 -59922 8 VDD
port 41 nsew
rlabel nwell s 85717 -59929 86326 -59922 8 VDD
port 41 nsew
rlabel nwell s 85717 -59922 88011 -59374 8 VDD
port 41 nsew
rlabel nwell s 85717 -59374 88043 -59180 8 VDD
port 41 nsew
rlabel nwell s 83496 -60303 84343 -59898 8 VDD
port 41 nsew
rlabel nwell s 82049 -60092 82571 -59898 8 VDD
port 41 nsew
rlabel nwell s 83278 -59898 84343 -59891 8 VDD
port 41 nsew
rlabel nwell s 82049 -59898 82658 -59891 8 VDD
port 41 nsew
rlabel nwell s 82049 -59891 84343 -59343 8 VDD
port 41 nsew
rlabel nwell s 77800 -60372 78647 -59967 8 VDD
port 41 nsew
rlabel nwell s 76353 -60161 76875 -59967 8 VDD
port 41 nsew
rlabel nwell s 77582 -59967 78647 -59960 8 VDD
port 41 nsew
rlabel nwell s 76353 -59967 76962 -59960 8 VDD
port 41 nsew
rlabel nwell s 76353 -59960 78647 -59412 8 VDD
port 41 nsew
rlabel nwell s 85743 -59180 88043 -59000 8 VDD
port 41 nsew
rlabel nwell s 85743 -59000 87325 -58993 8 VDD
port 41 nsew
rlabel nwell s 85743 -58993 87238 -58814 8 VDD
port 41 nsew
rlabel nwell s 82049 -59343 84375 -59149 8 VDD
port 41 nsew
rlabel nwell s 76353 -59412 78679 -59218 8 VDD
port 41 nsew
rlabel nwell s 74132 -60341 74979 -59936 8 VDD
port 41 nsew
rlabel nwell s 72685 -60130 73207 -59936 8 VDD
port 41 nsew
rlabel nwell s 73914 -59936 74979 -59929 8 VDD
port 41 nsew
rlabel nwell s 72685 -59936 73294 -59929 8 VDD
port 41 nsew
rlabel nwell s 72685 -59929 74979 -59381 8 VDD
port 41 nsew
rlabel nwell s 68647 -60389 69494 -59984 8 VDD
port 41 nsew
rlabel nwell s 67200 -60178 67722 -59984 8 VDD
port 41 nsew
rlabel nwell s 68429 -59984 69494 -59977 8 VDD
port 41 nsew
rlabel nwell s 67200 -59984 67809 -59977 8 VDD
port 41 nsew
rlabel nwell s 67200 -59977 69494 -59429 8 VDD
port 41 nsew
rlabel nwell s 82075 -59149 84375 -58969 8 VDD
port 41 nsew
rlabel nwell s 76379 -59218 78679 -59038 8 VDD
port 41 nsew
rlabel nwell s 76379 -59038 77961 -59031 8 VDD
port 41 nsew
rlabel nwell s 82075 -58969 83657 -58962 8 VDD
port 41 nsew
rlabel nwell s 86716 -58814 87238 -58799 8 VDD
port 41 nsew
rlabel nwell s 85743 -58814 86461 -58770 8 VDD
port 41 nsew
rlabel nwell s 82075 -58962 83570 -58783 8 VDD
port 41 nsew
rlabel nwell s 76379 -59031 77874 -58852 8 VDD
port 41 nsew
rlabel nwell s 72685 -59381 75011 -59187 8 VDD
port 41 nsew
rlabel nwell s 67200 -59429 69526 -59235 8 VDD
port 41 nsew
rlabel nwell s 64979 -60358 65826 -59953 8 VDD
port 41 nsew
rlabel nwell s 63532 -60147 64054 -59953 8 VDD
port 41 nsew
rlabel nwell s 64761 -59953 65826 -59946 8 VDD
port 41 nsew
rlabel nwell s 63532 -59953 64141 -59946 8 VDD
port 41 nsew
rlabel nwell s 63532 -59946 65826 -59398 8 VDD
port 41 nsew
rlabel nwell s 59893 -60455 60740 -60050 8 VDD
port 41 nsew
rlabel nwell s 58446 -60244 58968 -60050 8 VDD
port 41 nsew
rlabel nwell s 59675 -60050 60740 -60043 8 VDD
port 41 nsew
rlabel nwell s 58446 -60050 59055 -60043 8 VDD
port 41 nsew
rlabel nwell s 58446 -60043 60740 -59495 8 VDD
port 41 nsew
rlabel nwell s 72711 -59187 75011 -59007 8 VDD
port 41 nsew
rlabel nwell s 67226 -59235 69526 -59055 8 VDD
port 41 nsew
rlabel nwell s 67226 -59055 68808 -59048 8 VDD
port 41 nsew
rlabel nwell s 72711 -59007 74293 -59000 8 VDD
port 41 nsew
rlabel nwell s 77352 -58852 77874 -58837 8 VDD
port 41 nsew
rlabel nwell s 76379 -58852 77097 -58808 8 VDD
port 41 nsew
rlabel nwell s 72711 -59000 74206 -58821 8 VDD
port 41 nsew
rlabel nwell s 67226 -59048 68721 -58869 8 VDD
port 41 nsew
rlabel nwell s 63532 -59398 65858 -59204 8 VDD
port 41 nsew
rlabel nwell s 58446 -59495 60772 -59301 8 VDD
port 41 nsew
rlabel nwell s 56225 -60424 57072 -60019 8 VDD
port 41 nsew
rlabel nwell s 54778 -60213 55300 -60019 8 VDD
port 41 nsew
rlabel nwell s 56007 -60019 57072 -60012 8 VDD
port 41 nsew
rlabel nwell s 54778 -60019 55387 -60012 8 VDD
port 41 nsew
rlabel nwell s 54778 -60012 57072 -59464 8 VDD
port 41 nsew
rlabel nwell s 50695 -60489 51542 -60084 8 VDD
port 41 nsew
rlabel nwell s 49248 -60278 49770 -60084 8 VDD
port 41 nsew
rlabel nwell s 50477 -60084 51542 -60077 8 VDD
port 41 nsew
rlabel nwell s 49248 -60084 49857 -60077 8 VDD
port 41 nsew
rlabel nwell s 49248 -60077 51542 -59529 8 VDD
port 41 nsew
rlabel nwell s 63558 -59204 65858 -59024 8 VDD
port 41 nsew
rlabel nwell s 58472 -59301 60772 -59121 8 VDD
port 41 nsew
rlabel nwell s 58472 -59121 60054 -59114 8 VDD
port 41 nsew
rlabel nwell s 63558 -59024 65140 -59017 8 VDD
port 41 nsew
rlabel nwell s 68199 -58869 68721 -58854 8 VDD
port 41 nsew
rlabel nwell s 67226 -58869 67944 -58825 8 VDD
port 41 nsew
rlabel nwell s 63558 -59017 65053 -58838 8 VDD
port 41 nsew
rlabel nwell s 58472 -59114 59967 -58935 8 VDD
port 41 nsew
rlabel nwell s 54778 -59464 57104 -59270 8 VDD
port 41 nsew
rlabel nwell s 49248 -59529 51574 -59335 8 VDD
port 41 nsew
rlabel nwell s 47027 -60458 47874 -60053 8 VDD
port 41 nsew
rlabel nwell s 45580 -60247 46102 -60053 8 VDD
port 41 nsew
rlabel nwell s 46809 -60053 47874 -60046 8 VDD
port 41 nsew
rlabel nwell s 45580 -60053 46189 -60046 8 VDD
port 41 nsew
rlabel nwell s 45580 -60046 47874 -59498 8 VDD
port 41 nsew
rlabel nwell s 54804 -59270 57104 -59090 8 VDD
port 41 nsew
rlabel nwell s 49274 -59335 51574 -59155 8 VDD
port 41 nsew
rlabel nwell s 49274 -59155 50856 -59148 8 VDD
port 41 nsew
rlabel nwell s 54804 -59090 56386 -59083 8 VDD
port 41 nsew
rlabel nwell s 59445 -58935 59967 -58920 8 VDD
port 41 nsew
rlabel nwell s 58472 -58935 59190 -58891 8 VDD
port 41 nsew
rlabel nwell s 54804 -59083 56299 -58904 8 VDD
port 41 nsew
rlabel nwell s 49274 -59148 50769 -58969 8 VDD
port 41 nsew
rlabel nwell s 45580 -59498 47906 -59304 8 VDD
port 41 nsew
rlabel nwell s 41832 -60450 42679 -60045 8 VDD
port 41 nsew
rlabel nwell s 40385 -60239 40907 -60045 8 VDD
port 41 nsew
rlabel nwell s 41614 -60045 42679 -60038 8 VDD
port 41 nsew
rlabel nwell s 40385 -60045 40994 -60038 8 VDD
port 41 nsew
rlabel nwell s 40385 -60038 42679 -59490 8 VDD
port 41 nsew
rlabel nwell s 45606 -59304 47906 -59124 8 VDD
port 41 nsew
rlabel nwell s 45606 -59124 47188 -59117 8 VDD
port 41 nsew
rlabel nwell s 50247 -58969 50769 -58954 8 VDD
port 41 nsew
rlabel nwell s 49274 -58969 49992 -58925 8 VDD
port 41 nsew
rlabel nwell s 45606 -59117 47101 -58938 8 VDD
port 41 nsew
rlabel nwell s 40385 -59490 42711 -59296 8 VDD
port 41 nsew
rlabel nwell s 38164 -60419 39011 -60014 8 VDD
port 41 nsew
rlabel nwell s 36717 -60208 37239 -60014 8 VDD
port 41 nsew
rlabel nwell s 37946 -60014 39011 -60007 8 VDD
port 41 nsew
rlabel nwell s 36717 -60014 37326 -60007 8 VDD
port 41 nsew
rlabel nwell s 36717 -60007 39011 -59459 8 VDD
port 41 nsew
rlabel nwell s 33392 -60439 34239 -60034 8 VDD
port 41 nsew
rlabel nwell s 31945 -60228 32467 -60034 8 VDD
port 41 nsew
rlabel nwell s 33174 -60034 34239 -60027 8 VDD
port 41 nsew
rlabel nwell s 31945 -60034 32554 -60027 8 VDD
port 41 nsew
rlabel nwell s 31945 -60027 34239 -59479 8 VDD
port 41 nsew
rlabel nwell s 40411 -59296 42711 -59116 8 VDD
port 41 nsew
rlabel nwell s 40411 -59116 41993 -59109 8 VDD
port 41 nsew
rlabel nwell s 46579 -58938 47101 -58923 8 VDD
port 41 nsew
rlabel nwell s 55777 -58904 56299 -58889 8 VDD
port 41 nsew
rlabel nwell s 54804 -58904 55522 -58860 8 VDD
port 41 nsew
rlabel nwell s 45606 -58938 46324 -58894 8 VDD
port 41 nsew
rlabel nwell s 40411 -59109 41906 -58930 8 VDD
port 41 nsew
rlabel nwell s 36717 -59459 39043 -59265 8 VDD
port 41 nsew
rlabel nwell s 31945 -59479 34271 -59285 8 VDD
port 41 nsew
rlabel nwell s 29724 -60408 30571 -60003 8 VDD
port 41 nsew
rlabel nwell s 28277 -60197 28799 -60003 8 VDD
port 41 nsew
rlabel nwell s 11925 -60624 17883 -60171 8 VDD
port 41 nsew
rlabel nwell s 15147 -60171 17883 -60170 8 VDD
port 41 nsew
rlabel nwell s -17750 -60657 -15456 -60109 2 VDD
port 41 nsew
rlabel nwell s -16521 -60109 -15456 -60102 2 VDD
port 41 nsew
rlabel nwell s -17750 -60109 -17141 -60102 2 VDD
port 41 nsew
rlabel nwell s 29506 -60003 30571 -59996 8 VDD
port 41 nsew
rlabel nwell s 28277 -60003 28886 -59996 8 VDD
port 41 nsew
rlabel nwell s 28277 -59996 30571 -59448 8 VDD
port 41 nsew
rlabel nwell s 20589 -59781 22014 -59780 8 VDD
port 41 nsew
rlabel nwell s 36743 -59265 39043 -59085 8 VDD
port 41 nsew
rlabel nwell s 31971 -59285 34271 -59105 8 VDD
port 41 nsew
rlabel nwell s 31971 -59105 33553 -59098 8 VDD
port 41 nsew
rlabel nwell s 36743 -59085 38325 -59078 8 VDD
port 41 nsew
rlabel nwell s 41384 -58930 41906 -58915 8 VDD
port 41 nsew
rlabel nwell s 40411 -58930 41129 -58886 8 VDD
port 41 nsew
rlabel nwell s 36743 -59078 38238 -58899 8 VDD
port 41 nsew
rlabel nwell s 31971 -59098 33466 -58919 8 VDD
port 41 nsew
rlabel nwell s 28277 -59448 30603 -59254 8 VDD
port 41 nsew
rlabel nwell s 28303 -59254 30603 -59074 8 VDD
port 41 nsew
rlabel nwell s 28303 -59074 29885 -59067 8 VDD
port 41 nsew
rlabel nwell s 32944 -58919 33466 -58904 8 VDD
port 41 nsew
rlabel nwell s 37716 -58899 38238 -58884 8 VDD
port 41 nsew
rlabel nwell s 36743 -58899 37461 -58855 8 VDD
port 41 nsew
rlabel nwell s 31971 -58919 32689 -58875 8 VDD
port 41 nsew
rlabel nwell s 28303 -59067 29798 -58888 8 VDD
port 41 nsew
rlabel nwell s 29276 -58888 29798 -58873 8 VDD
port 41 nsew
rlabel nwell s 28303 -58888 29021 -58844 8 VDD
port 41 nsew
rlabel nwell s 64531 -58838 65053 -58823 8 VDD
port 41 nsew
rlabel nwell s 73684 -58821 74206 -58806 8 VDD
port 41 nsew
rlabel nwell s 83048 -58783 83570 -58768 8 VDD
port 41 nsew
rlabel nwell s 82075 -58783 82793 -58739 8 VDD
port 41 nsew
rlabel nwell s 72711 -58821 73429 -58777 8 VDD
port 41 nsew
rlabel nwell s 63558 -58838 64276 -58794 8 VDD
port 41 nsew
rlabel nwell s 23328 -59776 26054 -58744 8 VDD
port 41 nsew
rlabel nwell s 22448 -59768 23068 -59315 8 VDD
port 41 nsew
rlabel nwell s 20589 -59780 22045 -59322 8 VDD
port 41 nsew
rlabel nwell s 19673 -59769 20308 -59088 8 VDD
port 41 nsew
rlabel nwell s 18727 -59769 19362 -59088 8 VDD
port 41 nsew
rlabel nwell s -5925 -60005 8835 -59619 8 VDD
port 41 nsew
rlabel nwell s -13799 -59736 -11063 -59735 2 VDD
port 41 nsew
rlabel nwell s 2696 -59619 8835 -59617 8 VDD
port 41 nsew
rlabel nwell s 4301 -59617 8835 -59610 8 VDD
port 41 nsew
rlabel nwell s 2696 -59617 3305 -59612 8 VDD
port 41 nsew
rlabel nwell s 4388 -59610 8835 -59530 8 VDD
port 41 nsew
rlabel nwell s 4388 -59530 4910 -59416 8 VDD
port 41 nsew
rlabel nwell s 2783 -59612 3305 -59418 8 VDD
port 41 nsew
rlabel nwell s -5925 -59619 1701 -59549 2 VDD
port 41 nsew
rlabel nwell s -285 -59549 1701 -59532 8 VDD
port 41 nsew
rlabel nwell s -912 -59549 -571 -59538 2 VDD
port 41 nsew
rlabel nwell s -13799 -59735 -7841 -59282 2 VDD
port 41 nsew
rlabel nwell s -16303 -60102 -15456 -59697 2 VDD
port 41 nsew
rlabel nwell s -17750 -60102 -17228 -59908 2 VDD
port 41 nsew
rlabel nwell s -8786 -59282 -8445 -59271 2 VDD
port 41 nsew
rlabel nwell s -19152 -59503 -18517 -58822 2 VDD
port 41 nsew
rlabel nwell s -20057 -59502 -19422 -58821 2 VDD
port 41 nsew
rlabel nwell s -21263 -59773 -20318 -58828 2 VDD
port 41 nsew
rlabel nwell s -3211 -58561 -2370 -58555 2 VDD
port 41 nsew
rlabel nwell s 22498 -58338 23020 -57784 8 VDD
port 41 nsew
rlabel nwell s -5912 -58555 -850 -58102 2 VDD
port 41 nsew
rlabel nwell s -5912 -58102 -3176 -58101 2 VDD
port 41 nsew
rlabel nwell s -7495 -58705 -6648 -57828 2 VDD
port 41 nsew
rlabel nwell s -11085 -58294 -10244 -58288 2 VDD
port 41 nsew
rlabel nwell s -13786 -58288 -8724 -57835 2 VDD
port 41 nsew
rlabel nwell s -13786 -57835 -11050 -57834 2 VDD
port 41 nsew
rlabel nwell s 23275 -57516 26011 -57515 8 VDD
port 41 nsew
rlabel nwell s 22487 -57784 23020 -57515 8 VDD
port 41 nsew
rlabel nwell s 18731 -57515 26011 -57062 8 VDD
port 41 nsew
rlabel nwell s -5912 -57247 -3176 -57246 2 VDD
port 41 nsew
rlabel nwell s 20657 -57062 20998 -57051 8 VDD
port 41 nsew
rlabel nwell s 85496 -56608 86973 -55735 8 VDD
port 41 nsew
rlabel nwell s 83504 -56850 84351 -56445 8 VDD
port 41 nsew
rlabel nwell s 82057 -56639 82579 -56445 8 VDD
port 41 nsew
rlabel nwell s 83286 -56445 84351 -56438 8 VDD
port 41 nsew
rlabel nwell s 82057 -56445 82666 -56438 8 VDD
port 41 nsew
rlabel nwell s 82057 -56438 84351 -55890 8 VDD
port 41 nsew
rlabel nwell s 82057 -55890 84383 -55696 8 VDD
port 41 nsew
rlabel nwell s 76132 -56646 77609 -55773 8 VDD
port 41 nsew
rlabel nwell s 74140 -56888 74987 -56483 8 VDD
port 41 nsew
rlabel nwell s 72693 -56677 73215 -56483 8 VDD
port 41 nsew
rlabel nwell s 73922 -56483 74987 -56476 8 VDD
port 41 nsew
rlabel nwell s 72693 -56483 73302 -56476 8 VDD
port 41 nsew
rlabel nwell s 72693 -56476 74987 -55928 8 VDD
port 41 nsew
rlabel nwell s 72693 -55928 75019 -55734 8 VDD
port 41 nsew
rlabel nwell s 66979 -56663 68456 -55790 8 VDD
port 41 nsew
rlabel nwell s 64987 -56905 65834 -56500 8 VDD
port 41 nsew
rlabel nwell s 63540 -56694 64062 -56500 8 VDD
port 41 nsew
rlabel nwell s 64769 -56500 65834 -56493 8 VDD
port 41 nsew
rlabel nwell s 63540 -56500 64149 -56493 8 VDD
port 41 nsew
rlabel nwell s 63540 -56493 65834 -55945 8 VDD
port 41 nsew
rlabel nwell s 63540 -55945 65866 -55751 8 VDD
port 41 nsew
rlabel nwell s 58225 -56729 59702 -55856 8 VDD
port 41 nsew
rlabel nwell s 56233 -56971 57080 -56566 8 VDD
port 41 nsew
rlabel nwell s 54786 -56760 55308 -56566 8 VDD
port 41 nsew
rlabel nwell s 56015 -56566 57080 -56559 8 VDD
port 41 nsew
rlabel nwell s 54786 -56566 55395 -56559 8 VDD
port 41 nsew
rlabel nwell s 54786 -56559 57080 -56011 8 VDD
port 41 nsew
rlabel nwell s 54786 -56011 57112 -55817 8 VDD
port 41 nsew
rlabel nwell s 49027 -56763 50504 -55890 8 VDD
port 41 nsew
rlabel nwell s 47035 -57005 47882 -56600 8 VDD
port 41 nsew
rlabel nwell s 45588 -56794 46110 -56600 8 VDD
port 41 nsew
rlabel nwell s 46817 -56600 47882 -56593 8 VDD
port 41 nsew
rlabel nwell s 45588 -56600 46197 -56593 8 VDD
port 41 nsew
rlabel nwell s 45588 -56593 47882 -56045 8 VDD
port 41 nsew
rlabel nwell s 45588 -56045 47914 -55851 8 VDD
port 41 nsew
rlabel nwell s 40164 -56724 41641 -55851 8 VDD
port 41 nsew
rlabel nwell s 38172 -56966 39019 -56561 8 VDD
port 41 nsew
rlabel nwell s 36725 -56755 37247 -56561 8 VDD
port 41 nsew
rlabel nwell s 37954 -56561 39019 -56554 8 VDD
port 41 nsew
rlabel nwell s 36725 -56561 37334 -56554 8 VDD
port 41 nsew
rlabel nwell s 36725 -56554 39019 -56006 8 VDD
port 41 nsew
rlabel nwell s 82083 -55696 84383 -55516 8 VDD
port 41 nsew
rlabel nwell s 72719 -55734 75019 -55554 8 VDD
port 41 nsew
rlabel nwell s 63566 -55751 65866 -55571 8 VDD
port 41 nsew
rlabel nwell s 54812 -55817 57112 -55637 8 VDD
port 41 nsew
rlabel nwell s 45614 -55851 47914 -55671 8 VDD
port 41 nsew
rlabel nwell s 45614 -55671 47196 -55664 8 VDD
port 41 nsew
rlabel nwell s 54812 -55637 56394 -55630 8 VDD
port 41 nsew
rlabel nwell s 63566 -55571 65148 -55564 8 VDD
port 41 nsew
rlabel nwell s 72719 -55554 74301 -55547 8 VDD
port 41 nsew
rlabel nwell s 82083 -55516 83665 -55509 8 VDD
port 41 nsew
rlabel nwell s 82083 -55509 83578 -55330 8 VDD
port 41 nsew
rlabel nwell s 72719 -55547 74214 -55368 8 VDD
port 41 nsew
rlabel nwell s 63566 -55564 65061 -55385 8 VDD
port 41 nsew
rlabel nwell s 54812 -55630 56307 -55451 8 VDD
port 41 nsew
rlabel nwell s 45614 -55664 47109 -55485 8 VDD
port 41 nsew
rlabel nwell s 36725 -56006 39051 -55812 8 VDD
port 41 nsew
rlabel nwell s 31724 -56713 33201 -55840 8 VDD
port 41 nsew
rlabel nwell s 29732 -56955 30579 -56550 8 VDD
port 41 nsew
rlabel nwell s 28285 -56744 28807 -56550 8 VDD
port 41 nsew
rlabel nwell s 29514 -56550 30579 -56543 8 VDD
port 41 nsew
rlabel nwell s 28285 -56550 28894 -56543 8 VDD
port 41 nsew
rlabel nwell s 28285 -56543 30579 -55995 8 VDD
port 41 nsew
rlabel nwell s 18732 -57062 19677 -56542 8 VDD
port 41 nsew
rlabel nwell s -5912 -57246 -850 -56793 2 VDD
port 41 nsew
rlabel nwell s -11762 -57208 -11240 -57193 2 VDD
port 41 nsew
rlabel nwell s -12735 -57237 -12017 -57193 2 VDD
port 41 nsew
rlabel nwell s -12735 -57193 -11240 -57014 2 VDD
port 41 nsew
rlabel nwell s -12735 -57014 -11153 -57007 2 VDD
port 41 nsew
rlabel nwell s -12735 -57007 -10435 -56827 2 VDD
port 41 nsew
rlabel nwell s -3211 -56793 -2370 -56787 2 VDD
port 41 nsew
rlabel nwell s -12761 -56827 -10435 -56633 2 VDD
port 41 nsew
rlabel nwell s -12761 -56633 -10467 -56085 2 VDD
port 41 nsew
rlabel nwell s -11532 -56085 -10467 -56078 2 VDD
port 41 nsew
rlabel nwell s -12761 -56085 -12152 -56078 2 VDD
port 41 nsew
rlabel nwell s 22456 -56074 23297 -56068 8 VDD
port 41 nsew
rlabel nwell s 36751 -55812 39051 -55632 8 VDD
port 41 nsew
rlabel nwell s 36751 -55632 38333 -55625 8 VDD
port 41 nsew
rlabel nwell s 46587 -55485 47109 -55470 8 VDD
port 41 nsew
rlabel nwell s 55785 -55451 56307 -55436 8 VDD
port 41 nsew
rlabel nwell s 54812 -55451 55530 -55407 8 VDD
port 41 nsew
rlabel nwell s 45614 -55485 46332 -55441 8 VDD
port 41 nsew
rlabel nwell s 36751 -55625 38246 -55446 8 VDD
port 41 nsew
rlabel nwell s 28285 -55995 30611 -55801 8 VDD
port 41 nsew
rlabel nwell s 28311 -55801 30611 -55621 8 VDD
port 41 nsew
rlabel nwell s 28311 -55621 29893 -55614 8 VDD
port 41 nsew
rlabel nwell s 20936 -56068 25998 -55615 8 VDD
port 41 nsew
rlabel nwell s 4388 -55932 4910 -55818 8 VDD
port 41 nsew
rlabel nwell s 4388 -55818 8835 -55738 8 VDD
port 41 nsew
rlabel nwell s 4301 -55738 8835 -55731 8 VDD
port 41 nsew
rlabel nwell s 2783 -55930 3305 -55736 8 VDD
port 41 nsew
rlabel nwell s -285 -55816 1701 -55799 8 VDD
port 41 nsew
rlabel nwell s -912 -55810 -571 -55799 2 VDD
port 41 nsew
rlabel nwell s 2696 -55736 3305 -55731 8 VDD
port 41 nsew
rlabel nwell s 2696 -55731 8835 -55729 8 VDD
port 41 nsew
rlabel nwell s -5925 -55799 1701 -55729 2 VDD
port 41 nsew
rlabel nwell s 23262 -55615 25998 -55614 8 VDD
port 41 nsew
rlabel nwell s 37724 -55446 38246 -55431 8 VDD
port 41 nsew
rlabel nwell s 36751 -55446 37469 -55402 8 VDD
port 41 nsew
rlabel nwell s 28311 -55614 29806 -55435 8 VDD
port 41 nsew
rlabel nwell s 29284 -55435 29806 -55420 8 VDD
port 41 nsew
rlabel nwell s 28311 -55435 29029 -55391 8 VDD
port 41 nsew
rlabel nwell s 64539 -55385 65061 -55370 8 VDD
port 41 nsew
rlabel nwell s 73692 -55368 74214 -55353 8 VDD
port 41 nsew
rlabel nwell s 83056 -55330 83578 -55315 8 VDD
port 41 nsew
rlabel nwell s 82083 -55330 82801 -55286 8 VDD
port 41 nsew
rlabel nwell s 72719 -55368 73437 -55324 8 VDD
port 41 nsew
rlabel nwell s 63566 -55385 64284 -55341 8 VDD
port 41 nsew
rlabel nwell s -5925 -55729 8835 -55343 8 VDD
port 41 nsew
rlabel nwell s -11314 -56078 -10467 -55673 2 VDD
port 41 nsew
rlabel nwell s -12761 -56078 -12239 -55884 2 VDD
port 41 nsew
rlabel nwell s -16751 -56232 -16229 -56217 2 VDD
port 41 nsew
rlabel nwell s -17724 -56261 -17006 -56217 2 VDD
port 41 nsew
rlabel nwell s -17724 -56217 -16229 -56038 2 VDD
port 41 nsew
rlabel nwell s -21328 -56279 -20806 -56085 2 VDD
port 41 nsew
rlabel nwell s -17724 -56038 -16142 -56031 2 VDD
port 41 nsew
rlabel nwell s -17724 -56031 -15424 -55851 2 VDD
port 41 nsew
rlabel nwell s -17750 -55851 -15424 -55657 2 VDD
port 41 nsew
rlabel nwell s -17750 -55657 -15456 -55109 2 VDD
port 41 nsew
rlabel nwell s -19555 -56084 -18099 -55626 2 VDD
port 41 nsew
rlabel nwell s -21328 -56085 -20719 -56078 2 VDD
port 41 nsew
rlabel nwell s -21328 -56078 -20001 -55704 2 VDD
port 41 nsew
rlabel nwell s -19555 -55626 -18130 -55625 2 VDD
port 41 nsew
rlabel nwell s -16521 -55109 -15456 -55102 2 VDD
port 41 nsew
rlabel nwell s -17750 -55109 -17141 -55102 2 VDD
port 41 nsew
rlabel nwell s -5655 -55025 -5035 -54572 2 VDD
port 41 nsew
rlabel nwell s -13799 -54809 -11063 -54808 2 VDD
port 41 nsew
rlabel nwell s -13799 -54808 -7841 -54355 2 VDD
port 41 nsew
rlabel nwell s -16303 -55102 -15456 -54697 2 VDD
port 41 nsew
rlabel nwell s -17750 -55102 -17228 -54908 2 VDD
port 41 nsew
rlabel nwell s -8786 -54355 -8445 -54344 2 VDD
port 41 nsew
rlabel nwell s -19386 -54370 -18864 -54176 2 VDD
port 41 nsew
rlabel nwell s -19386 -54176 -18777 -54169 2 VDD
port 41 nsew
rlabel nwell s -19386 -54169 -18059 -53795 2 VDD
port 41 nsew
rlabel nwell s 6908 -53567 8825 -53494 8 VDD
port 41 nsew
rlabel nwell s 3908 -53567 5825 -53494 8 VDD
port 41 nsew
rlabel nwell s 1408 -53567 3325 -53494 8 VDD
port 41 nsew
rlabel nwell s -1092 -53567 825 -53494 2 VDD
port 41 nsew
rlabel nwell s -3592 -53567 -1675 -53494 2 VDD
port 41 nsew
rlabel nwell s -6092 -53567 -4175 -53494 2 VDD
port 41 nsew
rlabel nwell s 6907 -53494 8825 -53092 8 VDD
port 41 nsew
rlabel nwell s 3907 -53494 5825 -53092 8 VDD
port 41 nsew
rlabel nwell s 1407 -53494 3325 -53092 8 VDD
port 41 nsew
rlabel nwell s -1093 -53494 825 -53092 2 VDD
port 41 nsew
rlabel nwell s -3593 -53494 -1675 -53092 2 VDD
port 41 nsew
rlabel nwell s -6093 -53494 -4175 -53092 2 VDD
port 41 nsew
rlabel nwell s -7522 -53771 -6675 -52894 2 VDD
port 41 nsew
rlabel nwell s -21385 -54148 -19929 -53690 2 VDD
port 41 nsew
rlabel nwell s -21385 -53690 -19960 -53689 2 VDD
port 41 nsew
rlabel nwell s -11085 -53367 -10244 -53361 2 VDD
port 41 nsew
rlabel nwell s -13786 -53361 -8724 -52908 2 VDD
port 41 nsew
rlabel nwell s -13786 -52908 -11050 -52907 2 VDD
port 41 nsew
rlabel nwell s -27894 -59716 -27125 -52116 2 VDD
port 41 nsew
rlabel nwell s -22272 -44215 -20847 -44214 2 VDD
port 41 nsew
rlabel nwell s 14431 -43961 17167 -43960 8 VDD
port 41 nsew
rlabel nwell s 12105 -43960 17167 -43507 8 VDD
port 41 nsew
rlabel nwell s 6204 -44145 8122 -43743 8 VDD
port 41 nsew
rlabel nwell s 3204 -44145 5122 -43743 8 VDD
port 41 nsew
rlabel nwell s 704 -44145 2622 -43743 8 VDD
port 41 nsew
rlabel nwell s -1796 -44145 122 -43743 2 VDD
port 41 nsew
rlabel nwell s -4296 -44145 -2378 -43743 2 VDD
port 41 nsew
rlabel nwell s -6796 -44145 -4878 -43743 2 VDD
port 41 nsew
rlabel nwell s -22303 -44214 -20847 -43756 2 VDD
port 41 nsew
rlabel nwell s 6205 -43743 8122 -43670 8 VDD
port 41 nsew
rlabel nwell s 3205 -43743 5122 -43670 8 VDD
port 41 nsew
rlabel nwell s 705 -43743 2622 -43670 8 VDD
port 41 nsew
rlabel nwell s -1795 -43743 122 -43670 2 VDD
port 41 nsew
rlabel nwell s -4295 -43743 -2378 -43670 2 VDD
port 41 nsew
rlabel nwell s -6795 -43743 -4878 -43670 2 VDD
port 41 nsew
rlabel nwell s 13625 -43507 14466 -43501 8 VDD
port 41 nsew
rlabel nwell s -17454 -43121 -16932 -43106 2 VDD
port 41 nsew
rlabel nwell s -18427 -43150 -17709 -43106 2 VDD
port 41 nsew
rlabel nwell s -18427 -43106 -16932 -42927 2 VDD
port 41 nsew
rlabel nwell s -18427 -42927 -16845 -42920 2 VDD
port 41 nsew
rlabel nwell s -18427 -42920 -16127 -42740 2 VDD
port 41 nsew
rlabel nwell s -18453 -42740 -16127 -42546 2 VDD
port 41 nsew
rlabel nwell s 11826 -42524 12167 -42513 8 VDD
port 41 nsew
rlabel nwell s 86461 -42223 87308 -41818 8 VDD
port 41 nsew
rlabel nwell s 85014 -42012 85536 -41818 8 VDD
port 41 nsew
rlabel nwell s 86243 -41818 87308 -41811 8 VDD
port 41 nsew
rlabel nwell s 85014 -41818 85623 -41811 8 VDD
port 41 nsew
rlabel nwell s 85014 -41811 87308 -41263 8 VDD
port 41 nsew
rlabel nwell s 85014 -41263 87340 -41069 8 VDD
port 41 nsew
rlabel nwell s 82793 -42192 83640 -41787 8 VDD
port 41 nsew
rlabel nwell s 81346 -41981 81868 -41787 8 VDD
port 41 nsew
rlabel nwell s 82575 -41787 83640 -41780 8 VDD
port 41 nsew
rlabel nwell s 81346 -41787 81955 -41780 8 VDD
port 41 nsew
rlabel nwell s 81346 -41780 83640 -41232 8 VDD
port 41 nsew
rlabel nwell s 77097 -42261 77944 -41856 8 VDD
port 41 nsew
rlabel nwell s 75650 -42050 76172 -41856 8 VDD
port 41 nsew
rlabel nwell s 76879 -41856 77944 -41849 8 VDD
port 41 nsew
rlabel nwell s 75650 -41856 76259 -41849 8 VDD
port 41 nsew
rlabel nwell s 75650 -41849 77944 -41301 8 VDD
port 41 nsew
rlabel nwell s 85040 -41069 87340 -40889 8 VDD
port 41 nsew
rlabel nwell s 85040 -40889 86622 -40882 8 VDD
port 41 nsew
rlabel nwell s 85040 -40882 86535 -40703 8 VDD
port 41 nsew
rlabel nwell s 81346 -41232 83672 -41038 8 VDD
port 41 nsew
rlabel nwell s 75650 -41301 77976 -41107 8 VDD
port 41 nsew
rlabel nwell s 73429 -42230 74276 -41825 8 VDD
port 41 nsew
rlabel nwell s 71982 -42019 72504 -41825 8 VDD
port 41 nsew
rlabel nwell s 73211 -41825 74276 -41818 8 VDD
port 41 nsew
rlabel nwell s 71982 -41825 72591 -41818 8 VDD
port 41 nsew
rlabel nwell s 71982 -41818 74276 -41270 8 VDD
port 41 nsew
rlabel nwell s 67944 -42278 68791 -41873 8 VDD
port 41 nsew
rlabel nwell s 66497 -42067 67019 -41873 8 VDD
port 41 nsew
rlabel nwell s 67726 -41873 68791 -41866 8 VDD
port 41 nsew
rlabel nwell s 66497 -41873 67106 -41866 8 VDD
port 41 nsew
rlabel nwell s 66497 -41866 68791 -41318 8 VDD
port 41 nsew
rlabel nwell s 81372 -41038 83672 -40858 8 VDD
port 41 nsew
rlabel nwell s 75676 -41107 77976 -40927 8 VDD
port 41 nsew
rlabel nwell s 75676 -40927 77258 -40920 8 VDD
port 41 nsew
rlabel nwell s 81372 -40858 82954 -40851 8 VDD
port 41 nsew
rlabel nwell s 86013 -40703 86535 -40688 8 VDD
port 41 nsew
rlabel nwell s 85040 -40703 85758 -40659 8 VDD
port 41 nsew
rlabel nwell s 81372 -40851 82867 -40672 8 VDD
port 41 nsew
rlabel nwell s 75676 -40920 77171 -40741 8 VDD
port 41 nsew
rlabel nwell s 71982 -41270 74308 -41076 8 VDD
port 41 nsew
rlabel nwell s 66497 -41318 68823 -41124 8 VDD
port 41 nsew
rlabel nwell s 64276 -42247 65123 -41842 8 VDD
port 41 nsew
rlabel nwell s 62829 -42036 63351 -41842 8 VDD
port 41 nsew
rlabel nwell s 64058 -41842 65123 -41835 8 VDD
port 41 nsew
rlabel nwell s 62829 -41842 63438 -41835 8 VDD
port 41 nsew
rlabel nwell s 62829 -41835 65123 -41287 8 VDD
port 41 nsew
rlabel nwell s 59190 -42344 60037 -41939 8 VDD
port 41 nsew
rlabel nwell s 57743 -42133 58265 -41939 8 VDD
port 41 nsew
rlabel nwell s 58972 -41939 60037 -41932 8 VDD
port 41 nsew
rlabel nwell s 57743 -41939 58352 -41932 8 VDD
port 41 nsew
rlabel nwell s 57743 -41932 60037 -41384 8 VDD
port 41 nsew
rlabel nwell s 72008 -41076 74308 -40896 8 VDD
port 41 nsew
rlabel nwell s 66523 -41124 68823 -40944 8 VDD
port 41 nsew
rlabel nwell s 66523 -40944 68105 -40937 8 VDD
port 41 nsew
rlabel nwell s 72008 -40896 73590 -40889 8 VDD
port 41 nsew
rlabel nwell s 76649 -40741 77171 -40726 8 VDD
port 41 nsew
rlabel nwell s 75676 -40741 76394 -40697 8 VDD
port 41 nsew
rlabel nwell s 72008 -40889 73503 -40710 8 VDD
port 41 nsew
rlabel nwell s 66523 -40937 68018 -40758 8 VDD
port 41 nsew
rlabel nwell s 62829 -41287 65155 -41093 8 VDD
port 41 nsew
rlabel nwell s 57743 -41384 60069 -41190 8 VDD
port 41 nsew
rlabel nwell s 55522 -42313 56369 -41908 8 VDD
port 41 nsew
rlabel nwell s 54075 -42102 54597 -41908 8 VDD
port 41 nsew
rlabel nwell s 55304 -41908 56369 -41901 8 VDD
port 41 nsew
rlabel nwell s 54075 -41908 54684 -41901 8 VDD
port 41 nsew
rlabel nwell s 54075 -41901 56369 -41353 8 VDD
port 41 nsew
rlabel nwell s 49992 -42378 50839 -41973 8 VDD
port 41 nsew
rlabel nwell s 48545 -42167 49067 -41973 8 VDD
port 41 nsew
rlabel nwell s 49774 -41973 50839 -41966 8 VDD
port 41 nsew
rlabel nwell s 48545 -41973 49154 -41966 8 VDD
port 41 nsew
rlabel nwell s 48545 -41966 50839 -41418 8 VDD
port 41 nsew
rlabel nwell s 62855 -41093 65155 -40913 8 VDD
port 41 nsew
rlabel nwell s 57769 -41190 60069 -41010 8 VDD
port 41 nsew
rlabel nwell s 57769 -41010 59351 -41003 8 VDD
port 41 nsew
rlabel nwell s 62855 -40913 64437 -40906 8 VDD
port 41 nsew
rlabel nwell s 67496 -40758 68018 -40743 8 VDD
port 41 nsew
rlabel nwell s 66523 -40758 67241 -40714 8 VDD
port 41 nsew
rlabel nwell s 62855 -40906 64350 -40727 8 VDD
port 41 nsew
rlabel nwell s 57769 -41003 59264 -40824 8 VDD
port 41 nsew
rlabel nwell s 54075 -41353 56401 -41159 8 VDD
port 41 nsew
rlabel nwell s 48545 -41418 50871 -41224 8 VDD
port 41 nsew
rlabel nwell s 46324 -42347 47171 -41942 8 VDD
port 41 nsew
rlabel nwell s 44877 -42136 45399 -41942 8 VDD
port 41 nsew
rlabel nwell s 46106 -41942 47171 -41935 8 VDD
port 41 nsew
rlabel nwell s 44877 -41942 45486 -41935 8 VDD
port 41 nsew
rlabel nwell s 44877 -41935 47171 -41387 8 VDD
port 41 nsew
rlabel nwell s 54101 -41159 56401 -40979 8 VDD
port 41 nsew
rlabel nwell s 48571 -41224 50871 -41044 8 VDD
port 41 nsew
rlabel nwell s 48571 -41044 50153 -41037 8 VDD
port 41 nsew
rlabel nwell s 54101 -40979 55683 -40972 8 VDD
port 41 nsew
rlabel nwell s 58742 -40824 59264 -40809 8 VDD
port 41 nsew
rlabel nwell s 57769 -40824 58487 -40780 8 VDD
port 41 nsew
rlabel nwell s 54101 -40972 55596 -40793 8 VDD
port 41 nsew
rlabel nwell s 48571 -41037 50066 -40858 8 VDD
port 41 nsew
rlabel nwell s 44877 -41387 47203 -41193 8 VDD
port 41 nsew
rlabel nwell s 41129 -42339 41976 -41934 8 VDD
port 41 nsew
rlabel nwell s 39682 -42128 40204 -41934 8 VDD
port 41 nsew
rlabel nwell s 40911 -41934 41976 -41927 8 VDD
port 41 nsew
rlabel nwell s 39682 -41934 40291 -41927 8 VDD
port 41 nsew
rlabel nwell s 39682 -41927 41976 -41379 8 VDD
port 41 nsew
rlabel nwell s 44903 -41193 47203 -41013 8 VDD
port 41 nsew
rlabel nwell s 44903 -41013 46485 -41006 8 VDD
port 41 nsew
rlabel nwell s 49544 -40858 50066 -40843 8 VDD
port 41 nsew
rlabel nwell s 48571 -40858 49289 -40814 8 VDD
port 41 nsew
rlabel nwell s 44903 -41006 46398 -40827 8 VDD
port 41 nsew
rlabel nwell s 39682 -41379 42008 -41185 8 VDD
port 41 nsew
rlabel nwell s 37461 -42308 38308 -41903 8 VDD
port 41 nsew
rlabel nwell s 36014 -42097 36536 -41903 8 VDD
port 41 nsew
rlabel nwell s 37243 -41903 38308 -41896 8 VDD
port 41 nsew
rlabel nwell s 36014 -41903 36623 -41896 8 VDD
port 41 nsew
rlabel nwell s 36014 -41896 38308 -41348 8 VDD
port 41 nsew
rlabel nwell s 32689 -42328 33536 -41923 8 VDD
port 41 nsew
rlabel nwell s 31242 -42117 31764 -41923 8 VDD
port 41 nsew
rlabel nwell s 32471 -41923 33536 -41916 8 VDD
port 41 nsew
rlabel nwell s 31242 -41923 31851 -41916 8 VDD
port 41 nsew
rlabel nwell s 31242 -41916 33536 -41368 8 VDD
port 41 nsew
rlabel nwell s 39708 -41185 42008 -41005 8 VDD
port 41 nsew
rlabel nwell s 39708 -41005 41290 -40998 8 VDD
port 41 nsew
rlabel nwell s 45876 -40827 46398 -40812 8 VDD
port 41 nsew
rlabel nwell s 55074 -40793 55596 -40778 8 VDD
port 41 nsew
rlabel nwell s 54101 -40793 54819 -40749 8 VDD
port 41 nsew
rlabel nwell s 44903 -40827 45621 -40783 8 VDD
port 41 nsew
rlabel nwell s 39708 -40998 41203 -40819 8 VDD
port 41 nsew
rlabel nwell s 36014 -41348 38340 -41154 8 VDD
port 41 nsew
rlabel nwell s 31242 -41368 33568 -41174 8 VDD
port 41 nsew
rlabel nwell s 29021 -42297 29868 -41892 8 VDD
port 41 nsew
rlabel nwell s 27574 -42086 28096 -41892 8 VDD
port 41 nsew
rlabel nwell s 11222 -42513 17180 -42060 8 VDD
port 41 nsew
rlabel nwell s 14444 -42060 17180 -42059 8 VDD
port 41 nsew
rlabel nwell s -18453 -42546 -16159 -41998 2 VDD
port 41 nsew
rlabel nwell s -17224 -41998 -16159 -41991 2 VDD
port 41 nsew
rlabel nwell s -18453 -41998 -17844 -41991 2 VDD
port 41 nsew
rlabel nwell s 28803 -41892 29868 -41885 8 VDD
port 41 nsew
rlabel nwell s 27574 -41892 28183 -41885 8 VDD
port 41 nsew
rlabel nwell s 27574 -41885 29868 -41337 8 VDD
port 41 nsew
rlabel nwell s 19886 -41670 21311 -41669 8 VDD
port 41 nsew
rlabel nwell s 36040 -41154 38340 -40974 8 VDD
port 41 nsew
rlabel nwell s 31268 -41174 33568 -40994 8 VDD
port 41 nsew
rlabel nwell s 31268 -40994 32850 -40987 8 VDD
port 41 nsew
rlabel nwell s 36040 -40974 37622 -40967 8 VDD
port 41 nsew
rlabel nwell s 40681 -40819 41203 -40804 8 VDD
port 41 nsew
rlabel nwell s 39708 -40819 40426 -40775 8 VDD
port 41 nsew
rlabel nwell s 36040 -40967 37535 -40788 8 VDD
port 41 nsew
rlabel nwell s 31268 -40987 32763 -40808 8 VDD
port 41 nsew
rlabel nwell s 27574 -41337 29900 -41143 8 VDD
port 41 nsew
rlabel nwell s 27600 -41143 29900 -40963 8 VDD
port 41 nsew
rlabel nwell s 27600 -40963 29182 -40956 8 VDD
port 41 nsew
rlabel nwell s 32241 -40808 32763 -40793 8 VDD
port 41 nsew
rlabel nwell s 37013 -40788 37535 -40773 8 VDD
port 41 nsew
rlabel nwell s 36040 -40788 36758 -40744 8 VDD
port 41 nsew
rlabel nwell s 31268 -40808 31986 -40764 8 VDD
port 41 nsew
rlabel nwell s 27600 -40956 29095 -40777 8 VDD
port 41 nsew
rlabel nwell s 28573 -40777 29095 -40762 8 VDD
port 41 nsew
rlabel nwell s 27600 -40777 28318 -40733 8 VDD
port 41 nsew
rlabel nwell s 63828 -40727 64350 -40712 8 VDD
port 41 nsew
rlabel nwell s 72981 -40710 73503 -40695 8 VDD
port 41 nsew
rlabel nwell s 82345 -40672 82867 -40657 8 VDD
port 41 nsew
rlabel nwell s 81372 -40672 82090 -40628 8 VDD
port 41 nsew
rlabel nwell s 72008 -40710 72726 -40666 8 VDD
port 41 nsew
rlabel nwell s 62855 -40727 63573 -40683 8 VDD
port 41 nsew
rlabel nwell s 22625 -41665 25351 -40633 8 VDD
port 41 nsew
rlabel nwell s 21745 -41657 22365 -41204 8 VDD
port 41 nsew
rlabel nwell s 19886 -41669 21342 -41211 8 VDD
port 41 nsew
rlabel nwell s 18970 -41658 19605 -40977 8 VDD
port 41 nsew
rlabel nwell s 18024 -41658 18659 -40977 8 VDD
port 41 nsew
rlabel nwell s -6628 -41894 8132 -41508 8 VDD
port 41 nsew
rlabel nwell s -14502 -41625 -11766 -41624 2 VDD
port 41 nsew
rlabel nwell s 1993 -41508 8132 -41506 8 VDD
port 41 nsew
rlabel nwell s 3598 -41506 8132 -41499 8 VDD
port 41 nsew
rlabel nwell s 1993 -41506 2602 -41501 8 VDD
port 41 nsew
rlabel nwell s 3685 -41499 8132 -41419 8 VDD
port 41 nsew
rlabel nwell s 3685 -41419 4207 -41305 8 VDD
port 41 nsew
rlabel nwell s 2080 -41501 2602 -41307 8 VDD
port 41 nsew
rlabel nwell s -6628 -41508 998 -41438 2 VDD
port 41 nsew
rlabel nwell s -988 -41438 998 -41421 8 VDD
port 41 nsew
rlabel nwell s -1615 -41438 -1274 -41427 2 VDD
port 41 nsew
rlabel nwell s -14502 -41624 -8544 -41171 2 VDD
port 41 nsew
rlabel nwell s -17006 -41991 -16159 -41586 2 VDD
port 41 nsew
rlabel nwell s -18453 -41991 -17931 -41797 2 VDD
port 41 nsew
rlabel nwell s -9489 -41171 -9148 -41160 2 VDD
port 41 nsew
rlabel nwell s -19855 -41392 -19220 -40711 2 VDD
port 41 nsew
rlabel nwell s -20760 -41391 -20125 -40710 2 VDD
port 41 nsew
rlabel nwell s -21966 -41662 -21021 -40717 2 VDD
port 41 nsew
rlabel nwell s -3914 -40450 -3073 -40444 2 VDD
port 41 nsew
rlabel nwell s 21795 -40227 22317 -39673 8 VDD
port 41 nsew
rlabel nwell s -6615 -40444 -1553 -39991 2 VDD
port 41 nsew
rlabel nwell s -6615 -39991 -3879 -39990 2 VDD
port 41 nsew
rlabel nwell s -8198 -40594 -7351 -39717 2 VDD
port 41 nsew
rlabel nwell s -11788 -40183 -10947 -40177 2 VDD
port 41 nsew
rlabel nwell s -14489 -40177 -9427 -39724 2 VDD
port 41 nsew
rlabel nwell s -14489 -39724 -11753 -39723 2 VDD
port 41 nsew
rlabel nwell s 22572 -39405 25308 -39404 8 VDD
port 41 nsew
rlabel nwell s 21784 -39673 22317 -39404 8 VDD
port 41 nsew
rlabel nwell s 18028 -39404 25308 -38951 8 VDD
port 41 nsew
rlabel nwell s -6615 -39136 -3879 -39135 2 VDD
port 41 nsew
rlabel nwell s 19954 -38951 20295 -38940 8 VDD
port 41 nsew
rlabel nwell s 84793 -38497 86270 -37624 8 VDD
port 41 nsew
rlabel nwell s 82801 -38739 83648 -38334 8 VDD
port 41 nsew
rlabel nwell s 81354 -38528 81876 -38334 8 VDD
port 41 nsew
rlabel nwell s 82583 -38334 83648 -38327 8 VDD
port 41 nsew
rlabel nwell s 81354 -38334 81963 -38327 8 VDD
port 41 nsew
rlabel nwell s 81354 -38327 83648 -37779 8 VDD
port 41 nsew
rlabel nwell s 81354 -37779 83680 -37585 8 VDD
port 41 nsew
rlabel nwell s 75429 -38535 76906 -37662 8 VDD
port 41 nsew
rlabel nwell s 73437 -38777 74284 -38372 8 VDD
port 41 nsew
rlabel nwell s 71990 -38566 72512 -38372 8 VDD
port 41 nsew
rlabel nwell s 73219 -38372 74284 -38365 8 VDD
port 41 nsew
rlabel nwell s 71990 -38372 72599 -38365 8 VDD
port 41 nsew
rlabel nwell s 71990 -38365 74284 -37817 8 VDD
port 41 nsew
rlabel nwell s 71990 -37817 74316 -37623 8 VDD
port 41 nsew
rlabel nwell s 66276 -38552 67753 -37679 8 VDD
port 41 nsew
rlabel nwell s 64284 -38794 65131 -38389 8 VDD
port 41 nsew
rlabel nwell s 62837 -38583 63359 -38389 8 VDD
port 41 nsew
rlabel nwell s 64066 -38389 65131 -38382 8 VDD
port 41 nsew
rlabel nwell s 62837 -38389 63446 -38382 8 VDD
port 41 nsew
rlabel nwell s 62837 -38382 65131 -37834 8 VDD
port 41 nsew
rlabel nwell s 62837 -37834 65163 -37640 8 VDD
port 41 nsew
rlabel nwell s 57522 -38618 58999 -37745 8 VDD
port 41 nsew
rlabel nwell s 55530 -38860 56377 -38455 8 VDD
port 41 nsew
rlabel nwell s 54083 -38649 54605 -38455 8 VDD
port 41 nsew
rlabel nwell s 55312 -38455 56377 -38448 8 VDD
port 41 nsew
rlabel nwell s 54083 -38455 54692 -38448 8 VDD
port 41 nsew
rlabel nwell s 54083 -38448 56377 -37900 8 VDD
port 41 nsew
rlabel nwell s 54083 -37900 56409 -37706 8 VDD
port 41 nsew
rlabel nwell s 48324 -38652 49801 -37779 8 VDD
port 41 nsew
rlabel nwell s 46332 -38894 47179 -38489 8 VDD
port 41 nsew
rlabel nwell s 44885 -38683 45407 -38489 8 VDD
port 41 nsew
rlabel nwell s 46114 -38489 47179 -38482 8 VDD
port 41 nsew
rlabel nwell s 44885 -38489 45494 -38482 8 VDD
port 41 nsew
rlabel nwell s 44885 -38482 47179 -37934 8 VDD
port 41 nsew
rlabel nwell s 44885 -37934 47211 -37740 8 VDD
port 41 nsew
rlabel nwell s 39461 -38613 40938 -37740 8 VDD
port 41 nsew
rlabel nwell s 37469 -38855 38316 -38450 8 VDD
port 41 nsew
rlabel nwell s 36022 -38644 36544 -38450 8 VDD
port 41 nsew
rlabel nwell s 37251 -38450 38316 -38443 8 VDD
port 41 nsew
rlabel nwell s 36022 -38450 36631 -38443 8 VDD
port 41 nsew
rlabel nwell s 36022 -38443 38316 -37895 8 VDD
port 41 nsew
rlabel nwell s 81380 -37585 83680 -37405 8 VDD
port 41 nsew
rlabel nwell s 72016 -37623 74316 -37443 8 VDD
port 41 nsew
rlabel nwell s 62863 -37640 65163 -37460 8 VDD
port 41 nsew
rlabel nwell s 54109 -37706 56409 -37526 8 VDD
port 41 nsew
rlabel nwell s 44911 -37740 47211 -37560 8 VDD
port 41 nsew
rlabel nwell s 44911 -37560 46493 -37553 8 VDD
port 41 nsew
rlabel nwell s 54109 -37526 55691 -37519 8 VDD
port 41 nsew
rlabel nwell s 62863 -37460 64445 -37453 8 VDD
port 41 nsew
rlabel nwell s 72016 -37443 73598 -37436 8 VDD
port 41 nsew
rlabel nwell s 81380 -37405 82962 -37398 8 VDD
port 41 nsew
rlabel nwell s 81380 -37398 82875 -37219 8 VDD
port 41 nsew
rlabel nwell s 72016 -37436 73511 -37257 8 VDD
port 41 nsew
rlabel nwell s 62863 -37453 64358 -37274 8 VDD
port 41 nsew
rlabel nwell s 54109 -37519 55604 -37340 8 VDD
port 41 nsew
rlabel nwell s 44911 -37553 46406 -37374 8 VDD
port 41 nsew
rlabel nwell s 36022 -37895 38348 -37701 8 VDD
port 41 nsew
rlabel nwell s 31021 -38602 32498 -37729 8 VDD
port 41 nsew
rlabel nwell s 29029 -38844 29876 -38439 8 VDD
port 41 nsew
rlabel nwell s 27582 -38633 28104 -38439 8 VDD
port 41 nsew
rlabel nwell s 28811 -38439 29876 -38432 8 VDD
port 41 nsew
rlabel nwell s 27582 -38439 28191 -38432 8 VDD
port 41 nsew
rlabel nwell s 27582 -38432 29876 -37884 8 VDD
port 41 nsew
rlabel nwell s 18029 -38951 18974 -38431 8 VDD
port 41 nsew
rlabel nwell s -6615 -39135 -1553 -38682 2 VDD
port 41 nsew
rlabel nwell s -12465 -39097 -11943 -39082 2 VDD
port 41 nsew
rlabel nwell s -13438 -39126 -12720 -39082 2 VDD
port 41 nsew
rlabel nwell s -13438 -39082 -11943 -38903 2 VDD
port 41 nsew
rlabel nwell s -13438 -38903 -11856 -38896 2 VDD
port 41 nsew
rlabel nwell s -13438 -38896 -11138 -38716 2 VDD
port 41 nsew
rlabel nwell s -3914 -38682 -3073 -38676 2 VDD
port 41 nsew
rlabel nwell s -13464 -38716 -11138 -38522 2 VDD
port 41 nsew
rlabel nwell s -13464 -38522 -11170 -37974 2 VDD
port 41 nsew
rlabel nwell s -12235 -37974 -11170 -37967 2 VDD
port 41 nsew
rlabel nwell s -13464 -37974 -12855 -37967 2 VDD
port 41 nsew
rlabel nwell s 21753 -37963 22594 -37957 8 VDD
port 41 nsew
rlabel nwell s 36048 -37701 38348 -37521 8 VDD
port 41 nsew
rlabel nwell s 36048 -37521 37630 -37514 8 VDD
port 41 nsew
rlabel nwell s 45884 -37374 46406 -37359 8 VDD
port 41 nsew
rlabel nwell s 55082 -37340 55604 -37325 8 VDD
port 41 nsew
rlabel nwell s 54109 -37340 54827 -37296 8 VDD
port 41 nsew
rlabel nwell s 44911 -37374 45629 -37330 8 VDD
port 41 nsew
rlabel nwell s 36048 -37514 37543 -37335 8 VDD
port 41 nsew
rlabel nwell s 27582 -37884 29908 -37690 8 VDD
port 41 nsew
rlabel nwell s 27608 -37690 29908 -37510 8 VDD
port 41 nsew
rlabel nwell s 27608 -37510 29190 -37503 8 VDD
port 41 nsew
rlabel nwell s 20233 -37957 25295 -37504 8 VDD
port 41 nsew
rlabel nwell s 3685 -37821 4207 -37707 8 VDD
port 41 nsew
rlabel nwell s 3685 -37707 8132 -37627 8 VDD
port 41 nsew
rlabel nwell s 3598 -37627 8132 -37620 8 VDD
port 41 nsew
rlabel nwell s 2080 -37819 2602 -37625 8 VDD
port 41 nsew
rlabel nwell s -988 -37705 998 -37688 8 VDD
port 41 nsew
rlabel nwell s -1615 -37699 -1274 -37688 2 VDD
port 41 nsew
rlabel nwell s 1993 -37625 2602 -37620 8 VDD
port 41 nsew
rlabel nwell s 1993 -37620 8132 -37618 8 VDD
port 41 nsew
rlabel nwell s -6628 -37688 998 -37618 2 VDD
port 41 nsew
rlabel nwell s 22559 -37504 25295 -37503 8 VDD
port 41 nsew
rlabel nwell s 37021 -37335 37543 -37320 8 VDD
port 41 nsew
rlabel nwell s 36048 -37335 36766 -37291 8 VDD
port 41 nsew
rlabel nwell s 27608 -37503 29103 -37324 8 VDD
port 41 nsew
rlabel nwell s 28581 -37324 29103 -37309 8 VDD
port 41 nsew
rlabel nwell s 27608 -37324 28326 -37280 8 VDD
port 41 nsew
rlabel nwell s 63836 -37274 64358 -37259 8 VDD
port 41 nsew
rlabel nwell s 72989 -37257 73511 -37242 8 VDD
port 41 nsew
rlabel nwell s 82353 -37219 82875 -37204 8 VDD
port 41 nsew
rlabel nwell s 81380 -37219 82098 -37175 8 VDD
port 41 nsew
rlabel nwell s 72016 -37257 72734 -37213 8 VDD
port 41 nsew
rlabel nwell s 62863 -37274 63581 -37230 8 VDD
port 41 nsew
rlabel nwell s -6628 -37618 8132 -37232 8 VDD
port 41 nsew
rlabel nwell s -12017 -37967 -11170 -37562 2 VDD
port 41 nsew
rlabel nwell s -13464 -37967 -12942 -37773 2 VDD
port 41 nsew
rlabel nwell s -17454 -38121 -16932 -38106 2 VDD
port 41 nsew
rlabel nwell s -18427 -38150 -17709 -38106 2 VDD
port 41 nsew
rlabel nwell s -18427 -38106 -16932 -37927 2 VDD
port 41 nsew
rlabel nwell s -22031 -38168 -21509 -37974 2 VDD
port 41 nsew
rlabel nwell s -18427 -37927 -16845 -37920 2 VDD
port 41 nsew
rlabel nwell s -18427 -37920 -16127 -37740 2 VDD
port 41 nsew
rlabel nwell s -18453 -37740 -16127 -37546 2 VDD
port 41 nsew
rlabel nwell s -18453 -37546 -16159 -36998 2 VDD
port 41 nsew
rlabel nwell s -20258 -37973 -18802 -37515 2 VDD
port 41 nsew
rlabel nwell s -22031 -37974 -21422 -37967 2 VDD
port 41 nsew
rlabel nwell s -22031 -37967 -20704 -37593 2 VDD
port 41 nsew
rlabel nwell s -20258 -37515 -18833 -37514 2 VDD
port 41 nsew
rlabel nwell s -17224 -36998 -16159 -36991 2 VDD
port 41 nsew
rlabel nwell s -18453 -36998 -17844 -36991 2 VDD
port 41 nsew
rlabel nwell s -6358 -36914 -5738 -36461 2 VDD
port 41 nsew
rlabel nwell s -14502 -36698 -11766 -36697 2 VDD
port 41 nsew
rlabel nwell s -14502 -36697 -8544 -36244 2 VDD
port 41 nsew
rlabel nwell s -17006 -36991 -16159 -36586 2 VDD
port 41 nsew
rlabel nwell s -18453 -36991 -17931 -36797 2 VDD
port 41 nsew
rlabel nwell s -9489 -36244 -9148 -36233 2 VDD
port 41 nsew
rlabel nwell s -20089 -36259 -19567 -36065 2 VDD
port 41 nsew
rlabel nwell s -20089 -36065 -19480 -36058 2 VDD
port 41 nsew
rlabel nwell s -20089 -36058 -18762 -35684 2 VDD
port 41 nsew
rlabel nwell s 6205 -35456 8122 -35383 8 VDD
port 41 nsew
rlabel nwell s 3205 -35456 5122 -35383 8 VDD
port 41 nsew
rlabel nwell s 705 -35456 2622 -35383 8 VDD
port 41 nsew
rlabel nwell s -1795 -35456 122 -35383 2 VDD
port 41 nsew
rlabel nwell s -4295 -35456 -2378 -35383 2 VDD
port 41 nsew
rlabel nwell s -6795 -35456 -4878 -35383 2 VDD
port 41 nsew
rlabel nwell s 6204 -35383 8122 -34981 8 VDD
port 41 nsew
rlabel nwell s 3204 -35383 5122 -34981 8 VDD
port 41 nsew
rlabel nwell s 704 -35383 2622 -34981 8 VDD
port 41 nsew
rlabel nwell s -1796 -35383 122 -34981 2 VDD
port 41 nsew
rlabel nwell s -4296 -35383 -2378 -34981 2 VDD
port 41 nsew
rlabel nwell s -6796 -35383 -4878 -34981 2 VDD
port 41 nsew
rlabel nwell s -8225 -35660 -7378 -34783 2 VDD
port 41 nsew
rlabel nwell s -22088 -36037 -20632 -35579 2 VDD
port 41 nsew
rlabel nwell s -22088 -35579 -20663 -35578 2 VDD
port 41 nsew
rlabel nwell s -11788 -35256 -10947 -35250 2 VDD
port 41 nsew
rlabel nwell s -14489 -35250 -9427 -34797 2 VDD
port 41 nsew
rlabel nwell s -14489 -34797 -11753 -34796 2 VDD
port 41 nsew
rlabel nwell s -26074 -41571 -25305 -33971 2 VDD
port 41 nsew
rlabel nwell s -22970 -27624 -21545 -27623 2 VDD
port 41 nsew
rlabel nwell s 13733 -27370 16469 -27369 8 VDD
port 41 nsew
rlabel nwell s 11407 -27369 16469 -26916 8 VDD
port 41 nsew
rlabel nwell s 5506 -27554 7424 -27152 8 VDD
port 41 nsew
rlabel nwell s 2506 -27554 4424 -27152 8 VDD
port 41 nsew
rlabel nwell s 6 -27554 1924 -27152 8 VDD
port 41 nsew
rlabel nwell s -2494 -27554 -576 -27152 2 VDD
port 41 nsew
rlabel nwell s -4994 -27554 -3076 -27152 2 VDD
port 41 nsew
rlabel nwell s -7494 -27554 -5576 -27152 2 VDD
port 41 nsew
rlabel nwell s -23001 -27623 -21545 -27165 2 VDD
port 41 nsew
rlabel nwell s 5507 -27152 7424 -27079 8 VDD
port 41 nsew
rlabel nwell s 2507 -27152 4424 -27079 8 VDD
port 41 nsew
rlabel nwell s 7 -27152 1924 -27079 8 VDD
port 41 nsew
rlabel nwell s -2493 -27152 -576 -27079 2 VDD
port 41 nsew
rlabel nwell s -4993 -27152 -3076 -27079 2 VDD
port 41 nsew
rlabel nwell s -7493 -27152 -5576 -27079 2 VDD
port 41 nsew
rlabel nwell s 12927 -26916 13768 -26910 8 VDD
port 41 nsew
rlabel nwell s -18152 -26530 -17630 -26515 2 VDD
port 41 nsew
rlabel nwell s -19125 -26559 -18407 -26515 2 VDD
port 41 nsew
rlabel nwell s -19125 -26515 -17630 -26336 2 VDD
port 41 nsew
rlabel nwell s -19125 -26336 -17543 -26329 2 VDD
port 41 nsew
rlabel nwell s -19125 -26329 -16825 -26149 2 VDD
port 41 nsew
rlabel nwell s -19151 -26149 -16825 -25955 2 VDD
port 41 nsew
rlabel nwell s 11128 -25933 11469 -25922 8 VDD
port 41 nsew
rlabel nwell s 85763 -25632 86610 -25227 8 VDD
port 41 nsew
rlabel nwell s 84316 -25421 84838 -25227 8 VDD
port 41 nsew
rlabel nwell s 85545 -25227 86610 -25220 8 VDD
port 41 nsew
rlabel nwell s 84316 -25227 84925 -25220 8 VDD
port 41 nsew
rlabel nwell s 84316 -25220 86610 -24672 8 VDD
port 41 nsew
rlabel nwell s 84316 -24672 86642 -24478 8 VDD
port 41 nsew
rlabel nwell s 82095 -25601 82942 -25196 8 VDD
port 41 nsew
rlabel nwell s 80648 -25390 81170 -25196 8 VDD
port 41 nsew
rlabel nwell s 81877 -25196 82942 -25189 8 VDD
port 41 nsew
rlabel nwell s 80648 -25196 81257 -25189 8 VDD
port 41 nsew
rlabel nwell s 80648 -25189 82942 -24641 8 VDD
port 41 nsew
rlabel nwell s 76399 -25670 77246 -25265 8 VDD
port 41 nsew
rlabel nwell s 74952 -25459 75474 -25265 8 VDD
port 41 nsew
rlabel nwell s 76181 -25265 77246 -25258 8 VDD
port 41 nsew
rlabel nwell s 74952 -25265 75561 -25258 8 VDD
port 41 nsew
rlabel nwell s 74952 -25258 77246 -24710 8 VDD
port 41 nsew
rlabel nwell s 84342 -24478 86642 -24298 8 VDD
port 41 nsew
rlabel nwell s 84342 -24298 85924 -24291 8 VDD
port 41 nsew
rlabel nwell s 84342 -24291 85837 -24112 8 VDD
port 41 nsew
rlabel nwell s 80648 -24641 82974 -24447 8 VDD
port 41 nsew
rlabel nwell s 74952 -24710 77278 -24516 8 VDD
port 41 nsew
rlabel nwell s 72731 -25639 73578 -25234 8 VDD
port 41 nsew
rlabel nwell s 71284 -25428 71806 -25234 8 VDD
port 41 nsew
rlabel nwell s 72513 -25234 73578 -25227 8 VDD
port 41 nsew
rlabel nwell s 71284 -25234 71893 -25227 8 VDD
port 41 nsew
rlabel nwell s 71284 -25227 73578 -24679 8 VDD
port 41 nsew
rlabel nwell s 67246 -25687 68093 -25282 8 VDD
port 41 nsew
rlabel nwell s 65799 -25476 66321 -25282 8 VDD
port 41 nsew
rlabel nwell s 67028 -25282 68093 -25275 8 VDD
port 41 nsew
rlabel nwell s 65799 -25282 66408 -25275 8 VDD
port 41 nsew
rlabel nwell s 65799 -25275 68093 -24727 8 VDD
port 41 nsew
rlabel nwell s 80674 -24447 82974 -24267 8 VDD
port 41 nsew
rlabel nwell s 74978 -24516 77278 -24336 8 VDD
port 41 nsew
rlabel nwell s 74978 -24336 76560 -24329 8 VDD
port 41 nsew
rlabel nwell s 80674 -24267 82256 -24260 8 VDD
port 41 nsew
rlabel nwell s 85315 -24112 85837 -24097 8 VDD
port 41 nsew
rlabel nwell s 84342 -24112 85060 -24068 8 VDD
port 41 nsew
rlabel nwell s 80674 -24260 82169 -24081 8 VDD
port 41 nsew
rlabel nwell s 74978 -24329 76473 -24150 8 VDD
port 41 nsew
rlabel nwell s 71284 -24679 73610 -24485 8 VDD
port 41 nsew
rlabel nwell s 65799 -24727 68125 -24533 8 VDD
port 41 nsew
rlabel nwell s 63578 -25656 64425 -25251 8 VDD
port 41 nsew
rlabel nwell s 62131 -25445 62653 -25251 8 VDD
port 41 nsew
rlabel nwell s 63360 -25251 64425 -25244 8 VDD
port 41 nsew
rlabel nwell s 62131 -25251 62740 -25244 8 VDD
port 41 nsew
rlabel nwell s 62131 -25244 64425 -24696 8 VDD
port 41 nsew
rlabel nwell s 58492 -25753 59339 -25348 8 VDD
port 41 nsew
rlabel nwell s 57045 -25542 57567 -25348 8 VDD
port 41 nsew
rlabel nwell s 58274 -25348 59339 -25341 8 VDD
port 41 nsew
rlabel nwell s 57045 -25348 57654 -25341 8 VDD
port 41 nsew
rlabel nwell s 57045 -25341 59339 -24793 8 VDD
port 41 nsew
rlabel nwell s 71310 -24485 73610 -24305 8 VDD
port 41 nsew
rlabel nwell s 65825 -24533 68125 -24353 8 VDD
port 41 nsew
rlabel nwell s 65825 -24353 67407 -24346 8 VDD
port 41 nsew
rlabel nwell s 71310 -24305 72892 -24298 8 VDD
port 41 nsew
rlabel nwell s 75951 -24150 76473 -24135 8 VDD
port 41 nsew
rlabel nwell s 74978 -24150 75696 -24106 8 VDD
port 41 nsew
rlabel nwell s 71310 -24298 72805 -24119 8 VDD
port 41 nsew
rlabel nwell s 65825 -24346 67320 -24167 8 VDD
port 41 nsew
rlabel nwell s 62131 -24696 64457 -24502 8 VDD
port 41 nsew
rlabel nwell s 57045 -24793 59371 -24599 8 VDD
port 41 nsew
rlabel nwell s 54824 -25722 55671 -25317 8 VDD
port 41 nsew
rlabel nwell s 53377 -25511 53899 -25317 8 VDD
port 41 nsew
rlabel nwell s 54606 -25317 55671 -25310 8 VDD
port 41 nsew
rlabel nwell s 53377 -25317 53986 -25310 8 VDD
port 41 nsew
rlabel nwell s 53377 -25310 55671 -24762 8 VDD
port 41 nsew
rlabel nwell s 49294 -25787 50141 -25382 8 VDD
port 41 nsew
rlabel nwell s 47847 -25576 48369 -25382 8 VDD
port 41 nsew
rlabel nwell s 49076 -25382 50141 -25375 8 VDD
port 41 nsew
rlabel nwell s 47847 -25382 48456 -25375 8 VDD
port 41 nsew
rlabel nwell s 47847 -25375 50141 -24827 8 VDD
port 41 nsew
rlabel nwell s 62157 -24502 64457 -24322 8 VDD
port 41 nsew
rlabel nwell s 57071 -24599 59371 -24419 8 VDD
port 41 nsew
rlabel nwell s 57071 -24419 58653 -24412 8 VDD
port 41 nsew
rlabel nwell s 62157 -24322 63739 -24315 8 VDD
port 41 nsew
rlabel nwell s 66798 -24167 67320 -24152 8 VDD
port 41 nsew
rlabel nwell s 65825 -24167 66543 -24123 8 VDD
port 41 nsew
rlabel nwell s 62157 -24315 63652 -24136 8 VDD
port 41 nsew
rlabel nwell s 57071 -24412 58566 -24233 8 VDD
port 41 nsew
rlabel nwell s 53377 -24762 55703 -24568 8 VDD
port 41 nsew
rlabel nwell s 47847 -24827 50173 -24633 8 VDD
port 41 nsew
rlabel nwell s 45626 -25756 46473 -25351 8 VDD
port 41 nsew
rlabel nwell s 44179 -25545 44701 -25351 8 VDD
port 41 nsew
rlabel nwell s 45408 -25351 46473 -25344 8 VDD
port 41 nsew
rlabel nwell s 44179 -25351 44788 -25344 8 VDD
port 41 nsew
rlabel nwell s 44179 -25344 46473 -24796 8 VDD
port 41 nsew
rlabel nwell s 53403 -24568 55703 -24388 8 VDD
port 41 nsew
rlabel nwell s 47873 -24633 50173 -24453 8 VDD
port 41 nsew
rlabel nwell s 47873 -24453 49455 -24446 8 VDD
port 41 nsew
rlabel nwell s 53403 -24388 54985 -24381 8 VDD
port 41 nsew
rlabel nwell s 58044 -24233 58566 -24218 8 VDD
port 41 nsew
rlabel nwell s 57071 -24233 57789 -24189 8 VDD
port 41 nsew
rlabel nwell s 53403 -24381 54898 -24202 8 VDD
port 41 nsew
rlabel nwell s 47873 -24446 49368 -24267 8 VDD
port 41 nsew
rlabel nwell s 44179 -24796 46505 -24602 8 VDD
port 41 nsew
rlabel nwell s 40431 -25748 41278 -25343 8 VDD
port 41 nsew
rlabel nwell s 38984 -25537 39506 -25343 8 VDD
port 41 nsew
rlabel nwell s 40213 -25343 41278 -25336 8 VDD
port 41 nsew
rlabel nwell s 38984 -25343 39593 -25336 8 VDD
port 41 nsew
rlabel nwell s 38984 -25336 41278 -24788 8 VDD
port 41 nsew
rlabel nwell s 44205 -24602 46505 -24422 8 VDD
port 41 nsew
rlabel nwell s 44205 -24422 45787 -24415 8 VDD
port 41 nsew
rlabel nwell s 48846 -24267 49368 -24252 8 VDD
port 41 nsew
rlabel nwell s 47873 -24267 48591 -24223 8 VDD
port 41 nsew
rlabel nwell s 44205 -24415 45700 -24236 8 VDD
port 41 nsew
rlabel nwell s 38984 -24788 41310 -24594 8 VDD
port 41 nsew
rlabel nwell s 36763 -25717 37610 -25312 8 VDD
port 41 nsew
rlabel nwell s 35316 -25506 35838 -25312 8 VDD
port 41 nsew
rlabel nwell s 36545 -25312 37610 -25305 8 VDD
port 41 nsew
rlabel nwell s 35316 -25312 35925 -25305 8 VDD
port 41 nsew
rlabel nwell s 35316 -25305 37610 -24757 8 VDD
port 41 nsew
rlabel nwell s 31991 -25737 32838 -25332 8 VDD
port 41 nsew
rlabel nwell s 30544 -25526 31066 -25332 8 VDD
port 41 nsew
rlabel nwell s 31773 -25332 32838 -25325 8 VDD
port 41 nsew
rlabel nwell s 30544 -25332 31153 -25325 8 VDD
port 41 nsew
rlabel nwell s 30544 -25325 32838 -24777 8 VDD
port 41 nsew
rlabel nwell s 39010 -24594 41310 -24414 8 VDD
port 41 nsew
rlabel nwell s 39010 -24414 40592 -24407 8 VDD
port 41 nsew
rlabel nwell s 45178 -24236 45700 -24221 8 VDD
port 41 nsew
rlabel nwell s 54376 -24202 54898 -24187 8 VDD
port 41 nsew
rlabel nwell s 53403 -24202 54121 -24158 8 VDD
port 41 nsew
rlabel nwell s 44205 -24236 44923 -24192 8 VDD
port 41 nsew
rlabel nwell s 39010 -24407 40505 -24228 8 VDD
port 41 nsew
rlabel nwell s 35316 -24757 37642 -24563 8 VDD
port 41 nsew
rlabel nwell s 30544 -24777 32870 -24583 8 VDD
port 41 nsew
rlabel nwell s 28323 -25706 29170 -25301 8 VDD
port 41 nsew
rlabel nwell s 26876 -25495 27398 -25301 8 VDD
port 41 nsew
rlabel nwell s 10524 -25922 16482 -25469 8 VDD
port 41 nsew
rlabel nwell s 13746 -25469 16482 -25468 8 VDD
port 41 nsew
rlabel nwell s -19151 -25955 -16857 -25407 2 VDD
port 41 nsew
rlabel nwell s -17922 -25407 -16857 -25400 2 VDD
port 41 nsew
rlabel nwell s -19151 -25407 -18542 -25400 2 VDD
port 41 nsew
rlabel nwell s 28105 -25301 29170 -25294 8 VDD
port 41 nsew
rlabel nwell s 26876 -25301 27485 -25294 8 VDD
port 41 nsew
rlabel nwell s 26876 -25294 29170 -24746 8 VDD
port 41 nsew
rlabel nwell s 19188 -25079 20613 -25078 8 VDD
port 41 nsew
rlabel nwell s 35342 -24563 37642 -24383 8 VDD
port 41 nsew
rlabel nwell s 30570 -24583 32870 -24403 8 VDD
port 41 nsew
rlabel nwell s 30570 -24403 32152 -24396 8 VDD
port 41 nsew
rlabel nwell s 35342 -24383 36924 -24376 8 VDD
port 41 nsew
rlabel nwell s 39983 -24228 40505 -24213 8 VDD
port 41 nsew
rlabel nwell s 39010 -24228 39728 -24184 8 VDD
port 41 nsew
rlabel nwell s 35342 -24376 36837 -24197 8 VDD
port 41 nsew
rlabel nwell s 30570 -24396 32065 -24217 8 VDD
port 41 nsew
rlabel nwell s 26876 -24746 29202 -24552 8 VDD
port 41 nsew
rlabel nwell s 26902 -24552 29202 -24372 8 VDD
port 41 nsew
rlabel nwell s 26902 -24372 28484 -24365 8 VDD
port 41 nsew
rlabel nwell s 31543 -24217 32065 -24202 8 VDD
port 41 nsew
rlabel nwell s 36315 -24197 36837 -24182 8 VDD
port 41 nsew
rlabel nwell s 35342 -24197 36060 -24153 8 VDD
port 41 nsew
rlabel nwell s 30570 -24217 31288 -24173 8 VDD
port 41 nsew
rlabel nwell s 26902 -24365 28397 -24186 8 VDD
port 41 nsew
rlabel nwell s 27875 -24186 28397 -24171 8 VDD
port 41 nsew
rlabel nwell s 26902 -24186 27620 -24142 8 VDD
port 41 nsew
rlabel nwell s 63130 -24136 63652 -24121 8 VDD
port 41 nsew
rlabel nwell s 72283 -24119 72805 -24104 8 VDD
port 41 nsew
rlabel nwell s 81647 -24081 82169 -24066 8 VDD
port 41 nsew
rlabel nwell s 80674 -24081 81392 -24037 8 VDD
port 41 nsew
rlabel nwell s 71310 -24119 72028 -24075 8 VDD
port 41 nsew
rlabel nwell s 62157 -24136 62875 -24092 8 VDD
port 41 nsew
rlabel nwell s 21927 -25074 24653 -24042 8 VDD
port 41 nsew
rlabel nwell s 21047 -25066 21667 -24613 8 VDD
port 41 nsew
rlabel nwell s 19188 -25078 20644 -24620 8 VDD
port 41 nsew
rlabel nwell s 18272 -25067 18907 -24386 8 VDD
port 41 nsew
rlabel nwell s 17326 -25067 17961 -24386 8 VDD
port 41 nsew
rlabel nwell s -7326 -25303 7434 -24917 8 VDD
port 41 nsew
rlabel nwell s -15200 -25034 -12464 -25033 2 VDD
port 41 nsew
rlabel nwell s 1295 -24917 7434 -24915 8 VDD
port 41 nsew
rlabel nwell s 2900 -24915 7434 -24908 8 VDD
port 41 nsew
rlabel nwell s 1295 -24915 1904 -24910 8 VDD
port 41 nsew
rlabel nwell s 2987 -24908 7434 -24828 8 VDD
port 41 nsew
rlabel nwell s 2987 -24828 3509 -24714 8 VDD
port 41 nsew
rlabel nwell s 1382 -24910 1904 -24716 8 VDD
port 41 nsew
rlabel nwell s -7326 -24917 300 -24847 2 VDD
port 41 nsew
rlabel nwell s -1686 -24847 300 -24830 2 VDD
port 41 nsew
rlabel nwell s -2313 -24847 -1972 -24836 2 VDD
port 41 nsew
rlabel nwell s -15200 -25033 -9242 -24580 2 VDD
port 41 nsew
rlabel nwell s -17704 -25400 -16857 -24995 2 VDD
port 41 nsew
rlabel nwell s -19151 -25400 -18629 -25206 2 VDD
port 41 nsew
rlabel nwell s -10187 -24580 -9846 -24569 2 VDD
port 41 nsew
rlabel nwell s -20553 -24801 -19918 -24120 2 VDD
port 41 nsew
rlabel nwell s -21458 -24800 -20823 -24119 2 VDD
port 41 nsew
rlabel nwell s -22664 -25071 -21719 -24126 2 VDD
port 41 nsew
rlabel nwell s -4612 -23859 -3771 -23853 2 VDD
port 41 nsew
rlabel nwell s 21097 -23636 21619 -23082 8 VDD
port 41 nsew
rlabel nwell s -7313 -23853 -2251 -23400 2 VDD
port 41 nsew
rlabel nwell s -7313 -23400 -4577 -23399 2 VDD
port 41 nsew
rlabel nwell s -8896 -24003 -8049 -23126 2 VDD
port 41 nsew
rlabel nwell s -12486 -23592 -11645 -23586 2 VDD
port 41 nsew
rlabel nwell s -15187 -23586 -10125 -23133 2 VDD
port 41 nsew
rlabel nwell s -15187 -23133 -12451 -23132 2 VDD
port 41 nsew
rlabel nwell s 21874 -22814 24610 -22813 8 VDD
port 41 nsew
rlabel nwell s 21086 -23082 21619 -22813 8 VDD
port 41 nsew
rlabel nwell s 17330 -22813 24610 -22360 8 VDD
port 41 nsew
rlabel nwell s -7313 -22545 -4577 -22544 2 VDD
port 41 nsew
rlabel nwell s 19256 -22360 19597 -22349 8 VDD
port 41 nsew
rlabel nwell s 84095 -21906 85572 -21033 8 VDD
port 41 nsew
rlabel nwell s 82103 -22148 82950 -21743 8 VDD
port 41 nsew
rlabel nwell s 80656 -21937 81178 -21743 8 VDD
port 41 nsew
rlabel nwell s 81885 -21743 82950 -21736 8 VDD
port 41 nsew
rlabel nwell s 80656 -21743 81265 -21736 8 VDD
port 41 nsew
rlabel nwell s 80656 -21736 82950 -21188 8 VDD
port 41 nsew
rlabel nwell s 80656 -21188 82982 -20994 8 VDD
port 41 nsew
rlabel nwell s 74731 -21944 76208 -21071 8 VDD
port 41 nsew
rlabel nwell s 72739 -22186 73586 -21781 8 VDD
port 41 nsew
rlabel nwell s 71292 -21975 71814 -21781 8 VDD
port 41 nsew
rlabel nwell s 72521 -21781 73586 -21774 8 VDD
port 41 nsew
rlabel nwell s 71292 -21781 71901 -21774 8 VDD
port 41 nsew
rlabel nwell s 71292 -21774 73586 -21226 8 VDD
port 41 nsew
rlabel nwell s 71292 -21226 73618 -21032 8 VDD
port 41 nsew
rlabel nwell s 65578 -21961 67055 -21088 8 VDD
port 41 nsew
rlabel nwell s 63586 -22203 64433 -21798 8 VDD
port 41 nsew
rlabel nwell s 62139 -21992 62661 -21798 8 VDD
port 41 nsew
rlabel nwell s 63368 -21798 64433 -21791 8 VDD
port 41 nsew
rlabel nwell s 62139 -21798 62748 -21791 8 VDD
port 41 nsew
rlabel nwell s 62139 -21791 64433 -21243 8 VDD
port 41 nsew
rlabel nwell s 62139 -21243 64465 -21049 8 VDD
port 41 nsew
rlabel nwell s 56824 -22027 58301 -21154 8 VDD
port 41 nsew
rlabel nwell s 54832 -22269 55679 -21864 8 VDD
port 41 nsew
rlabel nwell s 53385 -22058 53907 -21864 8 VDD
port 41 nsew
rlabel nwell s 54614 -21864 55679 -21857 8 VDD
port 41 nsew
rlabel nwell s 53385 -21864 53994 -21857 8 VDD
port 41 nsew
rlabel nwell s 53385 -21857 55679 -21309 8 VDD
port 41 nsew
rlabel nwell s 53385 -21309 55711 -21115 8 VDD
port 41 nsew
rlabel nwell s 47626 -22061 49103 -21188 8 VDD
port 41 nsew
rlabel nwell s 45634 -22303 46481 -21898 8 VDD
port 41 nsew
rlabel nwell s 44187 -22092 44709 -21898 8 VDD
port 41 nsew
rlabel nwell s 45416 -21898 46481 -21891 8 VDD
port 41 nsew
rlabel nwell s 44187 -21898 44796 -21891 8 VDD
port 41 nsew
rlabel nwell s 44187 -21891 46481 -21343 8 VDD
port 41 nsew
rlabel nwell s 44187 -21343 46513 -21149 8 VDD
port 41 nsew
rlabel nwell s 38763 -22022 40240 -21149 8 VDD
port 41 nsew
rlabel nwell s 36771 -22264 37618 -21859 8 VDD
port 41 nsew
rlabel nwell s 35324 -22053 35846 -21859 8 VDD
port 41 nsew
rlabel nwell s 36553 -21859 37618 -21852 8 VDD
port 41 nsew
rlabel nwell s 35324 -21859 35933 -21852 8 VDD
port 41 nsew
rlabel nwell s 35324 -21852 37618 -21304 8 VDD
port 41 nsew
rlabel nwell s 80682 -20994 82982 -20814 8 VDD
port 41 nsew
rlabel nwell s 71318 -21032 73618 -20852 8 VDD
port 41 nsew
rlabel nwell s 62165 -21049 64465 -20869 8 VDD
port 41 nsew
rlabel nwell s 53411 -21115 55711 -20935 8 VDD
port 41 nsew
rlabel nwell s 44213 -21149 46513 -20969 8 VDD
port 41 nsew
rlabel nwell s 44213 -20969 45795 -20962 8 VDD
port 41 nsew
rlabel nwell s 53411 -20935 54993 -20928 8 VDD
port 41 nsew
rlabel nwell s 62165 -20869 63747 -20862 8 VDD
port 41 nsew
rlabel nwell s 71318 -20852 72900 -20845 8 VDD
port 41 nsew
rlabel nwell s 80682 -20814 82264 -20807 8 VDD
port 41 nsew
rlabel nwell s 80682 -20807 82177 -20628 8 VDD
port 41 nsew
rlabel nwell s 71318 -20845 72813 -20666 8 VDD
port 41 nsew
rlabel nwell s 62165 -20862 63660 -20683 8 VDD
port 41 nsew
rlabel nwell s 53411 -20928 54906 -20749 8 VDD
port 41 nsew
rlabel nwell s 44213 -20962 45708 -20783 8 VDD
port 41 nsew
rlabel nwell s 35324 -21304 37650 -21110 8 VDD
port 41 nsew
rlabel nwell s 30323 -22011 31800 -21138 8 VDD
port 41 nsew
rlabel nwell s 28331 -22253 29178 -21848 8 VDD
port 41 nsew
rlabel nwell s 26884 -22042 27406 -21848 8 VDD
port 41 nsew
rlabel nwell s 28113 -21848 29178 -21841 8 VDD
port 41 nsew
rlabel nwell s 26884 -21848 27493 -21841 8 VDD
port 41 nsew
rlabel nwell s 26884 -21841 29178 -21293 8 VDD
port 41 nsew
rlabel nwell s 17331 -22360 18276 -21840 8 VDD
port 41 nsew
rlabel nwell s -7313 -22544 -2251 -22091 2 VDD
port 41 nsew
rlabel nwell s -13163 -22506 -12641 -22491 2 VDD
port 41 nsew
rlabel nwell s -14136 -22535 -13418 -22491 2 VDD
port 41 nsew
rlabel nwell s -14136 -22491 -12641 -22312 2 VDD
port 41 nsew
rlabel nwell s -14136 -22312 -12554 -22305 2 VDD
port 41 nsew
rlabel nwell s -14136 -22305 -11836 -22125 2 VDD
port 41 nsew
rlabel nwell s -4612 -22091 -3771 -22085 2 VDD
port 41 nsew
rlabel nwell s -14162 -22125 -11836 -21931 2 VDD
port 41 nsew
rlabel nwell s -14162 -21931 -11868 -21383 2 VDD
port 41 nsew
rlabel nwell s -12933 -21383 -11868 -21376 2 VDD
port 41 nsew
rlabel nwell s -14162 -21383 -13553 -21376 2 VDD
port 41 nsew
rlabel nwell s 21055 -21372 21896 -21366 8 VDD
port 41 nsew
rlabel nwell s 35350 -21110 37650 -20930 8 VDD
port 41 nsew
rlabel nwell s 35350 -20930 36932 -20923 8 VDD
port 41 nsew
rlabel nwell s 45186 -20783 45708 -20768 8 VDD
port 41 nsew
rlabel nwell s 54384 -20749 54906 -20734 8 VDD
port 41 nsew
rlabel nwell s 53411 -20749 54129 -20705 8 VDD
port 41 nsew
rlabel nwell s 44213 -20783 44931 -20739 8 VDD
port 41 nsew
rlabel nwell s 35350 -20923 36845 -20744 8 VDD
port 41 nsew
rlabel nwell s 26884 -21293 29210 -21099 8 VDD
port 41 nsew
rlabel nwell s 26910 -21099 29210 -20919 8 VDD
port 41 nsew
rlabel nwell s 26910 -20919 28492 -20912 8 VDD
port 41 nsew
rlabel nwell s 19535 -21366 24597 -20913 8 VDD
port 41 nsew
rlabel nwell s 2987 -21230 3509 -21116 8 VDD
port 41 nsew
rlabel nwell s 2987 -21116 7434 -21036 8 VDD
port 41 nsew
rlabel nwell s 2900 -21036 7434 -21029 8 VDD
port 41 nsew
rlabel nwell s 1382 -21228 1904 -21034 8 VDD
port 41 nsew
rlabel nwell s -1686 -21114 300 -21097 2 VDD
port 41 nsew
rlabel nwell s -2313 -21108 -1972 -21097 2 VDD
port 41 nsew
rlabel nwell s 1295 -21034 1904 -21029 8 VDD
port 41 nsew
rlabel nwell s 1295 -21029 7434 -21027 8 VDD
port 41 nsew
rlabel nwell s -7326 -21097 300 -21027 2 VDD
port 41 nsew
rlabel nwell s 21861 -20913 24597 -20912 8 VDD
port 41 nsew
rlabel nwell s 36323 -20744 36845 -20729 8 VDD
port 41 nsew
rlabel nwell s 35350 -20744 36068 -20700 8 VDD
port 41 nsew
rlabel nwell s 26910 -20912 28405 -20733 8 VDD
port 41 nsew
rlabel nwell s 27883 -20733 28405 -20718 8 VDD
port 41 nsew
rlabel nwell s 26910 -20733 27628 -20689 8 VDD
port 41 nsew
rlabel nwell s 63138 -20683 63660 -20668 8 VDD
port 41 nsew
rlabel nwell s 72291 -20666 72813 -20651 8 VDD
port 41 nsew
rlabel nwell s 81655 -20628 82177 -20613 8 VDD
port 41 nsew
rlabel nwell s 80682 -20628 81400 -20584 8 VDD
port 41 nsew
rlabel nwell s 71318 -20666 72036 -20622 8 VDD
port 41 nsew
rlabel nwell s 62165 -20683 62883 -20639 8 VDD
port 41 nsew
rlabel nwell s -7326 -21027 7434 -20641 8 VDD
port 41 nsew
rlabel nwell s -12715 -21376 -11868 -20971 2 VDD
port 41 nsew
rlabel nwell s -14162 -21376 -13640 -21182 2 VDD
port 41 nsew
rlabel nwell s -18152 -21530 -17630 -21515 2 VDD
port 41 nsew
rlabel nwell s -19125 -21559 -18407 -21515 2 VDD
port 41 nsew
rlabel nwell s -19125 -21515 -17630 -21336 2 VDD
port 41 nsew
rlabel nwell s -22729 -21577 -22207 -21383 2 VDD
port 41 nsew
rlabel nwell s -19125 -21336 -17543 -21329 2 VDD
port 41 nsew
rlabel nwell s -19125 -21329 -16825 -21149 2 VDD
port 41 nsew
rlabel nwell s -19151 -21149 -16825 -20955 2 VDD
port 41 nsew
rlabel nwell s -19151 -20955 -16857 -20407 2 VDD
port 41 nsew
rlabel nwell s -20956 -21382 -19500 -20924 2 VDD
port 41 nsew
rlabel nwell s -22729 -21383 -22120 -21376 2 VDD
port 41 nsew
rlabel nwell s -22729 -21376 -21402 -21002 2 VDD
port 41 nsew
rlabel nwell s -20956 -20924 -19531 -20923 2 VDD
port 41 nsew
rlabel nwell s -17922 -20407 -16857 -20400 2 VDD
port 41 nsew
rlabel nwell s -19151 -20407 -18542 -20400 2 VDD
port 41 nsew
rlabel nwell s -7056 -20323 -6436 -19870 2 VDD
port 41 nsew
rlabel nwell s -15200 -20107 -12464 -20106 2 VDD
port 41 nsew
rlabel nwell s -15200 -20106 -9242 -19653 2 VDD
port 41 nsew
rlabel nwell s -17704 -20400 -16857 -19995 2 VDD
port 41 nsew
rlabel nwell s -19151 -20400 -18629 -20206 2 VDD
port 41 nsew
rlabel nwell s -10187 -19653 -9846 -19642 2 VDD
port 41 nsew
rlabel nwell s -20787 -19668 -20265 -19474 2 VDD
port 41 nsew
rlabel nwell s -20787 -19474 -20178 -19467 2 VDD
port 41 nsew
rlabel nwell s -20787 -19467 -19460 -19093 2 VDD
port 41 nsew
rlabel nwell s 5507 -18865 7424 -18792 8 VDD
port 41 nsew
rlabel nwell s 2507 -18865 4424 -18792 8 VDD
port 41 nsew
rlabel nwell s 7 -18865 1924 -18792 8 VDD
port 41 nsew
rlabel nwell s -2493 -18865 -576 -18792 2 VDD
port 41 nsew
rlabel nwell s -4993 -18865 -3076 -18792 2 VDD
port 41 nsew
rlabel nwell s -7493 -18865 -5576 -18792 2 VDD
port 41 nsew
rlabel nwell s 5506 -18792 7424 -18390 8 VDD
port 41 nsew
rlabel nwell s 2506 -18792 4424 -18390 8 VDD
port 41 nsew
rlabel nwell s 6 -18792 1924 -18390 8 VDD
port 41 nsew
rlabel nwell s -2494 -18792 -576 -18390 2 VDD
port 41 nsew
rlabel nwell s -4994 -18792 -3076 -18390 2 VDD
port 41 nsew
rlabel nwell s -7494 -18792 -5576 -18390 2 VDD
port 41 nsew
rlabel nwell s -8923 -19069 -8076 -18192 2 VDD
port 41 nsew
rlabel nwell s -22786 -19446 -21330 -18988 2 VDD
port 41 nsew
rlabel nwell s -22786 -18988 -21361 -18987 2 VDD
port 41 nsew
rlabel nwell s -12486 -18665 -11645 -18659 2 VDD
port 41 nsew
rlabel nwell s -15187 -18659 -10125 -18206 2 VDD
port 41 nsew
rlabel nwell s -15187 -18206 -12451 -18205 2 VDD
port 41 nsew
rlabel nwell s -15097 -16843 -7497 -16074 2 VDD
port 41 nsew
rlabel nwell s 63195 -4347 64755 -3851 8 VDD
port 41 nsew
rlabel nwell s 62345 -3100 64755 -2604 8 VDD
port 41 nsew
rlabel nwell s 50645 -3386 58245 -2617 8 VDD
port 41 nsew
rlabel nwell s 5332 -1986 6892 -1490 8 VDD
port 41 nsew
rlabel nwell s 20768 -1481 22328 -985 8 VDD
port 41 nsew
rlabel nwell s -4250 -1844 -2690 -1348 2 VDD
port 41 nsew
rlabel nwell s 50645 -339 58245 430 6 VDD
port 41 nsew
rlabel nwell s 19918 -234 22328 262 6 VDD
port 41 nsew
rlabel nwell s 7529 -961 15129 -192 8 VDD
port 41 nsew
rlabel nwell s 4482 -739 6892 -243 8 VDD
port 41 nsew
rlabel nwell s -5100 -597 -2690 -101 2 VDD
port 41 nsew
rlabel nwell s 42347 1225 45083 1226 6 VDD
port 41 nsew
rlabel nwell s 45531 1316 46151 1769 6 VDD
port 41 nsew
rlabel nwell s 40021 1226 45083 1679 6 VDD
port 41 nsew
rlabel nwell s 41541 1679 42382 1685 6 VDD
port 41 nsew
rlabel nwell s 36738 444 38132 1881 6 VDD
port 41 nsew
rlabel nwell s 35017 401 36411 1924 6 VDD
port 41 nsew
rlabel nwell s 34124 1398 34412 1399 6 VDD
port 41 nsew
rlabel nwell s 32528 1399 34412 2046 6 VDD
port 41 nsew
rlabel nwell s 30282 378 31676 1902 6 VDD
port 41 nsew
rlabel nwell s 5317 704 6877 1200 6 VDD
port 41 nsew
rlabel nwell s 1717 935 1921 979 6 VDD
port 41 nsew
rlabel nwell s 1717 979 2979 981 6 VDD
port 41 nsew
rlabel nwell s 577 979 913 981 6 VDD
port 41 nsew
rlabel nwell s 29269 1405 29557 1406 6 VDD
port 41 nsew
rlabel nwell s 32916 2046 34412 2117 6 VDD
port 41 nsew
rlabel nwell s 32916 2117 34125 2375 6 VDD
port 41 nsew
rlabel nwell s 27673 1406 29557 2053 6 VDD
port 41 nsew
rlabel nwell s 28061 2053 29557 2124 6 VDD
port 41 nsew
rlabel nwell s 28061 2124 29270 2382 6 VDD
port 41 nsew
rlabel nwell s 20596 1869 22156 2365 6 VDD
port 41 nsew
rlabel nwell s 7570 1795 15170 2564 6 VDD
port 41 nsew
rlabel nwell s 577 981 2979 1881 6 VDD
port 41 nsew
rlabel nwell s -2782 528 -1222 1024 4 VDD
port 41 nsew
rlabel nwell s 1717 1881 2979 1883 6 VDD
port 41 nsew
rlabel nwell s 577 1881 913 1883 6 VDD
port 41 nsew
rlabel nwell s 1717 1883 1921 1927 6 VDD
port 41 nsew
rlabel nwell s 4467 1951 6877 2447 6 VDD
port 41 nsew
rlabel nwell s -3632 1775 -1222 2271 4 VDD
port 41 nsew
rlabel nwell s -13457 1513 -5857 2282 4 VDD
port 41 nsew
rlabel nwell s 50848 2572 58448 3341 6 VDD
port 41 nsew
rlabel nwell s 39742 2662 40083 2673 6 VDD
port 41 nsew
rlabel nwell s 39138 2673 45096 3126 6 VDD
port 41 nsew
rlabel nwell s 42360 3126 45096 3127 6 VDD
port 41 nsew
rlabel nwell s 19746 3116 22156 3612 6 VDD
port 41 nsew
rlabel nwell s 8190 6589 12714 6634 6 VDD
port 41 nsew
rlabel nwell s 8096 6634 12765 7919 6 VDD
port 41 nsew
rlabel nwell s 15664 8806 15948 9053 6 VDD
port 41 nsew
rlabel nwell s 14469 9053 15950 10215 6 VDD
port 41 nsew
rlabel nwell s -14092 10312 -13634 10343 4 VDD
port 41 nsew
rlabel nwell s -5915 10527 -5456 11952 4 VDD
port 41 nsew
rlabel nwell s -8046 10584 -7471 11106 4 VDD
port 41 nsew
rlabel nwell s -7852 11106 -7471 11193 4 VDD
port 41 nsew
rlabel nwell s -7845 11193 -7471 11911 4 VDD
port 41 nsew
rlabel nwell s -11540 10649 -10595 11594 4 VDD
port 41 nsew
rlabel nwell s -14093 10343 -13634 11768 4 VDD
port 41 nsew
rlabel nwell s -5915 11952 -5457 11983 4 VDD
port 41 nsew
rlabel nwell s -6137 12526 -5562 13048 4 VDD
port 41 nsew
rlabel nwell s -5943 13048 -5562 13135 4 VDD
port 41 nsew
rlabel nwell s -5936 13135 -5562 13853 4 VDD
port 41 nsew
rlabel nwell s -7851 12357 -7392 13782 4 VDD
port 41 nsew
rlabel nwell s -11269 11855 -10588 12490 4 VDD
port 41 nsew
rlabel nwell s -11270 12760 -10589 13395 4 VDD
port 41 nsew
rlabel nwell s -7851 13782 -7393 13813 4 VDD
port 41 nsew
rlabel nwell s -7618 14162 -6675 14188 4 VDD
port 41 nsew
rlabel nwell s -12618 14162 -11675 14188 4 VDD
port 41 nsew
rlabel nwell s -8028 14188 -6675 14684 4 VDD
port 41 nsew
rlabel nwell s -13028 14188 -11675 14684 4 VDD
port 41 nsew
rlabel nwell s -8028 14684 -6869 14771 4 VDD
port 41 nsew
rlabel nwell s -13028 14684 -11869 14771 4 VDD
port 41 nsew
rlabel nwell s -8028 14771 -6876 14906 4 VDD
port 41 nsew
rlabel nwell s -13028 14771 -11876 14906 4 VDD
port 41 nsew
rlabel nwell s -7984 14906 -6876 15161 4 VDD
port 41 nsew
rlabel nwell s -12984 14906 -11876 15161 4 VDD
port 41 nsew
rlabel nwell s -7999 15161 -6876 15391 4 VDD
port 41 nsew
rlabel nwell s -12999 15161 -11876 15391 4 VDD
port 41 nsew
rlabel nwell s -7999 15391 -6869 15609 4 VDD
port 41 nsew
rlabel nwell s -12999 15391 -11869 15609 4 VDD
port 41 nsew
rlabel nwell s -7999 15609 -6464 15683 4 VDD
port 41 nsew
rlabel nwell s -12999 15609 -11464 15683 4 VDD
port 41 nsew
rlabel nwell s -7805 15683 -6464 15770 4 VDD
port 41 nsew
rlabel nwell s -12805 15683 -11464 15770 4 VDD
port 41 nsew
rlabel nwell s -7798 15770 -6464 16456 4 VDD
port 41 nsew
rlabel nwell s -12798 15770 -11464 16456 4 VDD
port 41 nsew
rlabel nwell s -7798 16456 -7424 16488 4 VDD
port 41 nsew
rlabel nwell s -12798 16456 -12424 16488 4 VDD
port 41 nsew
rlabel nwell s -5128 18126 -4674 20827 4 VDD
port 41 nsew
rlabel nwell s -5134 20827 -4674 20862 4 VDD
port 41 nsew
rlabel nwell s -5134 20862 -4675 21668 4 VDD
port 41 nsew
rlabel nwell s -6576 18113 -6122 20849 4 VDD
port 41 nsew
rlabel nwell s -8594 19151 -7651 19177 4 VDD
port 41 nsew
rlabel nwell s -9004 19177 -7651 19673 4 VDD
port 41 nsew
rlabel nwell s -9004 19673 -7845 19760 4 VDD
port 41 nsew
rlabel nwell s -9004 19760 -7852 19895 4 VDD
port 41 nsew
rlabel nwell s -8960 19895 -7852 20150 4 VDD
port 41 nsew
rlabel nwell s -8975 20150 -7852 20380 4 VDD
port 41 nsew
rlabel nwell s -8975 20380 -7845 20598 4 VDD
port 41 nsew
rlabel nwell s -8975 20598 -7440 20672 4 VDD
port 41 nsew
rlabel nwell s -8781 20672 -7440 20759 4 VDD
port 41 nsew
rlabel nwell s -5128 21668 -4675 23188 4 VDD
port 41 nsew
rlabel nwell s -6575 20849 -6122 23126 4 VDD
port 41 nsew
rlabel nwell s -8774 20759 -7440 21445 4 VDD
port 41 nsew
rlabel nwell s -10055 18126 -9601 20827 4 VDD
port 41 nsew
rlabel nwell s -10061 20827 -9601 20862 4 VDD
port 41 nsew
rlabel nwell s -8774 21445 -8400 21477 4 VDD
port 41 nsew
rlabel nwell s -6575 23126 -6111 23467 4 VDD
port 41 nsew
rlabel nwell s -10061 20862 -9602 21668 4 VDD
port 41 nsew
rlabel nwell s -11503 18113 -11049 20849 4 VDD
port 41 nsew
rlabel nwell s -10055 21668 -9602 23188 4 VDD
port 41 nsew
rlabel nwell s -11502 20849 -11049 23126 4 VDD
port 41 nsew
rlabel nwell s -11502 23126 -11038 23467 4 VDD
port 41 nsew
rlabel nwell s -6575 23467 -6122 24071 4 VDD
port 41 nsew
rlabel nwell s -11502 23467 -11049 24071 4 VDD
port 41 nsew
rlabel nwell s -5538 24390 -4661 25237 4 VDD
port 41 nsew
rlabel nwell s -10472 24417 -9595 25264 4 VDD
port 41 nsew
rlabel nwell s -5261 25819 -4859 25820 4 VDD
port 41 nsew
rlabel nwell s -14023 25819 -13621 25820 4 VDD
port 41 nsew
rlabel nwell s -5334 25820 -4859 27737 4 VDD
port 41 nsew
rlabel nwell s -6792 26257 -6339 26877 4 VDD
port 41 nsew
rlabel nwell s -5261 28319 -4859 28320 4 VDD
port 41 nsew
rlabel nwell s -5334 28320 -4859 30237 4 VDD
port 41 nsew
rlabel nwell s -5261 30819 -4859 30820 4 VDD
port 41 nsew
rlabel nwell s -5334 30820 -4859 32737 4 VDD
port 41 nsew
rlabel nwell s -7566 25987 -7110 31000 4 VDD
port 41 nsew
rlabel nwell s -9014 26000 -8560 28701 4 VDD
port 41 nsew
rlabel nwell s -9014 28701 -8554 28736 4 VDD
port 41 nsew
rlabel nwell s -10322 26000 -9868 28701 4 VDD
port 41 nsew
rlabel nwell s -10328 28701 -9868 28736 4 VDD
port 41 nsew
rlabel nwell s -9013 28736 -8554 29542 4 VDD
port 41 nsew
rlabel nwell s -7577 31000 -7110 31341 4 VDD
port 41 nsew
rlabel nwell s -9013 29542 -8560 31062 4 VDD
port 41 nsew
rlabel nwell s -10328 28736 -9869 29542 4 VDD
port 41 nsew
rlabel nwell s -10322 29542 -9869 31062 4 VDD
port 41 nsew
rlabel nwell s -11772 25987 -11316 31000 4 VDD
port 41 nsew
rlabel nwell s -14023 25820 -13548 27737 4 VDD
port 41 nsew
rlabel nwell s -14023 28319 -13621 28320 4 VDD
port 41 nsew
rlabel nwell s -14023 28320 -13548 30237 4 VDD
port 41 nsew
rlabel nwell s -14023 30819 -13621 30820 4 VDD
port 41 nsew
rlabel nwell s -11772 31000 -11305 31341 4 VDD
port 41 nsew
rlabel nwell s -7566 31341 -7110 31627 4 VDD
port 41 nsew
rlabel nwell s -11772 31341 -11316 31627 4 VDD
port 41 nsew
rlabel nwell s -5261 33319 -4859 33320 4 VDD
port 41 nsew
rlabel nwell s -5334 33320 -4859 35237 4 VDD
port 41 nsew
rlabel nwell s -7583 31627 -7110 33613 4 VDD
port 41 nsew
rlabel nwell s -11772 31627 -11299 33613 4 VDD
port 41 nsew
rlabel nwell s -14023 30820 -13548 32737 4 VDD
port 41 nsew
rlabel nwell s -14023 33319 -13621 33320 4 VDD
port 41 nsew
rlabel nwell s -7496 33613 -7110 34608 4 VDD
port 41 nsew
rlabel nwell s -11772 33613 -11386 34608 4 VDD
port 41 nsew
rlabel nwell s -7503 34608 -7110 34695 4 VDD
port 41 nsew
rlabel nwell s -11772 34608 -11379 34695 4 VDD
port 41 nsew
rlabel nwell s -7697 34695 -7110 35217 4 VDD
port 41 nsew
rlabel nwell s -11772 34695 -11185 35217 4 VDD
port 41 nsew
rlabel nwell s -5261 35819 -4859 35820 4 VDD
port 41 nsew
rlabel nwell s -5334 35820 -4859 37737 4 VDD
port 41 nsew
rlabel nwell s -7498 35217 -7110 36213 4 VDD
port 41 nsew
rlabel nwell s -11772 35217 -11384 36213 4 VDD
port 41 nsew
rlabel nwell s -14023 33320 -13548 35237 4 VDD
port 41 nsew
rlabel nwell s -14023 35819 -13621 35820 4 VDD
port 41 nsew
rlabel nwell s -7505 36213 -7110 36300 4 VDD
port 41 nsew
rlabel nwell s -11772 36213 -11377 36300 4 VDD
port 41 nsew
rlabel nwell s -7699 36300 -7110 36822 4 VDD
port 41 nsew
rlabel nwell s -11772 36300 -11183 36822 4 VDD
port 41 nsew
rlabel nwell s -5261 38819 -4859 38820 4 VDD
port 41 nsew
rlabel nwell s -5334 38820 -4859 40737 4 VDD
port 41 nsew
rlabel nwell s -7585 36822 -7110 40747 4 VDD
port 41 nsew
rlabel nwell s -11772 36822 -11297 40747 4 VDD
port 41 nsew
rlabel nwell s -14023 35820 -13548 37737 4 VDD
port 41 nsew
rlabel nwell s -14023 38819 -13621 38820 4 VDD
port 41 nsew
rlabel nwell s -14023 38820 -13548 40737 4 VDD
port 41 nsew
rlabel nwell s -12391 43837 -11938 44441 4 VDD
port 41 nsew
rlabel nwell s -12402 44441 -11938 44782 4 VDD
port 41 nsew
rlabel nwell s -12391 44782 -11938 47059 4 VDD
port 41 nsew
rlabel nwell s -13838 44720 -13385 46240 4 VDD
port 41 nsew
rlabel nwell s -12391 47059 -11937 49795 4 VDD
port 41 nsew
rlabel nwell s -13838 46240 -13379 47046 4 VDD
port 41 nsew
rlabel nwell s -13839 47046 -13379 47081 4 VDD
port 41 nsew
rlabel nwell s -13839 47081 -13385 49782 4 VDD
port 41 nsew
rlabel nwell s -9282 50643 -8829 50644 4 VDD
port 41 nsew
rlabel nwell s -9282 50644 -8309 51589 4 VDD
port 41 nsew
rlabel nwell s -11536 50639 -10855 51274 4 VDD
port 41 nsew
rlabel nwell s -9282 51589 -8829 52569 4 VDD
port 41 nsew
rlabel nwell s -11536 51585 -10855 52220 4 VDD
port 41 nsew
rlabel nwell s -7835 52848 -7382 54368 4 VDD
port 41 nsew
rlabel nwell s -9282 52569 -8818 52910 4 VDD
port 41 nsew
rlabel nwell s -7841 54368 -7382 55174 4 VDD
port 41 nsew
rlabel nwell s -7841 55174 -7381 55209 4 VDD
port 41 nsew
rlabel nwell s -9282 52910 -8829 54399 4 VDD
port 41 nsew
rlabel nwell s -11548 52501 -11089 53926 4 VDD
port 41 nsew
rlabel nwell s -11547 53926 -11089 53957 4 VDD
port 41 nsew
rlabel nwell s -9551 54399 -8829 54410 4 VDD
port 41 nsew
rlabel nwell s -10105 54410 -8829 54932 4 VDD
port 41 nsew
rlabel nwell s -9282 54932 -8829 55187 4 VDD
port 41 nsew
rlabel nwell s -11535 54360 -11082 54980 4 VDD
port 41 nsew
rlabel nwell s -7835 55209 -7381 57910 4 VDD
port 41 nsew
rlabel nwell s -9283 55187 -8829 57923 4 VDD
port 41 nsew
rlabel nwell s -11543 55240 -10511 57966 4 VDD
port 41 nsew
rlabel nwell s -8511 60197 -7568 60223 4 VDD
port 41 nsew
rlabel nwell s -11964 60189 -11021 60215 4 VDD
port 41 nsew
rlabel nwell s -8511 60223 -7158 60719 4 VDD
port 41 nsew
rlabel nwell s -11964 60215 -10611 60711 4 VDD
port 41 nsew
rlabel nwell s -8317 60719 -7158 60806 4 VDD
port 41 nsew
rlabel nwell s -11770 60711 -10611 60798 4 VDD
port 41 nsew
rlabel nwell s -8310 60806 -7158 60941 4 VDD
port 41 nsew
rlabel nwell s -11763 60798 -10611 60933 4 VDD
port 41 nsew
rlabel nwell s -8310 60941 -7202 61196 4 VDD
port 41 nsew
rlabel nwell s -11763 60933 -10655 61188 4 VDD
port 41 nsew
rlabel nwell s -8310 61196 -7187 61426 4 VDD
port 41 nsew
rlabel nwell s -11763 61188 -10640 61418 4 VDD
port 41 nsew
rlabel nwell s -8317 61426 -7187 61644 4 VDD
port 41 nsew
rlabel nwell s -11770 61418 -10640 61636 4 VDD
port 41 nsew
rlabel nwell s -8722 61644 -7187 61718 4 VDD
port 41 nsew
rlabel nwell s -12175 61636 -10640 61710 4 VDD
port 41 nsew
rlabel nwell s -8722 61718 -7381 61805 4 VDD
port 41 nsew
rlabel nwell s -12175 61710 -10834 61797 4 VDD
port 41 nsew
rlabel nwell s -8722 61805 -7388 62491 4 VDD
port 41 nsew
rlabel nwell s -12175 61797 -10841 62483 4 VDD
port 41 nsew
rlabel nwell s -7762 62491 -7388 62523 4 VDD
port 41 nsew
rlabel nwell s -11215 62483 -10841 62515 4 VDD
port 41 nsew
rlabel nwell s -8480 63636 -7607 65113 4 VDD
port 41 nsew
rlabel nwell s -11995 63857 -11052 63883 4 VDD
port 41 nsew
rlabel nwell s -11995 63883 -10642 64379 4 VDD
port 41 nsew
rlabel nwell s -11801 64379 -10642 64466 4 VDD
port 41 nsew
rlabel nwell s -11794 64466 -10642 64601 4 VDD
port 41 nsew
rlabel nwell s -11794 64601 -10686 64856 4 VDD
port 41 nsew
rlabel nwell s -11794 64856 -10671 65086 4 VDD
port 41 nsew
rlabel nwell s -11801 65086 -10671 65304 4 VDD
port 41 nsew
rlabel nwell s -12206 65304 -10671 65378 4 VDD
port 41 nsew
rlabel nwell s -12206 65378 -10865 65465 4 VDD
port 41 nsew
rlabel nwell s -12206 65465 -10872 66151 4 VDD
port 41 nsew
rlabel nwell s -11246 66151 -10872 66183 4 VDD
port 41 nsew
rlabel nwell s -8522 68637 -7579 68663 4 VDD
port 41 nsew
rlabel nwell s -11975 68629 -11032 68655 4 VDD
port 41 nsew
rlabel nwell s -8522 68663 -7169 69159 4 VDD
port 41 nsew
rlabel nwell s -11975 68655 -10622 69151 4 VDD
port 41 nsew
rlabel nwell s -8328 69159 -7169 69246 4 VDD
port 41 nsew
rlabel nwell s -11781 69151 -10622 69238 4 VDD
port 41 nsew
rlabel nwell s -8321 69246 -7169 69381 4 VDD
port 41 nsew
rlabel nwell s -11774 69238 -10622 69373 4 VDD
port 41 nsew
rlabel nwell s -8321 69381 -7213 69636 4 VDD
port 41 nsew
rlabel nwell s -11774 69373 -10666 69628 4 VDD
port 41 nsew
rlabel nwell s -8321 69636 -7198 69866 4 VDD
port 41 nsew
rlabel nwell s -11774 69628 -10651 69858 4 VDD
port 41 nsew
rlabel nwell s -8328 69866 -7198 70084 4 VDD
port 41 nsew
rlabel nwell s -11781 69858 -10651 70076 4 VDD
port 41 nsew
rlabel nwell s -8733 70084 -7198 70158 4 VDD
port 41 nsew
rlabel nwell s -12186 70076 -10651 70150 4 VDD
port 41 nsew
rlabel nwell s -8733 70158 -7392 70245 4 VDD
port 41 nsew
rlabel nwell s -12186 70150 -10845 70237 4 VDD
port 41 nsew
rlabel nwell s -8733 70245 -7399 70931 4 VDD
port 41 nsew
rlabel nwell s -12186 70237 -10852 70923 4 VDD
port 41 nsew
rlabel nwell s -7773 70931 -7399 70963 4 VDD
port 41 nsew
rlabel nwell s -11226 70923 -10852 70955 4 VDD
port 41 nsew
rlabel nwell s -8491 72076 -7618 73553 4 VDD
port 41 nsew
rlabel nwell s -12006 72297 -11063 72323 4 VDD
port 41 nsew
rlabel nwell s -12006 72323 -10653 72819 4 VDD
port 41 nsew
rlabel nwell s -11812 72819 -10653 72906 4 VDD
port 41 nsew
rlabel nwell s -11805 72906 -10653 73041 4 VDD
port 41 nsew
rlabel nwell s -11805 73041 -10697 73296 4 VDD
port 41 nsew
rlabel nwell s -11805 73296 -10682 73526 4 VDD
port 41 nsew
rlabel nwell s -11812 73526 -10682 73744 4 VDD
port 41 nsew
rlabel nwell s -12217 73744 -10682 73818 4 VDD
port 41 nsew
rlabel nwell s -12217 73818 -10876 73905 4 VDD
port 41 nsew
rlabel nwell s -12217 73905 -10883 74591 4 VDD
port 41 nsew
rlabel nwell s -11257 74591 -10883 74623 4 VDD
port 41 nsew
rlabel nwell s -8561 77500 -7618 77526 4 VDD
port 41 nsew
rlabel nwell s -12014 77492 -11071 77518 4 VDD
port 41 nsew
rlabel nwell s -8561 77526 -7208 78022 4 VDD
port 41 nsew
rlabel nwell s -12014 77518 -10661 78014 4 VDD
port 41 nsew
rlabel nwell s -8367 78022 -7208 78109 4 VDD
port 41 nsew
rlabel nwell s -11820 78014 -10661 78101 4 VDD
port 41 nsew
rlabel nwell s -8360 78109 -7208 78244 4 VDD
port 41 nsew
rlabel nwell s -11813 78101 -10661 78236 4 VDD
port 41 nsew
rlabel nwell s -8360 78244 -7252 78499 4 VDD
port 41 nsew
rlabel nwell s -11813 78236 -10705 78491 4 VDD
port 41 nsew
rlabel nwell s -8360 78499 -7237 78729 4 VDD
port 41 nsew
rlabel nwell s -11813 78491 -10690 78721 4 VDD
port 41 nsew
rlabel nwell s -8367 78729 -7237 78947 4 VDD
port 41 nsew
rlabel nwell s -11820 78721 -10690 78939 4 VDD
port 41 nsew
rlabel nwell s -8772 78947 -7237 79021 4 VDD
port 41 nsew
rlabel nwell s -12225 78939 -10690 79013 4 VDD
port 41 nsew
rlabel nwell s -8772 79021 -7431 79108 4 VDD
port 41 nsew
rlabel nwell s -12225 79013 -10884 79100 4 VDD
port 41 nsew
rlabel nwell s -8772 79108 -7438 79794 4 VDD
port 41 nsew
rlabel nwell s -12225 79100 -10891 79786 4 VDD
port 41 nsew
rlabel nwell s -7812 79794 -7438 79826 4 VDD
port 41 nsew
rlabel nwell s -11265 79786 -10891 79818 4 VDD
port 41 nsew
rlabel nwell s -8530 80939 -7657 82416 4 VDD
port 41 nsew
rlabel nwell s -12045 81160 -11102 81186 4 VDD
port 41 nsew
rlabel nwell s -12045 81186 -10692 81682 4 VDD
port 41 nsew
rlabel nwell s -11851 81682 -10692 81769 4 VDD
port 41 nsew
rlabel nwell s -11844 81769 -10692 81904 4 VDD
port 41 nsew
rlabel nwell s -11844 81904 -10736 82159 4 VDD
port 41 nsew
rlabel nwell s -11844 82159 -10721 82389 4 VDD
port 41 nsew
rlabel nwell s -11851 82389 -10721 82607 4 VDD
port 41 nsew
rlabel nwell s -12256 82607 -10721 82681 4 VDD
port 41 nsew
rlabel nwell s -12256 82681 -10915 82768 4 VDD
port 41 nsew
rlabel nwell s -12256 82768 -10922 83454 4 VDD
port 41 nsew
rlabel nwell s -11296 83454 -10922 83486 4 VDD
port 41 nsew
rlabel nwell s -8527 86698 -7584 86724 4 VDD
port 41 nsew
rlabel nwell s -11980 86690 -11037 86716 4 VDD
port 41 nsew
rlabel nwell s -8527 86724 -7174 87220 4 VDD
port 41 nsew
rlabel nwell s -11980 86716 -10627 87212 4 VDD
port 41 nsew
rlabel nwell s -8333 87220 -7174 87307 4 VDD
port 41 nsew
rlabel nwell s -11786 87212 -10627 87299 4 VDD
port 41 nsew
rlabel nwell s -8326 87307 -7174 87442 4 VDD
port 41 nsew
rlabel nwell s -11779 87299 -10627 87434 4 VDD
port 41 nsew
rlabel nwell s -8326 87442 -7218 87697 4 VDD
port 41 nsew
rlabel nwell s -11779 87434 -10671 87689 4 VDD
port 41 nsew
rlabel nwell s -8326 87697 -7203 87927 4 VDD
port 41 nsew
rlabel nwell s -11779 87689 -10656 87919 4 VDD
port 41 nsew
rlabel nwell s -8333 87927 -7203 88145 4 VDD
port 41 nsew
rlabel nwell s -11786 87919 -10656 88137 4 VDD
port 41 nsew
rlabel nwell s -8738 88145 -7203 88219 4 VDD
port 41 nsew
rlabel nwell s -12191 88137 -10656 88211 4 VDD
port 41 nsew
rlabel nwell s -8738 88219 -7397 88306 4 VDD
port 41 nsew
rlabel nwell s -12191 88211 -10850 88298 4 VDD
port 41 nsew
rlabel nwell s -8738 88306 -7404 88992 4 VDD
port 41 nsew
rlabel nwell s -12191 88298 -10857 88984 4 VDD
port 41 nsew
rlabel nwell s -7778 88992 -7404 89024 4 VDD
port 41 nsew
rlabel nwell s -11231 88984 -10857 89016 4 VDD
port 41 nsew
rlabel nwell s -8496 90137 -7623 91614 4 VDD
port 41 nsew
rlabel nwell s -12011 90358 -11068 90384 4 VDD
port 41 nsew
rlabel nwell s -12011 90384 -10658 90880 4 VDD
port 41 nsew
rlabel nwell s -11817 90880 -10658 90967 4 VDD
port 41 nsew
rlabel nwell s -11810 90967 -10658 91102 4 VDD
port 41 nsew
rlabel nwell s -11810 91102 -10702 91357 4 VDD
port 41 nsew
rlabel nwell s -11810 91357 -10687 91587 4 VDD
port 41 nsew
rlabel nwell s -11817 91587 -10687 91805 4 VDD
port 41 nsew
rlabel nwell s -12222 91805 -10687 91879 4 VDD
port 41 nsew
rlabel nwell s -12222 91879 -10881 91966 4 VDD
port 41 nsew
rlabel nwell s -12222 91966 -10888 92652 4 VDD
port 41 nsew
rlabel nwell s -11262 92652 -10888 92684 4 VDD
port 41 nsew
rlabel nwell s -8461 95452 -7518 95478 4 VDD
port 41 nsew
rlabel nwell s -11914 95444 -10971 95470 4 VDD
port 41 nsew
rlabel nwell s -8461 95478 -7108 95974 4 VDD
port 41 nsew
rlabel nwell s -11914 95470 -10561 95966 4 VDD
port 41 nsew
rlabel nwell s -8267 95974 -7108 96061 4 VDD
port 41 nsew
rlabel nwell s -11720 95966 -10561 96053 4 VDD
port 41 nsew
rlabel nwell s -8260 96061 -7108 96196 4 VDD
port 41 nsew
rlabel nwell s -11713 96053 -10561 96188 4 VDD
port 41 nsew
rlabel nwell s -8260 96196 -7152 96451 4 VDD
port 41 nsew
rlabel nwell s -11713 96188 -10605 96443 4 VDD
port 41 nsew
rlabel nwell s -8260 96451 -7137 96681 4 VDD
port 41 nsew
rlabel nwell s -11713 96443 -10590 96673 4 VDD
port 41 nsew
rlabel nwell s -8267 96681 -7137 96899 4 VDD
port 41 nsew
rlabel nwell s -11720 96673 -10590 96891 4 VDD
port 41 nsew
rlabel nwell s -8672 96899 -7137 96973 4 VDD
port 41 nsew
rlabel nwell s -12125 96891 -10590 96965 4 VDD
port 41 nsew
rlabel nwell s -8672 96973 -7331 97060 4 VDD
port 41 nsew
rlabel nwell s -12125 96965 -10784 97052 4 VDD
port 41 nsew
rlabel nwell s -8672 97060 -7338 97746 4 VDD
port 41 nsew
rlabel nwell s -12125 97052 -10791 97738 4 VDD
port 41 nsew
rlabel nwell s -7712 97746 -7338 97778 4 VDD
port 41 nsew
rlabel nwell s -11165 97738 -10791 97770 4 VDD
port 41 nsew
rlabel nwell s -8430 98891 -7557 100368 4 VDD
port 41 nsew
rlabel nwell s -11945 99112 -11002 99138 4 VDD
port 41 nsew
rlabel nwell s -11945 99138 -10592 99634 4 VDD
port 41 nsew
rlabel nwell s -11751 99634 -10592 99721 4 VDD
port 41 nsew
rlabel nwell s -11744 99721 -10592 99856 4 VDD
port 41 nsew
rlabel nwell s -11744 99856 -10636 100111 4 VDD
port 41 nsew
rlabel nwell s -11744 100111 -10621 100341 4 VDD
port 41 nsew
rlabel nwell s -11751 100341 -10621 100559 4 VDD
port 41 nsew
rlabel nwell s -12156 100559 -10621 100633 4 VDD
port 41 nsew
rlabel nwell s -12156 100633 -10815 100720 4 VDD
port 41 nsew
rlabel nwell s -12156 100720 -10822 101406 4 VDD
port 41 nsew
rlabel nwell s -11196 101406 -10822 101438 4 VDD
port 41 nsew
rlabel nwell s -8444 104605 -7501 104631 4 VDD
port 41 nsew
rlabel nwell s -11897 104597 -10954 104623 4 VDD
port 41 nsew
rlabel nwell s -8444 104631 -7091 105127 4 VDD
port 41 nsew
rlabel nwell s -11897 104623 -10544 105119 4 VDD
port 41 nsew
rlabel nwell s -8250 105127 -7091 105214 4 VDD
port 41 nsew
rlabel nwell s -11703 105119 -10544 105206 4 VDD
port 41 nsew
rlabel nwell s -8243 105214 -7091 105349 4 VDD
port 41 nsew
rlabel nwell s -11696 105206 -10544 105341 4 VDD
port 41 nsew
rlabel nwell s -8243 105349 -7135 105604 4 VDD
port 41 nsew
rlabel nwell s -11696 105341 -10588 105596 4 VDD
port 41 nsew
rlabel nwell s -8243 105604 -7120 105834 4 VDD
port 41 nsew
rlabel nwell s -11696 105596 -10573 105826 4 VDD
port 41 nsew
rlabel nwell s -8250 105834 -7120 106052 4 VDD
port 41 nsew
rlabel nwell s -11703 105826 -10573 106044 4 VDD
port 41 nsew
rlabel nwell s -8655 106052 -7120 106126 4 VDD
port 41 nsew
rlabel nwell s -12108 106044 -10573 106118 4 VDD
port 41 nsew
rlabel nwell s -8655 106126 -7314 106213 4 VDD
port 41 nsew
rlabel nwell s -12108 106118 -10767 106205 4 VDD
port 41 nsew
rlabel nwell s -8655 106213 -7321 106899 4 VDD
port 41 nsew
rlabel nwell s -12108 106205 -10774 106891 4 VDD
port 41 nsew
rlabel nwell s -7695 106899 -7321 106931 4 VDD
port 41 nsew
rlabel nwell s -11148 106891 -10774 106923 4 VDD
port 41 nsew
rlabel nwell s -8413 108044 -7540 109521 4 VDD
port 41 nsew
rlabel nwell s -11928 108265 -10985 108291 4 VDD
port 41 nsew
rlabel nwell s -11928 108291 -10575 108787 4 VDD
port 41 nsew
rlabel nwell s -11734 108787 -10575 108874 4 VDD
port 41 nsew
rlabel nwell s -11727 108874 -10575 109009 4 VDD
port 41 nsew
rlabel nwell s -11727 109009 -10619 109264 4 VDD
port 41 nsew
rlabel nwell s -11727 109264 -10604 109494 4 VDD
port 41 nsew
rlabel nwell s -11734 109494 -10604 109712 4 VDD
port 41 nsew
rlabel nwell s -12139 109712 -10604 109786 4 VDD
port 41 nsew
rlabel nwell s -12139 109786 -10798 109873 4 VDD
port 41 nsew
rlabel nwell s -12139 109873 -10805 110559 4 VDD
port 41 nsew
rlabel nwell s -11179 110559 -10805 110591 4 VDD
port 41 nsew
rlabel nwell s -8406 113969 -7463 113995 4 VDD
port 41 nsew
rlabel nwell s -11859 113961 -10916 113987 4 VDD
port 41 nsew
rlabel nwell s -8406 113995 -7053 114491 4 VDD
port 41 nsew
rlabel nwell s -11859 113987 -10506 114483 4 VDD
port 41 nsew
rlabel nwell s -8212 114491 -7053 114578 4 VDD
port 41 nsew
rlabel nwell s -11665 114483 -10506 114570 4 VDD
port 41 nsew
rlabel nwell s -8205 114578 -7053 114713 4 VDD
port 41 nsew
rlabel nwell s -11658 114570 -10506 114705 4 VDD
port 41 nsew
rlabel nwell s -8205 114713 -7097 114968 4 VDD
port 41 nsew
rlabel nwell s -11658 114705 -10550 114960 4 VDD
port 41 nsew
rlabel nwell s -8205 114968 -7082 115198 4 VDD
port 41 nsew
rlabel nwell s -11658 114960 -10535 115190 4 VDD
port 41 nsew
rlabel nwell s -8212 115198 -7082 115416 4 VDD
port 41 nsew
rlabel nwell s -11665 115190 -10535 115408 4 VDD
port 41 nsew
rlabel nwell s -8617 115416 -7082 115490 4 VDD
port 41 nsew
rlabel nwell s -12070 115408 -10535 115482 4 VDD
port 41 nsew
rlabel nwell s -8617 115490 -7276 115577 4 VDD
port 41 nsew
rlabel nwell s -12070 115482 -10729 115569 4 VDD
port 41 nsew
rlabel nwell s -8617 115577 -7283 116263 4 VDD
port 41 nsew
rlabel nwell s -12070 115569 -10736 116255 4 VDD
port 41 nsew
rlabel nwell s -7657 116263 -7283 116295 4 VDD
port 41 nsew
rlabel nwell s -11110 116255 -10736 116287 4 VDD
port 41 nsew
rlabel nwell s -8375 117408 -7502 118885 4 VDD
port 41 nsew
rlabel nwell s -11890 117629 -10947 117655 4 VDD
port 41 nsew
rlabel nwell s -11890 117655 -10537 118151 4 VDD
port 41 nsew
rlabel nwell s -11696 118151 -10537 118238 4 VDD
port 41 nsew
rlabel nwell s -11689 118238 -10537 118373 4 VDD
port 41 nsew
rlabel nwell s -11689 118373 -10581 118628 4 VDD
port 41 nsew
rlabel nwell s -11689 118628 -10566 118858 4 VDD
port 41 nsew
rlabel nwell s -11696 118858 -10566 119076 4 VDD
port 41 nsew
rlabel nwell s -12101 119076 -10566 119150 4 VDD
port 41 nsew
rlabel nwell s -12101 119150 -10760 119237 4 VDD
port 41 nsew
rlabel nwell s -12101 119237 -10767 119923 4 VDD
port 41 nsew
rlabel nwell s -11141 119923 -10767 119955 4 VDD
port 41 nsew
rlabel metal4 s 16812 11245 17392 11509 6 VSS
port 42 nsew
rlabel metal4 s 16812 11509 18030 13083 6 VSS
port 42 nsew
rlabel metal4 s 197 13083 18030 13187 6 VSS
port 42 nsew
rlabel metal4 s 16812 13187 18030 15695 6 VSS
port 42 nsew
rlabel metal4 s 197 15695 18030 15799 6 VSS
port 42 nsew
rlabel metal4 s 16812 15799 18030 16176 6 VSS
port 42 nsew
rlabel metal4 s 16812 16176 92620 16280 6 VSS
port 42 nsew
rlabel metal4 s 16812 16280 18030 18307 6 VSS
port 42 nsew
rlabel metal4 s 197 18307 18030 18411 6 VSS
port 42 nsew
rlabel metal4 s 16812 18411 18030 20919 6 VSS
port 42 nsew
rlabel metal4 s 197 20919 18030 21023 6 VSS
port 42 nsew
rlabel metal4 s 16812 21023 18030 21788 6 VSS
port 42 nsew
rlabel metal4 s 16812 21788 92620 21892 6 VSS
port 42 nsew
rlabel metal4 s 16812 21892 18030 23531 6 VSS
port 42 nsew
rlabel metal4 s 197 23531 18030 23635 6 VSS
port 42 nsew
rlabel metal4 s 16812 23635 18030 26143 6 VSS
port 42 nsew
rlabel metal4 s 197 26143 18030 26247 6 VSS
port 42 nsew
rlabel metal4 s 16812 26247 18030 27400 6 VSS
port 42 nsew
rlabel metal4 s 16812 27400 92620 27504 6 VSS
port 42 nsew
rlabel metal4 s 16812 27504 18030 28755 6 VSS
port 42 nsew
rlabel metal4 s 197 28755 18030 28859 6 VSS
port 42 nsew
rlabel metal4 s 17174 28859 18030 33012 6 VSS
port 42 nsew
rlabel metal4 s 17174 33012 92620 33116 6 VSS
port 42 nsew
rlabel metal4 s 17174 33116 18030 38624 6 VSS
port 42 nsew
rlabel metal4 s 17174 38624 92620 38728 6 VSS
port 42 nsew
rlabel metal4 s 17174 38728 18030 44236 6 VSS
port 42 nsew
rlabel metal4 s 17174 44236 92620 44340 6 VSS
port 42 nsew
rlabel metal4 s 17174 44340 18030 49848 6 VSS
port 42 nsew
rlabel metal4 s 17174 49848 92620 49952 6 VSS
port 42 nsew
rlabel metal4 s 17174 49952 18030 55460 6 VSS
port 42 nsew
rlabel metal4 s 17174 55460 92620 55564 6 VSS
port 42 nsew
rlabel metal4 s 17174 55564 18030 61072 6 VSS
port 42 nsew
rlabel metal4 s 17174 61072 92620 61176 6 VSS
port 42 nsew
rlabel metal4 s 17174 61176 18030 66684 6 VSS
port 42 nsew
rlabel metal4 s 17174 66684 92620 66788 6 VSS
port 42 nsew
rlabel metal4 s 17174 66788 18030 72296 6 VSS
port 42 nsew
rlabel metal4 s 17174 72296 92620 72400 6 VSS
port 42 nsew
rlabel metal4 s 17174 72400 18030 77908 6 VSS
port 42 nsew
rlabel metal4 s 17174 77908 92620 78012 6 VSS
port 42 nsew
rlabel metal4 s 17174 78012 18030 83520 6 VSS
port 42 nsew
rlabel metal4 s 17174 83520 92620 83624 6 VSS
port 42 nsew
rlabel metal4 s 17174 83624 18030 89132 6 VSS
port 42 nsew
rlabel metal4 s 17174 89132 92620 89236 6 VSS
port 42 nsew
rlabel metal4 s 17174 89236 18030 89308 6 VSS
port 42 nsew
rlabel metal3 s 87420 10908 92500 16280 6 VSS
port 42 nsew
rlabel metal3 s 82100 10908 87180 16280 6 VSS
port 42 nsew
rlabel metal3 s 76780 10908 81860 16280 6 VSS
port 42 nsew
rlabel metal3 s 71460 10908 76540 16280 6 VSS
port 42 nsew
rlabel metal3 s 66140 10908 71220 16280 6 VSS
port 42 nsew
rlabel metal3 s 60820 10908 65900 16280 6 VSS
port 42 nsew
rlabel metal3 s 55500 10908 60580 16280 6 VSS
port 42 nsew
rlabel metal3 s 50180 10908 55260 16280 6 VSS
port 42 nsew
rlabel metal3 s 44860 10908 49940 16280 6 VSS
port 42 nsew
rlabel metal3 s 39540 10908 44620 16280 6 VSS
port 42 nsew
rlabel metal3 s 34220 10908 39300 16280 6 VSS
port 42 nsew
rlabel metal3 s 28900 10908 33980 16280 6 VSS
port 42 nsew
rlabel metal3 s 23580 10908 28660 16280 6 VSS
port 42 nsew
rlabel metal3 s 18260 10908 23340 16280 6 VSS
port 42 nsew
rlabel metal3 s 87420 16520 92500 21892 6 VSS
port 42 nsew
rlabel metal3 s 82100 16520 87180 21892 6 VSS
port 42 nsew
rlabel metal3 s 76780 16520 81860 21892 6 VSS
port 42 nsew
rlabel metal3 s 71460 16520 76540 21892 6 VSS
port 42 nsew
rlabel metal3 s 66140 16520 71220 21892 6 VSS
port 42 nsew
rlabel metal3 s 60820 16520 65900 21892 6 VSS
port 42 nsew
rlabel metal3 s 55500 16520 60580 21892 6 VSS
port 42 nsew
rlabel metal3 s 50180 16520 55260 21892 6 VSS
port 42 nsew
rlabel metal3 s 44860 16520 49940 21892 6 VSS
port 42 nsew
rlabel metal3 s 39540 16520 44620 21892 6 VSS
port 42 nsew
rlabel metal3 s 34220 16520 39300 21892 6 VSS
port 42 nsew
rlabel metal3 s 28900 16520 33980 21892 6 VSS
port 42 nsew
rlabel metal3 s 23580 16520 28660 21892 6 VSS
port 42 nsew
rlabel metal3 s 18260 16520 23340 21892 6 VSS
port 42 nsew
rlabel metal3 s 16949 11350 17282 16839 6 VSS
port 42 nsew
rlabel metal3 s 14237 10815 16317 13187 6 VSS
port 42 nsew
rlabel metal3 s 11917 10815 13997 13187 6 VSS
port 42 nsew
rlabel metal3 s 9597 10815 11677 13187 6 VSS
port 42 nsew
rlabel metal3 s 7277 10815 9357 13187 6 VSS
port 42 nsew
rlabel metal3 s 4957 10815 7037 13187 6 VSS
port 42 nsew
rlabel metal3 s 2637 10815 4717 13187 6 VSS
port 42 nsew
rlabel metal3 s 317 10815 2397 13187 6 VSS
port 42 nsew
rlabel metal3 s 14237 13427 16317 15799 6 VSS
port 42 nsew
rlabel metal3 s 11917 13427 13997 15799 6 VSS
port 42 nsew
rlabel metal3 s 9597 13427 11677 15799 6 VSS
port 42 nsew
rlabel metal3 s 7277 13427 9357 15799 6 VSS
port 42 nsew
rlabel metal3 s 4957 13427 7037 15799 6 VSS
port 42 nsew
rlabel metal3 s 2637 13427 4717 15799 6 VSS
port 42 nsew
rlabel metal3 s 317 13427 2397 15799 6 VSS
port 42 nsew
rlabel metal3 s 14237 16039 16317 18411 6 VSS
port 42 nsew
rlabel metal3 s 11917 16039 13997 18411 6 VSS
port 42 nsew
rlabel metal3 s 9597 16039 11677 18411 6 VSS
port 42 nsew
rlabel metal3 s 7277 16039 9357 18411 6 VSS
port 42 nsew
rlabel metal3 s 4957 16039 7037 18411 6 VSS
port 42 nsew
rlabel metal3 s 2637 16039 4717 18411 6 VSS
port 42 nsew
rlabel metal3 s 317 16039 2397 18411 6 VSS
port 42 nsew
rlabel metal3 s 14237 18651 16317 21023 6 VSS
port 42 nsew
rlabel metal3 s 11917 18651 13997 21023 6 VSS
port 42 nsew
rlabel metal3 s 9597 18651 11677 21023 6 VSS
port 42 nsew
rlabel metal3 s 7277 18651 9357 21023 6 VSS
port 42 nsew
rlabel metal3 s 4957 18651 7037 21023 6 VSS
port 42 nsew
rlabel metal3 s 2637 18651 4717 21023 6 VSS
port 42 nsew
rlabel metal3 s 317 18651 2397 21023 6 VSS
port 42 nsew
rlabel metal3 s 87420 22132 92500 27504 6 VSS
port 42 nsew
rlabel metal3 s 82100 22132 87180 27504 6 VSS
port 42 nsew
rlabel metal3 s 76780 22132 81860 27504 6 VSS
port 42 nsew
rlabel metal3 s 71460 22132 76540 27504 6 VSS
port 42 nsew
rlabel metal3 s 66140 22132 71220 27504 6 VSS
port 42 nsew
rlabel metal3 s 60820 22132 65900 27504 6 VSS
port 42 nsew
rlabel metal3 s 55500 22132 60580 27504 6 VSS
port 42 nsew
rlabel metal3 s 50180 22132 55260 27504 6 VSS
port 42 nsew
rlabel metal3 s 44860 22132 49940 27504 6 VSS
port 42 nsew
rlabel metal3 s 39540 22132 44620 27504 6 VSS
port 42 nsew
rlabel metal3 s 34220 22132 39300 27504 6 VSS
port 42 nsew
rlabel metal3 s 28900 22132 33980 27504 6 VSS
port 42 nsew
rlabel metal3 s 23580 22132 28660 27504 6 VSS
port 42 nsew
rlabel metal3 s 18260 22132 23340 27504 6 VSS
port 42 nsew
rlabel metal3 s 14237 21263 16317 23635 6 VSS
port 42 nsew
rlabel metal3 s 11917 21263 13997 23635 6 VSS
port 42 nsew
rlabel metal3 s 9597 21263 11677 23635 6 VSS
port 42 nsew
rlabel metal3 s 7277 21263 9357 23635 6 VSS
port 42 nsew
rlabel metal3 s 4957 21263 7037 23635 6 VSS
port 42 nsew
rlabel metal3 s 2637 21263 4717 23635 6 VSS
port 42 nsew
rlabel metal3 s 317 21263 2397 23635 6 VSS
port 42 nsew
rlabel metal3 s 14237 23875 16317 26247 6 VSS
port 42 nsew
rlabel metal3 s 11917 23875 13997 26247 6 VSS
port 42 nsew
rlabel metal3 s 9597 23875 11677 26247 6 VSS
port 42 nsew
rlabel metal3 s 7277 23875 9357 26247 6 VSS
port 42 nsew
rlabel metal3 s 4957 23875 7037 26247 6 VSS
port 42 nsew
rlabel metal3 s 2637 23875 4717 26247 6 VSS
port 42 nsew
rlabel metal3 s 317 23875 2397 26247 6 VSS
port 42 nsew
rlabel metal3 s 87420 27744 92500 33116 6 VSS
port 42 nsew
rlabel metal3 s 82100 27744 87180 33116 6 VSS
port 42 nsew
rlabel metal3 s 76780 27744 81860 33116 6 VSS
port 42 nsew
rlabel metal3 s 71460 27744 76540 33116 6 VSS
port 42 nsew
rlabel metal3 s 66140 27744 71220 33116 6 VSS
port 42 nsew
rlabel metal3 s 60820 27744 65900 33116 6 VSS
port 42 nsew
rlabel metal3 s 55500 27744 60580 33116 6 VSS
port 42 nsew
rlabel metal3 s 50180 27744 55260 33116 6 VSS
port 42 nsew
rlabel metal3 s 44860 27744 49940 33116 6 VSS
port 42 nsew
rlabel metal3 s 39540 27744 44620 33116 6 VSS
port 42 nsew
rlabel metal3 s 34220 27744 39300 33116 6 VSS
port 42 nsew
rlabel metal3 s 28900 27744 33980 33116 6 VSS
port 42 nsew
rlabel metal3 s 23580 27744 28660 33116 6 VSS
port 42 nsew
rlabel metal3 s 18260 27744 23340 33116 6 VSS
port 42 nsew
rlabel metal3 s 14237 26487 16317 28859 6 VSS
port 42 nsew
rlabel metal3 s 11917 26487 13997 28859 6 VSS
port 42 nsew
rlabel metal3 s 9597 26487 11677 28859 6 VSS
port 42 nsew
rlabel metal3 s 7277 26487 9357 28859 6 VSS
port 42 nsew
rlabel metal3 s 4957 26487 7037 28859 6 VSS
port 42 nsew
rlabel metal3 s 2637 26487 4717 28859 6 VSS
port 42 nsew
rlabel metal3 s 317 26487 2397 28859 6 VSS
port 42 nsew
rlabel metal3 s 87420 33356 92500 38728 6 VSS
port 42 nsew
rlabel metal3 s 82100 33356 87180 38728 6 VSS
port 42 nsew
rlabel metal3 s 76780 33356 81860 38728 6 VSS
port 42 nsew
rlabel metal3 s 71460 33356 76540 38728 6 VSS
port 42 nsew
rlabel metal3 s 66140 33356 71220 38728 6 VSS
port 42 nsew
rlabel metal3 s 60820 33356 65900 38728 6 VSS
port 42 nsew
rlabel metal3 s 55500 33356 60580 38728 6 VSS
port 42 nsew
rlabel metal3 s 50180 33356 55260 38728 6 VSS
port 42 nsew
rlabel metal3 s 44860 33356 49940 38728 6 VSS
port 42 nsew
rlabel metal3 s 39540 33356 44620 38728 6 VSS
port 42 nsew
rlabel metal3 s 34220 33356 39300 38728 6 VSS
port 42 nsew
rlabel metal3 s 28900 33356 33980 38728 6 VSS
port 42 nsew
rlabel metal3 s 23580 33356 28660 38728 6 VSS
port 42 nsew
rlabel metal3 s 18260 33356 23340 38728 6 VSS
port 42 nsew
rlabel metal3 s 87420 38968 92500 44340 6 VSS
port 42 nsew
rlabel metal3 s 82100 38968 87180 44340 6 VSS
port 42 nsew
rlabel metal3 s 76780 38968 81860 44340 6 VSS
port 42 nsew
rlabel metal3 s 71460 38968 76540 44340 6 VSS
port 42 nsew
rlabel metal3 s 66140 38968 71220 44340 6 VSS
port 42 nsew
rlabel metal3 s 60820 38968 65900 44340 6 VSS
port 42 nsew
rlabel metal3 s 55500 38968 60580 44340 6 VSS
port 42 nsew
rlabel metal3 s 50180 38968 55260 44340 6 VSS
port 42 nsew
rlabel metal3 s 44860 38968 49940 44340 6 VSS
port 42 nsew
rlabel metal3 s 39540 38968 44620 44340 6 VSS
port 42 nsew
rlabel metal3 s 34220 38968 39300 44340 6 VSS
port 42 nsew
rlabel metal3 s 28900 38968 33980 44340 6 VSS
port 42 nsew
rlabel metal3 s 23580 38968 28660 44340 6 VSS
port 42 nsew
rlabel metal3 s 18260 38968 23340 44340 6 VSS
port 42 nsew
rlabel metal3 s 87420 44580 92500 49952 6 VSS
port 42 nsew
rlabel metal3 s 82100 44580 87180 49952 6 VSS
port 42 nsew
rlabel metal3 s 76780 44580 81860 49952 6 VSS
port 42 nsew
rlabel metal3 s 71460 44580 76540 49952 6 VSS
port 42 nsew
rlabel metal3 s 66140 44580 71220 49952 6 VSS
port 42 nsew
rlabel metal3 s 60820 44580 65900 49952 6 VSS
port 42 nsew
rlabel metal3 s 55500 44580 60580 49952 6 VSS
port 42 nsew
rlabel metal3 s 50180 44580 55260 49952 6 VSS
port 42 nsew
rlabel metal3 s 44860 44580 49940 49952 6 VSS
port 42 nsew
rlabel metal3 s 39540 44580 44620 49952 6 VSS
port 42 nsew
rlabel metal3 s 34220 44580 39300 49952 6 VSS
port 42 nsew
rlabel metal3 s 28900 44580 33980 49952 6 VSS
port 42 nsew
rlabel metal3 s 23580 44580 28660 49952 6 VSS
port 42 nsew
rlabel metal3 s 18260 44580 23340 49952 6 VSS
port 42 nsew
rlabel metal3 s 87420 50192 92500 55564 6 VSS
port 42 nsew
rlabel metal3 s 82100 50192 87180 55564 6 VSS
port 42 nsew
rlabel metal3 s 76780 50192 81860 55564 6 VSS
port 42 nsew
rlabel metal3 s 71460 50192 76540 55564 6 VSS
port 42 nsew
rlabel metal3 s 66140 50192 71220 55564 6 VSS
port 42 nsew
rlabel metal3 s 60820 50192 65900 55564 6 VSS
port 42 nsew
rlabel metal3 s 55500 50192 60580 55564 6 VSS
port 42 nsew
rlabel metal3 s 50180 50192 55260 55564 6 VSS
port 42 nsew
rlabel metal3 s 44860 50192 49940 55564 6 VSS
port 42 nsew
rlabel metal3 s 39540 50192 44620 55564 6 VSS
port 42 nsew
rlabel metal3 s 34220 50192 39300 55564 6 VSS
port 42 nsew
rlabel metal3 s 28900 50192 33980 55564 6 VSS
port 42 nsew
rlabel metal3 s 23580 50192 28660 55564 6 VSS
port 42 nsew
rlabel metal3 s 18260 50192 23340 55564 6 VSS
port 42 nsew
rlabel metal3 s 87420 55804 92500 61176 6 VSS
port 42 nsew
rlabel metal3 s 82100 55804 87180 61176 6 VSS
port 42 nsew
rlabel metal3 s 76780 55804 81860 61176 6 VSS
port 42 nsew
rlabel metal3 s 71460 55804 76540 61176 6 VSS
port 42 nsew
rlabel metal3 s 66140 55804 71220 61176 6 VSS
port 42 nsew
rlabel metal3 s 60820 55804 65900 61176 6 VSS
port 42 nsew
rlabel metal3 s 55500 55804 60580 61176 6 VSS
port 42 nsew
rlabel metal3 s 50180 55804 55260 61176 6 VSS
port 42 nsew
rlabel metal3 s 44860 55804 49940 61176 6 VSS
port 42 nsew
rlabel metal3 s 39540 55804 44620 61176 6 VSS
port 42 nsew
rlabel metal3 s 34220 55804 39300 61176 6 VSS
port 42 nsew
rlabel metal3 s 28900 55804 33980 61176 6 VSS
port 42 nsew
rlabel metal3 s 23580 55804 28660 61176 6 VSS
port 42 nsew
rlabel metal3 s 18260 55804 23340 61176 6 VSS
port 42 nsew
rlabel metal3 s 87420 61416 92500 66788 6 VSS
port 42 nsew
rlabel metal3 s 82100 61416 87180 66788 6 VSS
port 42 nsew
rlabel metal3 s 76780 61416 81860 66788 6 VSS
port 42 nsew
rlabel metal3 s 71460 61416 76540 66788 6 VSS
port 42 nsew
rlabel metal3 s 66140 61416 71220 66788 6 VSS
port 42 nsew
rlabel metal3 s 60820 61416 65900 66788 6 VSS
port 42 nsew
rlabel metal3 s 55500 61416 60580 66788 6 VSS
port 42 nsew
rlabel metal3 s 50180 61416 55260 66788 6 VSS
port 42 nsew
rlabel metal3 s 44860 61416 49940 66788 6 VSS
port 42 nsew
rlabel metal3 s 39540 61416 44620 66788 6 VSS
port 42 nsew
rlabel metal3 s 34220 61416 39300 66788 6 VSS
port 42 nsew
rlabel metal3 s 28900 61416 33980 66788 6 VSS
port 42 nsew
rlabel metal3 s 23580 61416 28660 66788 6 VSS
port 42 nsew
rlabel metal3 s 18260 61416 23340 66788 6 VSS
port 42 nsew
rlabel metal3 s 87420 67028 92500 72400 6 VSS
port 42 nsew
rlabel metal3 s 82100 67028 87180 72400 6 VSS
port 42 nsew
rlabel metal3 s 76780 67028 81860 72400 6 VSS
port 42 nsew
rlabel metal3 s 71460 67028 76540 72400 6 VSS
port 42 nsew
rlabel metal3 s 66140 67028 71220 72400 6 VSS
port 42 nsew
rlabel metal3 s 60820 67028 65900 72400 6 VSS
port 42 nsew
rlabel metal3 s 55500 67028 60580 72400 6 VSS
port 42 nsew
rlabel metal3 s 50180 67028 55260 72400 6 VSS
port 42 nsew
rlabel metal3 s 44860 67028 49940 72400 6 VSS
port 42 nsew
rlabel metal3 s 39540 67028 44620 72400 6 VSS
port 42 nsew
rlabel metal3 s 34220 67028 39300 72400 6 VSS
port 42 nsew
rlabel metal3 s 28900 67028 33980 72400 6 VSS
port 42 nsew
rlabel metal3 s 23580 67028 28660 72400 6 VSS
port 42 nsew
rlabel metal3 s 18260 67028 23340 72400 6 VSS
port 42 nsew
rlabel metal3 s 87420 72640 92500 78012 6 VSS
port 42 nsew
rlabel metal3 s 82100 72640 87180 78012 6 VSS
port 42 nsew
rlabel metal3 s 76780 72640 81860 78012 6 VSS
port 42 nsew
rlabel metal3 s 71460 72640 76540 78012 6 VSS
port 42 nsew
rlabel metal3 s 66140 72640 71220 78012 6 VSS
port 42 nsew
rlabel metal3 s 60820 72640 65900 78012 6 VSS
port 42 nsew
rlabel metal3 s 55500 72640 60580 78012 6 VSS
port 42 nsew
rlabel metal3 s 50180 72640 55260 78012 6 VSS
port 42 nsew
rlabel metal3 s 44860 72640 49940 78012 6 VSS
port 42 nsew
rlabel metal3 s 39540 72640 44620 78012 6 VSS
port 42 nsew
rlabel metal3 s 34220 72640 39300 78012 6 VSS
port 42 nsew
rlabel metal3 s 28900 72640 33980 78012 6 VSS
port 42 nsew
rlabel metal3 s 23580 72640 28660 78012 6 VSS
port 42 nsew
rlabel metal3 s 18260 72640 23340 78012 6 VSS
port 42 nsew
rlabel metal3 s 87420 78252 92500 83624 6 VSS
port 42 nsew
rlabel metal3 s 82100 78252 87180 83624 6 VSS
port 42 nsew
rlabel metal3 s 76780 78252 81860 83624 6 VSS
port 42 nsew
rlabel metal3 s 71460 78252 76540 83624 6 VSS
port 42 nsew
rlabel metal3 s 66140 78252 71220 83624 6 VSS
port 42 nsew
rlabel metal3 s 60820 78252 65900 83624 6 VSS
port 42 nsew
rlabel metal3 s 55500 78252 60580 83624 6 VSS
port 42 nsew
rlabel metal3 s 50180 78252 55260 83624 6 VSS
port 42 nsew
rlabel metal3 s 44860 78252 49940 83624 6 VSS
port 42 nsew
rlabel metal3 s 39540 78252 44620 83624 6 VSS
port 42 nsew
rlabel metal3 s 34220 78252 39300 83624 6 VSS
port 42 nsew
rlabel metal3 s 28900 78252 33980 83624 6 VSS
port 42 nsew
rlabel metal3 s 23580 78252 28660 83624 6 VSS
port 42 nsew
rlabel metal3 s 18260 78252 23340 83624 6 VSS
port 42 nsew
rlabel metal3 s 87420 83864 92500 89236 6 VSS
port 42 nsew
rlabel metal3 s 82100 83864 87180 89236 6 VSS
port 42 nsew
rlabel metal3 s 76780 83864 81860 89236 6 VSS
port 42 nsew
rlabel metal3 s 71460 83864 76540 89236 6 VSS
port 42 nsew
rlabel metal3 s 66140 83864 71220 89236 6 VSS
port 42 nsew
rlabel metal3 s 60820 83864 65900 89236 6 VSS
port 42 nsew
rlabel metal3 s 55500 83864 60580 89236 6 VSS
port 42 nsew
rlabel metal3 s 50180 83864 55260 89236 6 VSS
port 42 nsew
rlabel metal3 s 44860 83864 49940 89236 6 VSS
port 42 nsew
rlabel metal3 s 39540 83864 44620 89236 6 VSS
port 42 nsew
rlabel metal3 s 34220 83864 39300 89236 6 VSS
port 42 nsew
rlabel metal3 s 28900 83864 33980 89236 6 VSS
port 42 nsew
rlabel metal3 s 23580 83864 28660 89236 6 VSS
port 42 nsew
rlabel metal3 s 18260 83864 23340 89236 6 VSS
port 42 nsew
rlabel metal2 s 16949 11350 17282 16839 6 VSS
port 42 nsew
rlabel metal1 s 90119 -54278 92731 -7667 8 VSS
port 42 nsew
rlabel metal1 s 89990 -7667 92959 -4698 8 VSS
port 42 nsew
rlabel metal1 s 61261 -5041 61482 -4779 8 VSS
port 42 nsew
rlabel metal1 s 63629 -3733 63675 -3633 8 VSS
port 42 nsew
rlabel metal1 s 63433 -3733 63479 -3633 8 VSS
port 42 nsew
rlabel metal1 s 63237 -3733 63283 -3633 8 VSS
port 42 nsew
rlabel metal1 s 62387 -3431 62910 -3425 8 VSS
port 42 nsew
rlabel metal1 s 62111 -3425 62910 -3360 8 VSS
port 42 nsew
rlabel metal1 s 63629 -3318 63675 -3218 8 VSS
port 42 nsew
rlabel metal1 s 63433 -3318 63479 -3218 8 VSS
port 42 nsew
rlabel metal1 s 63237 -3318 63283 -3218 8 VSS
port 42 nsew
rlabel metal1 s 62779 -3318 62825 -3218 8 VSS
port 42 nsew
rlabel metal1 s 62583 -3318 62629 -3218 8 VSS
port 42 nsew
rlabel metal1 s 62387 -3318 62433 -3218 8 VSS
port 42 nsew
rlabel metal1 s 62111 -3360 62176 -3293 8 VSS
port 42 nsew
rlabel metal1 s 61353 -4779 61418 -3293 8 VSS
port 42 nsew
rlabel metal1 s 46778 -5304 47412 -4670 8 VSS
port 42 nsew
rlabel metal1 s 58059 -4132 58105 -3732 8 VSS
port 42 nsew
rlabel metal1 s 57941 -4132 57987 -3732 8 VSS
port 42 nsew
rlabel metal1 s 57823 -4132 57869 -3732 8 VSS
port 42 nsew
rlabel metal1 s 57705 -4132 57751 -3732 8 VSS
port 42 nsew
rlabel metal1 s 57587 -4132 57633 -3732 8 VSS
port 42 nsew
rlabel metal1 s 57469 -4132 57515 -3732 8 VSS
port 42 nsew
rlabel metal1 s 57351 -4132 57397 -3732 8 VSS
port 42 nsew
rlabel metal1 s 57233 -4132 57279 -3732 8 VSS
port 42 nsew
rlabel metal1 s 57115 -4132 57161 -3732 8 VSS
port 42 nsew
rlabel metal1 s 56997 -4132 57043 -3732 8 VSS
port 42 nsew
rlabel metal1 s 56879 -4132 56925 -3732 8 VSS
port 42 nsew
rlabel metal1 s 56761 -4132 56807 -3732 8 VSS
port 42 nsew
rlabel metal1 s 56643 -4132 56689 -3732 8 VSS
port 42 nsew
rlabel metal1 s 56525 -4132 56571 -3732 8 VSS
port 42 nsew
rlabel metal1 s 56407 -4132 56453 -3732 8 VSS
port 42 nsew
rlabel metal1 s 56289 -4132 56335 -3732 8 VSS
port 42 nsew
rlabel metal1 s 56171 -4132 56217 -3732 8 VSS
port 42 nsew
rlabel metal1 s 56053 -4132 56099 -3732 8 VSS
port 42 nsew
rlabel metal1 s 55935 -4132 55981 -3732 8 VSS
port 42 nsew
rlabel metal1 s 55817 -4132 55863 -3732 8 VSS
port 42 nsew
rlabel metal1 s 55699 -4132 55745 -3732 8 VSS
port 42 nsew
rlabel metal1 s 55581 -4132 55627 -3732 8 VSS
port 42 nsew
rlabel metal1 s 55463 -4132 55509 -3732 8 VSS
port 42 nsew
rlabel metal1 s 55345 -4132 55391 -3732 8 VSS
port 42 nsew
rlabel metal1 s 55227 -4132 55273 -3732 8 VSS
port 42 nsew
rlabel metal1 s 55109 -4132 55155 -3732 8 VSS
port 42 nsew
rlabel metal1 s 54991 -4132 55037 -3732 8 VSS
port 42 nsew
rlabel metal1 s 54873 -4132 54919 -3732 8 VSS
port 42 nsew
rlabel metal1 s 54755 -4132 54801 -3732 8 VSS
port 42 nsew
rlabel metal1 s 54637 -4132 54683 -3732 8 VSS
port 42 nsew
rlabel metal1 s 54519 -4132 54565 -3732 8 VSS
port 42 nsew
rlabel metal1 s 54283 -4132 54329 -3732 8 VSS
port 42 nsew
rlabel metal1 s 54047 -4132 54093 -3732 8 VSS
port 42 nsew
rlabel metal1 s 53811 -4132 53857 -3732 8 VSS
port 42 nsew
rlabel metal1 s 53575 -4132 53621 -3732 8 VSS
port 42 nsew
rlabel metal1 s 53339 -4132 53385 -3732 8 VSS
port 42 nsew
rlabel metal1 s 53103 -4132 53149 -3732 8 VSS
port 42 nsew
rlabel metal1 s 52867 -4132 52913 -3732 8 VSS
port 42 nsew
rlabel metal1 s 52631 -4132 52677 -3732 8 VSS
port 42 nsew
rlabel metal1 s 52395 -4132 52441 -3732 8 VSS
port 42 nsew
rlabel metal1 s 52159 -4132 52205 -3732 8 VSS
port 42 nsew
rlabel metal1 s 51923 -4132 51969 -3732 8 VSS
port 42 nsew
rlabel metal1 s 51687 -4132 51733 -3732 8 VSS
port 42 nsew
rlabel metal1 s 51451 -4132 51497 -3732 8 VSS
port 42 nsew
rlabel metal1 s 51215 -4132 51261 -3732 8 VSS
port 42 nsew
rlabel metal1 s 50979 -4132 51025 -3732 8 VSS
port 42 nsew
rlabel metal1 s 61353 -3293 62176 -3228 8 VSS
port 42 nsew
rlabel metal1 s 46850 -4670 47412 -1960 8 VSS
port 42 nsew
rlabel metal1 s 14943 -1707 14989 -1307 8 VSS
port 42 nsew
rlabel metal1 s 14825 -1707 14871 -1307 8 VSS
port 42 nsew
rlabel metal1 s 14707 -1707 14753 -1307 8 VSS
port 42 nsew
rlabel metal1 s 14589 -1707 14635 -1307 8 VSS
port 42 nsew
rlabel metal1 s 14471 -1707 14517 -1307 8 VSS
port 42 nsew
rlabel metal1 s 14353 -1707 14399 -1307 8 VSS
port 42 nsew
rlabel metal1 s 14235 -1707 14281 -1307 8 VSS
port 42 nsew
rlabel metal1 s 14117 -1707 14163 -1307 8 VSS
port 42 nsew
rlabel metal1 s 13999 -1707 14045 -1307 8 VSS
port 42 nsew
rlabel metal1 s 13881 -1707 13927 -1307 8 VSS
port 42 nsew
rlabel metal1 s 13763 -1707 13809 -1307 8 VSS
port 42 nsew
rlabel metal1 s 13645 -1707 13691 -1307 8 VSS
port 42 nsew
rlabel metal1 s 13527 -1707 13573 -1307 8 VSS
port 42 nsew
rlabel metal1 s 13409 -1707 13455 -1307 8 VSS
port 42 nsew
rlabel metal1 s 13291 -1707 13337 -1307 8 VSS
port 42 nsew
rlabel metal1 s 13173 -1707 13219 -1307 8 VSS
port 42 nsew
rlabel metal1 s 13055 -1707 13101 -1307 8 VSS
port 42 nsew
rlabel metal1 s 12937 -1707 12983 -1307 8 VSS
port 42 nsew
rlabel metal1 s 12819 -1707 12865 -1307 8 VSS
port 42 nsew
rlabel metal1 s 12701 -1707 12747 -1307 8 VSS
port 42 nsew
rlabel metal1 s 12583 -1707 12629 -1307 8 VSS
port 42 nsew
rlabel metal1 s 12465 -1707 12511 -1307 8 VSS
port 42 nsew
rlabel metal1 s 12347 -1707 12393 -1307 8 VSS
port 42 nsew
rlabel metal1 s 12229 -1707 12275 -1307 8 VSS
port 42 nsew
rlabel metal1 s 12111 -1707 12157 -1307 8 VSS
port 42 nsew
rlabel metal1 s 11993 -1707 12039 -1307 8 VSS
port 42 nsew
rlabel metal1 s 11875 -1707 11921 -1307 8 VSS
port 42 nsew
rlabel metal1 s 11757 -1707 11803 -1307 8 VSS
port 42 nsew
rlabel metal1 s 11639 -1707 11685 -1307 8 VSS
port 42 nsew
rlabel metal1 s 11521 -1707 11567 -1307 8 VSS
port 42 nsew
rlabel metal1 s 11403 -1707 11449 -1307 8 VSS
port 42 nsew
rlabel metal1 s 11167 -1707 11213 -1307 8 VSS
port 42 nsew
rlabel metal1 s 10931 -1707 10977 -1307 8 VSS
port 42 nsew
rlabel metal1 s 10695 -1707 10741 -1307 8 VSS
port 42 nsew
rlabel metal1 s 10459 -1707 10505 -1307 8 VSS
port 42 nsew
rlabel metal1 s 10223 -1707 10269 -1307 8 VSS
port 42 nsew
rlabel metal1 s 9987 -1707 10033 -1307 8 VSS
port 42 nsew
rlabel metal1 s 9751 -1707 9797 -1307 8 VSS
port 42 nsew
rlabel metal1 s 9515 -1707 9561 -1307 8 VSS
port 42 nsew
rlabel metal1 s 9279 -1707 9325 -1307 8 VSS
port 42 nsew
rlabel metal1 s 9043 -1707 9089 -1307 8 VSS
port 42 nsew
rlabel metal1 s 8807 -1707 8853 -1307 8 VSS
port 42 nsew
rlabel metal1 s 8571 -1707 8617 -1307 8 VSS
port 42 nsew
rlabel metal1 s 8335 -1707 8381 -1307 8 VSS
port 42 nsew
rlabel metal1 s 8099 -1707 8145 -1307 8 VSS
port 42 nsew
rlabel metal1 s 7863 -1707 7909 -1307 8 VSS
port 42 nsew
rlabel metal1 s 5766 -1372 5812 -1272 8 VSS
port 42 nsew
rlabel metal1 s 5570 -1372 5616 -1272 8 VSS
port 42 nsew
rlabel metal1 s 5374 -1372 5420 -1272 8 VSS
port 42 nsew
rlabel metal1 s 58059 -1085 58105 -685 8 VSS
port 42 nsew
rlabel metal1 s 57941 -1085 57987 -685 8 VSS
port 42 nsew
rlabel metal1 s 57823 -1085 57869 -685 8 VSS
port 42 nsew
rlabel metal1 s 57705 -1085 57751 -685 8 VSS
port 42 nsew
rlabel metal1 s 57587 -1085 57633 -685 8 VSS
port 42 nsew
rlabel metal1 s 57469 -1085 57515 -685 8 VSS
port 42 nsew
rlabel metal1 s 57351 -1085 57397 -685 8 VSS
port 42 nsew
rlabel metal1 s 57233 -1085 57279 -685 8 VSS
port 42 nsew
rlabel metal1 s 57115 -1085 57161 -685 8 VSS
port 42 nsew
rlabel metal1 s 56997 -1085 57043 -685 8 VSS
port 42 nsew
rlabel metal1 s 56879 -1085 56925 -685 8 VSS
port 42 nsew
rlabel metal1 s 56761 -1085 56807 -685 8 VSS
port 42 nsew
rlabel metal1 s 56643 -1085 56689 -685 8 VSS
port 42 nsew
rlabel metal1 s 56525 -1085 56571 -685 8 VSS
port 42 nsew
rlabel metal1 s 56407 -1085 56453 -685 8 VSS
port 42 nsew
rlabel metal1 s 56289 -1085 56335 -685 8 VSS
port 42 nsew
rlabel metal1 s 56171 -1085 56217 -685 8 VSS
port 42 nsew
rlabel metal1 s 56053 -1085 56099 -685 8 VSS
port 42 nsew
rlabel metal1 s 55935 -1085 55981 -685 8 VSS
port 42 nsew
rlabel metal1 s 55817 -1085 55863 -685 8 VSS
port 42 nsew
rlabel metal1 s 55699 -1085 55745 -685 8 VSS
port 42 nsew
rlabel metal1 s 55581 -1085 55627 -685 8 VSS
port 42 nsew
rlabel metal1 s 55463 -1085 55509 -685 8 VSS
port 42 nsew
rlabel metal1 s 55345 -1085 55391 -685 8 VSS
port 42 nsew
rlabel metal1 s 55227 -1085 55273 -685 8 VSS
port 42 nsew
rlabel metal1 s 55109 -1085 55155 -685 8 VSS
port 42 nsew
rlabel metal1 s 54991 -1085 55037 -685 8 VSS
port 42 nsew
rlabel metal1 s 54873 -1085 54919 -685 8 VSS
port 42 nsew
rlabel metal1 s 54755 -1085 54801 -685 8 VSS
port 42 nsew
rlabel metal1 s 54637 -1085 54683 -685 8 VSS
port 42 nsew
rlabel metal1 s 54519 -1085 54565 -685 8 VSS
port 42 nsew
rlabel metal1 s 54283 -1085 54329 -685 8 VSS
port 42 nsew
rlabel metal1 s 54047 -1085 54093 -685 8 VSS
port 42 nsew
rlabel metal1 s 53811 -1085 53857 -685 8 VSS
port 42 nsew
rlabel metal1 s 53575 -1085 53621 -685 8 VSS
port 42 nsew
rlabel metal1 s 53339 -1085 53385 -685 8 VSS
port 42 nsew
rlabel metal1 s 53103 -1085 53149 -685 8 VSS
port 42 nsew
rlabel metal1 s 52867 -1085 52913 -685 8 VSS
port 42 nsew
rlabel metal1 s 52631 -1085 52677 -685 8 VSS
port 42 nsew
rlabel metal1 s 52395 -1085 52441 -685 8 VSS
port 42 nsew
rlabel metal1 s 52159 -1085 52205 -685 8 VSS
port 42 nsew
rlabel metal1 s 51923 -1085 51969 -685 8 VSS
port 42 nsew
rlabel metal1 s 51687 -1085 51733 -685 8 VSS
port 42 nsew
rlabel metal1 s 51451 -1085 51497 -685 8 VSS
port 42 nsew
rlabel metal1 s 51215 -1085 51261 -685 8 VSS
port 42 nsew
rlabel metal1 s 50979 -1085 51025 -685 8 VSS
port 42 nsew
rlabel metal1 s 3841 -1069 4601 -1066 8 VSS
port 42 nsew
rlabel metal1 s 3841 -1066 4999 -1011 8 VSS
port 42 nsew
rlabel metal1 s 21202 -867 21248 -767 8 VSS
port 42 nsew
rlabel metal1 s 21006 -867 21052 -767 8 VSS
port 42 nsew
rlabel metal1 s 20810 -867 20856 -767 8 VSS
port 42 nsew
rlabel metal1 s 5766 -957 5812 -857 8 VSS
port 42 nsew
rlabel metal1 s 5570 -957 5616 -857 8 VSS
port 42 nsew
rlabel metal1 s 5374 -957 5420 -857 8 VSS
port 42 nsew
rlabel metal1 s 4916 -957 4962 -857 8 VSS
port 42 nsew
rlabel metal1 s 4720 -957 4766 -857 8 VSS
port 42 nsew
rlabel metal1 s 4524 -957 4570 -857 8 VSS
port 42 nsew
rlabel metal1 s 19472 -566 20517 -496 8 VSS
port 42 nsew
rlabel metal1 s 21202 -452 21248 -352 8 VSS
port 42 nsew
rlabel metal1 s 21006 -452 21052 -352 8 VSS
port 42 nsew
rlabel metal1 s 20810 -452 20856 -352 8 VSS
port 42 nsew
rlabel metal1 s 20352 -452 20398 -352 8 VSS
port 42 nsew
rlabel metal1 s 20156 -452 20202 -352 8 VSS
port 42 nsew
rlabel metal1 s 19960 -452 20006 -352 8 VSS
port 42 nsew
rlabel metal1 s 38044 -150 38090 250 6 VSS
port 42 nsew
rlabel metal1 s 37886 -150 37932 250 6 VSS
port 42 nsew
rlabel metal1 s 37728 -150 37774 250 6 VSS
port 42 nsew
rlabel metal1 s 37570 -150 37616 250 6 VSS
port 42 nsew
rlabel metal1 s 37412 -150 37458 250 6 VSS
port 42 nsew
rlabel metal1 s 37096 -150 37142 250 6 VSS
port 42 nsew
rlabel metal1 s 36780 -150 36826 250 6 VSS
port 42 nsew
rlabel metal1 s 36323 -193 36369 207 6 VSS
port 42 nsew
rlabel metal1 s 36165 -193 36211 207 6 VSS
port 42 nsew
rlabel metal1 s 36007 -193 36053 207 6 VSS
port 42 nsew
rlabel metal1 s 35849 -193 35895 207 6 VSS
port 42 nsew
rlabel metal1 s 35691 -193 35737 207 6 VSS
port 42 nsew
rlabel metal1 s 35375 -193 35421 207 6 VSS
port 42 nsew
rlabel metal1 s 35059 -193 35105 207 6 VSS
port 42 nsew
rlabel metal1 s 34513 -28 34559 172 6 VSS
port 42 nsew
rlabel metal1 s 34355 -28 34401 316 6 VSS
port 42 nsew
rlabel metal1 s 34080 -28 34126 172 6 VSS
port 42 nsew
rlabel metal1 s 33764 -28 33810 172 6 VSS
port 42 nsew
rlabel metal1 s 33448 -28 33494 172 6 VSS
port 42 nsew
rlabel metal1 s 33132 -28 33178 172 6 VSS
port 42 nsew
rlabel metal1 s 32816 -28 32862 172 6 VSS
port 42 nsew
rlabel metal1 s 34128 316 34401 362 6 VSS
port 42 nsew
rlabel metal1 s 32544 -30 32590 345 6 VSS
port 42 nsew
rlabel metal1 s 32386 -30 32432 170 6 VSS
port 42 nsew
rlabel metal1 s 31588 -216 31634 184 8 VSS
port 42 nsew
rlabel metal1 s 31430 -216 31476 184 8 VSS
port 42 nsew
rlabel metal1 s 31272 -216 31318 184 8 VSS
port 42 nsew
rlabel metal1 s 31114 -216 31160 184 8 VSS
port 42 nsew
rlabel metal1 s 30956 -216 31002 184 8 VSS
port 42 nsew
rlabel metal1 s 30640 -216 30686 184 8 VSS
port 42 nsew
rlabel metal1 s 30324 -216 30370 184 8 VSS
port 42 nsew
rlabel metal1 s 29658 -21 29704 179 6 VSS
port 42 nsew
rlabel metal1 s 34128 362 34174 682 6 VSS
port 42 nsew
rlabel metal1 s 32544 345 32711 391 6 VSS
port 42 nsew
rlabel metal1 s 29500 -21 29546 323 6 VSS
port 42 nsew
rlabel metal1 s 29225 -21 29271 179 6 VSS
port 42 nsew
rlabel metal1 s 28909 -21 28955 179 6 VSS
port 42 nsew
rlabel metal1 s 28593 -21 28639 179 6 VSS
port 42 nsew
rlabel metal1 s 28277 -21 28323 179 6 VSS
port 42 nsew
rlabel metal1 s 27961 -21 28007 179 6 VSS
port 42 nsew
rlabel metal1 s 29273 323 29546 369 6 VSS
port 42 nsew
rlabel metal1 s 27689 -23 27735 352 6 VSS
port 42 nsew
rlabel metal1 s 27531 -23 27577 177 6 VSS
port 42 nsew
rlabel metal1 s 33970 482 34016 682 6 VSS
port 42 nsew
rlabel metal1 s 34129 930 34175 1130 6 VSS
port 42 nsew
rlabel metal1 s 33971 930 34017 1130 6 VSS
port 42 nsew
rlabel metal1 s 32823 482 32869 1134 6 VSS
port 42 nsew
rlabel metal1 s 32665 391 32711 1134 6 VSS
port 42 nsew
rlabel metal1 s 29273 369 29319 689 6 VSS
port 42 nsew
rlabel metal1 s 27689 352 27856 398 6 VSS
port 42 nsew
rlabel metal1 s 29115 489 29161 689 6 VSS
port 42 nsew
rlabel metal1 s 29274 937 29320 1137 6 VSS
port 42 nsew
rlabel metal1 s 29116 937 29162 1137 6 VSS
port 42 nsew
rlabel metal1 s 27968 489 28014 1141 6 VSS
port 42 nsew
rlabel metal1 s 27810 398 27856 1141 6 VSS
port 42 nsew
rlabel metal1 s 22436 895 22925 943 6 VSS
port 42 nsew
rlabel metal1 s 19472 -496 19542 943 6 VSS
port 42 nsew
rlabel metal1 s 19472 943 22925 1241 6 VSS
port 42 nsew
rlabel metal1 s 22436 1241 22925 1317 6 VSS
port 42 nsew
rlabel metal1 s 14984 1049 15030 1449 6 VSS
port 42 nsew
rlabel metal1 s 14866 1049 14912 1449 6 VSS
port 42 nsew
rlabel metal1 s 14748 1049 14794 1449 6 VSS
port 42 nsew
rlabel metal1 s 14630 1049 14676 1449 6 VSS
port 42 nsew
rlabel metal1 s 14512 1049 14558 1449 6 VSS
port 42 nsew
rlabel metal1 s 14394 1049 14440 1449 6 VSS
port 42 nsew
rlabel metal1 s 14276 1049 14322 1449 6 VSS
port 42 nsew
rlabel metal1 s 14158 1049 14204 1449 6 VSS
port 42 nsew
rlabel metal1 s 14040 1049 14086 1449 6 VSS
port 42 nsew
rlabel metal1 s 13922 1049 13968 1449 6 VSS
port 42 nsew
rlabel metal1 s 13804 1049 13850 1449 6 VSS
port 42 nsew
rlabel metal1 s 13686 1049 13732 1449 6 VSS
port 42 nsew
rlabel metal1 s 13568 1049 13614 1449 6 VSS
port 42 nsew
rlabel metal1 s 13450 1049 13496 1449 6 VSS
port 42 nsew
rlabel metal1 s 13332 1049 13378 1449 6 VSS
port 42 nsew
rlabel metal1 s 13214 1049 13260 1449 6 VSS
port 42 nsew
rlabel metal1 s 13096 1049 13142 1449 6 VSS
port 42 nsew
rlabel metal1 s 12978 1049 13024 1449 6 VSS
port 42 nsew
rlabel metal1 s 12860 1049 12906 1449 6 VSS
port 42 nsew
rlabel metal1 s 12742 1049 12788 1449 6 VSS
port 42 nsew
rlabel metal1 s 12624 1049 12670 1449 6 VSS
port 42 nsew
rlabel metal1 s 12506 1049 12552 1449 6 VSS
port 42 nsew
rlabel metal1 s 12388 1049 12434 1449 6 VSS
port 42 nsew
rlabel metal1 s 12270 1049 12316 1449 6 VSS
port 42 nsew
rlabel metal1 s 12152 1049 12198 1449 6 VSS
port 42 nsew
rlabel metal1 s 12034 1049 12080 1449 6 VSS
port 42 nsew
rlabel metal1 s 11916 1049 11962 1449 6 VSS
port 42 nsew
rlabel metal1 s 11798 1049 11844 1449 6 VSS
port 42 nsew
rlabel metal1 s 11680 1049 11726 1449 6 VSS
port 42 nsew
rlabel metal1 s 11562 1049 11608 1449 6 VSS
port 42 nsew
rlabel metal1 s 11444 1049 11490 1449 6 VSS
port 42 nsew
rlabel metal1 s 11208 1049 11254 1449 6 VSS
port 42 nsew
rlabel metal1 s 10972 1049 11018 1449 6 VSS
port 42 nsew
rlabel metal1 s 10736 1049 10782 1449 6 VSS
port 42 nsew
rlabel metal1 s 10500 1049 10546 1449 6 VSS
port 42 nsew
rlabel metal1 s 10264 1049 10310 1449 6 VSS
port 42 nsew
rlabel metal1 s 10028 1049 10074 1449 6 VSS
port 42 nsew
rlabel metal1 s 9792 1049 9838 1449 6 VSS
port 42 nsew
rlabel metal1 s 9556 1049 9602 1449 6 VSS
port 42 nsew
rlabel metal1 s 9320 1049 9366 1449 6 VSS
port 42 nsew
rlabel metal1 s 9084 1049 9130 1449 6 VSS
port 42 nsew
rlabel metal1 s 8848 1049 8894 1449 6 VSS
port 42 nsew
rlabel metal1 s 8612 1049 8658 1449 6 VSS
port 42 nsew
rlabel metal1 s 8376 1049 8422 1449 6 VSS
port 42 nsew
rlabel metal1 s 8140 1049 8186 1449 6 VSS
port 42 nsew
rlabel metal1 s 7904 1049 7950 1449 6 VSS
port 42 nsew
rlabel metal1 s 3841 -1011 3899 1101 6 VSS
port 42 nsew
rlabel metal1 s 2794 355 3099 439 6 VSS
port 42 nsew
rlabel metal1 s 2794 439 3235 470 6 VSS
port 42 nsew
rlabel metal1 s 2391 470 3235 506 6 VSS
port 42 nsew
rlabel metal1 s 2794 506 3235 589 6 VSS
port 42 nsew
rlabel metal1 s 3061 589 3235 1101 6 VSS
port 42 nsew
rlabel metal1 s 2803 777 2849 892 6 VSS
port 42 nsew
rlabel metal1 s 2494 777 2540 861 6 VSS
port 42 nsew
rlabel metal1 s 2391 506 2427 892 6 VSS
port 42 nsew
rlabel metal1 s 2177 740 2223 892 6 VSS
port 42 nsew
rlabel metal1 s 1941 740 1987 892 6 VSS
port 42 nsew
rlabel metal1 s 1509 747 1555 867 6 VSS
port 42 nsew
rlabel metal1 s 1219 752 1265 872 6 VSS
port 42 nsew
rlabel metal1 s 707 777 753 861 6 VSS
port 42 nsew
rlabel metal1 s 1941 892 2849 928 6 VSS
port 42 nsew
rlabel metal1 s 3061 1101 3899 1159 6 VSS
port 42 nsew
rlabel metal1 s 5751 1318 5797 1418 6 VSS
port 42 nsew
rlabel metal1 s 5555 1318 5601 1418 6 VSS
port 42 nsew
rlabel metal1 s 5359 1318 5405 1418 6 VSS
port 42 nsew
rlabel metal1 s 4580 1384 4827 1385 6 VSS
port 42 nsew
rlabel metal1 s 4186 1385 4963 1519 6 VSS
port 42 nsew
rlabel metal1 s 58262 1826 58308 2226 6 VSS
port 42 nsew
rlabel metal1 s 58144 1826 58190 2226 6 VSS
port 42 nsew
rlabel metal1 s 58026 1826 58072 2226 6 VSS
port 42 nsew
rlabel metal1 s 57908 1826 57954 2226 6 VSS
port 42 nsew
rlabel metal1 s 57790 1826 57836 2226 6 VSS
port 42 nsew
rlabel metal1 s 57672 1826 57718 2226 6 VSS
port 42 nsew
rlabel metal1 s 57554 1826 57600 2226 6 VSS
port 42 nsew
rlabel metal1 s 57436 1826 57482 2226 6 VSS
port 42 nsew
rlabel metal1 s 57318 1826 57364 2226 6 VSS
port 42 nsew
rlabel metal1 s 57200 1826 57246 2226 6 VSS
port 42 nsew
rlabel metal1 s 57082 1826 57128 2226 6 VSS
port 42 nsew
rlabel metal1 s 56964 1826 57010 2226 6 VSS
port 42 nsew
rlabel metal1 s 56846 1826 56892 2226 6 VSS
port 42 nsew
rlabel metal1 s 56728 1826 56774 2226 6 VSS
port 42 nsew
rlabel metal1 s 56610 1826 56656 2226 6 VSS
port 42 nsew
rlabel metal1 s 56492 1826 56538 2226 6 VSS
port 42 nsew
rlabel metal1 s 56374 1826 56420 2226 6 VSS
port 42 nsew
rlabel metal1 s 56256 1826 56302 2226 6 VSS
port 42 nsew
rlabel metal1 s 56138 1826 56184 2226 6 VSS
port 42 nsew
rlabel metal1 s 56020 1826 56066 2226 6 VSS
port 42 nsew
rlabel metal1 s 55902 1826 55948 2226 6 VSS
port 42 nsew
rlabel metal1 s 55784 1826 55830 2226 6 VSS
port 42 nsew
rlabel metal1 s 55666 1826 55712 2226 6 VSS
port 42 nsew
rlabel metal1 s 55548 1826 55594 2226 6 VSS
port 42 nsew
rlabel metal1 s 55430 1826 55476 2226 6 VSS
port 42 nsew
rlabel metal1 s 55312 1826 55358 2226 6 VSS
port 42 nsew
rlabel metal1 s 55194 1826 55240 2226 6 VSS
port 42 nsew
rlabel metal1 s 55076 1826 55122 2226 6 VSS
port 42 nsew
rlabel metal1 s 54958 1826 55004 2226 6 VSS
port 42 nsew
rlabel metal1 s 54840 1826 54886 2226 6 VSS
port 42 nsew
rlabel metal1 s 54722 1826 54768 2226 6 VSS
port 42 nsew
rlabel metal1 s 54486 1826 54532 2226 6 VSS
port 42 nsew
rlabel metal1 s 54250 1826 54296 2226 6 VSS
port 42 nsew
rlabel metal1 s 54014 1826 54060 2226 6 VSS
port 42 nsew
rlabel metal1 s 53778 1826 53824 2226 6 VSS
port 42 nsew
rlabel metal1 s 53542 1826 53588 2226 6 VSS
port 42 nsew
rlabel metal1 s 53306 1826 53352 2226 6 VSS
port 42 nsew
rlabel metal1 s 53070 1826 53116 2226 6 VSS
port 42 nsew
rlabel metal1 s 52834 1826 52880 2226 6 VSS
port 42 nsew
rlabel metal1 s 52598 1826 52644 2226 6 VSS
port 42 nsew
rlabel metal1 s 52362 1826 52408 2226 6 VSS
port 42 nsew
rlabel metal1 s 52126 1826 52172 2226 6 VSS
port 42 nsew
rlabel metal1 s 51890 1826 51936 2226 6 VSS
port 42 nsew
rlabel metal1 s 51654 1826 51700 2226 6 VSS
port 42 nsew
rlabel metal1 s 51418 1826 51464 2226 6 VSS
port 42 nsew
rlabel metal1 s 51182 1826 51228 2226 6 VSS
port 42 nsew
rlabel metal1 s 45965 1887 46011 1987 6 VSS
port 42 nsew
rlabel metal1 s 45769 1887 45815 1987 6 VSS
port 42 nsew
rlabel metal1 s 45573 1887 45619 1987 6 VSS
port 42 nsew
rlabel metal1 s 44995 1797 45041 1897 6 VSS
port 42 nsew
rlabel metal1 s 44799 1797 44845 1897 6 VSS
port 42 nsew
rlabel metal1 s 44603 1797 44649 1897 6 VSS
port 42 nsew
rlabel metal1 s 44158 1797 44204 1897 6 VSS
port 42 nsew
rlabel metal1 s 43962 1797 44008 1897 6 VSS
port 42 nsew
rlabel metal1 s 43766 1797 43812 1897 6 VSS
port 42 nsew
rlabel metal1 s 42295 1797 42341 1897 6 VSS
port 42 nsew
rlabel metal1 s 42099 1797 42145 1897 6 VSS
port 42 nsew
rlabel metal1 s 41903 1797 41949 1897 6 VSS
port 42 nsew
rlabel metal1 s 41458 1797 41504 1897 6 VSS
port 42 nsew
rlabel metal1 s 41262 1797 41308 1897 6 VSS
port 42 nsew
rlabel metal1 s 41066 1797 41112 1897 6 VSS
port 42 nsew
rlabel metal1 s 5751 1733 5797 1833 6 VSS
port 42 nsew
rlabel metal1 s 5555 1733 5601 1833 6 VSS
port 42 nsew
rlabel metal1 s 5359 1733 5405 1833 6 VSS
port 42 nsew
rlabel metal1 s 4901 1733 4947 1833 6 VSS
port 42 nsew
rlabel metal1 s 4705 1733 4751 1833 6 VSS
port 42 nsew
rlabel metal1 s 4509 1733 4555 1833 6 VSS
port 42 nsew
rlabel metal1 s 44670 2060 44807 2120 6 VSS
port 42 nsew
rlabel metal1 s 45804 2255 45950 2335 6 VSS
port 42 nsew
rlabel metal1 s 44697 2120 44792 2335 6 VSS
port 42 nsew
rlabel metal1 s 42073 2066 42210 2126 6 VSS
port 42 nsew
rlabel metal1 s 39440 2066 39572 2126 6 VSS
port 42 nsew
rlabel metal1 s 42104 2126 42199 2334 6 VSS
port 42 nsew
rlabel metal1 s 39460 2126 39555 2193 6 VSS
port 42 nsew
rlabel metal1 s 38780 2149 38972 2193 6 VSS
port 42 nsew
rlabel metal1 s 38780 2193 39555 2288 6 VSS
port 42 nsew
rlabel metal1 s 44697 2335 45950 2338 6 VSS
port 42 nsew
rlabel metal1 s 44684 2338 45950 2379 6 VSS
port 42 nsew
rlabel metal1 s 45804 2379 45950 2441 6 VSS
port 42 nsew
rlabel metal1 s 44684 2379 44816 2398 6 VSS
port 42 nsew
rlabel metal1 s 42080 2334 42217 2394 6 VSS
port 42 nsew
rlabel metal1 s 39460 2288 39555 2335 6 VSS
port 42 nsew
rlabel metal1 s 39453 2335 39590 2395 6 VSS
port 42 nsew
rlabel metal1 s 38780 2288 38972 2407 6 VSS
port 42 nsew
rlabel metal1 s 38805 2407 38941 2408 6 VSS
port 42 nsew
rlabel metal1 s 44897 2455 44943 2555 6 VSS
port 42 nsew
rlabel metal1 s 44701 2455 44747 2555 6 VSS
port 42 nsew
rlabel metal1 s 44505 2455 44551 2555 6 VSS
port 42 nsew
rlabel metal1 s 43154 2455 43200 2555 6 VSS
port 42 nsew
rlabel metal1 s 42958 2455 43004 2555 6 VSS
port 42 nsew
rlabel metal1 s 42762 2455 42808 2555 6 VSS
port 42 nsew
rlabel metal1 s 42197 2455 42243 2555 6 VSS
port 42 nsew
rlabel metal1 s 42001 2455 42047 2555 6 VSS
port 42 nsew
rlabel metal1 s 41805 2455 41851 2555 6 VSS
port 42 nsew
rlabel metal1 s 40454 2455 40500 2555 6 VSS
port 42 nsew
rlabel metal1 s 40258 2455 40304 2555 6 VSS
port 42 nsew
rlabel metal1 s 40062 2455 40108 2555 6 VSS
port 42 nsew
rlabel metal1 s 39572 2455 39618 2555 6 VSS
port 42 nsew
rlabel metal1 s 39376 2455 39422 2555 6 VSS
port 42 nsew
rlabel metal1 s 39180 2455 39226 2555 6 VSS
port 42 nsew
rlabel metal1 s 38044 2075 38090 2475 6 VSS
port 42 nsew
rlabel metal1 s 37886 2075 37932 2475 6 VSS
port 42 nsew
rlabel metal1 s 37728 2075 37774 2475 6 VSS
port 42 nsew
rlabel metal1 s 37570 2075 37616 2475 6 VSS
port 42 nsew
rlabel metal1 s 37412 2075 37458 2475 6 VSS
port 42 nsew
rlabel metal1 s 37096 2075 37142 2475 6 VSS
port 42 nsew
rlabel metal1 s 36780 2075 36826 2475 6 VSS
port 42 nsew
rlabel metal1 s 36323 2118 36369 2518 6 VSS
port 42 nsew
rlabel metal1 s 36165 2118 36211 2518 6 VSS
port 42 nsew
rlabel metal1 s 36007 2118 36053 2518 6 VSS
port 42 nsew
rlabel metal1 s 35849 2118 35895 2518 6 VSS
port 42 nsew
rlabel metal1 s 35691 2118 35737 2518 6 VSS
port 42 nsew
rlabel metal1 s 35375 2118 35421 2518 6 VSS
port 42 nsew
rlabel metal1 s 35059 2118 35105 2518 6 VSS
port 42 nsew
rlabel metal1 s 31588 2096 31634 2496 6 VSS
port 42 nsew
rlabel metal1 s 31430 2096 31476 2496 6 VSS
port 42 nsew
rlabel metal1 s 31272 2096 31318 2496 6 VSS
port 42 nsew
rlabel metal1 s 31114 2096 31160 2496 6 VSS
port 42 nsew
rlabel metal1 s 30956 2096 31002 2496 6 VSS
port 42 nsew
rlabel metal1 s 30640 2096 30686 2496 6 VSS
port 42 nsew
rlabel metal1 s 30324 2096 30370 2496 6 VSS
port 42 nsew
rlabel metal1 s 3061 1159 3235 2272 6 VSS
port 42 nsew
rlabel metal1 s 1941 1934 2849 1970 6 VSS
port 42 nsew
rlabel metal1 s 2803 1970 2849 2085 6 VSS
port 42 nsew
rlabel metal1 s 2494 2001 2540 2085 6 VSS
port 42 nsew
rlabel metal1 s 2809 2272 3235 2356 6 VSS
port 42 nsew
rlabel metal1 s 2391 1970 2427 2356 6 VSS
port 42 nsew
rlabel metal1 s 2177 1970 2223 2122 6 VSS
port 42 nsew
rlabel metal1 s 1941 1970 1987 2122 6 VSS
port 42 nsew
rlabel metal1 s 1509 1995 1555 2115 6 VSS
port 42 nsew
rlabel metal1 s 1219 1990 1265 2110 6 VSS
port 42 nsew
rlabel metal1 s 707 2001 753 2085 6 VSS
port 42 nsew
rlabel metal1 s 2391 2356 3235 2392 6 VSS
port 42 nsew
rlabel metal1 s 21030 2483 21076 2583 6 VSS
port 42 nsew
rlabel metal1 s 20834 2483 20880 2583 6 VSS
port 42 nsew
rlabel metal1 s 20638 2483 20684 2583 6 VSS
port 42 nsew
rlabel metal1 s 2809 2392 3235 2508 6 VSS
port 42 nsew
rlabel metal1 s 19552 2787 20314 2858 6 VSS
port 42 nsew
rlabel metal1 s 19552 2858 19659 2862 6 VSS
port 42 nsew
rlabel metal1 s 19552 2862 19650 2892 6 VSS
port 42 nsew
rlabel metal1 s 21030 2898 21076 2998 6 VSS
port 42 nsew
rlabel metal1 s 20834 2898 20880 2998 6 VSS
port 42 nsew
rlabel metal1 s 20638 2898 20684 2998 6 VSS
port 42 nsew
rlabel metal1 s 20180 2898 20226 2998 6 VSS
port 42 nsew
rlabel metal1 s 19984 2898 20030 2998 6 VSS
port 42 nsew
rlabel metal1 s 19788 2898 19834 2998 6 VSS
port 42 nsew
rlabel metal1 s 26583 3483 38866 3886 6 VSS
port 42 nsew
rlabel metal1 s 36381 3886 37574 7623 6 VSS
port 42 nsew
rlabel metal1 s 33884 3886 35077 7623 6 VSS
port 42 nsew
rlabel metal1 s 31275 3886 32468 7623 6 VSS
port 42 nsew
rlabel metal1 s 29111 3886 30304 7623 6 VSS
port 42 nsew
rlabel metal1 s 26836 3886 28029 7623 6 VSS
port 42 nsew
rlabel metal1 s 3061 2508 3235 4116 6 VSS
port 42 nsew
rlabel metal1 s 2866 4116 3250 4560 6 VSS
port 42 nsew
rlabel metal1 s 11606 4643 11652 5443 6 VSS
port 42 nsew
rlabel metal1 s 9890 4643 9936 5443 6 VSS
port 42 nsew
rlabel metal1 s 8174 4643 8220 5443 6 VSS
port 42 nsew
rlabel metal1 s 11606 5643 11652 6443 6 VSS
port 42 nsew
rlabel metal1 s 9890 5643 9936 6443 6 VSS
port 42 nsew
rlabel metal1 s 8174 5643 8220 6443 6 VSS
port 42 nsew
rlabel metal1 s 26753 7623 38073 8844 6 VSS
port 42 nsew
rlabel metal1 s -6540 7273 -5433 8032 4 VSS
port 42 nsew
rlabel metal1 s -16277 8032 -5433 8494 4 VSS
port 42 nsew
rlabel metal1 s -16277 8494 -5438 8555 4 VSS
port 42 nsew
rlabel metal1 s 17202 8956 17318 8966 6 VSS
port 42 nsew
rlabel metal1 s 16033 8966 17318 9012 6 VSS
port 42 nsew
rlabel metal1 s 17131 9012 17318 9181 6 VSS
port 42 nsew
rlabel metal1 s 16043 9012 16101 9100 6 VSS
port 42 nsew
rlabel metal1 s 16818 9100 17018 9146 6 VSS
port 42 nsew
rlabel metal1 s 15933 9100 16218 9146 6 VSS
port 42 nsew
rlabel metal1 s 15933 9146 15979 9616 6 VSS
port 42 nsew
rlabel metal1 s 16818 9616 17018 9662 6 VSS
port 42 nsew
rlabel metal1 s 15933 9616 16218 9662 6 VSS
port 42 nsew
rlabel metal1 s 15933 9662 16018 9663 6 VSS
port 42 nsew
rlabel metal1 s 15933 9663 15979 10132 6 VSS
port 42 nsew
rlabel metal1 s -15400 9872 -15366 9873 4 VSS
port 42 nsew
rlabel metal1 s -15485 9873 -15366 9941 4 VSS
port 42 nsew
rlabel metal1 s -15485 9941 -6799 10002 4 VSS
port 42 nsew
rlabel metal1 s -15485 10002 -15367 10003 4 VSS
port 42 nsew
rlabel metal1 s -15790 10032 -15666 10053 4 VSS
port 42 nsew
rlabel metal1 s -15790 10053 -15494 10055 4 VSS
port 42 nsew
rlabel metal1 s -15790 10055 -8271 10119 4 VSS
port 42 nsew
rlabel metal1 s 16818 10132 17018 10178 6 VSS
port 42 nsew
rlabel metal1 s 15933 10132 16218 10178 6 VSS
port 42 nsew
rlabel metal1 s -15790 10119 -15667 10155 4 VSS
port 42 nsew
rlabel metal1 s 15933 10178 16018 10179 6 VSS
port 42 nsew
rlabel metal1 s -16157 10183 -16034 10200 4 VSS
port 42 nsew
rlabel metal1 s -16157 10200 -7840 10260 4 VSS
port 42 nsew
rlabel metal1 s -16157 10260 -16034 10306 4 VSS
port 42 nsew
rlabel metal1 s -12288 10655 -12138 10667 4 VSS
port 42 nsew
rlabel metal1 s -12815 10442 -12700 10667 4 VSS
port 42 nsew
rlabel metal1 s -13188 10550 -12988 10596 4 VSS
port 42 nsew
rlabel metal1 s -6560 10667 -6260 10713 4 VSS
port 42 nsew
rlabel metal1 s -8521 10724 -8221 10770 4 VSS
port 42 nsew
rlabel metal1 s -12815 10667 -12138 10754 4 VSS
port 42 nsew
rlabel metal1 s -12042 10789 -11842 10835 4 VSS
port 42 nsew
rlabel metal1 s -12288 10754 -12138 10847 4 VSS
port 42 nsew
rlabel metal1 s -12815 10754 -12700 10847 4 VSS
port 42 nsew
rlabel metal1 s -12815 10847 -12138 10934 4 VSS
port 42 nsew
rlabel metal1 s -12042 10985 -11842 11031 4 VSS
port 42 nsew
rlabel metal1 s -12288 10934 -12138 11020 4 VSS
port 42 nsew
rlabel metal1 s -12815 10934 -12700 11020 4 VSS
port 42 nsew
rlabel metal1 s -12815 11020 -12138 11107 4 VSS
port 42 nsew
rlabel metal1 s -12288 11107 -12138 11204 4 VSS
port 42 nsew
rlabel metal1 s -12815 11107 -12700 11204 4 VSS
port 42 nsew
rlabel metal1 s -12815 11204 -12138 11291 4 VSS
port 42 nsew
rlabel metal1 s -12288 11291 -12138 11329 4 VSS
port 42 nsew
rlabel metal1 s -12815 11291 -12700 11329 4 VSS
port 42 nsew
rlabel metal1 s 16949 11350 17282 16839 6 VSS
port 42 nsew
rlabel metal1 s -8014 11333 -7914 11379 4 VSS
port 42 nsew
rlabel metal1 s -12815 11329 -12138 11416 4 VSS
port 42 nsew
rlabel metal1 s -12288 11416 -12138 11459 4 VSS
port 42 nsew
rlabel metal1 s -12815 11416 -12700 11425 4 VSS
port 42 nsew
rlabel metal1 s -8014 11529 -7914 11575 4 VSS
port 42 nsew
rlabel metal1 s -13289 11582 -12989 11628 4 VSS
port 42 nsew
rlabel metal1 s -6561 11699 -6361 11745 4 VSS
port 42 nsew
rlabel metal1 s -12494 11796 -12357 11797 4 VSS
port 42 nsew
rlabel metal1 s -12494 11797 -11407 11798 4 VSS
port 42 nsew
rlabel metal1 s -12494 11798 -11403 11840 4 VSS
port 42 nsew
rlabel metal1 s -11540 11840 -11403 11856 4 VSS
port 42 nsew
rlabel metal1 s -12494 11840 -12357 11854 4 VSS
port 42 nsew
rlabel metal1 s -11699 11995 -11499 12041 4 VSS
port 42 nsew
rlabel metal1 s -7013 12229 -6881 12231 4 VSS
port 42 nsew
rlabel metal1 s -7013 12231 -6130 12259 4 VSS
port 42 nsew
rlabel metal1 s -11699 12191 -11499 12237 4 VSS
port 42 nsew
rlabel metal1 s -7013 12259 -6113 12267 4 VSS
port 42 nsew
rlabel metal1 s -6171 12267 -6113 12396 4 VSS
port 42 nsew
rlabel metal1 s -7013 12267 -6881 12282 4 VSS
port 42 nsew
rlabel metal1 s -8496 12497 -8196 12543 4 VSS
port 42 nsew
rlabel metal1 s -12573 12617 -12436 12639 4 VSS
port 42 nsew
rlabel metal1 s -6612 12666 -6312 12712 4 VSS
port 42 nsew
rlabel metal1 s -12573 12639 -11233 12674 4 VSS
port 42 nsew
rlabel metal1 s -11370 12674 -11233 12697 4 VSS
port 42 nsew
rlabel metal1 s -12573 12674 -12436 12675 4 VSS
port 42 nsew
rlabel metal1 s -12650 12710 -12513 12716 4 VSS
port 42 nsew
rlabel metal1 s -12650 12716 -11405 12751 4 VSS
port 42 nsew
rlabel metal1 s -11542 12751 -11405 12774 4 VSS
port 42 nsew
rlabel metal1 s -12650 12751 -12513 12768 4 VSS
port 42 nsew
rlabel metal1 s -11700 12900 -11500 12946 4 VSS
port 42 nsew
rlabel metal1 s -11700 13096 -11500 13142 4 VSS
port 42 nsew
rlabel metal1 s -6105 13275 -6005 13321 4 VSS
port 42 nsew
rlabel metal1 s -6105 13471 -6005 13517 4 VSS
port 42 nsew
rlabel metal1 s -8497 13529 -8297 13575 4 VSS
port 42 nsew
rlabel metal1 s -6500 14302 -6200 14348 4 VSS
port 42 nsew
rlabel metal1 s -8296 14328 -8096 14374 4 VSS
port 42 nsew
rlabel metal1 s -11500 14302 -11200 14348 4 VSS
port 42 nsew
rlabel metal1 s -13296 14328 -13096 14374 4 VSS
port 42 nsew
rlabel metal1 s -8296 14524 -8096 14570 4 VSS
port 42 nsew
rlabel metal1 s -13296 14524 -13096 14570 4 VSS
port 42 nsew
rlabel metal1 s -6807 14911 -6707 14957 4 VSS
port 42 nsew
rlabel metal1 s -11807 14911 -11707 14957 4 VSS
port 42 nsew
rlabel metal1 s -6807 15107 -6707 15153 4 VSS
port 42 nsew
rlabel metal1 s -11807 15107 -11707 15153 4 VSS
port 42 nsew
rlabel metal1 s -8474 15301 -8174 15347 4 VSS
port 42 nsew
rlabel metal1 s -13474 15301 -13174 15347 4 VSS
port 42 nsew
rlabel metal1 s -6214 15749 -5914 15795 4 VSS
port 42 nsew
rlabel metal1 s -11214 15749 -10914 15795 4 VSS
port 42 nsew
rlabel metal1 s -6214 15945 -5914 15991 4 VSS
port 42 nsew
rlabel metal1 s -7967 15910 -7867 15956 4 VSS
port 42 nsew
rlabel metal1 s -11214 15945 -10914 15991 4 VSS
port 42 nsew
rlabel metal1 s -12967 15910 -12867 15956 4 VSS
port 42 nsew
rlabel metal1 s -7967 16106 -7867 16152 4 VSS
port 42 nsew
rlabel metal1 s -12967 16106 -12867 16152 4 VSS
port 42 nsew
rlabel metal1 s -6214 16187 -5914 16233 4 VSS
port 42 nsew
rlabel metal1 s -11214 16187 -10914 16233 4 VSS
port 42 nsew
rlabel metal1 s -5806 16328 -5693 16709 4 VSS
port 42 nsew
rlabel metal1 s -5806 16709 -4414 16892 4 VSS
port 42 nsew
rlabel metal1 s -8115 16297 -8002 16892 4 VSS
port 42 nsew
rlabel metal1 s -10806 16328 -10693 16892 4 VSS
port 42 nsew
rlabel metal1 s -13115 16297 -13002 16892 4 VSS
port 42 nsew
rlabel metal1 s -13115 16892 -4414 16899 4 VSS
port 42 nsew
rlabel metal1 s -4604 16899 -4414 24189 4 VSS
port 42 nsew
rlabel metal1 s -13115 16899 -5693 17005 4 VSS
port 42 nsew
rlabel metal1 s -5346 18168 -5246 18214 4 VSS
port 42 nsew
rlabel metal1 s -10273 18168 -10173 18214 4 VSS
port 42 nsew
rlabel metal1 s -6004 18266 -5904 18312 4 VSS
port 42 nsew
rlabel metal1 s -10931 18266 -10831 18312 4 VSS
port 42 nsew
rlabel metal1 s -5346 18364 -5246 18410 4 VSS
port 42 nsew
rlabel metal1 s -5569 18402 -5509 18417 4 VSS
port 42 nsew
rlabel metal1 s -5847 18393 -5787 18417 4 VSS
port 42 nsew
rlabel metal1 s -10273 18364 -10173 18410 4 VSS
port 42 nsew
rlabel metal1 s -5847 18417 -5509 18512 4 VSS
port 42 nsew
rlabel metal1 s -10496 18402 -10436 18417 4 VSS
port 42 nsew
rlabel metal1 s -10774 18393 -10714 18417 4 VSS
port 42 nsew
rlabel metal1 s -6004 18462 -5904 18508 4 VSS
port 42 nsew
rlabel metal1 s -5569 18512 -5509 18539 4 VSS
port 42 nsew
rlabel metal1 s -5847 18512 -5787 18525 4 VSS
port 42 nsew
rlabel metal1 s -10774 18417 -10436 18512 4 VSS
port 42 nsew
rlabel metal1 s -10931 18462 -10831 18508 4 VSS
port 42 nsew
rlabel metal1 s -10496 18512 -10436 18539 4 VSS
port 42 nsew
rlabel metal1 s -10774 18512 -10714 18525 4 VSS
port 42 nsew
rlabel metal1 s -5346 18560 -5246 18606 4 VSS
port 42 nsew
rlabel metal1 s -10273 18560 -10173 18606 4 VSS
port 42 nsew
rlabel metal1 s -6004 18658 -5904 18704 4 VSS
port 42 nsew
rlabel metal1 s -10931 18658 -10831 18704 4 VSS
port 42 nsew
rlabel metal1 s -5346 19005 -5246 19051 4 VSS
port 42 nsew
rlabel metal1 s -10273 19005 -10173 19051 4 VSS
port 42 nsew
rlabel metal1 s -5346 19201 -5246 19247 4 VSS
port 42 nsew
rlabel metal1 s -10273 19201 -10173 19247 4 VSS
port 42 nsew
rlabel metal1 s -7476 19291 -7176 19337 4 VSS
port 42 nsew
rlabel metal1 s -9272 19317 -9072 19363 4 VSS
port 42 nsew
rlabel metal1 s -5346 19397 -5246 19443 4 VSS
port 42 nsew
rlabel metal1 s -10273 19397 -10173 19443 4 VSS
port 42 nsew
rlabel metal1 s -9272 19513 -9072 19559 4 VSS
port 42 nsew
rlabel metal1 s -7783 19900 -7683 19946 4 VSS
port 42 nsew
rlabel metal1 s -6004 20009 -5904 20055 4 VSS
port 42 nsew
rlabel metal1 s -10931 20009 -10831 20055 4 VSS
port 42 nsew
rlabel metal1 s -7783 20096 -7683 20142 4 VSS
port 42 nsew
rlabel metal1 s -6004 20205 -5904 20251 4 VSS
port 42 nsew
rlabel metal1 s -10931 20205 -10831 20251 4 VSS
port 42 nsew
rlabel metal1 s -9450 20290 -9150 20336 4 VSS
port 42 nsew
rlabel metal1 s -6004 20401 -5904 20447 4 VSS
port 42 nsew
rlabel metal1 s -10931 20401 -10831 20447 4 VSS
port 42 nsew
rlabel metal1 s -7190 20738 -6890 20784 4 VSS
port 42 nsew
rlabel metal1 s -5346 20868 -5246 20914 4 VSS
port 42 nsew
rlabel metal1 s -5575 20999 -5515 21010 4 VSS
port 42 nsew
rlabel metal1 s -5843 20992 -5783 21010 4 VSS
port 42 nsew
rlabel metal1 s -5346 21064 -5246 21110 4 VSS
port 42 nsew
rlabel metal1 s -5843 21010 -5515 21105 4 VSS
port 42 nsew
rlabel metal1 s -6004 20966 -5904 21012 4 VSS
port 42 nsew
rlabel metal1 s -7190 20934 -6890 20980 4 VSS
port 42 nsew
rlabel metal1 s -8943 20899 -8843 20945 4 VSS
port 42 nsew
rlabel metal1 s -10273 20868 -10173 20914 4 VSS
port 42 nsew
rlabel metal1 s -10502 20999 -10442 21010 4 VSS
port 42 nsew
rlabel metal1 s -10770 20992 -10710 21010 4 VSS
port 42 nsew
rlabel metal1 s -5575 21105 -5515 21136 4 VSS
port 42 nsew
rlabel metal1 s -5843 21105 -5783 21129 4 VSS
port 42 nsew
rlabel metal1 s -8943 21095 -8843 21141 4 VSS
port 42 nsew
rlabel metal1 s -10273 21064 -10173 21110 4 VSS
port 42 nsew
rlabel metal1 s -10770 21010 -10442 21105 4 VSS
port 42 nsew
rlabel metal1 s -10931 20966 -10831 21012 4 VSS
port 42 nsew
rlabel metal1 s -10502 21105 -10442 21136 4 VSS
port 42 nsew
rlabel metal1 s -10770 21105 -10710 21129 4 VSS
port 42 nsew
rlabel metal1 s -6004 21162 -5904 21208 4 VSS
port 42 nsew
rlabel metal1 s -7190 21176 -6890 21222 4 VSS
port 42 nsew
rlabel metal1 s -10931 21162 -10831 21208 4 VSS
port 42 nsew
rlabel metal1 s -5346 21260 -5246 21306 4 VSS
port 42 nsew
rlabel metal1 s -6004 21358 -5904 21404 4 VSS
port 42 nsew
rlabel metal1 s -5346 21705 -5246 21751 4 VSS
port 42 nsew
rlabel metal1 s -6782 21317 -6669 21881 4 VSS
port 42 nsew
rlabel metal1 s -9091 21286 -8978 21881 4 VSS
port 42 nsew
rlabel metal1 s -10273 21260 -10173 21306 4 VSS
port 42 nsew
rlabel metal1 s -10931 21358 -10831 21404 4 VSS
port 42 nsew
rlabel metal1 s -10273 21705 -10173 21751 4 VSS
port 42 nsew
rlabel metal1 s -5346 21901 -5246 21947 4 VSS
port 42 nsew
rlabel metal1 s -9091 21881 -6669 21994 4 VSS
port 42 nsew
rlabel metal1 s -10273 21901 -10173 21947 4 VSS
port 42 nsew
rlabel metal1 s -5346 22097 -5246 22143 4 VSS
port 42 nsew
rlabel metal1 s -6004 22709 -5904 22755 4 VSS
port 42 nsew
rlabel metal1 s -6004 22905 -5904 22951 4 VSS
port 42 nsew
rlabel metal1 s -6004 23101 -5904 23147 4 VSS
port 42 nsew
rlabel metal1 s -5575 23637 -5515 23654 4 VSS
port 42 nsew
rlabel metal1 s -5844 23619 -5784 23654 4 VSS
port 42 nsew
rlabel metal1 s -6004 23591 -5904 23637 4 VSS
port 42 nsew
rlabel metal1 s -5844 23654 -5515 23749 4 VSS
port 42 nsew
rlabel metal1 s -5575 23749 -5515 23769 4 VSS
port 42 nsew
rlabel metal1 s -5735 23749 -5640 24189 4 VSS
port 42 nsew
rlabel metal1 s -5844 23749 -5784 23756 4 VSS
port 42 nsew
rlabel metal1 s -6782 21994 -6669 23654 4 VSS
port 42 nsew
rlabel metal1 s -10273 22097 -10173 22143 4 VSS
port 42 nsew
rlabel metal1 s -10931 22709 -10831 22755 4 VSS
port 42 nsew
rlabel metal1 s -10931 22905 -10831 22951 4 VSS
port 42 nsew
rlabel metal1 s -10931 23101 -10831 23147 4 VSS
port 42 nsew
rlabel metal1 s -10502 23637 -10442 23654 4 VSS
port 42 nsew
rlabel metal1 s -10771 23619 -10711 23654 4 VSS
port 42 nsew
rlabel metal1 s -10931 23591 -10831 23637 4 VSS
port 42 nsew
rlabel metal1 s -10771 23654 -6669 23749 4 VSS
port 42 nsew
rlabel metal1 s -6004 23787 -5904 23833 4 VSS
port 42 nsew
rlabel metal1 s -6004 23983 -5904 24029 4 VSS
port 42 nsew
rlabel metal1 s -6782 23749 -6669 24189 4 VSS
port 42 nsew
rlabel metal1 s -10502 23749 -10442 23769 4 VSS
port 42 nsew
rlabel metal1 s -10771 23749 -10711 23756 4 VSS
port 42 nsew
rlabel metal1 s -10931 23787 -10831 23833 4 VSS
port 42 nsew
rlabel metal1 s -10931 23983 -10831 24029 4 VSS
port 42 nsew
rlabel metal1 s -6782 24189 -4414 24284 4 VSS
port 42 nsew
rlabel metal1 s -4604 24284 -4414 41117 4 VSS
port 42 nsew
rlabel metal1 s -6782 24284 -6669 24285 4 VSS
port 42 nsew
rlabel metal1 s -6088 24613 -5788 24659 4 VSS
port 42 nsew
rlabel metal1 s -11022 24640 -10722 24686 4 VSS
port 42 nsew
rlabel metal1 s -6088 24855 -5788 24901 4 VSS
port 42 nsew
rlabel metal1 s -11022 24882 -10722 24928 4 VSS
port 42 nsew
rlabel metal1 s -6088 25051 -5788 25097 4 VSS
port 42 nsew
rlabel metal1 s -11022 25078 -10722 25124 4 VSS
port 42 nsew
rlabel metal1 s -11220 25589 -11125 25804 4 VSS
port 42 nsew
rlabel metal1 s -5878 25862 -5678 25908 4 VSS
port 42 nsew
rlabel metal1 s -11220 25804 -10951 25899 4 VSS
port 42 nsew
rlabel metal1 s -8442 26042 -8342 26088 4 VSS
port 42 nsew
rlabel metal1 s -10540 26042 -10440 26088 4 VSS
port 42 nsew
rlabel metal1 s -7784 26140 -7684 26186 4 VSS
port 42 nsew
rlabel metal1 s -5878 26276 -5678 26322 4 VSS
port 42 nsew
rlabel metal1 s -7901 26267 -7841 26291 4 VSS
port 42 nsew
rlabel metal1 s -8179 26276 -8119 26291 4 VSS
port 42 nsew
rlabel metal1 s -8442 26238 -8342 26284 4 VSS
port 42 nsew
rlabel metal1 s -10540 26238 -10440 26284 4 VSS
port 42 nsew
rlabel metal1 s -6221 26299 -6121 26345 4 VSS
port 42 nsew
rlabel metal1 s -7784 26336 -7684 26382 4 VSS
port 42 nsew
rlabel metal1 s -8179 26291 -7841 26386 4 VSS
port 42 nsew
rlabel metal1 s -7901 26386 -7841 26399 4 VSS
port 42 nsew
rlabel metal1 s -8179 26386 -8119 26413 4 VSS
port 42 nsew
rlabel metal1 s -10763 26276 -10703 26291 4 VSS
port 42 nsew
rlabel metal1 s -11046 25899 -10951 26291 4 VSS
port 42 nsew
rlabel metal1 s -13204 25862 -13004 25908 4 VSS
port 42 nsew
rlabel metal1 s -11198 26140 -11098 26186 4 VSS
port 42 nsew
rlabel metal1 s -11046 26291 -10703 26386 4 VSS
port 42 nsew
rlabel metal1 s -13204 26276 -13004 26322 4 VSS
port 42 nsew
rlabel metal1 s -11198 26336 -11098 26382 4 VSS
port 42 nsew
rlabel metal1 s -10763 26386 -10703 26413 4 VSS
port 42 nsew
rlabel metal1 s -11041 26386 -10981 26399 4 VSS
port 42 nsew
rlabel metal1 s -8442 26434 -8342 26480 4 VSS
port 42 nsew
rlabel metal1 s -10540 26434 -10440 26480 4 VSS
port 42 nsew
rlabel metal1 s -6221 26495 -6121 26541 4 VSS
port 42 nsew
rlabel metal1 s -7784 26532 -7684 26578 4 VSS
port 42 nsew
rlabel metal1 s -11198 26532 -11098 26578 4 VSS
port 42 nsew
rlabel metal1 s -6221 26691 -6121 26737 4 VSS
port 42 nsew
rlabel metal1 s -8442 26879 -8342 26925 4 VSS
port 42 nsew
rlabel metal1 s -10540 26879 -10440 26925 4 VSS
port 42 nsew
rlabel metal1 s -8442 27075 -8342 27121 4 VSS
port 42 nsew
rlabel metal1 s -10540 27075 -10440 27121 4 VSS
port 42 nsew
rlabel metal1 s -8442 27271 -8342 27317 4 VSS
port 42 nsew
rlabel metal1 s -10540 27271 -10440 27317 4 VSS
port 42 nsew
rlabel metal1 s -5878 27340 -5678 27386 4 VSS
port 42 nsew
rlabel metal1 s -13204 27340 -13004 27386 4 VSS
port 42 nsew
rlabel metal1 s -5878 27649 -5678 27695 4 VSS
port 42 nsew
rlabel metal1 s -13204 27649 -13004 27695 4 VSS
port 42 nsew
rlabel metal1 s -7784 27883 -7684 27929 4 VSS
port 42 nsew
rlabel metal1 s -11198 27883 -11098 27929 4 VSS
port 42 nsew
rlabel metal1 s -7784 28079 -7684 28125 4 VSS
port 42 nsew
rlabel metal1 s -11198 28079 -11098 28125 4 VSS
port 42 nsew
rlabel metal1 s -7784 28275 -7684 28321 4 VSS
port 42 nsew
rlabel metal1 s -11198 28275 -11098 28321 4 VSS
port 42 nsew
rlabel metal1 s -5878 28362 -5678 28408 4 VSS
port 42 nsew
rlabel metal1 s -13204 28362 -13004 28408 4 VSS
port 42 nsew
rlabel metal1 s -5584 28749 -5530 28888 4 VSS
port 42 nsew
rlabel metal1 s -5878 28776 -5678 28822 4 VSS
port 42 nsew
rlabel metal1 s -8442 28742 -8342 28788 4 VSS
port 42 nsew
rlabel metal1 s -10540 28742 -10440 28788 4 VSS
port 42 nsew
rlabel metal1 s -13204 28776 -13004 28822 4 VSS
port 42 nsew
rlabel metal1 s -7784 28840 -7684 28886 4 VSS
port 42 nsew
rlabel metal1 s -7905 28866 -7845 28884 4 VSS
port 42 nsew
rlabel metal1 s -8173 28873 -8113 28884 4 VSS
port 42 nsew
rlabel metal1 s -5567 28888 -5539 29827 4 VSS
port 42 nsew
rlabel metal1 s -8173 28884 -7845 28979 4 VSS
port 42 nsew
rlabel metal1 s -10769 28873 -10709 28884 4 VSS
port 42 nsew
rlabel metal1 s -11037 28866 -10977 28884 4 VSS
port 42 nsew
rlabel metal1 s -7905 28979 -7845 29003 4 VSS
port 42 nsew
rlabel metal1 s -8173 28979 -8113 29010 4 VSS
port 42 nsew
rlabel metal1 s -8442 28938 -8342 28984 4 VSS
port 42 nsew
rlabel metal1 s -10540 28938 -10440 28984 4 VSS
port 42 nsew
rlabel metal1 s -11037 28884 -10709 28979 4 VSS
port 42 nsew
rlabel metal1 s -11198 28840 -11098 28886 4 VSS
port 42 nsew
rlabel metal1 s -13352 28749 -13298 28888 4 VSS
port 42 nsew
rlabel metal1 s -10769 28979 -10709 29010 4 VSS
port 42 nsew
rlabel metal1 s -11037 28979 -10977 29003 4 VSS
port 42 nsew
rlabel metal1 s -7784 29036 -7684 29082 4 VSS
port 42 nsew
rlabel metal1 s -11198 29036 -11098 29082 4 VSS
port 42 nsew
rlabel metal1 s -8442 29134 -8342 29180 4 VSS
port 42 nsew
rlabel metal1 s -10540 29134 -10440 29180 4 VSS
port 42 nsew
rlabel metal1 s -7784 29232 -7684 29278 4 VSS
port 42 nsew
rlabel metal1 s -11198 29232 -11098 29278 4 VSS
port 42 nsew
rlabel metal1 s -8442 29579 -8342 29625 4 VSS
port 42 nsew
rlabel metal1 s -10540 29579 -10440 29625 4 VSS
port 42 nsew
rlabel metal1 s -8442 29775 -8342 29821 4 VSS
port 42 nsew
rlabel metal1 s -10540 29775 -10440 29821 4 VSS
port 42 nsew
rlabel metal1 s -13343 28888 -13315 29827 4 VSS
port 42 nsew
rlabel metal1 s -5590 29827 -5536 29966 4 VSS
port 42 nsew
rlabel metal1 s -5878 29840 -5678 29886 4 VSS
port 42 nsew
rlabel metal1 s -13204 29840 -13004 29886 4 VSS
port 42 nsew
rlabel metal1 s -13346 29827 -13292 29966 4 VSS
port 42 nsew
rlabel metal1 s -5565 29966 -5537 30387 4 VSS
port 42 nsew
rlabel metal1 s -8442 29971 -8342 30017 4 VSS
port 42 nsew
rlabel metal1 s -10540 29971 -10440 30017 4 VSS
port 42 nsew
rlabel metal1 s -5878 30149 -5678 30195 4 VSS
port 42 nsew
rlabel metal1 s -13204 30149 -13004 30195 4 VSS
port 42 nsew
rlabel metal1 s -13345 29966 -13317 30387 4 VSS
port 42 nsew
rlabel metal1 s -6605 30387 -5537 30415 4 VSS
port 42 nsew
rlabel metal1 s -5878 30862 -5678 30908 4 VSS
port 42 nsew
rlabel metal1 s -5584 31249 -5530 31388 4 VSS
port 42 nsew
rlabel metal1 s -5878 31276 -5678 31322 4 VSS
port 42 nsew
rlabel metal1 s -5567 31388 -5539 32327 4 VSS
port 42 nsew
rlabel metal1 s -5590 32327 -5536 32466 4 VSS
port 42 nsew
rlabel metal1 s -5878 32340 -5678 32386 4 VSS
port 42 nsew
rlabel metal1 s -5565 32466 -5537 32871 4 VSS
port 42 nsew
rlabel metal1 s -5878 32649 -5678 32695 4 VSS
port 42 nsew
rlabel metal1 s -6458 32871 -5537 32899 4 VSS
port 42 nsew
rlabel metal1 s -5878 33362 -5678 33408 4 VSS
port 42 nsew
rlabel metal1 s -5584 33749 -5530 33888 4 VSS
port 42 nsew
rlabel metal1 s -5878 33776 -5678 33822 4 VSS
port 42 nsew
rlabel metal1 s -5567 33888 -5539 34827 4 VSS
port 42 nsew
rlabel metal1 s -5590 34827 -5536 34966 4 VSS
port 42 nsew
rlabel metal1 s -5878 34840 -5678 34886 4 VSS
port 42 nsew
rlabel metal1 s -5565 34966 -5537 35337 4 VSS
port 42 nsew
rlabel metal1 s -5878 35149 -5678 35195 4 VSS
port 42 nsew
rlabel metal1 s -6338 35337 -5537 35365 4 VSS
port 42 nsew
rlabel metal1 s -5878 35862 -5678 35908 4 VSS
port 42 nsew
rlabel metal1 s -5878 36276 -5678 36322 4 VSS
port 42 nsew
rlabel metal1 s -5878 37340 -5678 37386 4 VSS
port 42 nsew
rlabel metal1 s -5878 37649 -5678 37695 4 VSS
port 42 nsew
rlabel metal1 s -5878 38862 -5678 38908 4 VSS
port 42 nsew
rlabel metal1 s -5878 39276 -5678 39322 4 VSS
port 42 nsew
rlabel metal1 s -5878 40340 -5678 40386 4 VSS
port 42 nsew
rlabel metal1 s -5878 40649 -5678 40695 4 VSS
port 42 nsew
rlabel metal1 s -1993 42470 -862 42503 4 VSS
port 42 nsew
rlabel metal1 s -4820 42470 -3786 42503 4 VSS
port 42 nsew
rlabel metal1 s -4820 42503 -797 44054 4 VSS
port 42 nsew
rlabel metal1 s -6338 35365 -6310 42498 4 VSS
port 42 nsew
rlabel metal1 s -6458 32899 -6430 42336 4 VSS
port 42 nsew
rlabel metal1 s -6605 30415 -6569 42169 4 VSS
port 42 nsew
rlabel metal1 s -13345 30387 -12277 30415 4 VSS
port 42 nsew
rlabel metal1 s -7784 30583 -7684 30629 4 VSS
port 42 nsew
rlabel metal1 s -11198 30583 -11098 30629 4 VSS
port 42 nsew
rlabel metal1 s -7784 30779 -7684 30825 4 VSS
port 42 nsew
rlabel metal1 s -11198 30779 -11098 30825 4 VSS
port 42 nsew
rlabel metal1 s -7784 30975 -7684 31021 4 VSS
port 42 nsew
rlabel metal1 s -11198 30975 -11098 31021 4 VSS
port 42 nsew
rlabel metal1 s -7784 31465 -7684 31511 4 VSS
port 42 nsew
rlabel metal1 s -10769 31511 -10709 31528 4 VSS
port 42 nsew
rlabel metal1 s -11038 31493 -10978 31528 4 VSS
port 42 nsew
rlabel metal1 s -11198 31465 -11098 31511 4 VSS
port 42 nsew
rlabel metal1 s -11038 31528 -10709 31623 4 VSS
port 42 nsew
rlabel metal1 s -7904 31623 -7844 31658 4 VSS
port 42 nsew
rlabel metal1 s -8173 31641 -8113 31658 4 VSS
port 42 nsew
rlabel metal1 s -10769 31623 -10709 31643 4 VSS
port 42 nsew
rlabel metal1 s -11038 31623 -10978 31630 4 VSS
port 42 nsew
rlabel metal1 s -7784 31661 -7684 31707 4 VSS
port 42 nsew
rlabel metal1 s -8173 31658 -7844 31753 4 VSS
port 42 nsew
rlabel metal1 s -11198 31661 -11098 31707 4 VSS
port 42 nsew
rlabel metal1 s -7904 31753 -7844 31760 4 VSS
port 42 nsew
rlabel metal1 s -8173 31753 -8113 31773 4 VSS
port 42 nsew
rlabel metal1 s -7784 31857 -7684 31903 4 VSS
port 42 nsew
rlabel metal1 s -11198 31857 -11098 31903 4 VSS
port 42 nsew
rlabel metal1 s -8229 32395 -8029 32441 4 VSS
port 42 nsew
rlabel metal1 s -10853 32395 -10653 32441 4 VSS
port 42 nsew
rlabel metal1 s -8228 33427 -7928 33473 4 VSS
port 42 nsew
rlabel metal1 s -10954 33427 -10654 33473 4 VSS
port 42 nsew
rlabel metal1 s -7665 34226 -7565 34272 4 VSS
port 42 nsew
rlabel metal1 s -11317 34226 -11217 34272 4 VSS
port 42 nsew
rlabel metal1 s -7665 34422 -7565 34468 4 VSS
port 42 nsew
rlabel metal1 s -11317 34422 -11217 34468 4 VSS
port 42 nsew
rlabel metal1 s -8172 35031 -7872 35077 4 VSS
port 42 nsew
rlabel metal1 s -11010 35031 -10710 35077 4 VSS
port 42 nsew
rlabel metal1 s -7667 35831 -7567 35877 4 VSS
port 42 nsew
rlabel metal1 s -11315 35831 -11215 35877 4 VSS
port 42 nsew
rlabel metal1 s -7667 36027 -7567 36073 4 VSS
port 42 nsew
rlabel metal1 s -11315 36027 -11215 36073 4 VSS
port 42 nsew
rlabel metal1 s -8174 36636 -7874 36682 4 VSS
port 42 nsew
rlabel metal1 s -11008 36636 -10708 36682 4 VSS
port 42 nsew
rlabel metal1 s -8220 37357 -8020 37403 4 VSS
port 42 nsew
rlabel metal1 s -10862 37357 -10662 37403 4 VSS
port 42 nsew
rlabel metal1 s -8219 38389 -7919 38435 4 VSS
port 42 nsew
rlabel metal1 s -10963 38389 -10663 38435 4 VSS
port 42 nsew
rlabel metal1 s -8129 38872 -7929 38918 4 VSS
port 42 nsew
rlabel metal1 s -10953 38872 -10753 38918 4 VSS
port 42 nsew
rlabel metal1 s -8129 39286 -7929 39332 4 VSS
port 42 nsew
rlabel metal1 s -10953 39286 -10753 39332 4 VSS
port 42 nsew
rlabel metal1 s -8129 40350 -7929 40396 4 VSS
port 42 nsew
rlabel metal1 s -10953 40350 -10753 40396 4 VSS
port 42 nsew
rlabel metal1 s -8129 40659 -7929 40705 4 VSS
port 42 nsew
rlabel metal1 s -10953 40659 -10753 40705 4 VSS
port 42 nsew
rlabel metal1 s -12313 30415 -12277 41898 4 VSS
port 42 nsew
rlabel metal1 s -13204 30862 -13004 30908 4 VSS
port 42 nsew
rlabel metal1 s -13204 31276 -13004 31322 4 VSS
port 42 nsew
rlabel metal1 s -13352 31249 -13298 31388 4 VSS
port 42 nsew
rlabel metal1 s -13343 31388 -13315 32327 4 VSS
port 42 nsew
rlabel metal1 s -13204 32340 -13004 32386 4 VSS
port 42 nsew
rlabel metal1 s -13346 32327 -13292 32466 4 VSS
port 42 nsew
rlabel metal1 s -13204 32649 -13004 32695 4 VSS
port 42 nsew
rlabel metal1 s -13345 32466 -13317 32871 4 VSS
port 42 nsew
rlabel metal1 s -13345 32871 -12424 32899 4 VSS
port 42 nsew
rlabel metal1 s -12452 32899 -12424 41738 4 VSS
port 42 nsew
rlabel metal1 s -13204 33362 -13004 33408 4 VSS
port 42 nsew
rlabel metal1 s -13204 33776 -13004 33822 4 VSS
port 42 nsew
rlabel metal1 s -13352 33749 -13298 33888 4 VSS
port 42 nsew
rlabel metal1 s -13343 33888 -13315 34827 4 VSS
port 42 nsew
rlabel metal1 s -13204 34840 -13004 34886 4 VSS
port 42 nsew
rlabel metal1 s -13346 34827 -13292 34966 4 VSS
port 42 nsew
rlabel metal1 s -13204 35149 -13004 35195 4 VSS
port 42 nsew
rlabel metal1 s -13345 34966 -13317 35337 4 VSS
port 42 nsew
rlabel metal1 s -13345 35337 -12544 35365 4 VSS
port 42 nsew
rlabel metal1 s -12572 35365 -12544 41612 4 VSS
port 42 nsew
rlabel metal1 s -13204 35862 -13004 35908 4 VSS
port 42 nsew
rlabel metal1 s -13204 36276 -13004 36322 4 VSS
port 42 nsew
rlabel metal1 s -13204 37340 -13004 37386 4 VSS
port 42 nsew
rlabel metal1 s -13204 37649 -13004 37695 4 VSS
port 42 nsew
rlabel metal1 s -13204 38862 -13004 38908 4 VSS
port 42 nsew
rlabel metal1 s -13204 39276 -13004 39322 4 VSS
port 42 nsew
rlabel metal1 s -13204 40340 -13004 40386 4 VSS
port 42 nsew
rlabel metal1 s -13204 40649 -13004 40695 4 VSS
port 42 nsew
rlabel metal1 s -15395 41511 -15361 41512 4 VSS
port 42 nsew
rlabel metal1 s -15480 41512 -15361 41580 4 VSS
port 42 nsew
rlabel metal1 s -12453 41738 -12406 41881 4 VSS
port 42 nsew
rlabel metal1 s -12584 41612 -12537 41756 4 VSS
port 42 nsew
rlabel metal1 s -15480 41580 -13984 41641 4 VSS
port 42 nsew
rlabel metal1 s -15480 41641 -15362 41642 4 VSS
port 42 nsew
rlabel metal1 s -15785 41671 -15661 41692 4 VSS
port 42 nsew
rlabel metal1 s -15785 41692 -15489 41694 4 VSS
port 42 nsew
rlabel metal1 s -12317 41898 -12269 42046 4 VSS
port 42 nsew
rlabel metal1 s -12313 42046 -12277 42169 4 VSS
port 42 nsew
rlabel metal1 s -12313 42169 -6569 42205 4 VSS
port 42 nsew
rlabel metal1 s -12452 41881 -12424 42336 4 VSS
port 42 nsew
rlabel metal1 s -12452 42336 -6430 42364 4 VSS
port 42 nsew
rlabel metal1 s -12572 41756 -12544 42498 4 VSS
port 42 nsew
rlabel metal1 s -15785 41694 -13980 41758 4 VSS
port 42 nsew
rlabel metal1 s -15785 41758 -15662 41794 4 VSS
port 42 nsew
rlabel metal1 s -16152 41822 -16029 41839 4 VSS
port 42 nsew
rlabel metal1 s -16152 41839 -13944 41899 4 VSS
port 42 nsew
rlabel metal1 s -16152 41899 -16029 41945 4 VSS
port 42 nsew
rlabel metal1 s -12572 42498 -6310 42526 4 VSS
port 42 nsew
rlabel metal1 s -12609 43879 -12509 43925 4 VSS
port 42 nsew
rlabel metal1 s -1993 44054 -862 44070 4 VSS
port 42 nsew
rlabel metal1 s -4820 44054 -3786 44102 4 VSS
port 42 nsew
rlabel metal1 s -12609 44075 -12509 44121 4 VSS
port 42 nsew
rlabel metal1 s -12729 44152 -12669 44159 4 VSS
port 42 nsew
rlabel metal1 s -12998 44139 -12938 44159 4 VSS
port 42 nsew
rlabel metal1 s -12998 44159 -12669 44254 4 VSS
port 42 nsew
rlabel metal1 s -12609 44271 -12509 44317 4 VSS
port 42 nsew
rlabel metal1 s -12729 44254 -12669 44289 4 VSS
port 42 nsew
rlabel metal1 s -12998 44254 -12938 44271 4 VSS
port 42 nsew
rlabel metal1 s -12609 44761 -12509 44807 4 VSS
port 42 nsew
rlabel metal1 s -12609 44957 -12509 45003 4 VSS
port 42 nsew
rlabel metal1 s -12609 45153 -12509 45199 4 VSS
port 42 nsew
rlabel metal1 s -13267 45765 -13167 45811 4 VSS
port 42 nsew
rlabel metal1 s -13267 45961 -13167 46007 4 VSS
port 42 nsew
rlabel metal1 s -13267 46157 -13167 46203 4 VSS
port 42 nsew
rlabel metal1 s -12609 46504 -12509 46550 4 VSS
port 42 nsew
rlabel metal1 s -13267 46602 -13167 46648 4 VSS
port 42 nsew
rlabel metal1 s -12609 46700 -12509 46746 4 VSS
port 42 nsew
rlabel metal1 s -12730 46779 -12670 46803 4 VSS
port 42 nsew
rlabel metal1 s -12998 46772 -12938 46803 4 VSS
port 42 nsew
rlabel metal1 s -12609 46896 -12509 46942 4 VSS
port 42 nsew
rlabel metal1 s -12998 46803 -12670 46898 4 VSS
port 42 nsew
rlabel metal1 s -13267 46798 -13167 46844 4 VSS
port 42 nsew
rlabel metal1 s -12730 46898 -12670 46916 4 VSS
port 42 nsew
rlabel metal1 s -12998 46898 -12938 46909 4 VSS
port 42 nsew
rlabel metal1 s -13267 46994 -13167 47040 4 VSS
port 42 nsew
rlabel metal1 s -12609 47461 -12509 47507 4 VSS
port 42 nsew
rlabel metal1 s -12609 47657 -12509 47703 4 VSS
port 42 nsew
rlabel metal1 s -12609 47853 -12509 47899 4 VSS
port 42 nsew
rlabel metal1 s -13267 48465 -13167 48511 4 VSS
port 42 nsew
rlabel metal1 s -13267 48661 -13167 48707 4 VSS
port 42 nsew
rlabel metal1 s -13267 48857 -13167 48903 4 VSS
port 42 nsew
rlabel metal1 s -12609 49204 -12509 49250 4 VSS
port 42 nsew
rlabel metal1 s -13267 49302 -13167 49348 4 VSS
port 42 nsew
rlabel metal1 s -12726 49383 -12666 49396 4 VSS
port 42 nsew
rlabel metal1 s -13004 49369 -12944 49396 4 VSS
port 42 nsew
rlabel metal1 s -12609 49400 -12509 49446 4 VSS
port 42 nsew
rlabel metal1 s -13004 49396 -12666 49491 4 VSS
port 42 nsew
rlabel metal1 s -12726 49491 -12666 49515 4 VSS
port 42 nsew
rlabel metal1 s -13004 49491 -12944 49506 4 VSS
port 42 nsew
rlabel metal1 s -13267 49498 -13167 49544 4 VSS
port 42 nsew
rlabel metal1 s -12609 49596 -12509 49642 4 VSS
port 42 nsew
rlabel metal1 s -13267 49694 -13167 49740 4 VSS
port 42 nsew
rlabel metal1 s -8007 50784 -7807 50830 4 VSS
port 42 nsew
rlabel metal1 s -10625 50779 -10425 50825 4 VSS
port 42 nsew
rlabel metal1 s -8007 50980 -7807 51026 4 VSS
port 42 nsew
rlabel metal1 s -10625 50975 -10425 51021 4 VSS
port 42 nsew
rlabel metal1 s -10625 51725 -10425 51771 4 VSS
port 42 nsew
rlabel metal1 s -10625 51921 -10425 51967 4 VSS
port 42 nsew
rlabel metal1 s -8711 52007 -8611 52053 4 VSS
port 42 nsew
rlabel metal1 s -8711 52203 -8611 52249 4 VSS
port 42 nsew
rlabel metal1 s -8282 52267 -8222 52287 4 VSS
port 42 nsew
rlabel metal1 s -8551 52280 -8491 52287 4 VSS
port 42 nsew
rlabel metal1 s -8551 52287 -8222 52382 4 VSS
port 42 nsew
rlabel metal1 s -8282 52382 -8222 52399 4 VSS
port 42 nsew
rlabel metal1 s -8551 52382 -8491 52417 4 VSS
port 42 nsew
rlabel metal1 s -8711 52399 -8611 52445 4 VSS
port 42 nsew
rlabel metal1 s -10744 52641 -10444 52687 4 VSS
port 42 nsew
rlabel metal1 s -8711 52889 -8611 52935 4 VSS
port 42 nsew
rlabel metal1 s -8711 53085 -8611 53131 4 VSS
port 42 nsew
rlabel metal1 s -8711 53281 -8611 53327 4 VSS
port 42 nsew
rlabel metal1 s -10643 53673 -10443 53719 4 VSS
port 42 nsew
rlabel metal1 s -8053 53893 -7953 53939 4 VSS
port 42 nsew
rlabel metal1 s -8053 54089 -7953 54135 4 VSS
port 42 nsew
rlabel metal1 s -8053 54285 -7953 54331 4 VSS
port 42 nsew
rlabel metal1 s -10964 54402 -10864 54448 4 VSS
port 42 nsew
rlabel metal1 s -10497 54452 -10297 54498 4 VSS
port 42 nsew
rlabel metal1 s -8711 54632 -8611 54678 4 VSS
port 42 nsew
rlabel metal1 s -10964 54598 -10864 54644 4 VSS
port 42 nsew
rlabel metal1 s -8053 54730 -7953 54776 4 VSS
port 42 nsew
rlabel metal1 s -8711 54828 -8611 54874 4 VSS
port 42 nsew
rlabel metal1 s -10964 54794 -10864 54840 4 VSS
port 42 nsew
rlabel metal1 s -8053 54926 -7953 54972 4 VSS
port 42 nsew
rlabel metal1 s -8282 54900 -8222 54931 4 VSS
port 42 nsew
rlabel metal1 s -8550 54907 -8490 54931 4 VSS
port 42 nsew
rlabel metal1 s -8550 54931 -8222 55026 4 VSS
port 42 nsew
rlabel metal1 s -8282 55026 -8222 55037 4 VSS
port 42 nsew
rlabel metal1 s -8550 55026 -8490 55044 4 VSS
port 42 nsew
rlabel metal1 s -8711 55024 -8611 55070 4 VSS
port 42 nsew
rlabel metal1 s -8053 55122 -7953 55168 4 VSS
port 42 nsew
rlabel metal1 s -10388 55282 -9688 55328 4 VSS
port 42 nsew
rlabel metal1 s -8711 55589 -8611 55635 4 VSS
port 42 nsew
rlabel metal1 s -10388 55682 -9688 55728 4 VSS
port 42 nsew
rlabel metal1 s -8711 55785 -8611 55831 4 VSS
port 42 nsew
rlabel metal1 s -8711 55981 -8611 56027 4 VSS
port 42 nsew
rlabel metal1 s -10388 56282 -9688 56328 4 VSS
port 42 nsew
rlabel metal1 s -8053 56593 -7953 56639 4 VSS
port 42 nsew
rlabel metal1 s -10388 56682 -9688 56728 4 VSS
port 42 nsew
rlabel metal1 s -8053 56789 -7953 56835 4 VSS
port 42 nsew
rlabel metal1 s -8053 56985 -7953 57031 4 VSS
port 42 nsew
rlabel metal1 s -10388 57282 -9688 57328 4 VSS
port 42 nsew
rlabel metal1 s -8711 57332 -8611 57378 4 VSS
port 42 nsew
rlabel metal1 s -8053 57430 -7953 57476 4 VSS
port 42 nsew
rlabel metal1 s -8276 57497 -8216 57524 4 VSS
port 42 nsew
rlabel metal1 s -8554 57511 -8494 57524 4 VSS
port 42 nsew
rlabel metal1 s -8554 57524 -8216 57619 4 VSS
port 42 nsew
rlabel metal1 s -8711 57528 -8611 57574 4 VSS
port 42 nsew
rlabel metal1 s -8053 57626 -7953 57672 4 VSS
port 42 nsew
rlabel metal1 s -8276 57619 -8216 57634 4 VSS
port 42 nsew
rlabel metal1 s -8554 57619 -8494 57643 4 VSS
port 42 nsew
rlabel metal1 s -8711 57724 -8611 57770 4 VSS
port 42 nsew
rlabel metal1 s -10388 57682 -9688 57728 4 VSS
port 42 nsew
rlabel metal1 s -8053 57822 -7953 57868 4 VSS
port 42 nsew
rlabel metal1 s -7090 60363 -6890 60409 4 VSS
port 42 nsew
rlabel metal1 s -8986 60337 -8686 60383 4 VSS
port 42 nsew
rlabel metal1 s -10543 60355 -10343 60401 4 VSS
port 42 nsew
rlabel metal1 s -12439 60329 -12139 60375 4 VSS
port 42 nsew
rlabel metal1 s -7090 60559 -6890 60605 4 VSS
port 42 nsew
rlabel metal1 s -10543 60551 -10343 60597 4 VSS
port 42 nsew
rlabel metal1 s -8479 60946 -8379 60992 4 VSS
port 42 nsew
rlabel metal1 s -11932 60938 -11832 60984 4 VSS
port 42 nsew
rlabel metal1 s -8479 61142 -8379 61188 4 VSS
port 42 nsew
rlabel metal1 s -11932 61134 -11832 61180 4 VSS
port 42 nsew
rlabel metal1 s -7012 61336 -6712 61382 4 VSS
port 42 nsew
rlabel metal1 s -10465 61328 -10165 61374 4 VSS
port 42 nsew
rlabel metal1 s -9272 61784 -8972 61830 4 VSS
port 42 nsew
rlabel metal1 s -12725 61776 -12425 61822 4 VSS
port 42 nsew
rlabel metal1 s -7319 61945 -7219 61991 4 VSS
port 42 nsew
rlabel metal1 s -9272 61980 -8972 62026 4 VSS
port 42 nsew
rlabel metal1 s -10772 61937 -10672 61983 4 VSS
port 42 nsew
rlabel metal1 s -12725 61972 -12425 62018 4 VSS
port 42 nsew
rlabel metal1 s -7319 62141 -7219 62187 4 VSS
port 42 nsew
rlabel metal1 s -10772 62133 -10672 62179 4 VSS
port 42 nsew
rlabel metal1 s -9272 62222 -8972 62268 4 VSS
port 42 nsew
rlabel metal1 s -12725 62214 -12425 62260 4 VSS
port 42 nsew
rlabel metal1 s -7184 62332 -7071 62927 4 VSS
port 42 nsew
rlabel metal1 s -9493 62363 -9380 62553 4 VSS
port 42 nsew
rlabel metal1 s -10637 62324 -10524 62553 4 VSS
port 42 nsew
rlabel metal1 s -10637 62553 -9379 62666 4 VSS
port 42 nsew
rlabel metal1 s -9493 62666 -9380 62927 4 VSS
port 42 nsew
rlabel metal1 s -9493 62927 -7071 63040 4 VSS
port 42 nsew
rlabel metal1 s -10637 62666 -10524 62919 4 VSS
port 42 nsew
rlabel metal1 s -12946 62355 -12833 62359 4 VSS
port 42 nsew
rlabel metal1 s -12977 62359 -12833 62919 4 VSS
port 42 nsew
rlabel metal1 s -12977 62919 -10524 63032 4 VSS
port 42 nsew
rlabel metal1 s -9214 63678 -8914 63724 4 VSS
port 42 nsew
rlabel metal1 s -10574 64023 -10374 64069 4 VSS
port 42 nsew
rlabel metal1 s -12470 63997 -12170 64043 4 VSS
port 42 nsew
rlabel metal1 s -10574 64219 -10374 64265 4 VSS
port 42 nsew
rlabel metal1 s -9214 64469 -8714 64515 4 VSS
port 42 nsew
rlabel metal1 s -9214 64599 -8714 64645 4 VSS
port 42 nsew
rlabel metal1 s -11963 64606 -11863 64652 4 VSS
port 42 nsew
rlabel metal1 s -11963 64802 -11863 64848 4 VSS
port 42 nsew
rlabel metal1 s -9214 64925 -8914 64971 4 VSS
port 42 nsew
rlabel metal1 s -10496 64996 -10196 65042 4 VSS
port 42 nsew
rlabel metal1 s -12756 65444 -12456 65490 4 VSS
port 42 nsew
rlabel metal1 s -10803 65605 -10703 65651 4 VSS
port 42 nsew
rlabel metal1 s -12756 65640 -12456 65686 4 VSS
port 42 nsew
rlabel metal1 s -10803 65801 -10703 65847 4 VSS
port 42 nsew
rlabel metal1 s -12756 65882 -12456 65928 4 VSS
port 42 nsew
rlabel metal1 s -10668 65992 -10555 66587 4 VSS
port 42 nsew
rlabel metal1 s -12977 63032 -12864 66587 4 VSS
port 42 nsew
rlabel metal1 s -12977 66587 -10555 66700 4 VSS
port 42 nsew
rlabel metal1 s -7101 68803 -6901 68849 4 VSS
port 42 nsew
rlabel metal1 s -8997 68777 -8697 68823 4 VSS
port 42 nsew
rlabel metal1 s -10554 68795 -10354 68841 4 VSS
port 42 nsew
rlabel metal1 s -12450 68769 -12150 68815 4 VSS
port 42 nsew
rlabel metal1 s -7101 68999 -6901 69045 4 VSS
port 42 nsew
rlabel metal1 s -10554 68991 -10354 69037 4 VSS
port 42 nsew
rlabel metal1 s -8490 69386 -8390 69432 4 VSS
port 42 nsew
rlabel metal1 s -11943 69378 -11843 69424 4 VSS
port 42 nsew
rlabel metal1 s -8490 69582 -8390 69628 4 VSS
port 42 nsew
rlabel metal1 s -11943 69574 -11843 69620 4 VSS
port 42 nsew
rlabel metal1 s -7023 69776 -6723 69822 4 VSS
port 42 nsew
rlabel metal1 s -10476 69768 -10176 69814 4 VSS
port 42 nsew
rlabel metal1 s -9283 70224 -8983 70270 4 VSS
port 42 nsew
rlabel metal1 s -12736 70216 -12436 70262 4 VSS
port 42 nsew
rlabel metal1 s -7330 70385 -7230 70431 4 VSS
port 42 nsew
rlabel metal1 s -9283 70420 -8983 70466 4 VSS
port 42 nsew
rlabel metal1 s -10783 70377 -10683 70423 4 VSS
port 42 nsew
rlabel metal1 s -12736 70412 -12436 70458 4 VSS
port 42 nsew
rlabel metal1 s -7330 70581 -7230 70627 4 VSS
port 42 nsew
rlabel metal1 s -10783 70573 -10683 70619 4 VSS
port 42 nsew
rlabel metal1 s -9283 70662 -8983 70708 4 VSS
port 42 nsew
rlabel metal1 s -12736 70654 -12436 70700 4 VSS
port 42 nsew
rlabel metal1 s -7195 70772 -7082 71367 4 VSS
port 42 nsew
rlabel metal1 s -9504 70803 -9391 70993 4 VSS
port 42 nsew
rlabel metal1 s -10648 70764 -10535 70993 4 VSS
port 42 nsew
rlabel metal1 s -10648 70993 -9390 71106 4 VSS
port 42 nsew
rlabel metal1 s -9504 71106 -9391 71367 4 VSS
port 42 nsew
rlabel metal1 s -9504 71367 -7082 71480 4 VSS
port 42 nsew
rlabel metal1 s -10648 71106 -10535 71359 4 VSS
port 42 nsew
rlabel metal1 s -12957 70795 -12844 70799 4 VSS
port 42 nsew
rlabel metal1 s -12988 70799 -12844 71359 4 VSS
port 42 nsew
rlabel metal1 s -12988 71359 -10535 71472 4 VSS
port 42 nsew
rlabel metal1 s -9225 72118 -8925 72164 4 VSS
port 42 nsew
rlabel metal1 s -10585 72463 -10385 72509 4 VSS
port 42 nsew
rlabel metal1 s -12481 72437 -12181 72483 4 VSS
port 42 nsew
rlabel metal1 s -10585 72659 -10385 72705 4 VSS
port 42 nsew
rlabel metal1 s -9225 72909 -8725 72955 4 VSS
port 42 nsew
rlabel metal1 s -9225 73039 -8725 73085 4 VSS
port 42 nsew
rlabel metal1 s -11974 73046 -11874 73092 4 VSS
port 42 nsew
rlabel metal1 s -11974 73242 -11874 73288 4 VSS
port 42 nsew
rlabel metal1 s -9225 73365 -8925 73411 4 VSS
port 42 nsew
rlabel metal1 s -10507 73436 -10207 73482 4 VSS
port 42 nsew
rlabel metal1 s -12767 73884 -12467 73930 4 VSS
port 42 nsew
rlabel metal1 s -10814 74045 -10714 74091 4 VSS
port 42 nsew
rlabel metal1 s -12767 74080 -12467 74126 4 VSS
port 42 nsew
rlabel metal1 s -10814 74241 -10714 74287 4 VSS
port 42 nsew
rlabel metal1 s -12767 74322 -12467 74368 4 VSS
port 42 nsew
rlabel metal1 s -10679 74432 -10566 75027 4 VSS
port 42 nsew
rlabel metal1 s -12988 71472 -12875 75027 4 VSS
port 42 nsew
rlabel metal1 s -12988 75027 -10566 75140 4 VSS
port 42 nsew
rlabel metal1 s -7140 77666 -6940 77712 4 VSS
port 42 nsew
rlabel metal1 s -9036 77640 -8736 77686 4 VSS
port 42 nsew
rlabel metal1 s -10593 77658 -10393 77704 4 VSS
port 42 nsew
rlabel metal1 s -12489 77632 -12189 77678 4 VSS
port 42 nsew
rlabel metal1 s -7140 77862 -6940 77908 4 VSS
port 42 nsew
rlabel metal1 s -10593 77854 -10393 77900 4 VSS
port 42 nsew
rlabel metal1 s -8529 78249 -8429 78295 4 VSS
port 42 nsew
rlabel metal1 s -11982 78241 -11882 78287 4 VSS
port 42 nsew
rlabel metal1 s -8529 78445 -8429 78491 4 VSS
port 42 nsew
rlabel metal1 s -11982 78437 -11882 78483 4 VSS
port 42 nsew
rlabel metal1 s -7062 78639 -6762 78685 4 VSS
port 42 nsew
rlabel metal1 s -10515 78631 -10215 78677 4 VSS
port 42 nsew
rlabel metal1 s -9322 79087 -9022 79133 4 VSS
port 42 nsew
rlabel metal1 s -12775 79079 -12475 79125 4 VSS
port 42 nsew
rlabel metal1 s -7369 79248 -7269 79294 4 VSS
port 42 nsew
rlabel metal1 s -9322 79283 -9022 79329 4 VSS
port 42 nsew
rlabel metal1 s -10822 79240 -10722 79286 4 VSS
port 42 nsew
rlabel metal1 s -12775 79275 -12475 79321 4 VSS
port 42 nsew
rlabel metal1 s -7369 79444 -7269 79490 4 VSS
port 42 nsew
rlabel metal1 s -10822 79436 -10722 79482 4 VSS
port 42 nsew
rlabel metal1 s -9322 79525 -9022 79571 4 VSS
port 42 nsew
rlabel metal1 s -12775 79517 -12475 79563 4 VSS
port 42 nsew
rlabel metal1 s -7234 79635 -7121 80230 4 VSS
port 42 nsew
rlabel metal1 s -9543 79666 -9430 79856 4 VSS
port 42 nsew
rlabel metal1 s -10687 79627 -10574 79856 4 VSS
port 42 nsew
rlabel metal1 s -10687 79856 -9429 79969 4 VSS
port 42 nsew
rlabel metal1 s -9543 79969 -9430 80230 4 VSS
port 42 nsew
rlabel metal1 s -9543 80230 -7121 80343 4 VSS
port 42 nsew
rlabel metal1 s -10687 79969 -10574 80222 4 VSS
port 42 nsew
rlabel metal1 s -12996 79658 -12883 79662 4 VSS
port 42 nsew
rlabel metal1 s -13027 79662 -12883 80222 4 VSS
port 42 nsew
rlabel metal1 s -13027 80222 -10574 80335 4 VSS
port 42 nsew
rlabel metal1 s -9264 80981 -8964 81027 4 VSS
port 42 nsew
rlabel metal1 s -10624 81326 -10424 81372 4 VSS
port 42 nsew
rlabel metal1 s -12520 81300 -12220 81346 4 VSS
port 42 nsew
rlabel metal1 s -10624 81522 -10424 81568 4 VSS
port 42 nsew
rlabel metal1 s -9264 81772 -8764 81818 4 VSS
port 42 nsew
rlabel metal1 s -9264 81902 -8764 81948 4 VSS
port 42 nsew
rlabel metal1 s -12013 81909 -11913 81955 4 VSS
port 42 nsew
rlabel metal1 s -12013 82105 -11913 82151 4 VSS
port 42 nsew
rlabel metal1 s -9264 82228 -8964 82274 4 VSS
port 42 nsew
rlabel metal1 s -10546 82299 -10246 82345 4 VSS
port 42 nsew
rlabel metal1 s -12806 82747 -12506 82793 4 VSS
port 42 nsew
rlabel metal1 s -10853 82908 -10753 82954 4 VSS
port 42 nsew
rlabel metal1 s -12806 82943 -12506 82989 4 VSS
port 42 nsew
rlabel metal1 s -10853 83104 -10753 83150 4 VSS
port 42 nsew
rlabel metal1 s -12806 83185 -12506 83231 4 VSS
port 42 nsew
rlabel metal1 s -10718 83295 -10605 83890 4 VSS
port 42 nsew
rlabel metal1 s -13027 80335 -12914 83890 4 VSS
port 42 nsew
rlabel metal1 s -13027 83890 -10605 84003 4 VSS
port 42 nsew
rlabel metal1 s -7106 86864 -6906 86910 4 VSS
port 42 nsew
rlabel metal1 s -9002 86838 -8702 86884 4 VSS
port 42 nsew
rlabel metal1 s -10559 86856 -10359 86902 4 VSS
port 42 nsew
rlabel metal1 s -12455 86830 -12155 86876 4 VSS
port 42 nsew
rlabel metal1 s -7106 87060 -6906 87106 4 VSS
port 42 nsew
rlabel metal1 s -10559 87052 -10359 87098 4 VSS
port 42 nsew
rlabel metal1 s -8495 87447 -8395 87493 4 VSS
port 42 nsew
rlabel metal1 s -11948 87439 -11848 87485 4 VSS
port 42 nsew
rlabel metal1 s -8495 87643 -8395 87689 4 VSS
port 42 nsew
rlabel metal1 s -11948 87635 -11848 87681 4 VSS
port 42 nsew
rlabel metal1 s -7028 87837 -6728 87883 4 VSS
port 42 nsew
rlabel metal1 s -10481 87829 -10181 87875 4 VSS
port 42 nsew
rlabel metal1 s -9288 88285 -8988 88331 4 VSS
port 42 nsew
rlabel metal1 s -12741 88277 -12441 88323 4 VSS
port 42 nsew
rlabel metal1 s -7335 88446 -7235 88492 4 VSS
port 42 nsew
rlabel metal1 s -9288 88481 -8988 88527 4 VSS
port 42 nsew
rlabel metal1 s -10788 88438 -10688 88484 4 VSS
port 42 nsew
rlabel metal1 s -12741 88473 -12441 88519 4 VSS
port 42 nsew
rlabel metal1 s -7335 88642 -7235 88688 4 VSS
port 42 nsew
rlabel metal1 s -10788 88634 -10688 88680 4 VSS
port 42 nsew
rlabel metal1 s -9288 88723 -8988 88769 4 VSS
port 42 nsew
rlabel metal1 s -12741 88715 -12441 88761 4 VSS
port 42 nsew
rlabel metal1 s -7200 88833 -7087 89428 4 VSS
port 42 nsew
rlabel metal1 s -9509 88864 -9396 89054 4 VSS
port 42 nsew
rlabel metal1 s -10653 88825 -10540 89054 4 VSS
port 42 nsew
rlabel metal1 s -10653 89054 -9395 89167 4 VSS
port 42 nsew
rlabel metal1 s -9509 89167 -9396 89428 4 VSS
port 42 nsew
rlabel metal1 s -9509 89428 -7087 89541 4 VSS
port 42 nsew
rlabel metal1 s -10653 89167 -10540 89420 4 VSS
port 42 nsew
rlabel metal1 s -12962 88856 -12849 88860 4 VSS
port 42 nsew
rlabel metal1 s -12993 88860 -12849 89420 4 VSS
port 42 nsew
rlabel metal1 s -12993 89420 -10540 89533 4 VSS
port 42 nsew
rlabel metal1 s -9230 90179 -8930 90225 4 VSS
port 42 nsew
rlabel metal1 s -10590 90524 -10390 90570 4 VSS
port 42 nsew
rlabel metal1 s -12486 90498 -12186 90544 4 VSS
port 42 nsew
rlabel metal1 s -10590 90720 -10390 90766 4 VSS
port 42 nsew
rlabel metal1 s -9230 90970 -8730 91016 4 VSS
port 42 nsew
rlabel metal1 s -9230 91100 -8730 91146 4 VSS
port 42 nsew
rlabel metal1 s -11979 91107 -11879 91153 4 VSS
port 42 nsew
rlabel metal1 s -11979 91303 -11879 91349 4 VSS
port 42 nsew
rlabel metal1 s -9230 91426 -8930 91472 4 VSS
port 42 nsew
rlabel metal1 s -10512 91497 -10212 91543 4 VSS
port 42 nsew
rlabel metal1 s -12772 91945 -12472 91991 4 VSS
port 42 nsew
rlabel metal1 s -10819 92106 -10719 92152 4 VSS
port 42 nsew
rlabel metal1 s -12772 92141 -12472 92187 4 VSS
port 42 nsew
rlabel metal1 s -10819 92302 -10719 92348 4 VSS
port 42 nsew
rlabel metal1 s -12772 92383 -12472 92429 4 VSS
port 42 nsew
rlabel metal1 s -10684 92493 -10571 93088 4 VSS
port 42 nsew
rlabel metal1 s -12993 89533 -12880 93088 4 VSS
port 42 nsew
rlabel metal1 s -12993 93088 -10571 93201 4 VSS
port 42 nsew
rlabel metal1 s -7040 95618 -6840 95664 4 VSS
port 42 nsew
rlabel metal1 s -8936 95592 -8636 95638 4 VSS
port 42 nsew
rlabel metal1 s -10493 95610 -10293 95656 4 VSS
port 42 nsew
rlabel metal1 s -12389 95584 -12089 95630 4 VSS
port 42 nsew
rlabel metal1 s -7040 95814 -6840 95860 4 VSS
port 42 nsew
rlabel metal1 s -10493 95806 -10293 95852 4 VSS
port 42 nsew
rlabel metal1 s -8429 96201 -8329 96247 4 VSS
port 42 nsew
rlabel metal1 s -11882 96193 -11782 96239 4 VSS
port 42 nsew
rlabel metal1 s -8429 96397 -8329 96443 4 VSS
port 42 nsew
rlabel metal1 s -11882 96389 -11782 96435 4 VSS
port 42 nsew
rlabel metal1 s -6962 96591 -6662 96637 4 VSS
port 42 nsew
rlabel metal1 s -10415 96583 -10115 96629 4 VSS
port 42 nsew
rlabel metal1 s -9222 97039 -8922 97085 4 VSS
port 42 nsew
rlabel metal1 s -12675 97031 -12375 97077 4 VSS
port 42 nsew
rlabel metal1 s -7269 97200 -7169 97246 4 VSS
port 42 nsew
rlabel metal1 s -9222 97235 -8922 97281 4 VSS
port 42 nsew
rlabel metal1 s -10722 97192 -10622 97238 4 VSS
port 42 nsew
rlabel metal1 s -12675 97227 -12375 97273 4 VSS
port 42 nsew
rlabel metal1 s -7269 97396 -7169 97442 4 VSS
port 42 nsew
rlabel metal1 s -10722 97388 -10622 97434 4 VSS
port 42 nsew
rlabel metal1 s -9222 97477 -8922 97523 4 VSS
port 42 nsew
rlabel metal1 s -12675 97469 -12375 97515 4 VSS
port 42 nsew
rlabel metal1 s -7134 97587 -7021 98182 4 VSS
port 42 nsew
rlabel metal1 s -9443 97618 -9330 97808 4 VSS
port 42 nsew
rlabel metal1 s -10587 97579 -10474 97808 4 VSS
port 42 nsew
rlabel metal1 s -10587 97808 -9329 97921 4 VSS
port 42 nsew
rlabel metal1 s -9443 97921 -9330 98182 4 VSS
port 42 nsew
rlabel metal1 s -9443 98182 -7021 98295 4 VSS
port 42 nsew
rlabel metal1 s -10587 97921 -10474 98174 4 VSS
port 42 nsew
rlabel metal1 s -12896 97610 -12783 97614 4 VSS
port 42 nsew
rlabel metal1 s -12927 97614 -12783 98174 4 VSS
port 42 nsew
rlabel metal1 s -12927 98174 -10474 98287 4 VSS
port 42 nsew
rlabel metal1 s -9164 98933 -8864 98979 4 VSS
port 42 nsew
rlabel metal1 s -10524 99278 -10324 99324 4 VSS
port 42 nsew
rlabel metal1 s -12420 99252 -12120 99298 4 VSS
port 42 nsew
rlabel metal1 s -10524 99474 -10324 99520 4 VSS
port 42 nsew
rlabel metal1 s -9164 99724 -8664 99770 4 VSS
port 42 nsew
rlabel metal1 s -9164 99854 -8664 99900 4 VSS
port 42 nsew
rlabel metal1 s -11913 99861 -11813 99907 4 VSS
port 42 nsew
rlabel metal1 s -11913 100057 -11813 100103 4 VSS
port 42 nsew
rlabel metal1 s -9164 100180 -8864 100226 4 VSS
port 42 nsew
rlabel metal1 s -10446 100251 -10146 100297 4 VSS
port 42 nsew
rlabel metal1 s -12706 100699 -12406 100745 4 VSS
port 42 nsew
rlabel metal1 s -10753 100860 -10653 100906 4 VSS
port 42 nsew
rlabel metal1 s -12706 100895 -12406 100941 4 VSS
port 42 nsew
rlabel metal1 s -10753 101056 -10653 101102 4 VSS
port 42 nsew
rlabel metal1 s -12706 101137 -12406 101183 4 VSS
port 42 nsew
rlabel metal1 s -10618 101247 -10505 101842 4 VSS
port 42 nsew
rlabel metal1 s -12927 98287 -12814 101842 4 VSS
port 42 nsew
rlabel metal1 s -12927 101842 -10505 101955 4 VSS
port 42 nsew
rlabel metal1 s -7023 104771 -6823 104817 4 VSS
port 42 nsew
rlabel metal1 s -8919 104745 -8619 104791 4 VSS
port 42 nsew
rlabel metal1 s -10476 104763 -10276 104809 4 VSS
port 42 nsew
rlabel metal1 s -12372 104737 -12072 104783 4 VSS
port 42 nsew
rlabel metal1 s -7023 104967 -6823 105013 4 VSS
port 42 nsew
rlabel metal1 s -10476 104959 -10276 105005 4 VSS
port 42 nsew
rlabel metal1 s -8412 105354 -8312 105400 4 VSS
port 42 nsew
rlabel metal1 s -11865 105346 -11765 105392 4 VSS
port 42 nsew
rlabel metal1 s -8412 105550 -8312 105596 4 VSS
port 42 nsew
rlabel metal1 s -11865 105542 -11765 105588 4 VSS
port 42 nsew
rlabel metal1 s -6945 105744 -6645 105790 4 VSS
port 42 nsew
rlabel metal1 s -10398 105736 -10098 105782 4 VSS
port 42 nsew
rlabel metal1 s -9205 106192 -8905 106238 4 VSS
port 42 nsew
rlabel metal1 s -12658 106184 -12358 106230 4 VSS
port 42 nsew
rlabel metal1 s -7252 106353 -7152 106399 4 VSS
port 42 nsew
rlabel metal1 s -9205 106388 -8905 106434 4 VSS
port 42 nsew
rlabel metal1 s -10705 106345 -10605 106391 4 VSS
port 42 nsew
rlabel metal1 s -12658 106380 -12358 106426 4 VSS
port 42 nsew
rlabel metal1 s -7252 106549 -7152 106595 4 VSS
port 42 nsew
rlabel metal1 s -10705 106541 -10605 106587 4 VSS
port 42 nsew
rlabel metal1 s -9205 106630 -8905 106676 4 VSS
port 42 nsew
rlabel metal1 s -12658 106622 -12358 106668 4 VSS
port 42 nsew
rlabel metal1 s -7117 106740 -7004 107335 4 VSS
port 42 nsew
rlabel metal1 s -9426 106771 -9313 106961 4 VSS
port 42 nsew
rlabel metal1 s -10570 106732 -10457 106961 4 VSS
port 42 nsew
rlabel metal1 s -10570 106961 -9312 107074 4 VSS
port 42 nsew
rlabel metal1 s -9426 107074 -9313 107335 4 VSS
port 42 nsew
rlabel metal1 s -9426 107335 -7004 107448 4 VSS
port 42 nsew
rlabel metal1 s -10570 107074 -10457 107327 4 VSS
port 42 nsew
rlabel metal1 s -12879 106763 -12766 106767 4 VSS
port 42 nsew
rlabel metal1 s -12910 106767 -12766 107327 4 VSS
port 42 nsew
rlabel metal1 s -12910 107327 -10457 107440 4 VSS
port 42 nsew
rlabel metal1 s -9147 108086 -8847 108132 4 VSS
port 42 nsew
rlabel metal1 s -10507 108431 -10307 108477 4 VSS
port 42 nsew
rlabel metal1 s -12403 108405 -12103 108451 4 VSS
port 42 nsew
rlabel metal1 s -10507 108627 -10307 108673 4 VSS
port 42 nsew
rlabel metal1 s -9147 108877 -8647 108923 4 VSS
port 42 nsew
rlabel metal1 s -9147 109007 -8647 109053 4 VSS
port 42 nsew
rlabel metal1 s -11896 109014 -11796 109060 4 VSS
port 42 nsew
rlabel metal1 s -11896 109210 -11796 109256 4 VSS
port 42 nsew
rlabel metal1 s -9147 109333 -8847 109379 4 VSS
port 42 nsew
rlabel metal1 s -10429 109404 -10129 109450 4 VSS
port 42 nsew
rlabel metal1 s -12689 109852 -12389 109898 4 VSS
port 42 nsew
rlabel metal1 s -10736 110013 -10636 110059 4 VSS
port 42 nsew
rlabel metal1 s -12689 110048 -12389 110094 4 VSS
port 42 nsew
rlabel metal1 s -10736 110209 -10636 110255 4 VSS
port 42 nsew
rlabel metal1 s -12689 110290 -12389 110336 4 VSS
port 42 nsew
rlabel metal1 s -10601 110400 -10488 110995 4 VSS
port 42 nsew
rlabel metal1 s -12910 107440 -12797 110995 4 VSS
port 42 nsew
rlabel metal1 s -12910 110995 -10488 111108 4 VSS
port 42 nsew
rlabel metal1 s -6985 114135 -6785 114181 4 VSS
port 42 nsew
rlabel metal1 s -8881 114109 -8581 114155 4 VSS
port 42 nsew
rlabel metal1 s -10438 114127 -10238 114173 4 VSS
port 42 nsew
rlabel metal1 s -12334 114101 -12034 114147 4 VSS
port 42 nsew
rlabel metal1 s -6985 114331 -6785 114377 4 VSS
port 42 nsew
rlabel metal1 s -10438 114323 -10238 114369 4 VSS
port 42 nsew
rlabel metal1 s -8374 114718 -8274 114764 4 VSS
port 42 nsew
rlabel metal1 s -11827 114710 -11727 114756 4 VSS
port 42 nsew
rlabel metal1 s -8374 114914 -8274 114960 4 VSS
port 42 nsew
rlabel metal1 s -11827 114906 -11727 114952 4 VSS
port 42 nsew
rlabel metal1 s -6907 115108 -6607 115154 4 VSS
port 42 nsew
rlabel metal1 s -10360 115100 -10060 115146 4 VSS
port 42 nsew
rlabel metal1 s -9167 115556 -8867 115602 4 VSS
port 42 nsew
rlabel metal1 s -12620 115548 -12320 115594 4 VSS
port 42 nsew
rlabel metal1 s -7214 115717 -7114 115763 4 VSS
port 42 nsew
rlabel metal1 s -9167 115752 -8867 115798 4 VSS
port 42 nsew
rlabel metal1 s -10667 115709 -10567 115755 4 VSS
port 42 nsew
rlabel metal1 s -12620 115744 -12320 115790 4 VSS
port 42 nsew
rlabel metal1 s -7214 115913 -7114 115959 4 VSS
port 42 nsew
rlabel metal1 s -10667 115905 -10567 115951 4 VSS
port 42 nsew
rlabel metal1 s -9167 115994 -8867 116040 4 VSS
port 42 nsew
rlabel metal1 s -12620 115986 -12320 116032 4 VSS
port 42 nsew
rlabel metal1 s -7079 116104 -6966 116699 4 VSS
port 42 nsew
rlabel metal1 s -9388 116135 -9275 116325 4 VSS
port 42 nsew
rlabel metal1 s -10532 116096 -10419 116325 4 VSS
port 42 nsew
rlabel metal1 s -10532 116325 -9274 116438 4 VSS
port 42 nsew
rlabel metal1 s -9388 116438 -9275 116699 4 VSS
port 42 nsew
rlabel metal1 s -9388 116699 -6966 116812 4 VSS
port 42 nsew
rlabel metal1 s -10532 116438 -10419 116691 4 VSS
port 42 nsew
rlabel metal1 s -12841 116127 -12728 116131 4 VSS
port 42 nsew
rlabel metal1 s -12872 116131 -12728 116691 4 VSS
port 42 nsew
rlabel metal1 s -12872 116691 -10419 116804 4 VSS
port 42 nsew
rlabel metal1 s -9109 117450 -8809 117496 4 VSS
port 42 nsew
rlabel metal1 s -10469 117795 -10269 117841 4 VSS
port 42 nsew
rlabel metal1 s -12365 117769 -12065 117815 4 VSS
port 42 nsew
rlabel metal1 s -10469 117991 -10269 118037 4 VSS
port 42 nsew
rlabel metal1 s -9109 118241 -8609 118287 4 VSS
port 42 nsew
rlabel metal1 s -9109 118371 -8609 118417 4 VSS
port 42 nsew
rlabel metal1 s -11858 118378 -11758 118424 4 VSS
port 42 nsew
rlabel metal1 s -11858 118574 -11758 118620 4 VSS
port 42 nsew
rlabel metal1 s -9109 118697 -8809 118743 4 VSS
port 42 nsew
rlabel metal1 s -10391 118768 -10091 118814 4 VSS
port 42 nsew
rlabel metal1 s -12651 119216 -12351 119262 4 VSS
port 42 nsew
rlabel metal1 s -10698 119377 -10598 119423 4 VSS
port 42 nsew
rlabel metal1 s -12651 119412 -12351 119458 4 VSS
port 42 nsew
rlabel metal1 s -10698 119573 -10598 119619 4 VSS
port 42 nsew
rlabel metal1 s -12651 119654 -12351 119700 4 VSS
port 42 nsew
rlabel metal1 s -10563 119764 -10450 120359 4 VSS
port 42 nsew
rlabel metal1 s -12872 116804 -12759 120359 4 VSS
port 42 nsew
rlabel metal1 s -12872 120359 -10450 120472 4 VSS
port 42 nsew
rlabel locali s 91309 -53546 92592 -53281 8 VSS
port 42 nsew
rlabel locali s 89400 -53281 92592 -52743 8 VSS
port 42 nsew
rlabel locali s 91309 -52743 92592 -52202 8 VSS
port 42 nsew
rlabel locali s 90604 -35414 92221 -35170 8 VSS
port 42 nsew
rlabel locali s 88763 -35170 92221 -34632 8 VSS
port 42 nsew
rlabel locali s 90604 -34632 92221 -33888 8 VSS
port 42 nsew
rlabel locali s 90329 -18877 91702 -18579 8 VSS
port 42 nsew
rlabel locali s 88428 -18579 91702 -18041 8 VSS
port 42 nsew
rlabel locali s 90329 -18041 91702 -17504 8 VSS
port 42 nsew
rlabel locali s 81551 -7803 84520 -7667 8 VSS
port 42 nsew
rlabel locali s 70077 -7803 73046 -7667 8 VSS
port 42 nsew
rlabel locali s 70077 -7667 92959 -5275 8 VSS
port 42 nsew
rlabel locali s 46778 -5304 47412 -5275 8 VSS
port 42 nsew
rlabel locali s 46778 -5275 92959 -4698 8 VSS
port 42 nsew
rlabel locali s 52571 -4698 53148 -4341 8 VSS
port 42 nsew
rlabel locali s 46778 -4698 47398 -4670 8 VSS
port 42 nsew
rlabel locali s 50943 -4341 58130 -4221 8 VSS
port 42 nsew
rlabel locali s 63635 -3737 63669 -3578 8 VSS
port 42 nsew
rlabel locali s 63439 -3737 63473 -3578 8 VSS
port 42 nsew
rlabel locali s 63243 -3737 63277 -3578 8 VSS
port 42 nsew
rlabel locali s 58065 -4136 58099 -3728 8 VSS
port 42 nsew
rlabel locali s 57947 -4136 57981 -3728 8 VSS
port 42 nsew
rlabel locali s 57829 -4136 57863 -3728 8 VSS
port 42 nsew
rlabel locali s 57711 -4136 57745 -3728 8 VSS
port 42 nsew
rlabel locali s 57593 -4136 57627 -3728 8 VSS
port 42 nsew
rlabel locali s 57475 -4136 57509 -3728 8 VSS
port 42 nsew
rlabel locali s 57357 -4136 57391 -3728 8 VSS
port 42 nsew
rlabel locali s 57239 -4136 57273 -3728 8 VSS
port 42 nsew
rlabel locali s 57121 -4136 57155 -3728 8 VSS
port 42 nsew
rlabel locali s 57003 -4136 57037 -3728 8 VSS
port 42 nsew
rlabel locali s 56885 -4136 56919 -3728 8 VSS
port 42 nsew
rlabel locali s 56767 -4136 56801 -3728 8 VSS
port 42 nsew
rlabel locali s 56649 -4136 56683 -3728 8 VSS
port 42 nsew
rlabel locali s 56531 -4136 56565 -3728 8 VSS
port 42 nsew
rlabel locali s 56413 -4136 56447 -3728 8 VSS
port 42 nsew
rlabel locali s 56295 -4136 56329 -3728 8 VSS
port 42 nsew
rlabel locali s 56177 -4136 56211 -3728 8 VSS
port 42 nsew
rlabel locali s 56059 -4136 56093 -3728 8 VSS
port 42 nsew
rlabel locali s 55941 -4136 55975 -3728 8 VSS
port 42 nsew
rlabel locali s 55823 -4136 55857 -3728 8 VSS
port 42 nsew
rlabel locali s 55705 -4136 55739 -3728 8 VSS
port 42 nsew
rlabel locali s 55587 -4136 55621 -3728 8 VSS
port 42 nsew
rlabel locali s 55469 -4136 55503 -3728 8 VSS
port 42 nsew
rlabel locali s 55351 -4136 55385 -3728 8 VSS
port 42 nsew
rlabel locali s 55233 -4136 55267 -3728 8 VSS
port 42 nsew
rlabel locali s 55115 -4136 55149 -3728 8 VSS
port 42 nsew
rlabel locali s 54997 -4136 55031 -3728 8 VSS
port 42 nsew
rlabel locali s 54879 -4136 54913 -3728 8 VSS
port 42 nsew
rlabel locali s 54761 -4136 54795 -3728 8 VSS
port 42 nsew
rlabel locali s 54643 -4136 54677 -3728 8 VSS
port 42 nsew
rlabel locali s 54525 -4221 54559 -3728 8 VSS
port 42 nsew
rlabel locali s 54289 -4221 54323 -3728 8 VSS
port 42 nsew
rlabel locali s 54053 -4221 54087 -3728 8 VSS
port 42 nsew
rlabel locali s 53817 -4221 53851 -3728 8 VSS
port 42 nsew
rlabel locali s 53581 -4221 53615 -3728 8 VSS
port 42 nsew
rlabel locali s 53345 -4221 53379 -3728 8 VSS
port 42 nsew
rlabel locali s 53109 -4221 53143 -3728 8 VSS
port 42 nsew
rlabel locali s 52873 -4221 52907 -3728 8 VSS
port 42 nsew
rlabel locali s 52637 -4221 52671 -3728 8 VSS
port 42 nsew
rlabel locali s 52401 -4221 52435 -3728 8 VSS
port 42 nsew
rlabel locali s 52165 -4221 52199 -3728 8 VSS
port 42 nsew
rlabel locali s 51929 -4221 51963 -3728 8 VSS
port 42 nsew
rlabel locali s 51693 -4221 51727 -3728 8 VSS
port 42 nsew
rlabel locali s 51457 -4221 51491 -3728 8 VSS
port 42 nsew
rlabel locali s 51221 -4221 51255 -3728 8 VSS
port 42 nsew
rlabel locali s 50985 -4221 51019 -3728 8 VSS
port 42 nsew
rlabel locali s 54495 -3728 58125 -3664 8 VSS
port 42 nsew
rlabel locali s 54643 -3664 58125 -3636 8 VSS
port 42 nsew
rlabel locali s 63234 -3578 63768 -3441 8 VSS
port 42 nsew
rlabel locali s 62384 -3441 63768 -3373 8 VSS
port 42 nsew
rlabel locali s 63635 -3373 63669 -3214 8 VSS
port 42 nsew
rlabel locali s 63439 -3373 63473 -3214 8 VSS
port 42 nsew
rlabel locali s 63243 -3373 63277 -3214 8 VSS
port 42 nsew
rlabel locali s 62785 -3373 62819 -3214 8 VSS
port 42 nsew
rlabel locali s 62589 -3373 62623 -3214 8 VSS
port 42 nsew
rlabel locali s 62393 -3373 62427 -3214 8 VSS
port 42 nsew
rlabel locali s 46864 -2515 47369 -2242 8 VSS
port 42 nsew
rlabel locali s 46864 -2242 52968 -1737 8 VSS
port 42 nsew
rlabel locali s 52463 -1737 52968 -1294 8 VSS
port 42 nsew
rlabel locali s 46864 -1737 47369 -1450 8 VSS
port 42 nsew
rlabel locali s 8168 -2323 26638 -1966 8 VSS
port 42 nsew
rlabel locali s 26281 -1966 26638 -1450 8 VSS
port 42 nsew
rlabel locali s 13931 -1966 14204 -1916 8 VSS
port 42 nsew
rlabel locali s 13206 -1966 13479 -1916 8 VSS
port 42 nsew
rlabel locali s 12412 -1966 12685 -1916 8 VSS
port 42 nsew
rlabel locali s 11457 -1966 11730 -1916 8 VSS
port 42 nsew
rlabel locali s 10255 -1966 10528 -1916 8 VSS
port 42 nsew
rlabel locali s 9274 -1966 9547 -1916 8 VSS
port 42 nsew
rlabel locali s 8336 -1966 8557 -1916 8 VSS
port 42 nsew
rlabel locali s 7827 -1916 15014 -1796 8 VSS
port 42 nsew
rlabel locali s 50943 -1294 58130 -1174 8 VSS
port 42 nsew
rlabel locali s 58065 -1089 58099 -681 8 VSS
port 42 nsew
rlabel locali s 57947 -1089 57981 -681 8 VSS
port 42 nsew
rlabel locali s 57829 -1089 57863 -681 8 VSS
port 42 nsew
rlabel locali s 57711 -1089 57745 -681 8 VSS
port 42 nsew
rlabel locali s 57593 -1089 57627 -681 8 VSS
port 42 nsew
rlabel locali s 57475 -1089 57509 -681 8 VSS
port 42 nsew
rlabel locali s 57357 -1089 57391 -681 8 VSS
port 42 nsew
rlabel locali s 57239 -1089 57273 -681 8 VSS
port 42 nsew
rlabel locali s 57121 -1089 57155 -681 8 VSS
port 42 nsew
rlabel locali s 57003 -1089 57037 -681 8 VSS
port 42 nsew
rlabel locali s 56885 -1089 56919 -681 8 VSS
port 42 nsew
rlabel locali s 56767 -1089 56801 -681 8 VSS
port 42 nsew
rlabel locali s 56649 -1089 56683 -681 8 VSS
port 42 nsew
rlabel locali s 56531 -1089 56565 -681 8 VSS
port 42 nsew
rlabel locali s 56413 -1089 56447 -681 8 VSS
port 42 nsew
rlabel locali s 56295 -1089 56329 -681 8 VSS
port 42 nsew
rlabel locali s 56177 -1089 56211 -681 8 VSS
port 42 nsew
rlabel locali s 56059 -1089 56093 -681 8 VSS
port 42 nsew
rlabel locali s 55941 -1089 55975 -681 8 VSS
port 42 nsew
rlabel locali s 55823 -1089 55857 -681 8 VSS
port 42 nsew
rlabel locali s 55705 -1089 55739 -681 8 VSS
port 42 nsew
rlabel locali s 55587 -1089 55621 -681 8 VSS
port 42 nsew
rlabel locali s 55469 -1089 55503 -681 8 VSS
port 42 nsew
rlabel locali s 55351 -1089 55385 -681 8 VSS
port 42 nsew
rlabel locali s 55233 -1089 55267 -681 8 VSS
port 42 nsew
rlabel locali s 55115 -1089 55149 -681 8 VSS
port 42 nsew
rlabel locali s 54997 -1089 55031 -681 8 VSS
port 42 nsew
rlabel locali s 54879 -1089 54913 -681 8 VSS
port 42 nsew
rlabel locali s 54761 -1089 54795 -681 8 VSS
port 42 nsew
rlabel locali s 54643 -1089 54677 -681 8 VSS
port 42 nsew
rlabel locali s 54525 -1174 54559 -681 8 VSS
port 42 nsew
rlabel locali s 54289 -1174 54323 -681 8 VSS
port 42 nsew
rlabel locali s 54053 -1174 54087 -681 8 VSS
port 42 nsew
rlabel locali s 53817 -1174 53851 -681 8 VSS
port 42 nsew
rlabel locali s 53581 -1174 53615 -681 8 VSS
port 42 nsew
rlabel locali s 53345 -1174 53379 -681 8 VSS
port 42 nsew
rlabel locali s 53109 -1174 53143 -681 8 VSS
port 42 nsew
rlabel locali s 52873 -1174 52907 -681 8 VSS
port 42 nsew
rlabel locali s 52637 -1174 52671 -681 8 VSS
port 42 nsew
rlabel locali s 52401 -1174 52435 -681 8 VSS
port 42 nsew
rlabel locali s 52165 -1174 52199 -681 8 VSS
port 42 nsew
rlabel locali s 51929 -1174 51963 -681 8 VSS
port 42 nsew
rlabel locali s 51693 -1174 51727 -681 8 VSS
port 42 nsew
rlabel locali s 51457 -1174 51491 -681 8 VSS
port 42 nsew
rlabel locali s 51221 -1174 51255 -681 8 VSS
port 42 nsew
rlabel locali s 50985 -1174 51019 -681 8 VSS
port 42 nsew
rlabel locali s 25573 -1450 47674 -1155 8 VSS
port 42 nsew
rlabel locali s 14949 -1711 14983 -1303 8 VSS
port 42 nsew
rlabel locali s 14831 -1711 14865 -1303 8 VSS
port 42 nsew
rlabel locali s 14713 -1711 14747 -1303 8 VSS
port 42 nsew
rlabel locali s 14595 -1711 14629 -1303 8 VSS
port 42 nsew
rlabel locali s 14477 -1711 14511 -1303 8 VSS
port 42 nsew
rlabel locali s 14359 -1711 14393 -1303 8 VSS
port 42 nsew
rlabel locali s 14241 -1711 14275 -1303 8 VSS
port 42 nsew
rlabel locali s 14123 -1711 14157 -1303 8 VSS
port 42 nsew
rlabel locali s 14005 -1711 14039 -1303 8 VSS
port 42 nsew
rlabel locali s 13887 -1711 13921 -1303 8 VSS
port 42 nsew
rlabel locali s 13769 -1711 13803 -1303 8 VSS
port 42 nsew
rlabel locali s 13651 -1711 13685 -1303 8 VSS
port 42 nsew
rlabel locali s 13533 -1711 13567 -1303 8 VSS
port 42 nsew
rlabel locali s 13415 -1711 13449 -1303 8 VSS
port 42 nsew
rlabel locali s 13297 -1711 13331 -1303 8 VSS
port 42 nsew
rlabel locali s 13179 -1711 13213 -1303 8 VSS
port 42 nsew
rlabel locali s 13061 -1711 13095 -1303 8 VSS
port 42 nsew
rlabel locali s 12943 -1711 12977 -1303 8 VSS
port 42 nsew
rlabel locali s 12825 -1711 12859 -1303 8 VSS
port 42 nsew
rlabel locali s 12707 -1711 12741 -1303 8 VSS
port 42 nsew
rlabel locali s 12589 -1711 12623 -1303 8 VSS
port 42 nsew
rlabel locali s 12471 -1711 12505 -1303 8 VSS
port 42 nsew
rlabel locali s 12353 -1711 12387 -1303 8 VSS
port 42 nsew
rlabel locali s 12235 -1711 12269 -1303 8 VSS
port 42 nsew
rlabel locali s 12117 -1711 12151 -1303 8 VSS
port 42 nsew
rlabel locali s 11999 -1711 12033 -1303 8 VSS
port 42 nsew
rlabel locali s 11881 -1711 11915 -1303 8 VSS
port 42 nsew
rlabel locali s 11763 -1711 11797 -1303 8 VSS
port 42 nsew
rlabel locali s 11645 -1711 11679 -1303 8 VSS
port 42 nsew
rlabel locali s 11527 -1711 11561 -1303 8 VSS
port 42 nsew
rlabel locali s 11409 -1796 11443 -1303 8 VSS
port 42 nsew
rlabel locali s 11173 -1796 11207 -1303 8 VSS
port 42 nsew
rlabel locali s 10937 -1796 10971 -1303 8 VSS
port 42 nsew
rlabel locali s 10701 -1796 10735 -1303 8 VSS
port 42 nsew
rlabel locali s 10465 -1796 10499 -1303 8 VSS
port 42 nsew
rlabel locali s 10229 -1796 10263 -1303 8 VSS
port 42 nsew
rlabel locali s 9993 -1796 10027 -1303 8 VSS
port 42 nsew
rlabel locali s 9757 -1796 9791 -1303 8 VSS
port 42 nsew
rlabel locali s 9521 -1796 9555 -1303 8 VSS
port 42 nsew
rlabel locali s 9285 -1796 9319 -1303 8 VSS
port 42 nsew
rlabel locali s 9049 -1796 9083 -1303 8 VSS
port 42 nsew
rlabel locali s 8813 -1796 8847 -1303 8 VSS
port 42 nsew
rlabel locali s 8577 -1796 8611 -1303 8 VSS
port 42 nsew
rlabel locali s 8341 -1796 8375 -1303 8 VSS
port 42 nsew
rlabel locali s 8105 -1796 8139 -1303 8 VSS
port 42 nsew
rlabel locali s 7869 -1796 7903 -1303 8 VSS
port 42 nsew
rlabel locali s 11379 -1303 15009 -1239 8 VSS
port 42 nsew
rlabel locali s 11527 -1239 15009 -1211 8 VSS
port 42 nsew
rlabel locali s 5772 -1376 5806 -1217 8 VSS
port 42 nsew
rlabel locali s 5576 -1376 5610 -1217 8 VSS
port 42 nsew
rlabel locali s 5380 -1376 5414 -1217 8 VSS
port 42 nsew
rlabel locali s 54495 -681 58125 -617 8 VSS
port 42 nsew
rlabel locali s 54643 -617 58125 -589 8 VSS
port 42 nsew
rlabel locali s 47379 -1155 47674 537 8 VSS
port 42 nsew
rlabel locali s 36761 -433 38097 -308 8 VSS
port 42 nsew
rlabel locali s 35040 -476 36376 -351 8 VSS
port 42 nsew
rlabel locali s 30305 -499 31641 -374 8 VSS
port 42 nsew
rlabel locali s 38050 -308 38084 272 8 VSS
port 42 nsew
rlabel locali s 37892 -154 37926 272 6 VSS
port 42 nsew
rlabel locali s 37734 -308 37768 272 8 VSS
port 42 nsew
rlabel locali s 37576 -154 37610 272 6 VSS
port 42 nsew
rlabel locali s 37418 -308 37452 254 8 VSS
port 42 nsew
rlabel locali s 37102 -308 37136 254 8 VSS
port 42 nsew
rlabel locali s 36786 -308 36820 -265 8 VSS
port 42 nsew
rlabel locali s 36329 -351 36363 -265 8 VSS
port 42 nsew
rlabel locali s 36329 -265 36820 -210 8 VSS
port 42 nsew
rlabel locali s 36786 -210 36820 254 6 VSS
port 42 nsew
rlabel locali s 36329 -210 36363 229 6 VSS
port 42 nsew
rlabel locali s 36171 -197 36205 229 6 VSS
port 42 nsew
rlabel locali s 36013 -351 36047 229 8 VSS
port 42 nsew
rlabel locali s 35855 -197 35889 229 6 VSS
port 42 nsew
rlabel locali s 35697 -351 35731 211 8 VSS
port 42 nsew
rlabel locali s 35381 -351 35415 211 8 VSS
port 42 nsew
rlabel locali s 35065 -351 35099 -294 8 VSS
port 42 nsew
rlabel locali s 31594 -374 31628 -307 8 VSS
port 42 nsew
rlabel locali s 34420 -294 35099 -260 8 VSS
port 42 nsew
rlabel locali s 35065 -260 35099 211 8 VSS
port 42 nsew
rlabel locali s 34420 -260 34502 -247 8 VSS
port 42 nsew
rlabel locali s 32636 -247 34502 -232 8 VSS
port 42 nsew
rlabel locali s 31594 -307 32499 -232 8 VSS
port 42 nsew
rlabel locali s 31594 -232 34502 -217 8 VSS
port 42 nsew
rlabel locali s 32392 -217 34502 -198 8 VSS
port 42 nsew
rlabel locali s 32636 -198 34502 -189 8 VSS
port 42 nsew
rlabel locali s 34444 -189 34502 -139 8 VSS
port 42 nsew
rlabel locali s 34361 -139 34553 -48 8 VSS
port 42 nsew
rlabel locali s 34519 -48 34553 176 6 VSS
port 42 nsew
rlabel locali s 34361 -48 34395 176 6 VSS
port 42 nsew
rlabel locali s 34086 -189 34120 176 8 VSS
port 42 nsew
rlabel locali s 33770 -189 33804 176 8 VSS
port 42 nsew
rlabel locali s 33454 -189 33488 176 8 VSS
port 42 nsew
rlabel locali s 33138 -189 33172 176 8 VSS
port 42 nsew
rlabel locali s 32822 -189 32856 176 8 VSS
port 42 nsew
rlabel locali s 32550 -34 32584 195 6 VSS
port 42 nsew
rlabel locali s 32392 -198 32426 195 8 VSS
port 42 nsew
rlabel locali s 35855 229 36363 263 6 VSS
port 42 nsew
rlabel locali s 37576 272 38084 306 6 VSS
port 42 nsew
rlabel locali s 37625 306 38028 359 6 VSS
port 42 nsew
rlabel locali s 35904 263 36307 316 6 VSS
port 42 nsew
rlabel locali s 32392 195 32584 267 6 VSS
port 42 nsew
rlabel locali s 31594 -217 31628 206 8 VSS
port 42 nsew
rlabel locali s 31436 -220 31470 206 8 VSS
port 42 nsew
rlabel locali s 31278 -374 31312 206 8 VSS
port 42 nsew
rlabel locali s 31120 -220 31154 206 8 VSS
port 42 nsew
rlabel locali s 30962 -374 30996 188 8 VSS
port 42 nsew
rlabel locali s 30646 -374 30680 188 8 VSS
port 42 nsew
rlabel locali s 30330 -374 30364 -291 8 VSS
port 42 nsew
rlabel locali s 29583 -291 30364 -240 8 VSS
port 42 nsew
rlabel locali s 27781 -240 30364 -225 8 VSS
port 42 nsew
rlabel locali s 27537 -1155 27726 -225 8 VSS
port 42 nsew
rlabel locali s 27537 -225 30364 -191 8 VSS
port 42 nsew
rlabel locali s 27781 -191 30364 -182 8 VSS
port 42 nsew
rlabel locali s 30330 -182 30364 188 6 VSS
port 42 nsew
rlabel locali s 29589 -182 29647 -132 8 VSS
port 42 nsew
rlabel locali s 29506 -132 29698 -41 8 VSS
port 42 nsew
rlabel locali s 29664 -41 29698 183 6 VSS
port 42 nsew
rlabel locali s 29506 -41 29540 183 6 VSS
port 42 nsew
rlabel locali s 29231 -182 29265 183 8 VSS
port 42 nsew
rlabel locali s 28915 -182 28949 183 8 VSS
port 42 nsew
rlabel locali s 28599 -182 28633 183 8 VSS
port 42 nsew
rlabel locali s 28283 -182 28317 183 8 VSS
port 42 nsew
rlabel locali s 27967 -182 28001 183 8 VSS
port 42 nsew
rlabel locali s 31120 206 31628 240 6 VSS
port 42 nsew
rlabel locali s 27695 -27 27729 202 6 VSS
port 42 nsew
rlabel locali s 27537 -191 27571 202 6 VSS
port 42 nsew
rlabel locali s 31169 240 31572 293 6 VSS
port 42 nsew
rlabel locali s 27537 202 27729 274 6 VSS
port 42 nsew
rlabel locali s 47379 537 52157 824 6 VSS
port 42 nsew
rlabel locali s 34134 478 34168 770 6 VSS
port 42 nsew
rlabel locali s 33976 478 34010 770 6 VSS
port 42 nsew
rlabel locali s 32671 396 32863 479 6 VSS
port 42 nsew
rlabel locali s 32829 479 32863 686 6 VSS
port 42 nsew
rlabel locali s 32671 479 32705 686 6 VSS
port 42 nsew
rlabel locali s 51870 824 52157 1617 6 VSS
port 42 nsew
rlabel locali s 51146 1617 58333 1737 6 VSS
port 42 nsew
rlabel locali s 58268 1822 58302 2230 6 VSS
port 42 nsew
rlabel locali s 58150 1822 58184 2230 6 VSS
port 42 nsew
rlabel locali s 58032 1822 58066 2230 6 VSS
port 42 nsew
rlabel locali s 57914 1822 57948 2230 6 VSS
port 42 nsew
rlabel locali s 57796 1822 57830 2230 6 VSS
port 42 nsew
rlabel locali s 57678 1822 57712 2230 6 VSS
port 42 nsew
rlabel locali s 57560 1822 57594 2230 6 VSS
port 42 nsew
rlabel locali s 57442 1822 57476 2230 6 VSS
port 42 nsew
rlabel locali s 57324 1822 57358 2230 6 VSS
port 42 nsew
rlabel locali s 57206 1822 57240 2230 6 VSS
port 42 nsew
rlabel locali s 57088 1822 57122 2230 6 VSS
port 42 nsew
rlabel locali s 56970 1822 57004 2230 6 VSS
port 42 nsew
rlabel locali s 56852 1822 56886 2230 6 VSS
port 42 nsew
rlabel locali s 56734 1822 56768 2230 6 VSS
port 42 nsew
rlabel locali s 56616 1822 56650 2230 6 VSS
port 42 nsew
rlabel locali s 56498 1822 56532 2230 6 VSS
port 42 nsew
rlabel locali s 56380 1822 56414 2230 6 VSS
port 42 nsew
rlabel locali s 56262 1822 56296 2230 6 VSS
port 42 nsew
rlabel locali s 56144 1822 56178 2230 6 VSS
port 42 nsew
rlabel locali s 56026 1822 56060 2230 6 VSS
port 42 nsew
rlabel locali s 55908 1822 55942 2230 6 VSS
port 42 nsew
rlabel locali s 55790 1822 55824 2230 6 VSS
port 42 nsew
rlabel locali s 55672 1822 55706 2230 6 VSS
port 42 nsew
rlabel locali s 55554 1822 55588 2230 6 VSS
port 42 nsew
rlabel locali s 55436 1822 55470 2230 6 VSS
port 42 nsew
rlabel locali s 55318 1822 55352 2230 6 VSS
port 42 nsew
rlabel locali s 55200 1822 55234 2230 6 VSS
port 42 nsew
rlabel locali s 55082 1822 55116 2230 6 VSS
port 42 nsew
rlabel locali s 54964 1822 54998 2230 6 VSS
port 42 nsew
rlabel locali s 54846 1822 54880 2230 6 VSS
port 42 nsew
rlabel locali s 54728 1737 54762 2230 6 VSS
port 42 nsew
rlabel locali s 54492 1737 54526 2230 6 VSS
port 42 nsew
rlabel locali s 54256 1737 54290 2230 6 VSS
port 42 nsew
rlabel locali s 54020 1737 54054 2230 6 VSS
port 42 nsew
rlabel locali s 53784 1737 53818 2230 6 VSS
port 42 nsew
rlabel locali s 53548 1737 53582 2230 6 VSS
port 42 nsew
rlabel locali s 53312 1737 53346 2230 6 VSS
port 42 nsew
rlabel locali s 53076 1737 53110 2230 6 VSS
port 42 nsew
rlabel locali s 52840 1737 52874 2230 6 VSS
port 42 nsew
rlabel locali s 52604 1737 52638 2230 6 VSS
port 42 nsew
rlabel locali s 52368 1737 52402 2230 6 VSS
port 42 nsew
rlabel locali s 52132 1737 52166 2230 6 VSS
port 42 nsew
rlabel locali s 51896 1737 51930 2230 6 VSS
port 42 nsew
rlabel locali s 51660 1737 51694 2230 6 VSS
port 42 nsew
rlabel locali s 51424 1737 51458 2230 6 VSS
port 42 nsew
rlabel locali s 51188 1737 51222 2230 6 VSS
port 42 nsew
rlabel locali s 54698 2230 58328 2294 6 VSS
port 42 nsew
rlabel locali s 54846 2294 58328 2322 6 VSS
port 42 nsew
rlabel locali s 47379 824 47674 3483 6 VSS
port 42 nsew
rlabel locali s 33956 770 34191 851 6 VSS
port 42 nsew
rlabel locali s 29279 485 29313 777 6 VSS
port 42 nsew
rlabel locali s 29121 485 29155 777 6 VSS
port 42 nsew
rlabel locali s 27816 403 28008 486 6 VSS
port 42 nsew
rlabel locali s 27974 486 28008 693 6 VSS
port 42 nsew
rlabel locali s 27816 486 27850 693 6 VSS
port 42 nsew
rlabel locali s 34135 851 34169 1134 6 VSS
port 42 nsew
rlabel locali s 33977 851 34011 1134 6 VSS
port 42 nsew
rlabel locali s 29101 777 29336 858 6 VSS
port 42 nsew
rlabel locali s 32829 930 32863 1138 6 VSS
port 42 nsew
rlabel locali s 32671 930 32705 1138 6 VSS
port 42 nsew
rlabel locali s 29280 858 29314 1141 6 VSS
port 42 nsew
rlabel locali s 29122 858 29156 1141 6 VSS
port 42 nsew
rlabel locali s 25573 -1155 25868 876 8 VSS
port 42 nsew
rlabel locali s 5371 -1217 5905 -1080 8 VSS
port 42 nsew
rlabel locali s 4521 -1080 5905 -1012 8 VSS
port 42 nsew
rlabel locali s 21208 -871 21242 -712 8 VSS
port 42 nsew
rlabel locali s 21012 -871 21046 -712 8 VSS
port 42 nsew
rlabel locali s 20816 -871 20850 -712 8 VSS
port 42 nsew
rlabel locali s 5772 -1012 5806 -853 8 VSS
port 42 nsew
rlabel locali s 5576 -1012 5610 -853 8 VSS
port 42 nsew
rlabel locali s 5380 -1012 5414 -853 8 VSS
port 42 nsew
rlabel locali s 4922 -1012 4956 -853 8 VSS
port 42 nsew
rlabel locali s 4726 -1012 4760 -853 8 VSS
port 42 nsew
rlabel locali s 4530 -1012 4564 -853 8 VSS
port 42 nsew
rlabel locali s 20807 -712 21341 -575 8 VSS
port 42 nsew
rlabel locali s 19957 -575 21341 -507 8 VSS
port 42 nsew
rlabel locali s 21208 -507 21242 -348 8 VSS
port 42 nsew
rlabel locali s 21012 -507 21046 -348 8 VSS
port 42 nsew
rlabel locali s 20816 -507 20850 -348 8 VSS
port 42 nsew
rlabel locali s 20358 -507 20392 -348 8 VSS
port 42 nsew
rlabel locali s 20162 -507 20196 -348 8 VSS
port 42 nsew
rlabel locali s 19966 -507 20000 -348 8 VSS
port 42 nsew
rlabel locali s 2764 336 3099 382 6 VSS
port 42 nsew
rlabel locali s 2764 382 19742 495 6 VSS
port 42 nsew
rlabel locali s 565 495 19742 590 6 VSS
port 42 nsew
rlabel locali s 2455 590 19742 593 6 VSS
port 42 nsew
rlabel locali s 3030 593 19742 595 6 VSS
port 42 nsew
rlabel locali s 8089 595 19742 744 6 VSS
port 42 nsew
rlabel locali s 27974 937 28008 1145 6 VSS
port 42 nsew
rlabel locali s 27816 937 27850 1145 6 VSS
port 42 nsew
rlabel locali s 22419 876 25868 1356 6 VSS
port 42 nsew
rlabel locali s 19404 744 19742 943 6 VSS
port 42 nsew
rlabel locali s 14498 744 14866 840 6 VSS
port 42 nsew
rlabel locali s 13329 744 13697 840 6 VSS
port 42 nsew
rlabel locali s 12204 744 12572 840 6 VSS
port 42 nsew
rlabel locali s 10640 744 11008 840 6 VSS
port 42 nsew
rlabel locali s 9394 744 9762 840 6 VSS
port 42 nsew
rlabel locali s 8203 744 8571 840 6 VSS
port 42 nsew
rlabel locali s 19404 943 19770 1241 6 VSS
port 42 nsew
rlabel locali s 7868 840 15055 960 6 VSS
port 42 nsew
rlabel locali s 19404 1241 19736 1242 6 VSS
port 42 nsew
rlabel locali s 45971 1883 46005 2042 6 VSS
port 42 nsew
rlabel locali s 45775 1883 45809 2042 6 VSS
port 42 nsew
rlabel locali s 45579 1883 45613 2042 6 VSS
port 42 nsew
rlabel locali s 45001 1793 45035 1952 6 VSS
port 42 nsew
rlabel locali s 44805 1793 44839 1952 6 VSS
port 42 nsew
rlabel locali s 44609 1793 44643 1952 6 VSS
port 42 nsew
rlabel locali s 44164 1793 44198 1952 6 VSS
port 42 nsew
rlabel locali s 43968 1793 44002 1952 6 VSS
port 42 nsew
rlabel locali s 43772 1793 43806 1952 6 VSS
port 42 nsew
rlabel locali s 42301 1793 42335 1952 6 VSS
port 42 nsew
rlabel locali s 42105 1793 42139 1952 6 VSS
port 42 nsew
rlabel locali s 41909 1793 41943 1952 6 VSS
port 42 nsew
rlabel locali s 41464 1793 41498 1952 6 VSS
port 42 nsew
rlabel locali s 41268 1793 41302 1952 6 VSS
port 42 nsew
rlabel locali s 41072 1793 41106 1952 6 VSS
port 42 nsew
rlabel locali s 43673 1952 45044 2020 6 VSS
port 42 nsew
rlabel locali s 41810 1952 42344 1954 6 VSS
port 42 nsew
rlabel locali s 40973 1952 41507 1954 6 VSS
port 42 nsew
rlabel locali s 40973 1954 42344 2020 6 VSS
port 42 nsew
rlabel locali s 37625 1966 38028 2019 6 VSS
port 42 nsew
rlabel locali s 45570 2042 46104 2110 6 VSS
port 42 nsew
rlabel locali s 44685 2020 44796 2060 6 VSS
port 42 nsew
rlabel locali s 44670 2060 44807 2068 6 VSS
port 42 nsew
rlabel locali s 43874 2020 43985 2068 6 VSS
port 42 nsew
rlabel locali s 42076 2020 42187 2066 6 VSS
port 42 nsew
rlabel locali s 41484 2020 42004 2022 6 VSS
port 42 nsew
rlabel locali s 42073 2066 42210 2068 6 VSS
port 42 nsew
rlabel locali s 41198 2020 41309 2068 6 VSS
port 42 nsew
rlabel locali s 37576 2019 38084 2053 6 VSS
port 42 nsew
rlabel locali s 39440 2066 39572 2068 6 VSS
port 42 nsew
rlabel locali s 39439 2068 44824 2107 6 VSS
port 42 nsew
rlabel locali s 45853 2110 45897 2255 6 VSS
port 42 nsew
rlabel locali s 44670 2107 44807 2120 6 VSS
port 42 nsew
rlabel locali s 42073 2107 42210 2126 6 VSS
port 42 nsew
rlabel locali s 39440 2107 39572 2126 6 VSS
port 42 nsew
rlabel locali s 45804 2255 45950 2441 6 VSS
port 42 nsew
rlabel locali s 44502 2332 45036 2400 6 VSS
port 42 nsew
rlabel locali s 41802 2332 43293 2400 6 VSS
port 42 nsew
rlabel locali s 39177 2332 40593 2400 6 VSS
port 42 nsew
rlabel locali s 44903 2400 44937 2559 6 VSS
port 42 nsew
rlabel locali s 44707 2400 44741 2559 6 VSS
port 42 nsew
rlabel locali s 44511 2400 44545 2559 6 VSS
port 42 nsew
rlabel locali s 43160 2400 43194 2559 6 VSS
port 42 nsew
rlabel locali s 42964 2400 42998 2559 6 VSS
port 42 nsew
rlabel locali s 42768 2400 42802 2559 6 VSS
port 42 nsew
rlabel locali s 42203 2400 42237 2559 6 VSS
port 42 nsew
rlabel locali s 42007 2400 42041 2559 6 VSS
port 42 nsew
rlabel locali s 41811 2400 41845 2559 6 VSS
port 42 nsew
rlabel locali s 40460 2400 40494 2559 6 VSS
port 42 nsew
rlabel locali s 40264 2400 40298 2559 6 VSS
port 42 nsew
rlabel locali s 40068 2400 40102 2559 6 VSS
port 42 nsew
rlabel locali s 39578 2400 39612 2559 6 VSS
port 42 nsew
rlabel locali s 39382 2400 39416 2559 6 VSS
port 42 nsew
rlabel locali s 39186 2400 39220 2559 6 VSS
port 42 nsew
rlabel locali s 38780 2149 38972 2407 6 VSS
port 42 nsew
rlabel locali s 38874 2407 38938 2548 6 VSS
port 42 nsew
rlabel locali s 38050 2053 38084 2548 6 VSS
port 42 nsew
rlabel locali s 37892 2053 37926 2479 6 VSS
port 42 nsew
rlabel locali s 38050 2548 38938 2633 6 VSS
port 42 nsew
rlabel locali s 37734 2053 37768 2633 6 VSS
port 42 nsew
rlabel locali s 37576 2053 37610 2479 6 VSS
port 42 nsew
rlabel locali s 35904 2009 36307 2062 6 VSS
port 42 nsew
rlabel locali s 31169 1987 31572 2040 6 VSS
port 42 nsew
rlabel locali s 37418 2071 37452 2633 6 VSS
port 42 nsew
rlabel locali s 37102 2071 37136 2633 6 VSS
port 42 nsew
rlabel locali s 36786 2071 36820 2548 6 VSS
port 42 nsew
rlabel locali s 35855 2062 36363 2096 6 VSS
port 42 nsew
rlabel locali s 36329 2096 36363 2548 6 VSS
port 42 nsew
rlabel locali s 36171 2096 36205 2522 6 VSS
port 42 nsew
rlabel locali s 36329 2548 36820 2633 6 VSS
port 42 nsew
rlabel locali s 36329 2633 38938 2641 6 VSS
port 42 nsew
rlabel locali s 36761 2641 38938 2644 6 VSS
port 42 nsew
rlabel locali s 36761 2644 38097 2758 6 VSS
port 42 nsew
rlabel locali s 36329 2641 36363 2676 6 VSS
port 42 nsew
rlabel locali s 36013 2096 36047 2676 6 VSS
port 42 nsew
rlabel locali s 35855 2096 35889 2522 6 VSS
port 42 nsew
rlabel locali s 31120 2040 31628 2074 6 VSS
port 42 nsew
rlabel locali s 35697 2114 35731 2676 6 VSS
port 42 nsew
rlabel locali s 35381 2114 35415 2676 6 VSS
port 42 nsew
rlabel locali s 35065 2114 35099 2564 6 VSS
port 42 nsew
rlabel locali s 31594 2074 31628 2564 6 VSS
port 42 nsew
rlabel locali s 31436 2074 31470 2500 6 VSS
port 42 nsew
rlabel locali s 31594 2564 35099 2654 6 VSS
port 42 nsew
rlabel locali s 31278 2074 31312 2654 6 VSS
port 42 nsew
rlabel locali s 31120 2074 31154 2500 6 VSS
port 42 nsew
rlabel locali s 30962 2092 30996 2654 6 VSS
port 42 nsew
rlabel locali s 30646 2092 30680 2654 6 VSS
port 42 nsew
rlabel locali s 30330 2092 30364 2654 6 VSS
port 42 nsew
rlabel locali s 30305 2654 35099 2676 6 VSS
port 42 nsew
rlabel locali s 30305 2676 36376 2689 6 VSS
port 42 nsew
rlabel locali s 35040 2689 36376 2801 6 VSS
port 42 nsew
rlabel locali s 33299 2689 33705 3483 6 VSS
port 42 nsew
rlabel locali s 30305 2689 31641 2779 6 VSS
port 42 nsew
rlabel locali s 26289 3483 47674 3484 6 VSS
port 42 nsew
rlabel locali s 25573 1356 25868 3484 6 VSS
port 42 nsew
rlabel locali s 21036 2479 21070 2638 6 VSS
port 42 nsew
rlabel locali s 20840 2479 20874 2638 6 VSS
port 42 nsew
rlabel locali s 20644 2479 20678 2638 6 VSS
port 42 nsew
rlabel locali s 20635 2638 21169 2775 6 VSS
port 42 nsew
rlabel locali s 19785 2775 21169 2843 6 VSS
port 42 nsew
rlabel locali s 19567 1242 19632 2800 6 VSS
port 42 nsew
rlabel locali s 14990 1045 15024 1453 6 VSS
port 42 nsew
rlabel locali s 14872 1045 14906 1453 6 VSS
port 42 nsew
rlabel locali s 14754 1045 14788 1453 6 VSS
port 42 nsew
rlabel locali s 14636 1045 14670 1453 6 VSS
port 42 nsew
rlabel locali s 14518 1045 14552 1453 6 VSS
port 42 nsew
rlabel locali s 14400 1045 14434 1453 6 VSS
port 42 nsew
rlabel locali s 14282 1045 14316 1453 6 VSS
port 42 nsew
rlabel locali s 14164 1045 14198 1453 6 VSS
port 42 nsew
rlabel locali s 14046 1045 14080 1453 6 VSS
port 42 nsew
rlabel locali s 13928 1045 13962 1453 6 VSS
port 42 nsew
rlabel locali s 13810 1045 13844 1453 6 VSS
port 42 nsew
rlabel locali s 13692 1045 13726 1453 6 VSS
port 42 nsew
rlabel locali s 13574 1045 13608 1453 6 VSS
port 42 nsew
rlabel locali s 13456 1045 13490 1453 6 VSS
port 42 nsew
rlabel locali s 13338 1045 13372 1453 6 VSS
port 42 nsew
rlabel locali s 13220 1045 13254 1453 6 VSS
port 42 nsew
rlabel locali s 13102 1045 13136 1453 6 VSS
port 42 nsew
rlabel locali s 12984 1045 13018 1453 6 VSS
port 42 nsew
rlabel locali s 12866 1045 12900 1453 6 VSS
port 42 nsew
rlabel locali s 12748 1045 12782 1453 6 VSS
port 42 nsew
rlabel locali s 12630 1045 12664 1453 6 VSS
port 42 nsew
rlabel locali s 12512 1045 12546 1453 6 VSS
port 42 nsew
rlabel locali s 12394 1045 12428 1453 6 VSS
port 42 nsew
rlabel locali s 12276 1045 12310 1453 6 VSS
port 42 nsew
rlabel locali s 12158 1045 12192 1453 6 VSS
port 42 nsew
rlabel locali s 12040 1045 12074 1453 6 VSS
port 42 nsew
rlabel locali s 11922 1045 11956 1453 6 VSS
port 42 nsew
rlabel locali s 11804 1045 11838 1453 6 VSS
port 42 nsew
rlabel locali s 11686 1045 11720 1453 6 VSS
port 42 nsew
rlabel locali s 11568 1045 11602 1453 6 VSS
port 42 nsew
rlabel locali s 11450 960 11484 1453 6 VSS
port 42 nsew
rlabel locali s 11214 960 11248 1453 6 VSS
port 42 nsew
rlabel locali s 10978 960 11012 1453 6 VSS
port 42 nsew
rlabel locali s 10742 960 10776 1453 6 VSS
port 42 nsew
rlabel locali s 10506 960 10540 1453 6 VSS
port 42 nsew
rlabel locali s 10270 960 10304 1453 6 VSS
port 42 nsew
rlabel locali s 10034 960 10068 1453 6 VSS
port 42 nsew
rlabel locali s 9798 960 9832 1453 6 VSS
port 42 nsew
rlabel locali s 9394 960 9762 971 6 VSS
port 42 nsew
rlabel locali s 9562 971 9596 1453 6 VSS
port 42 nsew
rlabel locali s 9326 960 9360 1453 6 VSS
port 42 nsew
rlabel locali s 9090 960 9124 1453 6 VSS
port 42 nsew
rlabel locali s 8854 960 8888 1453 6 VSS
port 42 nsew
rlabel locali s 8618 960 8652 1453 6 VSS
port 42 nsew
rlabel locali s 8382 960 8416 1453 6 VSS
port 42 nsew
rlabel locali s 8146 960 8180 1453 6 VSS
port 42 nsew
rlabel locali s 7910 960 7944 1453 6 VSS
port 42 nsew
rlabel locali s 11420 1453 15050 1517 6 VSS
port 42 nsew
rlabel locali s 5757 1314 5791 1473 6 VSS
port 42 nsew
rlabel locali s 5561 1314 5595 1473 6 VSS
port 42 nsew
rlabel locali s 5365 1314 5399 1473 6 VSS
port 42 nsew
rlabel locali s 11568 1517 15050 1545 6 VSS
port 42 nsew
rlabel locali s 5356 1473 5890 1610 6 VSS
port 42 nsew
rlabel locali s 4600 1392 4817 1517 6 VSS
port 42 nsew
rlabel locali s 4196 595 4326 1504 6 VSS
port 42 nsew
rlabel locali s 2455 593 2965 690 6 VSS
port 42 nsew
rlabel locali s 2809 690 2843 865 6 VSS
port 42 nsew
rlabel locali s 2500 690 2534 865 6 VSS
port 42 nsew
rlabel locali s 2183 736 2217 864 6 VSS
port 42 nsew
rlabel locali s 1947 736 1981 864 6 VSS
port 42 nsew
rlabel locali s 1515 590 1549 871 6 VSS
port 42 nsew
rlabel locali s 1225 590 1259 876 6 VSS
port 42 nsew
rlabel locali s 591 590 792 690 6 VSS
port 42 nsew
rlabel locali s 713 690 747 865 6 VSS
port 42 nsew
rlabel locali s 4626 1517 4768 1610 6 VSS
port 42 nsew
rlabel locali s 4506 1610 5890 1678 6 VSS
port 42 nsew
rlabel locali s 5757 1678 5791 1837 6 VSS
port 42 nsew
rlabel locali s 5561 1678 5595 1837 6 VSS
port 42 nsew
rlabel locali s 5365 1678 5399 1837 6 VSS
port 42 nsew
rlabel locali s 4907 1678 4941 1837 6 VSS
port 42 nsew
rlabel locali s 4711 1678 4745 1837 6 VSS
port 42 nsew
rlabel locali s 4515 1678 4549 1837 6 VSS
port 42 nsew
rlabel locali s 2809 1997 2843 2172 6 VSS
port 42 nsew
rlabel locali s 2500 1997 2534 2172 6 VSS
port 42 nsew
rlabel locali s 2183 1998 2217 2126 6 VSS
port 42 nsew
rlabel locali s 1947 1998 1981 2126 6 VSS
port 42 nsew
rlabel locali s 2455 2172 2965 2272 6 VSS
port 42 nsew
rlabel locali s 1515 1991 1549 2272 6 VSS
port 42 nsew
rlabel locali s 1225 1986 1259 2272 6 VSS
port 42 nsew
rlabel locali s 713 1997 747 2172 6 VSS
port 42 nsew
rlabel locali s 591 2172 792 2272 6 VSS
port 42 nsew
rlabel locali s 565 2272 2965 2274 6 VSS
port 42 nsew
rlabel locali s 565 2274 3099 2367 6 VSS
port 42 nsew
rlabel locali s 2820 2367 3099 2508 6 VSS
port 42 nsew
rlabel locali s 21036 2843 21070 3002 6 VSS
port 42 nsew
rlabel locali s 20840 2843 20874 3002 6 VSS
port 42 nsew
rlabel locali s 20644 2843 20678 3002 6 VSS
port 42 nsew
rlabel locali s 19794 2843 20301 2844 6 VSS
port 42 nsew
rlabel locali s 20186 2844 20220 3002 6 VSS
port 42 nsew
rlabel locali s 19990 2844 20024 3002 6 VSS
port 42 nsew
rlabel locali s 19794 2844 19828 3002 6 VSS
port 42 nsew
rlabel locali s 19563 2800 19636 2877 6 VSS
port 42 nsew
rlabel locali s 19567 2877 19632 2878 6 VSS
port 42 nsew
rlabel locali s 25573 3484 47674 3778 6 VSS
port 42 nsew
rlabel locali s 26583 3778 38866 3886 6 VSS
port 42 nsew
rlabel locali s 25573 3778 26392 3779 6 VSS
port 42 nsew
rlabel locali s -2197 4085 12654 4551 6 VSS
port 42 nsew
rlabel locali s 11612 4551 11647 4643 6 VSS
port 42 nsew
rlabel locali s 11612 4643 11646 6447 6 VSS
port 42 nsew
rlabel locali s 9896 4551 9930 6447 6 VSS
port 42 nsew
rlabel locali s 8180 4551 8214 6447 6 VSS
port 42 nsew
rlabel locali s 2866 4551 3250 4560 6 VSS
port 42 nsew
rlabel locali s -2105 4551 -746 7185 4 VSS
port 42 nsew
rlabel locali s 26753 7623 38073 7646 6 VSS
port 42 nsew
rlabel locali s 17671 7646 92311 8151 6 VSS
port 42 nsew
rlabel locali s 17125 8151 92311 8341 6 VSS
port 42 nsew
rlabel locali s 17671 8341 92311 8878 6 VSS
port 42 nsew
rlabel locali s 69243 8878 92311 9648 6 VSS
port 42 nsew
rlabel locali s 17125 8341 17315 8908 6 VSS
port 42 nsew
rlabel locali s -6647 7185 -745 8544 4 VSS
port 42 nsew
rlabel locali s -16182 8044 -15367 8210 4 VSS
port 42 nsew
rlabel locali s 69243 9648 92336 9668 6 VSS
port 42 nsew
rlabel locali s 17118 8908 17337 9106 6 VSS
port 42 nsew
rlabel locali s 16029 8972 16121 9006 6 VSS
port 42 nsew
rlabel locali s 16814 9106 17337 9140 6 VSS
port 42 nsew
rlabel locali s 16014 9106 16222 9140 6 VSS
port 42 nsew
rlabel locali s 17118 9140 17337 9622 6 VSS
port 42 nsew
rlabel locali s 16814 9622 17337 9656 6 VSS
port 42 nsew
rlabel locali s 16014 9622 16222 9656 6 VSS
port 42 nsew
rlabel locali s 69244 9668 92336 9682 6 VSS
port 42 nsew
rlabel locali s 92302 9682 92336 10012 6 VSS
port 42 nsew
rlabel locali s 69244 9682 69278 10012 6 VSS
port 42 nsew
rlabel locali s 69244 10012 92336 10046 6 VSS
port 42 nsew
rlabel locali s 17118 9656 17337 10138 6 VSS
port 42 nsew
rlabel locali s 16814 10138 17337 10172 6 VSS
port 42 nsew
rlabel locali s 16014 10138 16222 10172 6 VSS
port 42 nsew
rlabel locali s 17118 10172 17337 10250 6 VSS
port 42 nsew
rlabel locali s 17125 10250 17315 11350 6 VSS
port 42 nsew
rlabel locali s 16949 11350 17315 13005 6 VSS
port 42 nsew
rlabel locali s 16949 13005 17282 16839 6 VSS
port 42 nsew
rlabel locali s -2105 8544 -746 44258 4 VSS
port 42 nsew
rlabel locali s -16182 8210 -15355 8555 4 VSS
port 42 nsew
rlabel locali s -7015 9941 -6799 10002 4 VSS
port 42 nsew
rlabel locali s -12587 9941 -12450 9999 4 VSS
port 42 nsew
rlabel locali s -6818 10575 -6753 10673 4 VSS
port 42 nsew
rlabel locali s -6818 10673 -6256 10707 4 VSS
port 42 nsew
rlabel locali s -6818 10707 -6753 11520 4 VSS
port 42 nsew
rlabel locali s -6818 11520 -6664 11705 4 VSS
port 42 nsew
rlabel locali s -6818 11705 -6357 11739 4 VSS
port 42 nsew
rlabel locali s -6818 11739 -6664 11849 4 VSS
port 42 nsew
rlabel locali s -6171 12259 -6113 12396 4 VSS
port 42 nsew
rlabel locali s -6166 12396 -6130 12469 4 VSS
port 42 nsew
rlabel locali s -6168 12469 -6128 12489 4 VSS
port 42 nsew
rlabel locali s -6176 12489 -6122 12624 4 VSS
port 42 nsew
rlabel locali s -6816 11849 -6664 12671 4 VSS
port 42 nsew
rlabel locali s -7013 10002 -6977 12229 4 VSS
port 42 nsew
rlabel locali s -8515 10057 -8278 10074 4 VSS
port 42 nsew
rlabel locali s -8515 10074 -8133 10114 4 VSS
port 42 nsew
rlabel locali s -8077 10200 -7840 10260 4 VSS
port 42 nsew
rlabel locali s -8075 10260 -8039 10527 4 VSS
port 42 nsew
rlabel locali s -8077 10527 -8037 10547 4 VSS
port 42 nsew
rlabel locali s -8085 10547 -8031 10682 4 VSS
port 42 nsew
rlabel locali s -8173 10114 -8133 10600 4 VSS
port 42 nsew
rlabel locali s -8515 10114 -8278 10117 4 VSS
port 42 nsew
rlabel locali s -8175 10600 -8133 10601 4 VSS
port 42 nsew
rlabel locali s -8175 10601 -8135 10671 4 VSS
port 42 nsew
rlabel locali s -8174 10671 -8135 11012 4 VSS
port 42 nsew
rlabel locali s -8638 10612 -8577 10729 4 VSS
port 42 nsew
rlabel locali s -8638 10729 -8525 10730 4 VSS
port 42 nsew
rlabel locali s -8638 10730 -8217 10764 4 VSS
port 42 nsew
rlabel locali s -8180 11012 -8109 11086 4 VSS
port 42 nsew
rlabel locali s -8638 10764 -8577 11053 4 VSS
port 42 nsew
rlabel locali s -12288 10655 -12138 10790 4 VSS
port 42 nsew
rlabel locali s -12288 10790 -12009 10795 4 VSS
port 42 nsew
rlabel locali s -12288 10795 -11838 10829 4 VSS
port 42 nsew
rlabel locali s -12288 10829 -12009 10838 4 VSS
port 42 nsew
rlabel locali s -12288 10838 -12138 10984 4 VSS
port 42 nsew
rlabel locali s -12288 10984 -12006 10991 4 VSS
port 42 nsew
rlabel locali s -12288 10991 -11838 11025 4 VSS
port 42 nsew
rlabel locali s -12288 11025 -12006 11032 4 VSS
port 42 nsew
rlabel locali s -8674 11053 -8577 11054 4 VSS
port 42 nsew
rlabel locali s -8152 11199 -8066 11339 4 VSS
port 42 nsew
rlabel locali s -8152 11339 -7910 11373 4 VSS
port 42 nsew
rlabel locali s -8152 11373 -8066 11443 4 VSS
port 42 nsew
rlabel locali s -8674 11054 -8559 11443 4 VSS
port 42 nsew
rlabel locali s -12288 11032 -12138 11313 4 VSS
port 42 nsew
rlabel locali s -8674 11443 -8066 11504 4 VSS
port 42 nsew
rlabel locali s -8152 11504 -8066 11535 4 VSS
port 42 nsew
rlabel locali s -8152 11535 -7910 11569 4 VSS
port 42 nsew
rlabel locali s -8152 11569 -8066 11814 4 VSS
port 42 nsew
rlabel locali s -8674 11504 -8559 12108 4 VSS
port 42 nsew
rlabel locali s -12288 11313 -11841 11429 4 VSS
port 42 nsew
rlabel locali s -11540 11798 -11403 11856 4 VSS
port 42 nsew
rlabel locali s -11452 11856 -11416 11907 4 VSS
port 42 nsew
rlabel locali s -11957 11429 -11841 11868 4 VSS
port 42 nsew
rlabel locali s -12288 11429 -12138 11459 4 VSS
port 42 nsew
rlabel locali s -12261 11459 -12155 11543 4 VSS
port 42 nsew
rlabel locali s -12494 9999 -12453 11796 4 VSS
port 42 nsew
rlabel locali s -12668 10055 -12531 10113 4 VSS
port 42 nsew
rlabel locali s -12494 11796 -12357 11854 4 VSS
port 42 nsew
rlabel locali s -11460 11907 -11400 12053 4 VSS
port 42 nsew
rlabel locali s -11957 11868 -11806 11997 4 VSS
port 42 nsew
rlabel locali s -11957 11997 -11654 12001 4 VSS
port 42 nsew
rlabel locali s -11957 12001 -11495 12035 4 VSS
port 42 nsew
rlabel locali s -11957 12035 -11654 12041 4 VSS
port 42 nsew
rlabel locali s -8817 12108 -8559 12223 4 VSS
port 42 nsew
rlabel locali s -11957 12041 -11806 12191 4 VSS
port 42 nsew
rlabel locali s -11957 12191 -11655 12197 4 VSS
port 42 nsew
rlabel locali s -7013 12229 -6881 12282 4 VSS
port 42 nsew
rlabel locali s -8817 12223 -8692 12405 4 VSS
port 42 nsew
rlabel locali s -11957 12197 -11495 12231 4 VSS
port 42 nsew
rlabel locali s -11957 12231 -11655 12235 4 VSS
port 42 nsew
rlabel locali s -8817 12405 -8689 12503 4 VSS
port 42 nsew
rlabel locali s -11957 12235 -11806 12465 4 VSS
port 42 nsew
rlabel locali s -8817 12503 -8192 12537 4 VSS
port 42 nsew
rlabel locali s -6816 12671 -6616 12672 4 VSS
port 42 nsew
rlabel locali s -6816 12672 -6308 12706 4 VSS
port 42 nsew
rlabel locali s -6816 12706 -6664 12996 4 VSS
port 42 nsew
rlabel locali s -6243 13141 -6157 13281 4 VSS
port 42 nsew
rlabel locali s -6243 13281 -6001 13315 4 VSS
port 42 nsew
rlabel locali s -6243 13315 -6157 13385 4 VSS
port 42 nsew
rlabel locali s -6816 12996 -6650 13385 4 VSS
port 42 nsew
rlabel locali s -8817 12537 -8689 13334 4 VSS
port 42 nsew
rlabel locali s -11370 12639 -11233 12697 4 VSS
port 42 nsew
rlabel locali s -11364 12697 -11328 13035 4 VSS
port 42 nsew
rlabel locali s -11542 12716 -11405 12774 4 VSS
port 42 nsew
rlabel locali s -11957 12465 -11841 12773 4 VSS
port 42 nsew
rlabel locali s -12573 10113 -12532 12617 4 VSS
port 42 nsew
rlabel locali s -12573 12617 -12436 12675 4 VSS
port 42 nsew
rlabel locali s -12746 10200 -12609 10258 4 VSS
port 42 nsew
rlabel locali s -12650 10258 -12609 12710 4 VSS
port 42 nsew
rlabel locali s -15496 8555 -15355 10372 4 VSS
port 42 nsew
rlabel locali s -12815 10442 -12700 10556 4 VSS
port 42 nsew
rlabel locali s -13192 10556 -12700 10590 4 VSS
port 42 nsew
rlabel locali s -12815 10590 -12700 11425 4 VSS
port 42 nsew
rlabel locali s -12796 11425 -12731 11588 4 VSS
port 42 nsew
rlabel locali s -13293 11588 -12731 11622 4 VSS
port 42 nsew
rlabel locali s -12796 11622 -12731 11720 4 VSS
port 42 nsew
rlabel locali s -12650 12710 -12513 12768 4 VSS
port 42 nsew
rlabel locali s -11453 12774 -11417 12812 4 VSS
port 42 nsew
rlabel locali s -11461 12812 -11401 12958 4 VSS
port 42 nsew
rlabel locali s -11957 12773 -11807 12902 4 VSS
port 42 nsew
rlabel locali s -11957 12902 -11655 12906 4 VSS
port 42 nsew
rlabel locali s -11957 12906 -11496 12940 4 VSS
port 42 nsew
rlabel locali s -11957 12940 -11655 12946 4 VSS
port 42 nsew
rlabel locali s -11381 13035 -11321 13178 4 VSS
port 42 nsew
rlabel locali s -11957 12946 -11807 13096 4 VSS
port 42 nsew
rlabel locali s -11957 13096 -11656 13102 4 VSS
port 42 nsew
rlabel locali s -11957 13102 -11496 13136 4 VSS
port 42 nsew
rlabel locali s -11957 13136 -11656 13140 4 VSS
port 42 nsew
rlabel locali s -11957 13140 -11807 13154 4 VSS
port 42 nsew
rlabel locali s -11896 13154 -11807 13291 4 VSS
port 42 nsew
rlabel locali s -6816 13385 -6157 13446 4 VSS
port 42 nsew
rlabel locali s -6243 13446 -6157 13477 4 VSS
port 42 nsew
rlabel locali s -6816 13446 -6664 13476 4 VSS
port 42 nsew
rlabel locali s -6243 13477 -6001 13511 4 VSS
port 42 nsew
rlabel locali s -6243 13511 -6157 13714 4 VSS
port 42 nsew
rlabel locali s -8817 13334 -8662 13535 4 VSS
port 42 nsew
rlabel locali s -8817 13535 -8293 13569 4 VSS
port 42 nsew
rlabel locali s -6245 13714 -6101 13775 4 VSS
port 42 nsew
rlabel locali s -6162 13775 -6101 14190 4 VSS
port 42 nsew
rlabel locali s -6162 14190 -6083 14307 4 VSS
port 42 nsew
rlabel locali s -6196 14307 -6083 14308 4 VSS
port 42 nsew
rlabel locali s -6504 14308 -6083 14342 4 VSS
port 42 nsew
rlabel locali s -8434 14194 -8348 14334 4 VSS
port 42 nsew
rlabel locali s -6162 14342 -6083 14639 4 VSS
port 42 nsew
rlabel locali s -8434 14334 -8092 14368 4 VSS
port 42 nsew
rlabel locali s -8434 14368 -8348 14530 4 VSS
port 42 nsew
rlabel locali s -8434 14530 -8092 14564 4 VSS
port 42 nsew
rlabel locali s -6162 14639 -6101 15021 4 VSS
port 42 nsew
rlabel locali s -6655 14777 -6569 14917 4 VSS
port 42 nsew
rlabel locali s -6811 14917 -6569 14951 4 VSS
port 42 nsew
rlabel locali s -6655 14951 -6569 15021 4 VSS
port 42 nsew
rlabel locali s -6655 15021 -5693 15082 4 VSS
port 42 nsew
rlabel locali s -5806 15082 -5693 15748 4 VSS
port 42 nsew
rlabel locali s -6655 15082 -6569 15113 4 VSS
port 42 nsew
rlabel locali s -8434 14564 -8348 15046 4 VSS
port 42 nsew
rlabel locali s -8601 15046 -8348 15082 4 VSS
port 42 nsew
rlabel locali s -8817 13569 -8662 15082 4 VSS
port 42 nsew
rlabel locali s -11896 13291 -11520 13352 4 VSS
port 42 nsew
rlabel locali s -11581 13352 -11520 13678 4 VSS
port 42 nsew
rlabel locali s -11896 13352 -11807 13370 4 VSS
port 42 nsew
rlabel locali s -11581 13678 -11101 13739 4 VSS
port 42 nsew
rlabel locali s -11162 13739 -11101 14190 4 VSS
port 42 nsew
rlabel locali s -11162 14190 -11083 14307 4 VSS
port 42 nsew
rlabel locali s -11196 14307 -11083 14308 4 VSS
port 42 nsew
rlabel locali s -11504 14308 -11083 14342 4 VSS
port 42 nsew
rlabel locali s -13434 14194 -13348 14334 4 VSS
port 42 nsew
rlabel locali s -11162 14342 -11083 14639 4 VSS
port 42 nsew
rlabel locali s -13434 14334 -13092 14368 4 VSS
port 42 nsew
rlabel locali s -13434 14368 -13348 14530 4 VSS
port 42 nsew
rlabel locali s -13434 14530 -13092 14564 4 VSS
port 42 nsew
rlabel locali s -11162 14639 -11101 15021 4 VSS
port 42 nsew
rlabel locali s -11655 14777 -11569 14917 4 VSS
port 42 nsew
rlabel locali s -11811 14917 -11569 14951 4 VSS
port 42 nsew
rlabel locali s -11655 14951 -11569 15021 4 VSS
port 42 nsew
rlabel locali s -6811 15113 -6569 15147 4 VSS
port 42 nsew
rlabel locali s -8817 15082 -8348 15132 4 VSS
port 42 nsew
rlabel locali s -6655 15147 -6569 15392 4 VSS
port 42 nsew
rlabel locali s -8817 15132 -8515 15292 4 VSS
port 42 nsew
rlabel locali s -11655 15021 -10693 15082 4 VSS
port 42 nsew
rlabel locali s -8601 15292 -8515 15306 4 VSS
port 42 nsew
rlabel locali s -8601 15306 -8478 15307 4 VSS
port 42 nsew
rlabel locali s -8601 15307 -8170 15341 4 VSS
port 42 nsew
rlabel locali s -8601 15341 -8515 15631 4 VSS
port 42 nsew
rlabel locali s -8601 15631 -8512 15711 4 VSS
port 42 nsew
rlabel locali s -5924 15748 -5693 15755 4 VSS
port 42 nsew
rlabel locali s -6218 15755 -5693 15789 4 VSS
port 42 nsew
rlabel locali s -5924 15789 -5693 15795 4 VSS
port 42 nsew
rlabel locali s -5806 15795 -5693 15944 4 VSS
port 42 nsew
rlabel locali s -8105 15776 -8019 15916 4 VSS
port 42 nsew
rlabel locali s -5925 15944 -5693 15951 4 VSS
port 42 nsew
rlabel locali s -8105 15916 -7863 15950 4 VSS
port 42 nsew
rlabel locali s -6218 15951 -5693 15985 4 VSS
port 42 nsew
rlabel locali s -5925 15985 -5693 15991 4 VSS
port 42 nsew
rlabel locali s -5806 15991 -5693 16186 4 VSS
port 42 nsew
rlabel locali s -8105 15950 -8019 16020 4 VSS
port 42 nsew
rlabel locali s -8573 15711 -8512 16020 4 VSS
port 42 nsew
rlabel locali s -8573 16020 -8019 16081 4 VSS
port 42 nsew
rlabel locali s -10806 15082 -10693 15748 4 VSS
port 42 nsew
rlabel locali s -11655 15082 -11569 15113 4 VSS
port 42 nsew
rlabel locali s -13434 14564 -13348 15046 4 VSS
port 42 nsew
rlabel locali s -11811 15113 -11569 15147 4 VSS
port 42 nsew
rlabel locali s -13601 15046 -13348 15132 4 VSS
port 42 nsew
rlabel locali s -11655 15147 -11569 15392 4 VSS
port 42 nsew
rlabel locali s -13601 15132 -13515 15306 4 VSS
port 42 nsew
rlabel locali s -13601 15306 -13478 15307 4 VSS
port 42 nsew
rlabel locali s -13601 15307 -13170 15341 4 VSS
port 42 nsew
rlabel locali s -13601 15341 -13515 15631 4 VSS
port 42 nsew
rlabel locali s -13601 15631 -13512 15711 4 VSS
port 42 nsew
rlabel locali s -10924 15748 -10693 15755 4 VSS
port 42 nsew
rlabel locali s -11218 15755 -10693 15789 4 VSS
port 42 nsew
rlabel locali s -10924 15789 -10693 15795 4 VSS
port 42 nsew
rlabel locali s -10806 15795 -10693 15944 4 VSS
port 42 nsew
rlabel locali s -13105 15776 -13019 15916 4 VSS
port 42 nsew
rlabel locali s -10925 15944 -10693 15951 4 VSS
port 42 nsew
rlabel locali s -13105 15916 -12863 15950 4 VSS
port 42 nsew
rlabel locali s -11218 15951 -10693 15985 4 VSS
port 42 nsew
rlabel locali s -10925 15985 -10693 15991 4 VSS
port 42 nsew
rlabel locali s -8105 16081 -8019 16112 4 VSS
port 42 nsew
rlabel locali s -8105 16112 -7863 16146 4 VSS
port 42 nsew
rlabel locali s -5935 16186 -5693 16193 4 VSS
port 42 nsew
rlabel locali s -6218 16193 -5693 16227 4 VSS
port 42 nsew
rlabel locali s -5935 16227 -5693 16233 4 VSS
port 42 nsew
rlabel locali s -5806 16233 -5693 16498 4 VSS
port 42 nsew
rlabel locali s -8105 16146 -8019 16561 4 VSS
port 42 nsew
rlabel locali s -10806 15991 -10693 16186 4 VSS
port 42 nsew
rlabel locali s -13105 15950 -13019 16020 4 VSS
port 42 nsew
rlabel locali s -13573 15711 -13512 16020 4 VSS
port 42 nsew
rlabel locali s -13573 16020 -13019 16081 4 VSS
port 42 nsew
rlabel locali s -13105 16081 -13019 16112 4 VSS
port 42 nsew
rlabel locali s -13105 16112 -12863 16146 4 VSS
port 42 nsew
rlabel locali s -10935 16186 -10693 16193 4 VSS
port 42 nsew
rlabel locali s -11218 16193 -10693 16227 4 VSS
port 42 nsew
rlabel locali s -10935 16227 -10693 16233 4 VSS
port 42 nsew
rlabel locali s -10806 16233 -10693 16498 4 VSS
port 42 nsew
rlabel locali s -13105 16146 -13019 16561 4 VSS
port 42 nsew
rlabel locali s -5469 18165 -5401 18174 4 VSS
port 42 nsew
rlabel locali s -5469 18174 -5242 18208 4 VSS
port 42 nsew
rlabel locali s -5469 18208 -5401 18370 4 VSS
port 42 nsew
rlabel locali s -5469 18370 -5242 18404 4 VSS
port 42 nsew
rlabel locali s -5849 18173 -5781 18272 4 VSS
port 42 nsew
rlabel locali s -10396 18165 -10328 18174 4 VSS
port 42 nsew
rlabel locali s -10396 18174 -10169 18208 4 VSS
port 42 nsew
rlabel locali s -6008 18272 -5781 18306 4 VSS
port 42 nsew
rlabel locali s -5556 18385 -5517 18402 4 VSS
port 42 nsew
rlabel locali s -5469 18404 -5401 18413 4 VSS
port 42 nsew
rlabel locali s -5569 18402 -5509 18413 4 VSS
port 42 nsew
rlabel locali s -5569 18413 -5401 18524 4 VSS
port 42 nsew
rlabel locali s -5469 18524 -5401 18566 4 VSS
port 42 nsew
rlabel locali s -5569 18524 -5509 18539 4 VSS
port 42 nsew
rlabel locali s -5849 18306 -5781 18468 4 VSS
port 42 nsew
rlabel locali s -10396 18208 -10328 18370 4 VSS
port 42 nsew
rlabel locali s -10396 18370 -10169 18404 4 VSS
port 42 nsew
rlabel locali s -10776 18173 -10708 18272 4 VSS
port 42 nsew
rlabel locali s -10935 18272 -10708 18306 4 VSS
port 42 nsew
rlabel locali s -10483 18385 -10444 18402 4 VSS
port 42 nsew
rlabel locali s -10396 18404 -10328 18413 4 VSS
port 42 nsew
rlabel locali s -10496 18402 -10436 18413 4 VSS
port 42 nsew
rlabel locali s -6008 18468 -5781 18502 4 VSS
port 42 nsew
rlabel locali s -5469 18566 -5242 18600 4 VSS
port 42 nsew
rlabel locali s -5469 18600 -5401 19011 4 VSS
port 42 nsew
rlabel locali s -5469 19011 -5242 19045 4 VSS
port 42 nsew
rlabel locali s -5469 19045 -5401 19207 4 VSS
port 42 nsew
rlabel locali s -5469 19207 -5242 19224 4 VSS
port 42 nsew
rlabel locali s -5556 18539 -5517 19224 4 VSS
port 42 nsew
rlabel locali s -5849 18502 -5781 18664 4 VSS
port 42 nsew
rlabel locali s -10496 18413 -10328 18524 4 VSS
port 42 nsew
rlabel locali s -10396 18524 -10328 18566 4 VSS
port 42 nsew
rlabel locali s -10496 18524 -10436 18539 4 VSS
port 42 nsew
rlabel locali s -10776 18306 -10708 18468 4 VSS
port 42 nsew
rlabel locali s -10935 18468 -10708 18502 4 VSS
port 42 nsew
rlabel locali s -10396 18566 -10169 18600 4 VSS
port 42 nsew
rlabel locali s -6008 18664 -5781 18698 4 VSS
port 42 nsew
rlabel locali s -5849 18698 -5781 18707 4 VSS
port 42 nsew
rlabel locali s -10396 18600 -10328 19011 4 VSS
port 42 nsew
rlabel locali s -10396 19011 -10169 19045 4 VSS
port 42 nsew
rlabel locali s -5556 19224 -5242 19241 4 VSS
port 42 nsew
rlabel locali s -5556 19241 -5401 19335 4 VSS
port 42 nsew
rlabel locali s -5469 19335 -5401 19403 4 VSS
port 42 nsew
rlabel locali s -5469 19403 -5242 19437 4 VSS
port 42 nsew
rlabel locali s -5469 19437 -5401 19536 4 VSS
port 42 nsew
rlabel locali s -5469 20865 -5401 20874 4 VSS
port 42 nsew
rlabel locali s -5469 20874 -5242 20908 4 VSS
port 42 nsew
rlabel locali s -5469 20908 -5401 21022 4 VSS
port 42 nsew
rlabel locali s -5556 19335 -5517 20999 4 VSS
port 42 nsew
rlabel locali s -7120 19179 -7059 19296 4 VSS
port 42 nsew
rlabel locali s -7172 19296 -7059 19297 4 VSS
port 42 nsew
rlabel locali s -7480 19297 -7059 19331 4 VSS
port 42 nsew
rlabel locali s -9410 19183 -9324 19323 4 VSS
port 42 nsew
rlabel locali s -10396 19045 -10328 19207 4 VSS
port 42 nsew
rlabel locali s -10396 19207 -10169 19224 4 VSS
port 42 nsew
rlabel locali s -10483 18539 -10444 19224 4 VSS
port 42 nsew
rlabel locali s -10776 18502 -10708 18664 4 VSS
port 42 nsew
rlabel locali s -10935 18664 -10708 18698 4 VSS
port 42 nsew
rlabel locali s -10776 18698 -10708 18707 4 VSS
port 42 nsew
rlabel locali s -10483 19224 -10169 19241 4 VSS
port 42 nsew
rlabel locali s -7120 19331 -7059 19621 4 VSS
port 42 nsew
rlabel locali s -9410 19323 -9068 19357 4 VSS
port 42 nsew
rlabel locali s -9410 19357 -9324 19519 4 VSS
port 42 nsew
rlabel locali s -10483 19241 -10328 19335 4 VSS
port 42 nsew
rlabel locali s -10396 19335 -10328 19403 4 VSS
port 42 nsew
rlabel locali s -10396 19403 -10169 19437 4 VSS
port 42 nsew
rlabel locali s -9410 19519 -9068 19553 4 VSS
port 42 nsew
rlabel locali s -10396 19437 -10328 19536 4 VSS
port 42 nsew
rlabel locali s -7138 19621 -7059 19628 4 VSS
port 42 nsew
rlabel locali s -5849 19916 -5781 20015 4 VSS
port 42 nsew
rlabel locali s -7138 19628 -7077 20010 4 VSS
port 42 nsew
rlabel locali s -7631 19766 -7545 19906 4 VSS
port 42 nsew
rlabel locali s -7787 19906 -7545 19940 4 VSS
port 42 nsew
rlabel locali s -7631 19940 -7545 20010 4 VSS
port 42 nsew
rlabel locali s -6008 20015 -5781 20049 4 VSS
port 42 nsew
rlabel locali s -5849 20049 -5781 20211 4 VSS
port 42 nsew
rlabel locali s -7631 20010 -6669 20071 4 VSS
port 42 nsew
rlabel locali s -6008 20211 -5781 20245 4 VSS
port 42 nsew
rlabel locali s -5849 20245 -5781 20407 4 VSS
port 42 nsew
rlabel locali s -6008 20407 -5781 20441 4 VSS
port 42 nsew
rlabel locali s -5849 20441 -5781 20972 4 VSS
port 42 nsew
rlabel locali s -6782 20071 -6669 20737 4 VSS
port 42 nsew
rlabel locali s -7631 20071 -7545 20102 4 VSS
port 42 nsew
rlabel locali s -9410 19553 -9324 20035 4 VSS
port 42 nsew
rlabel locali s -7787 20102 -7545 20136 4 VSS
port 42 nsew
rlabel locali s -9577 20035 -9324 20121 4 VSS
port 42 nsew
rlabel locali s -7631 20136 -7545 20381 4 VSS
port 42 nsew
rlabel locali s -9577 20121 -9491 20295 4 VSS
port 42 nsew
rlabel locali s -9577 20295 -9454 20296 4 VSS
port 42 nsew
rlabel locali s -9577 20296 -9146 20330 4 VSS
port 42 nsew
rlabel locali s -9577 20330 -9491 20620 4 VSS
port 42 nsew
rlabel locali s -9577 20620 -9488 20700 4 VSS
port 42 nsew
rlabel locali s -6900 20737 -6669 20744 4 VSS
port 42 nsew
rlabel locali s -7194 20744 -6669 20778 4 VSS
port 42 nsew
rlabel locali s -6900 20778 -6669 20784 4 VSS
port 42 nsew
rlabel locali s -6782 20784 -6669 20933 4 VSS
port 42 nsew
rlabel locali s -9081 20765 -8995 20905 4 VSS
port 42 nsew
rlabel locali s -6901 20933 -6669 20940 4 VSS
port 42 nsew
rlabel locali s -9081 20905 -8839 20939 4 VSS
port 42 nsew
rlabel locali s -5575 20999 -5515 21022 4 VSS
port 42 nsew
rlabel locali s -5575 21022 -5401 21070 4 VSS
port 42 nsew
rlabel locali s -5575 21070 -5242 21104 4 VSS
port 42 nsew
rlabel locali s -5575 21104 -5401 21133 4 VSS
port 42 nsew
rlabel locali s -5469 21133 -5401 21205 4 VSS
port 42 nsew
rlabel locali s -5575 21133 -5515 21136 4 VSS
port 42 nsew
rlabel locali s -6008 20972 -5781 21006 4 VSS
port 42 nsew
rlabel locali s -7194 20940 -6669 20974 4 VSS
port 42 nsew
rlabel locali s -6901 20974 -6669 20980 4 VSS
port 42 nsew
rlabel locali s -5471 21205 -5401 21266 4 VSS
port 42 nsew
rlabel locali s -5471 21266 -5242 21300 4 VSS
port 42 nsew
rlabel locali s -5471 21300 -5401 21399 4 VSS
port 42 nsew
rlabel locali s -5471 21399 -5403 21702 4 VSS
port 42 nsew
rlabel locali s -5471 21702 -5401 21711 4 VSS
port 42 nsew
rlabel locali s -5471 21711 -5242 21725 4 VSS
port 42 nsew
rlabel locali s -5469 21725 -5242 21745 4 VSS
port 42 nsew
rlabel locali s -5469 21745 -5401 21900 4 VSS
port 42 nsew
rlabel locali s -5556 21136 -5517 21900 4 VSS
port 42 nsew
rlabel locali s -5849 21006 -5781 21168 4 VSS
port 42 nsew
rlabel locali s -6008 21168 -5781 21202 4 VSS
port 42 nsew
rlabel locali s -6782 20980 -6669 21175 4 VSS
port 42 nsew
rlabel locali s -9081 20939 -8995 21009 4 VSS
port 42 nsew
rlabel locali s -9549 20700 -9488 21009 4 VSS
port 42 nsew
rlabel locali s -10396 20865 -10328 20874 4 VSS
port 42 nsew
rlabel locali s -10396 20874 -10169 20908 4 VSS
port 42 nsew
rlabel locali s -9549 21009 -8995 21070 4 VSS
port 42 nsew
rlabel locali s -10396 20908 -10328 21022 4 VSS
port 42 nsew
rlabel locali s -10483 19335 -10444 20999 4 VSS
port 42 nsew
rlabel locali s -10776 19916 -10708 20015 4 VSS
port 42 nsew
rlabel locali s -10935 20015 -10708 20049 4 VSS
port 42 nsew
rlabel locali s -10776 20049 -10708 20211 4 VSS
port 42 nsew
rlabel locali s -10935 20211 -10708 20245 4 VSS
port 42 nsew
rlabel locali s -10776 20245 -10708 20407 4 VSS
port 42 nsew
rlabel locali s -10935 20407 -10708 20441 4 VSS
port 42 nsew
rlabel locali s -10776 20441 -10708 20972 4 VSS
port 42 nsew
rlabel locali s -10502 20999 -10442 21022 4 VSS
port 42 nsew
rlabel locali s -10502 21022 -10328 21070 4 VSS
port 42 nsew
rlabel locali s -9081 21070 -8995 21101 4 VSS
port 42 nsew
rlabel locali s -9081 21101 -8839 21135 4 VSS
port 42 nsew
rlabel locali s -10502 21070 -10169 21104 4 VSS
port 42 nsew
rlabel locali s -6911 21175 -6669 21182 4 VSS
port 42 nsew
rlabel locali s -5849 21202 -5781 21364 4 VSS
port 42 nsew
rlabel locali s -7194 21182 -6669 21216 4 VSS
port 42 nsew
rlabel locali s -6911 21216 -6669 21222 4 VSS
port 42 nsew
rlabel locali s -6008 21364 -5781 21398 4 VSS
port 42 nsew
rlabel locali s -5849 21398 -5781 21407 4 VSS
port 42 nsew
rlabel locali s -6782 21222 -6669 21487 4 VSS
port 42 nsew
rlabel locali s -9081 21135 -8995 21550 4 VSS
port 42 nsew
rlabel locali s -10502 21104 -10328 21133 4 VSS
port 42 nsew
rlabel locali s -10396 21133 -10328 21205 4 VSS
port 42 nsew
rlabel locali s -10502 21133 -10442 21136 4 VSS
port 42 nsew
rlabel locali s -10935 20972 -10708 21006 4 VSS
port 42 nsew
rlabel locali s -10398 21205 -10328 21266 4 VSS
port 42 nsew
rlabel locali s -10398 21266 -10169 21300 4 VSS
port 42 nsew
rlabel locali s -10398 21300 -10328 21399 4 VSS
port 42 nsew
rlabel locali s -10398 21399 -10330 21702 4 VSS
port 42 nsew
rlabel locali s -10398 21702 -10328 21711 4 VSS
port 42 nsew
rlabel locali s -10398 21711 -10169 21725 4 VSS
port 42 nsew
rlabel locali s -10396 21725 -10169 21745 4 VSS
port 42 nsew
rlabel locali s -5556 21900 -5401 21907 4 VSS
port 42 nsew
rlabel locali s -10396 21745 -10328 21900 4 VSS
port 42 nsew
rlabel locali s -10483 21136 -10444 21900 4 VSS
port 42 nsew
rlabel locali s -10776 21006 -10708 21168 4 VSS
port 42 nsew
rlabel locali s -10935 21168 -10708 21202 4 VSS
port 42 nsew
rlabel locali s -10776 21202 -10708 21364 4 VSS
port 42 nsew
rlabel locali s -10935 21364 -10708 21398 4 VSS
port 42 nsew
rlabel locali s -10776 21398 -10708 21407 4 VSS
port 42 nsew
rlabel locali s -10483 21900 -10328 21907 4 VSS
port 42 nsew
rlabel locali s -5556 21907 -5242 21941 4 VSS
port 42 nsew
rlabel locali s -10483 21907 -10169 21941 4 VSS
port 42 nsew
rlabel locali s -5556 21941 -5401 22011 4 VSS
port 42 nsew
rlabel locali s -5469 22011 -5401 22103 4 VSS
port 42 nsew
rlabel locali s -5469 22103 -5242 22137 4 VSS
port 42 nsew
rlabel locali s -5469 22137 -5401 22236 4 VSS
port 42 nsew
rlabel locali s -5556 22011 -5517 23637 4 VSS
port 42 nsew
rlabel locali s -10483 21941 -10328 22011 4 VSS
port 42 nsew
rlabel locali s -10396 22011 -10328 22103 4 VSS
port 42 nsew
rlabel locali s -10396 22103 -10169 22137 4 VSS
port 42 nsew
rlabel locali s -10396 22137 -10328 22236 4 VSS
port 42 nsew
rlabel locali s -5849 22616 -5781 22715 4 VSS
port 42 nsew
rlabel locali s -6008 22715 -5781 22749 4 VSS
port 42 nsew
rlabel locali s -5849 22749 -5781 22911 4 VSS
port 42 nsew
rlabel locali s -6008 22911 -5781 22945 4 VSS
port 42 nsew
rlabel locali s -5849 22945 -5781 23107 4 VSS
port 42 nsew
rlabel locali s -6008 23107 -5781 23141 4 VSS
port 42 nsew
rlabel locali s -5849 23141 -5781 23597 4 VSS
port 42 nsew
rlabel locali s -6008 23597 -5781 23631 4 VSS
port 42 nsew
rlabel locali s -5575 23637 -5515 23769 4 VSS
port 42 nsew
rlabel locali s -5556 23769 -5517 23770 4 VSS
port 42 nsew
rlabel locali s -5849 23631 -5781 23793 4 VSS
port 42 nsew
rlabel locali s -10483 22011 -10444 23637 4 VSS
port 42 nsew
rlabel locali s -10776 22616 -10708 22715 4 VSS
port 42 nsew
rlabel locali s -10935 22715 -10708 22749 4 VSS
port 42 nsew
rlabel locali s -10776 22749 -10708 22911 4 VSS
port 42 nsew
rlabel locali s -10935 22911 -10708 22945 4 VSS
port 42 nsew
rlabel locali s -10776 22945 -10708 23107 4 VSS
port 42 nsew
rlabel locali s -10935 23107 -10708 23141 4 VSS
port 42 nsew
rlabel locali s -10776 23141 -10708 23597 4 VSS
port 42 nsew
rlabel locali s -10935 23597 -10708 23631 4 VSS
port 42 nsew
rlabel locali s -10502 23637 -10442 23769 4 VSS
port 42 nsew
rlabel locali s -10483 23769 -10444 23770 4 VSS
port 42 nsew
rlabel locali s -10776 23631 -10708 23793 4 VSS
port 42 nsew
rlabel locali s -6008 23793 -5781 23827 4 VSS
port 42 nsew
rlabel locali s -10935 23793 -10708 23827 4 VSS
port 42 nsew
rlabel locali s -5849 23827 -5781 23989 4 VSS
port 42 nsew
rlabel locali s -10776 23827 -10708 23989 4 VSS
port 42 nsew
rlabel locali s -6008 23989 -5781 24023 4 VSS
port 42 nsew
rlabel locali s -10935 23989 -10708 24023 4 VSS
port 42 nsew
rlabel locali s -5849 24023 -5781 24032 4 VSS
port 42 nsew
rlabel locali s -10776 24023 -10708 24032 4 VSS
port 42 nsew
rlabel locali s -6279 24189 -6196 24467 4 VSS
port 42 nsew
rlabel locali s -6279 24467 -6197 24613 4 VSS
port 42 nsew
rlabel locali s -6279 24613 -6067 24619 4 VSS
port 42 nsew
rlabel locali s -6279 24619 -5784 24653 4 VSS
port 42 nsew
rlabel locali s -11213 24460 -11131 24640 4 VSS
port 42 nsew
rlabel locali s -11213 24640 -11001 24646 4 VSS
port 42 nsew
rlabel locali s -6279 24653 -6067 24660 4 VSS
port 42 nsew
rlabel locali s -6279 24660 -6197 24855 4 VSS
port 42 nsew
rlabel locali s -11213 24646 -10718 24680 4 VSS
port 42 nsew
rlabel locali s -11213 24680 -11001 24687 4 VSS
port 42 nsew
rlabel locali s -6279 24855 -6077 24861 4 VSS
port 42 nsew
rlabel locali s -6279 24861 -5784 24895 4 VSS
port 42 nsew
rlabel locali s -11213 24687 -11131 24882 4 VSS
port 42 nsew
rlabel locali s -11213 24882 -11011 24888 4 VSS
port 42 nsew
rlabel locali s -6279 24895 -6077 24902 4 VSS
port 42 nsew
rlabel locali s -6279 24902 -6197 25051 4 VSS
port 42 nsew
rlabel locali s -11213 24888 -10718 24922 4 VSS
port 42 nsew
rlabel locali s -11213 24922 -11011 24929 4 VSS
port 42 nsew
rlabel locali s -6279 25051 -6078 25057 4 VSS
port 42 nsew
rlabel locali s -6279 25057 -5784 25091 4 VSS
port 42 nsew
rlabel locali s -11213 24929 -11131 25078 4 VSS
port 42 nsew
rlabel locali s -11213 25078 -11012 25084 4 VSS
port 42 nsew
rlabel locali s -6279 25091 -6078 25098 4 VSS
port 42 nsew
rlabel locali s -6279 25098 -6197 25180 4 VSS
port 42 nsew
rlabel locali s -11213 25084 -10718 25118 4 VSS
port 42 nsew
rlabel locali s -11213 25118 -11012 25125 4 VSS
port 42 nsew
rlabel locali s -11213 25125 -11131 25589 4 VSS
port 42 nsew
rlabel locali s -11220 25589 -11125 25694 4 VSS
port 42 nsew
rlabel locali s -5681 25866 -5561 25868 4 VSS
port 42 nsew
rlabel locali s -6046 25864 -5870 25868 4 VSS
port 42 nsew
rlabel locali s -6046 25868 -5561 25902 4 VSS
port 42 nsew
rlabel locali s -5681 25902 -5561 25903 4 VSS
port 42 nsew
rlabel locali s -6046 25902 -5870 25903 4 VSS
port 42 nsew
rlabel locali s -5598 25903 -5561 26160 4 VSS
port 42 nsew
rlabel locali s -5659 26160 -5561 26197 4 VSS
port 42 nsew
rlabel locali s -5659 26197 -5622 26279 4 VSS
port 42 nsew
rlabel locali s -5680 26279 -5622 26282 4 VSS
port 42 nsew
rlabel locali s -5882 26282 -5622 26316 4 VSS
port 42 nsew
rlabel locali s -6046 25903 -5993 26296 4 VSS
port 42 nsew
rlabel locali s -13012 25864 -12836 25868 4 VSS
port 42 nsew
rlabel locali s -13321 25866 -13201 25868 4 VSS
port 42 nsew
rlabel locali s -13321 25868 -12836 25902 4 VSS
port 42 nsew
rlabel locali s -13012 25902 -12836 25903 4 VSS
port 42 nsew
rlabel locali s -13321 25902 -13201 25903 4 VSS
port 42 nsew
rlabel locali s -7907 26047 -7839 26146 4 VSS
port 42 nsew
rlabel locali s -7907 26146 -7680 26180 4 VSS
port 42 nsew
rlabel locali s -6066 26296 -5993 26305 4 VSS
port 42 nsew
rlabel locali s -6225 26305 -5993 26339 4 VSS
port 42 nsew
rlabel locali s -6066 26339 -5993 26501 4 VSS
port 42 nsew
rlabel locali s -7907 26180 -7839 26342 4 VSS
port 42 nsew
rlabel locali s -8287 26039 -8219 26048 4 VSS
port 42 nsew
rlabel locali s -10663 26039 -10595 26048 4 VSS
port 42 nsew
rlabel locali s -8446 26048 -8219 26082 4 VSS
port 42 nsew
rlabel locali s -10663 26048 -10436 26082 4 VSS
port 42 nsew
rlabel locali s -8287 26082 -8219 26244 4 VSS
port 42 nsew
rlabel locali s -10663 26082 -10595 26244 4 VSS
port 42 nsew
rlabel locali s -8171 26259 -8132 26276 4 VSS
port 42 nsew
rlabel locali s -7907 26342 -7680 26376 4 VSS
port 42 nsew
rlabel locali s -6225 26501 -5993 26535 4 VSS
port 42 nsew
rlabel locali s -6066 26535 -5993 26697 4 VSS
port 42 nsew
rlabel locali s -7907 26376 -7839 26538 4 VSS
port 42 nsew
rlabel locali s -8179 26276 -8119 26287 4 VSS
port 42 nsew
rlabel locali s -8446 26244 -8219 26278 4 VSS
port 42 nsew
rlabel locali s -10663 26244 -10436 26278 4 VSS
port 42 nsew
rlabel locali s -11043 26047 -10975 26146 4 VSS
port 42 nsew
rlabel locali s -11202 26146 -10975 26180 4 VSS
port 42 nsew
rlabel locali s -10750 26259 -10711 26276 4 VSS
port 42 nsew
rlabel locali s -8287 26278 -8219 26287 4 VSS
port 42 nsew
rlabel locali s -8287 26287 -8119 26398 4 VSS
port 42 nsew
rlabel locali s -8179 26398 -8119 26413 4 VSS
port 42 nsew
rlabel locali s -7907 26538 -7680 26572 4 VSS
port 42 nsew
rlabel locali s -7907 26572 -7839 26581 4 VSS
port 42 nsew
rlabel locali s -6225 26697 -5993 26731 4 VSS
port 42 nsew
rlabel locali s -6066 26731 -5993 26830 4 VSS
port 42 nsew
rlabel locali s -6046 26830 -5993 27065 4 VSS
port 42 nsew
rlabel locali s -6055 27065 -5959 27341 4 VSS
port 42 nsew
rlabel locali s -6055 27341 -5875 27346 4 VSS
port 42 nsew
rlabel locali s -6055 27346 -5674 27380 4 VSS
port 42 nsew
rlabel locali s -6055 27380 -5875 27384 4 VSS
port 42 nsew
rlabel locali s -6055 27384 -5959 27576 4 VSS
port 42 nsew
rlabel locali s -6055 27576 -5958 27650 4 VSS
port 42 nsew
rlabel locali s -6055 27650 -5873 27655 4 VSS
port 42 nsew
rlabel locali s -6055 27655 -5674 27689 4 VSS
port 42 nsew
rlabel locali s -6055 27689 -5873 27693 4 VSS
port 42 nsew
rlabel locali s -6055 27693 -5958 27697 4 VSS
port 42 nsew
rlabel locali s -8171 26413 -8132 27098 4 VSS
port 42 nsew
rlabel locali s -8287 26398 -8219 26440 4 VSS
port 42 nsew
rlabel locali s -10663 26278 -10595 26287 4 VSS
port 42 nsew
rlabel locali s -10763 26276 -10703 26287 4 VSS
port 42 nsew
rlabel locali s -10763 26287 -10595 26398 4 VSS
port 42 nsew
rlabel locali s -10663 26398 -10595 26440 4 VSS
port 42 nsew
rlabel locali s -10763 26398 -10703 26413 4 VSS
port 42 nsew
rlabel locali s -11043 26180 -10975 26342 4 VSS
port 42 nsew
rlabel locali s -11202 26342 -10975 26376 4 VSS
port 42 nsew
rlabel locali s -8446 26440 -8219 26474 4 VSS
port 42 nsew
rlabel locali s -10663 26440 -10436 26474 4 VSS
port 42 nsew
rlabel locali s -8287 26474 -8219 26885 4 VSS
port 42 nsew
rlabel locali s -10663 26474 -10595 26885 4 VSS
port 42 nsew
rlabel locali s -8446 26885 -8219 26919 4 VSS
port 42 nsew
rlabel locali s -10663 26885 -10436 26919 4 VSS
port 42 nsew
rlabel locali s -8287 26919 -8219 27081 4 VSS
port 42 nsew
rlabel locali s -10663 26919 -10595 27081 4 VSS
port 42 nsew
rlabel locali s -8446 27081 -8219 27098 4 VSS
port 42 nsew
rlabel locali s -8446 27098 -8132 27115 4 VSS
port 42 nsew
rlabel locali s -10663 27081 -10436 27098 4 VSS
port 42 nsew
rlabel locali s -10750 26413 -10711 27098 4 VSS
port 42 nsew
rlabel locali s -11043 26376 -10975 26538 4 VSS
port 42 nsew
rlabel locali s -11202 26538 -10975 26572 4 VSS
port 42 nsew
rlabel locali s -11043 26572 -10975 26581 4 VSS
port 42 nsew
rlabel locali s -12889 25903 -12836 27065 4 VSS
port 42 nsew
rlabel locali s -13321 25903 -13284 26160 4 VSS
port 42 nsew
rlabel locali s -13321 26160 -13223 26197 4 VSS
port 42 nsew
rlabel locali s -13260 26197 -13223 26279 4 VSS
port 42 nsew
rlabel locali s -13260 26279 -13202 26282 4 VSS
port 42 nsew
rlabel locali s -13260 26282 -13000 26316 4 VSS
port 42 nsew
rlabel locali s -10750 27098 -10436 27115 4 VSS
port 42 nsew
rlabel locali s -8287 27115 -8132 27209 4 VSS
port 42 nsew
rlabel locali s -6045 27697 -5958 28364 4 VSS
port 42 nsew
rlabel locali s -7907 27790 -7839 27889 4 VSS
port 42 nsew
rlabel locali s -7907 27889 -7680 27923 4 VSS
port 42 nsew
rlabel locali s -7907 27923 -7839 28085 4 VSS
port 42 nsew
rlabel locali s -7907 28085 -7680 28119 4 VSS
port 42 nsew
rlabel locali s -7907 28119 -7839 28281 4 VSS
port 42 nsew
rlabel locali s -7907 28281 -7680 28315 4 VSS
port 42 nsew
rlabel locali s -5681 28366 -5561 28368 4 VSS
port 42 nsew
rlabel locali s -6046 28364 -5870 28368 4 VSS
port 42 nsew
rlabel locali s -6046 28368 -5561 28402 4 VSS
port 42 nsew
rlabel locali s -5681 28402 -5561 28403 4 VSS
port 42 nsew
rlabel locali s -6046 28402 -5870 28403 4 VSS
port 42 nsew
rlabel locali s -5598 28403 -5561 28660 4 VSS
port 42 nsew
rlabel locali s -5659 28660 -5561 28697 4 VSS
port 42 nsew
rlabel locali s -5584 28749 -5530 28888 4 VSS
port 42 nsew
rlabel locali s -5659 28697 -5622 28779 4 VSS
port 42 nsew
rlabel locali s -5680 28779 -5622 28782 4 VSS
port 42 nsew
rlabel locali s -5882 28782 -5622 28816 4 VSS
port 42 nsew
rlabel locali s -6046 28403 -5993 29565 4 VSS
port 42 nsew
rlabel locali s -7907 28315 -7839 28846 4 VSS
port 42 nsew
rlabel locali s -7907 28846 -7680 28880 4 VSS
port 42 nsew
rlabel locali s -8171 27209 -8132 28873 4 VSS
port 42 nsew
rlabel locali s -8287 27209 -8219 27277 4 VSS
port 42 nsew
rlabel locali s -10750 27115 -10595 27209 4 VSS
port 42 nsew
rlabel locali s -10663 27209 -10595 27277 4 VSS
port 42 nsew
rlabel locali s -8446 27277 -8219 27311 4 VSS
port 42 nsew
rlabel locali s -10663 27277 -10436 27311 4 VSS
port 42 nsew
rlabel locali s -8287 27311 -8219 27410 4 VSS
port 42 nsew
rlabel locali s -10663 27311 -10595 27410 4 VSS
port 42 nsew
rlabel locali s -8287 28739 -8219 28748 4 VSS
port 42 nsew
rlabel locali s -10663 28739 -10595 28748 4 VSS
port 42 nsew
rlabel locali s -8446 28748 -8219 28782 4 VSS
port 42 nsew
rlabel locali s -10663 28748 -10436 28782 4 VSS
port 42 nsew
rlabel locali s -7907 28880 -7839 29042 4 VSS
port 42 nsew
rlabel locali s -8173 28873 -8113 28896 4 VSS
port 42 nsew
rlabel locali s -8287 28782 -8219 28896 4 VSS
port 42 nsew
rlabel locali s -8287 28896 -8113 28944 4 VSS
port 42 nsew
rlabel locali s -10663 28782 -10595 28896 4 VSS
port 42 nsew
rlabel locali s -10750 27209 -10711 28873 4 VSS
port 42 nsew
rlabel locali s -12923 27065 -12827 27341 4 VSS
port 42 nsew
rlabel locali s -13007 27341 -12827 27346 4 VSS
port 42 nsew
rlabel locali s -13208 27346 -12827 27380 4 VSS
port 42 nsew
rlabel locali s -13007 27380 -12827 27384 4 VSS
port 42 nsew
rlabel locali s -12923 27384 -12827 27576 4 VSS
port 42 nsew
rlabel locali s -12924 27576 -12827 27650 4 VSS
port 42 nsew
rlabel locali s -13009 27650 -12827 27655 4 VSS
port 42 nsew
rlabel locali s -13208 27655 -12827 27689 4 VSS
port 42 nsew
rlabel locali s -13009 27689 -12827 27693 4 VSS
port 42 nsew
rlabel locali s -12924 27693 -12827 27697 4 VSS
port 42 nsew
rlabel locali s -11043 27790 -10975 27889 4 VSS
port 42 nsew
rlabel locali s -11202 27889 -10975 27923 4 VSS
port 42 nsew
rlabel locali s -11043 27923 -10975 28085 4 VSS
port 42 nsew
rlabel locali s -11202 28085 -10975 28119 4 VSS
port 42 nsew
rlabel locali s -11043 28119 -10975 28281 4 VSS
port 42 nsew
rlabel locali s -11202 28281 -10975 28315 4 VSS
port 42 nsew
rlabel locali s -11043 28315 -10975 28846 4 VSS
port 42 nsew
rlabel locali s -12924 27697 -12837 28364 4 VSS
port 42 nsew
rlabel locali s -13012 28364 -12836 28368 4 VSS
port 42 nsew
rlabel locali s -13321 28366 -13201 28368 4 VSS
port 42 nsew
rlabel locali s -13321 28368 -12836 28402 4 VSS
port 42 nsew
rlabel locali s -13012 28402 -12836 28403 4 VSS
port 42 nsew
rlabel locali s -13321 28402 -13201 28403 4 VSS
port 42 nsew
rlabel locali s -10769 28873 -10709 28896 4 VSS
port 42 nsew
rlabel locali s -10769 28896 -10595 28944 4 VSS
port 42 nsew
rlabel locali s -8446 28944 -8113 28978 4 VSS
port 42 nsew
rlabel locali s -10769 28944 -10436 28978 4 VSS
port 42 nsew
rlabel locali s -8287 28978 -8113 29007 4 VSS
port 42 nsew
rlabel locali s -8173 29007 -8113 29010 4 VSS
port 42 nsew
rlabel locali s -7907 29042 -7680 29076 4 VSS
port 42 nsew
rlabel locali s -7907 29076 -7839 29238 4 VSS
port 42 nsew
rlabel locali s -7907 29238 -7680 29272 4 VSS
port 42 nsew
rlabel locali s -7907 29272 -7839 29281 4 VSS
port 42 nsew
rlabel locali s -5590 29827 -5536 29966 4 VSS
port 42 nsew
rlabel locali s -6055 29565 -5959 29841 4 VSS
port 42 nsew
rlabel locali s -6055 29841 -5875 29846 4 VSS
port 42 nsew
rlabel locali s -6055 29846 -5674 29880 4 VSS
port 42 nsew
rlabel locali s -6055 29880 -5875 29884 4 VSS
port 42 nsew
rlabel locali s -6055 29884 -5959 30150 4 VSS
port 42 nsew
rlabel locali s -6055 30150 -5873 30155 4 VSS
port 42 nsew
rlabel locali s -6055 30155 -5674 30189 4 VSS
port 42 nsew
rlabel locali s -6055 30189 -5873 30193 4 VSS
port 42 nsew
rlabel locali s -6055 30193 -5959 30197 4 VSS
port 42 nsew
rlabel locali s -8171 29010 -8132 29774 4 VSS
port 42 nsew
rlabel locali s -8287 29007 -8219 29079 4 VSS
port 42 nsew
rlabel locali s -8287 29079 -8217 29140 4 VSS
port 42 nsew
rlabel locali s -10769 28978 -10595 29007 4 VSS
port 42 nsew
rlabel locali s -10663 29007 -10595 29079 4 VSS
port 42 nsew
rlabel locali s -10769 29007 -10709 29010 4 VSS
port 42 nsew
rlabel locali s -11202 28846 -10975 28880 4 VSS
port 42 nsew
rlabel locali s -10665 29079 -10595 29140 4 VSS
port 42 nsew
rlabel locali s -8446 29140 -8217 29174 4 VSS
port 42 nsew
rlabel locali s -10665 29140 -10436 29174 4 VSS
port 42 nsew
rlabel locali s -8287 29174 -8217 29273 4 VSS
port 42 nsew
rlabel locali s -10665 29174 -10595 29273 4 VSS
port 42 nsew
rlabel locali s -8285 29273 -8217 29576 4 VSS
port 42 nsew
rlabel locali s -10665 29273 -10597 29576 4 VSS
port 42 nsew
rlabel locali s -8287 29576 -8217 29585 4 VSS
port 42 nsew
rlabel locali s -10665 29576 -10595 29585 4 VSS
port 42 nsew
rlabel locali s -8446 29585 -8217 29599 4 VSS
port 42 nsew
rlabel locali s -8446 29599 -8219 29619 4 VSS
port 42 nsew
rlabel locali s -10665 29585 -10436 29599 4 VSS
port 42 nsew
rlabel locali s -10663 29599 -10436 29619 4 VSS
port 42 nsew
rlabel locali s -8287 29619 -8219 29774 4 VSS
port 42 nsew
rlabel locali s -8287 29774 -8132 29781 4 VSS
port 42 nsew
rlabel locali s -10663 29619 -10595 29774 4 VSS
port 42 nsew
rlabel locali s -10750 29010 -10711 29774 4 VSS
port 42 nsew
rlabel locali s -11043 28880 -10975 29042 4 VSS
port 42 nsew
rlabel locali s -11202 29042 -10975 29076 4 VSS
port 42 nsew
rlabel locali s -11043 29076 -10975 29238 4 VSS
port 42 nsew
rlabel locali s -11202 29238 -10975 29272 4 VSS
port 42 nsew
rlabel locali s -11043 29272 -10975 29281 4 VSS
port 42 nsew
rlabel locali s -12889 28403 -12836 29565 4 VSS
port 42 nsew
rlabel locali s -13321 28403 -13284 28660 4 VSS
port 42 nsew
rlabel locali s -13321 28660 -13223 28697 4 VSS
port 42 nsew
rlabel locali s -13260 28697 -13223 28779 4 VSS
port 42 nsew
rlabel locali s -13260 28779 -13202 28782 4 VSS
port 42 nsew
rlabel locali s -13260 28782 -13000 28816 4 VSS
port 42 nsew
rlabel locali s -13352 28749 -13298 28888 4 VSS
port 42 nsew
rlabel locali s -10750 29774 -10595 29781 4 VSS
port 42 nsew
rlabel locali s -8446 29781 -8132 29815 4 VSS
port 42 nsew
rlabel locali s -10750 29781 -10436 29815 4 VSS
port 42 nsew
rlabel locali s -8287 29815 -8132 29885 4 VSS
port 42 nsew
rlabel locali s -6046 30197 -5993 30864 4 VSS
port 42 nsew
rlabel locali s -7907 30490 -7839 30589 4 VSS
port 42 nsew
rlabel locali s -7907 30589 -7680 30623 4 VSS
port 42 nsew
rlabel locali s -7907 30623 -7839 30785 4 VSS
port 42 nsew
rlabel locali s -7907 30785 -7680 30819 4 VSS
port 42 nsew
rlabel locali s -5681 30866 -5561 30868 4 VSS
port 42 nsew
rlabel locali s -6046 30864 -5870 30868 4 VSS
port 42 nsew
rlabel locali s -6046 30868 -5561 30902 4 VSS
port 42 nsew
rlabel locali s -5681 30902 -5561 30903 4 VSS
port 42 nsew
rlabel locali s -6046 30902 -5870 30903 4 VSS
port 42 nsew
rlabel locali s -5598 30903 -5561 31160 4 VSS
port 42 nsew
rlabel locali s -5659 31160 -5561 31197 4 VSS
port 42 nsew
rlabel locali s -5584 31249 -5530 31388 4 VSS
port 42 nsew
rlabel locali s -5659 31197 -5622 31279 4 VSS
port 42 nsew
rlabel locali s -5680 31279 -5622 31282 4 VSS
port 42 nsew
rlabel locali s -5882 31282 -5622 31316 4 VSS
port 42 nsew
rlabel locali s -6046 30903 -5993 32065 4 VSS
port 42 nsew
rlabel locali s -7907 30819 -7839 30981 4 VSS
port 42 nsew
rlabel locali s -7907 30981 -7680 31015 4 VSS
port 42 nsew
rlabel locali s -7907 31015 -7839 31471 4 VSS
port 42 nsew
rlabel locali s -7907 31471 -7680 31505 4 VSS
port 42 nsew
rlabel locali s -7907 31505 -7839 31667 4 VSS
port 42 nsew
rlabel locali s -8171 29885 -8132 31258 4 VSS
port 42 nsew
rlabel locali s -8287 29885 -8219 29977 4 VSS
port 42 nsew
rlabel locali s -10750 29815 -10595 29885 4 VSS
port 42 nsew
rlabel locali s -10663 29885 -10595 29977 4 VSS
port 42 nsew
rlabel locali s -8446 29977 -8219 30011 4 VSS
port 42 nsew
rlabel locali s -10663 29977 -10436 30011 4 VSS
port 42 nsew
rlabel locali s -8287 30011 -8219 30110 4 VSS
port 42 nsew
rlabel locali s -10663 30011 -10595 30110 4 VSS
port 42 nsew
rlabel locali s -10750 29885 -10711 31258 4 VSS
port 42 nsew
rlabel locali s -12923 29565 -12827 29841 4 VSS
port 42 nsew
rlabel locali s -13007 29841 -12827 29846 4 VSS
port 42 nsew
rlabel locali s -13208 29846 -12827 29880 4 VSS
port 42 nsew
rlabel locali s -13007 29880 -12827 29884 4 VSS
port 42 nsew
rlabel locali s -12923 29884 -12827 30150 4 VSS
port 42 nsew
rlabel locali s -13346 29827 -13292 29966 4 VSS
port 42 nsew
rlabel locali s -13009 30150 -12827 30155 4 VSS
port 42 nsew
rlabel locali s -13208 30155 -12827 30189 4 VSS
port 42 nsew
rlabel locali s -13009 30189 -12827 30193 4 VSS
port 42 nsew
rlabel locali s -12923 30193 -12827 30197 4 VSS
port 42 nsew
rlabel locali s -10750 31258 -8132 31511 4 VSS
port 42 nsew
rlabel locali s -11043 30490 -10975 30589 4 VSS
port 42 nsew
rlabel locali s -11202 30589 -10975 30623 4 VSS
port 42 nsew
rlabel locali s -11043 30623 -10975 30785 4 VSS
port 42 nsew
rlabel locali s -11202 30785 -10975 30819 4 VSS
port 42 nsew
rlabel locali s -11043 30819 -10975 30981 4 VSS
port 42 nsew
rlabel locali s -12889 30197 -12836 30864 4 VSS
port 42 nsew
rlabel locali s -13012 30864 -12836 30868 4 VSS
port 42 nsew
rlabel locali s -13321 30866 -13201 30868 4 VSS
port 42 nsew
rlabel locali s -13321 30868 -12836 30902 4 VSS
port 42 nsew
rlabel locali s -13012 30902 -12836 30903 4 VSS
port 42 nsew
rlabel locali s -13321 30902 -13201 30903 4 VSS
port 42 nsew
rlabel locali s -11202 30981 -10975 31015 4 VSS
port 42 nsew
rlabel locali s -11043 31015 -10975 31471 4 VSS
port 42 nsew
rlabel locali s -11202 31471 -10975 31505 4 VSS
port 42 nsew
rlabel locali s -10769 31511 -8132 31556 4 VSS
port 42 nsew
rlabel locali s -8171 31556 -8132 31641 4 VSS
port 42 nsew
rlabel locali s -7907 31667 -7680 31701 4 VSS
port 42 nsew
rlabel locali s -7907 31701 -7839 31863 4 VSS
port 42 nsew
rlabel locali s -8173 31641 -8113 31773 4 VSS
port 42 nsew
rlabel locali s -8171 31773 -8132 31774 4 VSS
port 42 nsew
rlabel locali s -7907 31863 -7680 31897 4 VSS
port 42 nsew
rlabel locali s -7907 31897 -7839 31906 4 VSS
port 42 nsew
rlabel locali s -5590 32327 -5536 32466 4 VSS
port 42 nsew
rlabel locali s -6055 32065 -5959 32341 4 VSS
port 42 nsew
rlabel locali s -6055 32341 -5875 32346 4 VSS
port 42 nsew
rlabel locali s -6055 32346 -5674 32380 4 VSS
port 42 nsew
rlabel locali s -6055 32380 -5875 32384 4 VSS
port 42 nsew
rlabel locali s -6055 32384 -5959 32650 4 VSS
port 42 nsew
rlabel locali s -8486 32291 -8421 32304 4 VSS
port 42 nsew
rlabel locali s -9012 31556 -8751 32304 4 VSS
port 42 nsew
rlabel locali s -9012 32304 -8421 32401 4 VSS
port 42 nsew
rlabel locali s -9012 32401 -8025 32434 4 VSS
port 42 nsew
rlabel locali s -8486 32434 -8025 32435 4 VSS
port 42 nsew
rlabel locali s -6055 32650 -5873 32655 4 VSS
port 42 nsew
rlabel locali s -6055 32655 -5674 32689 4 VSS
port 42 nsew
rlabel locali s -6055 32689 -5873 32693 4 VSS
port 42 nsew
rlabel locali s -6055 32693 -5959 32697 4 VSS
port 42 nsew
rlabel locali s -8486 32435 -8421 32610 4 VSS
port 42 nsew
rlabel locali s -9012 32434 -8751 32610 4 VSS
port 42 nsew
rlabel locali s -6046 32697 -5993 33364 4 VSS
port 42 nsew
rlabel locali s -5681 33366 -5561 33368 4 VSS
port 42 nsew
rlabel locali s -6046 33364 -5870 33368 4 VSS
port 42 nsew
rlabel locali s -6046 33368 -5561 33402 4 VSS
port 42 nsew
rlabel locali s -5681 33402 -5561 33403 4 VSS
port 42 nsew
rlabel locali s -6046 33402 -5870 33403 4 VSS
port 42 nsew
rlabel locali s -5598 33403 -5561 33660 4 VSS
port 42 nsew
rlabel locali s -5659 33660 -5561 33697 4 VSS
port 42 nsew
rlabel locali s -5584 33749 -5530 33888 4 VSS
port 42 nsew
rlabel locali s -5659 33697 -5622 33779 4 VSS
port 42 nsew
rlabel locali s -5680 33779 -5622 33782 4 VSS
port 42 nsew
rlabel locali s -5882 33782 -5622 33816 4 VSS
port 42 nsew
rlabel locali s -6046 33403 -5993 34565 4 VSS
port 42 nsew
rlabel locali s -9012 32610 -8421 32740 4 VSS
port 42 nsew
rlabel locali s -8486 32740 -8421 32927 4 VSS
port 42 nsew
rlabel locali s -9012 32740 -8751 32867 4 VSS
port 42 nsew
rlabel locali s -10131 31556 -9870 32304 4 VSS
port 42 nsew
rlabel locali s -10769 31556 -10709 31643 4 VSS
port 42 nsew
rlabel locali s -10750 31643 -10711 31644 4 VSS
port 42 nsew
rlabel locali s -11043 31505 -10975 31667 4 VSS
port 42 nsew
rlabel locali s -11202 31667 -10975 31701 4 VSS
port 42 nsew
rlabel locali s -11043 31701 -10975 31863 4 VSS
port 42 nsew
rlabel locali s -11202 31863 -10975 31897 4 VSS
port 42 nsew
rlabel locali s -11043 31897 -10975 31906 4 VSS
port 42 nsew
rlabel locali s -12889 30903 -12836 32065 4 VSS
port 42 nsew
rlabel locali s -13321 30903 -13284 31160 4 VSS
port 42 nsew
rlabel locali s -13321 31160 -13223 31197 4 VSS
port 42 nsew
rlabel locali s -13260 31197 -13223 31279 4 VSS
port 42 nsew
rlabel locali s -13260 31279 -13202 31282 4 VSS
port 42 nsew
rlabel locali s -13260 31282 -13000 31316 4 VSS
port 42 nsew
rlabel locali s -13352 31249 -13298 31388 4 VSS
port 42 nsew
rlabel locali s -10461 32291 -10396 32304 4 VSS
port 42 nsew
rlabel locali s -10461 32304 -9870 32401 4 VSS
port 42 nsew
rlabel locali s -12923 32065 -12827 32341 4 VSS
port 42 nsew
rlabel locali s -13007 32341 -12827 32346 4 VSS
port 42 nsew
rlabel locali s -13208 32346 -12827 32380 4 VSS
port 42 nsew
rlabel locali s -13007 32380 -12827 32384 4 VSS
port 42 nsew
rlabel locali s -10857 32401 -9870 32434 4 VSS
port 42 nsew
rlabel locali s -10131 32434 -9870 32610 4 VSS
port 42 nsew
rlabel locali s -10857 32434 -10396 32435 4 VSS
port 42 nsew
rlabel locali s -10461 32435 -10396 32610 4 VSS
port 42 nsew
rlabel locali s -10461 32610 -9870 32740 4 VSS
port 42 nsew
rlabel locali s -12923 32384 -12827 32650 4 VSS
port 42 nsew
rlabel locali s -13346 32327 -13292 32466 4 VSS
port 42 nsew
rlabel locali s -13009 32650 -12827 32655 4 VSS
port 42 nsew
rlabel locali s -13208 32655 -12827 32689 4 VSS
port 42 nsew
rlabel locali s -13009 32689 -12827 32693 4 VSS
port 42 nsew
rlabel locali s -12923 32693 -12827 32697 4 VSS
port 42 nsew
rlabel locali s -10131 32740 -9870 32867 4 VSS
port 42 nsew
rlabel locali s -10131 32867 -8751 32927 4 VSS
port 42 nsew
rlabel locali s -10461 32740 -10396 32927 4 VSS
port 42 nsew
rlabel locali s -10461 32927 -8421 33057 4 VSS
port 42 nsew
rlabel locali s -8486 33057 -8421 33373 4 VSS
port 42 nsew
rlabel locali s -10131 33057 -8751 33128 4 VSS
port 42 nsew
rlabel locali s -9012 33128 -8751 33373 4 VSS
port 42 nsew
rlabel locali s -9012 33373 -8421 33433 4 VSS
port 42 nsew
rlabel locali s -9012 33433 -7924 33467 4 VSS
port 42 nsew
rlabel locali s -9012 33467 -8421 33503 4 VSS
port 42 nsew
rlabel locali s -8486 33503 -8421 33565 4 VSS
port 42 nsew
rlabel locali s -9012 33503 -8751 33704 4 VSS
port 42 nsew
rlabel locali s -10131 33128 -9870 33373 4 VSS
port 42 nsew
rlabel locali s -10461 33057 -10396 33373 4 VSS
port 42 nsew
rlabel locali s -10461 33373 -9870 33433 4 VSS
port 42 nsew
rlabel locali s -12889 32697 -12836 33364 4 VSS
port 42 nsew
rlabel locali s -13012 33364 -12836 33368 4 VSS
port 42 nsew
rlabel locali s -13321 33366 -13201 33368 4 VSS
port 42 nsew
rlabel locali s -13321 33368 -12836 33402 4 VSS
port 42 nsew
rlabel locali s -13012 33402 -12836 33403 4 VSS
port 42 nsew
rlabel locali s -13321 33402 -13201 33403 4 VSS
port 42 nsew
rlabel locali s -10958 33433 -9870 33467 4 VSS
port 42 nsew
rlabel locali s -10461 33467 -9870 33503 4 VSS
port 42 nsew
rlabel locali s -10131 33503 -9870 33704 4 VSS
port 42 nsew
rlabel locali s -10461 33503 -10396 33565 4 VSS
port 42 nsew
rlabel locali s -10131 33704 -8751 33965 4 VSS
port 42 nsew
rlabel locali s -7803 33987 -7717 34232 4 VSS
port 42 nsew
rlabel locali s -7803 34232 -7561 34266 4 VSS
port 42 nsew
rlabel locali s -7803 34266 -7717 34297 4 VSS
port 42 nsew
rlabel locali s -9012 33965 -8751 34297 4 VSS
port 42 nsew
rlabel locali s -9012 34297 -7717 34358 4 VSS
port 42 nsew
rlabel locali s -7803 34358 -7717 34428 4 VSS
port 42 nsew
rlabel locali s -7803 34428 -7561 34462 4 VSS
port 42 nsew
rlabel locali s -5590 34827 -5536 34966 4 VSS
port 42 nsew
rlabel locali s -6055 34565 -5959 34841 4 VSS
port 42 nsew
rlabel locali s -7803 34462 -7717 34602 4 VSS
port 42 nsew
rlabel locali s -9012 34358 -8210 34448 4 VSS
port 42 nsew
rlabel locali s -8271 34448 -8210 34674 4 VSS
port 42 nsew
rlabel locali s -9012 34448 -8751 34674 4 VSS
port 42 nsew
rlabel locali s -9012 34674 -8210 34744 4 VSS
port 42 nsew
rlabel locali s -10131 33965 -9870 34297 4 VSS
port 42 nsew
rlabel locali s -11165 33987 -11079 34232 4 VSS
port 42 nsew
rlabel locali s -11321 34232 -11079 34266 4 VSS
port 42 nsew
rlabel locali s -11165 34266 -11079 34297 4 VSS
port 42 nsew
rlabel locali s -11165 34297 -9870 34358 4 VSS
port 42 nsew
rlabel locali s -10672 34358 -9870 34448 4 VSS
port 42 nsew
rlabel locali s -10131 34448 -9870 34674 4 VSS
port 42 nsew
rlabel locali s -10672 34448 -10611 34674 4 VSS
port 42 nsew
rlabel locali s -11165 34358 -11079 34428 4 VSS
port 42 nsew
rlabel locali s -11321 34428 -11079 34462 4 VSS
port 42 nsew
rlabel locali s -11165 34462 -11079 34602 4 VSS
port 42 nsew
rlabel locali s -12889 33403 -12836 34565 4 VSS
port 42 nsew
rlabel locali s -13321 33403 -13284 33660 4 VSS
port 42 nsew
rlabel locali s -13321 33660 -13223 33697 4 VSS
port 42 nsew
rlabel locali s -13260 33697 -13223 33779 4 VSS
port 42 nsew
rlabel locali s -13260 33779 -13202 33782 4 VSS
port 42 nsew
rlabel locali s -13260 33782 -13000 33816 4 VSS
port 42 nsew
rlabel locali s -13352 33749 -13298 33888 4 VSS
port 42 nsew
rlabel locali s -10672 34674 -9870 34744 4 VSS
port 42 nsew
rlabel locali s -10672 34744 -8210 34747 4 VSS
port 42 nsew
rlabel locali s -6055 34841 -5875 34846 4 VSS
port 42 nsew
rlabel locali s -6055 34846 -5674 34880 4 VSS
port 42 nsew
rlabel locali s -6055 34880 -5875 34884 4 VSS
port 42 nsew
rlabel locali s -6055 34884 -5959 35150 4 VSS
port 42 nsew
rlabel locali s -10654 34747 -8228 34798 4 VSS
port 42 nsew
rlabel locali s -8289 34798 -8228 35004 4 VSS
port 42 nsew
rlabel locali s -10131 34798 -8751 35004 4 VSS
port 42 nsew
rlabel locali s -10654 34798 -10593 35004 4 VSS
port 42 nsew
rlabel locali s -10654 35004 -8228 35005 4 VSS
port 42 nsew
rlabel locali s -9012 35005 -8228 35037 4 VSS
port 42 nsew
rlabel locali s -9012 35037 -7868 35071 4 VSS
port 42 nsew
rlabel locali s -9012 35071 -8176 35072 4 VSS
port 42 nsew
rlabel locali s -6055 35150 -5873 35155 4 VSS
port 42 nsew
rlabel locali s -6055 35155 -5674 35189 4 VSS
port 42 nsew
rlabel locali s -9012 35072 -8228 35128 4 VSS
port 42 nsew
rlabel locali s -8289 35128 -8228 35189 4 VSS
port 42 nsew
rlabel locali s -6055 35189 -5873 35193 4 VSS
port 42 nsew
rlabel locali s -6055 35193 -5959 35197 4 VSS
port 42 nsew
rlabel locali s -6046 35197 -5993 35864 4 VSS
port 42 nsew
rlabel locali s -7805 35592 -7719 35837 4 VSS
port 42 nsew
rlabel locali s -5681 35866 -5561 35868 4 VSS
port 42 nsew
rlabel locali s -6046 35864 -5870 35868 4 VSS
port 42 nsew
rlabel locali s -6046 35868 -5561 35902 4 VSS
port 42 nsew
rlabel locali s -7805 35837 -7563 35871 4 VSS
port 42 nsew
rlabel locali s -5681 35902 -5561 35903 4 VSS
port 42 nsew
rlabel locali s -6046 35902 -5870 35903 4 VSS
port 42 nsew
rlabel locali s -5598 35903 -5561 36160 4 VSS
port 42 nsew
rlabel locali s -5659 36160 -5561 36197 4 VSS
port 42 nsew
rlabel locali s -5659 36197 -5622 36279 4 VSS
port 42 nsew
rlabel locali s -5680 36279 -5622 36282 4 VSS
port 42 nsew
rlabel locali s -5882 36282 -5622 36316 4 VSS
port 42 nsew
rlabel locali s -6046 35903 -5993 37065 4 VSS
port 42 nsew
rlabel locali s -7805 35871 -7719 35902 4 VSS
port 42 nsew
rlabel locali s -9012 35128 -8751 35902 4 VSS
port 42 nsew
rlabel locali s -9012 35902 -7719 35963 4 VSS
port 42 nsew
rlabel locali s -7805 35963 -7719 36033 4 VSS
port 42 nsew
rlabel locali s -7805 36033 -7563 36067 4 VSS
port 42 nsew
rlabel locali s -7805 36067 -7719 36207 4 VSS
port 42 nsew
rlabel locali s -9012 35963 -8212 36053 4 VSS
port 42 nsew
rlabel locali s -8273 36053 -8212 36344 4 VSS
port 42 nsew
rlabel locali s -9012 36053 -8751 36202 4 VSS
port 42 nsew
rlabel locali s -10654 35005 -9870 35037 4 VSS
port 42 nsew
rlabel locali s -12923 34565 -12827 34841 4 VSS
port 42 nsew
rlabel locali s -13007 34841 -12827 34846 4 VSS
port 42 nsew
rlabel locali s -13208 34846 -12827 34880 4 VSS
port 42 nsew
rlabel locali s -13007 34880 -12827 34884 4 VSS
port 42 nsew
rlabel locali s -11014 35037 -9870 35071 4 VSS
port 42 nsew
rlabel locali s -10706 35071 -9870 35072 4 VSS
port 42 nsew
rlabel locali s -10654 35072 -9870 35128 4 VSS
port 42 nsew
rlabel locali s -10131 35128 -9870 35902 4 VSS
port 42 nsew
rlabel locali s -10654 35128 -10593 35189 4 VSS
port 42 nsew
rlabel locali s -12923 34884 -12827 35150 4 VSS
port 42 nsew
rlabel locali s -13346 34827 -13292 34966 4 VSS
port 42 nsew
rlabel locali s -13009 35150 -12827 35155 4 VSS
port 42 nsew
rlabel locali s -13208 35155 -12827 35189 4 VSS
port 42 nsew
rlabel locali s -13009 35189 -12827 35193 4 VSS
port 42 nsew
rlabel locali s -12923 35193 -12827 35197 4 VSS
port 42 nsew
rlabel locali s -11163 35592 -11077 35837 4 VSS
port 42 nsew
rlabel locali s -11319 35837 -11077 35871 4 VSS
port 42 nsew
rlabel locali s -12889 35197 -12836 35864 4 VSS
port 42 nsew
rlabel locali s -13012 35864 -12836 35868 4 VSS
port 42 nsew
rlabel locali s -13321 35866 -13201 35868 4 VSS
port 42 nsew
rlabel locali s -11163 35871 -11077 35902 4 VSS
port 42 nsew
rlabel locali s -11163 35902 -9870 35963 4 VSS
port 42 nsew
rlabel locali s -10670 35963 -9870 36053 4 VSS
port 42 nsew
rlabel locali s -10131 36053 -9870 36202 4 VSS
port 42 nsew
rlabel locali s -10131 36202 -8751 36344 4 VSS
port 42 nsew
rlabel locali s -10670 36053 -10609 36344 4 VSS
port 42 nsew
rlabel locali s -11163 35963 -11077 36033 4 VSS
port 42 nsew
rlabel locali s -13321 35868 -12836 35902 4 VSS
port 42 nsew
rlabel locali s -13012 35902 -12836 35903 4 VSS
port 42 nsew
rlabel locali s -13321 35902 -13201 35903 4 VSS
port 42 nsew
rlabel locali s -11319 36033 -11077 36067 4 VSS
port 42 nsew
rlabel locali s -11163 36067 -11077 36207 4 VSS
port 42 nsew
rlabel locali s -10670 36344 -8212 36352 4 VSS
port 42 nsew
rlabel locali s -10652 36352 -8230 36463 4 VSS
port 42 nsew
rlabel locali s -9012 36463 -8230 36495 4 VSS
port 42 nsew
rlabel locali s -8291 36495 -8230 36637 4 VSS
port 42 nsew
rlabel locali s -9012 36495 -8751 36637 4 VSS
port 42 nsew
rlabel locali s -9012 36637 -8230 36642 4 VSS
port 42 nsew
rlabel locali s -9012 36642 -7870 36676 4 VSS
port 42 nsew
rlabel locali s -9012 36676 -8178 36677 4 VSS
port 42 nsew
rlabel locali s -9012 36677 -8230 36788 4 VSS
port 42 nsew
rlabel locali s -8291 36788 -8230 36794 4 VSS
port 42 nsew
rlabel locali s -6055 37065 -5959 37341 4 VSS
port 42 nsew
rlabel locali s -6055 37341 -5875 37346 4 VSS
port 42 nsew
rlabel locali s -6055 37346 -5674 37380 4 VSS
port 42 nsew
rlabel locali s -8477 37253 -8412 37277 4 VSS
port 42 nsew
rlabel locali s -9012 36788 -8751 37277 4 VSS
port 42 nsew
rlabel locali s -9012 37277 -8412 37363 4 VSS
port 42 nsew
rlabel locali s -6055 37380 -5875 37384 4 VSS
port 42 nsew
rlabel locali s -6055 37384 -5959 37650 4 VSS
port 42 nsew
rlabel locali s -9012 37363 -8016 37397 4 VSS
port 42 nsew
rlabel locali s -6055 37650 -5873 37655 4 VSS
port 42 nsew
rlabel locali s -6055 37655 -5674 37689 4 VSS
port 42 nsew
rlabel locali s -6055 37689 -5873 37693 4 VSS
port 42 nsew
rlabel locali s -6055 37693 -5959 37697 4 VSS
port 42 nsew
rlabel locali s -9012 37397 -8412 37416 4 VSS
port 42 nsew
rlabel locali s -10652 36463 -9870 36495 4 VSS
port 42 nsew
rlabel locali s -10131 36495 -9870 36637 4 VSS
port 42 nsew
rlabel locali s -10652 36495 -10591 36637 4 VSS
port 42 nsew
rlabel locali s -10652 36637 -9870 36642 4 VSS
port 42 nsew
rlabel locali s -11012 36642 -9870 36676 4 VSS
port 42 nsew
rlabel locali s -10704 36676 -9870 36677 4 VSS
port 42 nsew
rlabel locali s -10652 36677 -9870 36788 4 VSS
port 42 nsew
rlabel locali s -10131 36788 -9870 37277 4 VSS
port 42 nsew
rlabel locali s -10652 36788 -10591 36794 4 VSS
port 42 nsew
rlabel locali s -12889 35903 -12836 37065 4 VSS
port 42 nsew
rlabel locali s -13321 35903 -13284 36160 4 VSS
port 42 nsew
rlabel locali s -13321 36160 -13223 36197 4 VSS
port 42 nsew
rlabel locali s -13260 36197 -13223 36279 4 VSS
port 42 nsew
rlabel locali s -13260 36279 -13202 36282 4 VSS
port 42 nsew
rlabel locali s -13260 36282 -13000 36316 4 VSS
port 42 nsew
rlabel locali s -10470 37253 -10405 37277 4 VSS
port 42 nsew
rlabel locali s -10470 37277 -9870 37363 4 VSS
port 42 nsew
rlabel locali s -12923 37065 -12827 37341 4 VSS
port 42 nsew
rlabel locali s -13007 37341 -12827 37346 4 VSS
port 42 nsew
rlabel locali s -10866 37363 -9870 37397 4 VSS
port 42 nsew
rlabel locali s -13208 37346 -12827 37380 4 VSS
port 42 nsew
rlabel locali s -13007 37380 -12827 37384 4 VSS
port 42 nsew
rlabel locali s -10470 37397 -9870 37416 4 VSS
port 42 nsew
rlabel locali s -10470 37416 -8412 37423 4 VSS
port 42 nsew
rlabel locali s -6046 37697 -5993 38864 4 VSS
port 42 nsew
rlabel locali s -8477 37423 -8412 37722 4 VSS
port 42 nsew
rlabel locali s -10131 37423 -8751 37677 4 VSS
port 42 nsew
rlabel locali s -9012 37677 -8751 37722 4 VSS
port 42 nsew
rlabel locali s -9012 37722 -8412 37868 4 VSS
port 42 nsew
rlabel locali s -8477 37868 -8412 37988 4 VSS
port 42 nsew
rlabel locali s -9012 37868 -8751 37988 4 VSS
port 42 nsew
rlabel locali s -9012 37988 -8412 38134 4 VSS
port 42 nsew
rlabel locali s -8477 38134 -8412 38348 4 VSS
port 42 nsew
rlabel locali s -9012 38134 -8751 38348 4 VSS
port 42 nsew
rlabel locali s -9012 38348 -8412 38395 4 VSS
port 42 nsew
rlabel locali s -9012 38395 -7915 38429 4 VSS
port 42 nsew
rlabel locali s -9012 38429 -8412 38494 4 VSS
port 42 nsew
rlabel locali s -8477 38494 -8412 38527 4 VSS
port 42 nsew
rlabel locali s -5681 38866 -5561 38868 4 VSS
port 42 nsew
rlabel locali s -6046 38864 -5870 38868 4 VSS
port 42 nsew
rlabel locali s -6046 38868 -5561 38902 4 VSS
port 42 nsew
rlabel locali s -5681 38902 -5561 38903 4 VSS
port 42 nsew
rlabel locali s -6046 38902 -5870 38903 4 VSS
port 42 nsew
rlabel locali s -5598 38903 -5561 39160 4 VSS
port 42 nsew
rlabel locali s -5659 39160 -5561 39197 4 VSS
port 42 nsew
rlabel locali s -5659 39197 -5622 39279 4 VSS
port 42 nsew
rlabel locali s -5680 39279 -5622 39282 4 VSS
port 42 nsew
rlabel locali s -5882 39282 -5622 39316 4 VSS
port 42 nsew
rlabel locali s -6046 38903 -5993 40049 4 VSS
port 42 nsew
rlabel locali s -7932 38876 -7812 38878 4 VSS
port 42 nsew
rlabel locali s -8297 38874 -8121 38878 4 VSS
port 42 nsew
rlabel locali s -8297 38878 -7812 38912 4 VSS
port 42 nsew
rlabel locali s -9012 38494 -8751 38912 4 VSS
port 42 nsew
rlabel locali s -7932 38912 -7812 38913 4 VSS
port 42 nsew
rlabel locali s -9012 38912 -8121 38913 4 VSS
port 42 nsew
rlabel locali s -7849 38913 -7812 39170 4 VSS
port 42 nsew
rlabel locali s -9012 38913 -8244 39109 4 VSS
port 42 nsew
rlabel locali s -7910 39170 -7812 39207 4 VSS
port 42 nsew
rlabel locali s -7910 39207 -7873 39289 4 VSS
port 42 nsew
rlabel locali s -7931 39289 -7873 39292 4 VSS
port 42 nsew
rlabel locali s -8133 39292 -7873 39326 4 VSS
port 42 nsew
rlabel locali s -8297 39109 -8244 39445 4 VSS
port 42 nsew
rlabel locali s -9012 39109 -8751 39362 4 VSS
port 42 nsew
rlabel locali s -10131 37677 -9870 37722 4 VSS
port 42 nsew
rlabel locali s -10470 37423 -10405 37722 4 VSS
port 42 nsew
rlabel locali s -12923 37384 -12827 37650 4 VSS
port 42 nsew
rlabel locali s -13009 37650 -12827 37655 4 VSS
port 42 nsew
rlabel locali s -13208 37655 -12827 37689 4 VSS
port 42 nsew
rlabel locali s -13009 37689 -12827 37693 4 VSS
port 42 nsew
rlabel locali s -12923 37693 -12827 37697 4 VSS
port 42 nsew
rlabel locali s -10470 37722 -9870 37868 4 VSS
port 42 nsew
rlabel locali s -10131 37868 -9870 37988 4 VSS
port 42 nsew
rlabel locali s -10470 37868 -10405 37988 4 VSS
port 42 nsew
rlabel locali s -10470 37988 -9870 38134 4 VSS
port 42 nsew
rlabel locali s -10131 38134 -9870 38348 4 VSS
port 42 nsew
rlabel locali s -10470 38134 -10405 38348 4 VSS
port 42 nsew
rlabel locali s -10470 38348 -9870 38395 4 VSS
port 42 nsew
rlabel locali s -10967 38395 -9870 38429 4 VSS
port 42 nsew
rlabel locali s -10470 38429 -9870 38494 4 VSS
port 42 nsew
rlabel locali s -10131 38494 -9870 38912 4 VSS
port 42 nsew
rlabel locali s -10470 38494 -10405 38527 4 VSS
port 42 nsew
rlabel locali s -12889 37697 -12836 38864 4 VSS
port 42 nsew
rlabel locali s -13012 38864 -12836 38868 4 VSS
port 42 nsew
rlabel locali s -13321 38866 -13201 38868 4 VSS
port 42 nsew
rlabel locali s -10761 38874 -10585 38878 4 VSS
port 42 nsew
rlabel locali s -11070 38876 -10950 38878 4 VSS
port 42 nsew
rlabel locali s -11070 38878 -10585 38912 4 VSS
port 42 nsew
rlabel locali s -10761 38912 -9870 38913 4 VSS
port 42 nsew
rlabel locali s -11070 38912 -10950 38913 4 VSS
port 42 nsew
rlabel locali s -10638 38913 -9870 39109 4 VSS
port 42 nsew
rlabel locali s -10131 39109 -9870 39362 4 VSS
port 42 nsew
rlabel locali s -10131 39362 -8751 39445 4 VSS
port 42 nsew
rlabel locali s -10638 39109 -10585 39445 4 VSS
port 42 nsew
rlabel locali s -11070 38913 -11033 39170 4 VSS
port 42 nsew
rlabel locali s -11070 39170 -10972 39207 4 VSS
port 42 nsew
rlabel locali s -13321 38868 -12836 38902 4 VSS
port 42 nsew
rlabel locali s -13012 38902 -12836 38903 4 VSS
port 42 nsew
rlabel locali s -13321 38902 -13201 38903 4 VSS
port 42 nsew
rlabel locali s -11009 39207 -10972 39289 4 VSS
port 42 nsew
rlabel locali s -11009 39289 -10951 39292 4 VSS
port 42 nsew
rlabel locali s -11009 39292 -10749 39326 4 VSS
port 42 nsew
rlabel locali s -10638 39445 -8244 39623 4 VSS
port 42 nsew
rlabel locali s -9012 39623 -8244 39642 4 VSS
port 42 nsew
rlabel locali s -8297 39642 -8244 39958 4 VSS
port 42 nsew
rlabel locali s -9012 39642 -8751 39958 4 VSS
port 42 nsew
rlabel locali s -6068 40049 -5941 40341 4 VSS
port 42 nsew
rlabel locali s -9012 39958 -8244 40075 4 VSS
port 42 nsew
rlabel locali s -6068 40341 -5875 40346 4 VSS
port 42 nsew
rlabel locali s -6068 40346 -5674 40380 4 VSS
port 42 nsew
rlabel locali s -9012 40075 -8210 40155 4 VSS
port 42 nsew
rlabel locali s -8306 40155 -8210 40351 4 VSS
port 42 nsew
rlabel locali s -8306 40351 -8126 40356 4 VSS
port 42 nsew
rlabel locali s -6068 40380 -5875 40384 4 VSS
port 42 nsew
rlabel locali s -6068 40384 -5941 40650 4 VSS
port 42 nsew
rlabel locali s -8306 40356 -7925 40390 4 VSS
port 42 nsew
rlabel locali s -8306 40390 -8126 40394 4 VSS
port 42 nsew
rlabel locali s -6068 40650 -5873 40655 4 VSS
port 42 nsew
rlabel locali s -6068 40655 -5674 40689 4 VSS
port 42 nsew
rlabel locali s -8306 40394 -8210 40461 4 VSS
port 42 nsew
rlabel locali s -9012 40155 -8751 40461 4 VSS
port 42 nsew
rlabel locali s -9012 40461 -8210 40658 4 VSS
port 42 nsew
rlabel locali s -8306 40658 -8210 40660 4 VSS
port 42 nsew
rlabel locali s -8306 40660 -8124 40665 4 VSS
port 42 nsew
rlabel locali s -6068 40689 -5873 40693 4 VSS
port 42 nsew
rlabel locali s -6068 40693 -5941 40856 4 VSS
port 42 nsew
rlabel locali s -8306 40665 -7925 40699 4 VSS
port 42 nsew
rlabel locali s -8306 40699 -8124 40703 4 VSS
port 42 nsew
rlabel locali s -8306 40703 -8210 40707 4 VSS
port 42 nsew
rlabel locali s -9012 40658 -8751 40856 4 VSS
port 42 nsew
rlabel locali s -10638 39623 -9870 39642 4 VSS
port 42 nsew
rlabel locali s -10131 39642 -9870 39958 4 VSS
port 42 nsew
rlabel locali s -10638 39642 -10585 39958 4 VSS
port 42 nsew
rlabel locali s -10638 39958 -9870 40075 4 VSS
port 42 nsew
rlabel locali s -12889 38903 -12836 40049 4 VSS
port 42 nsew
rlabel locali s -13321 38903 -13284 39160 4 VSS
port 42 nsew
rlabel locali s -13321 39160 -13223 39197 4 VSS
port 42 nsew
rlabel locali s -13260 39197 -13223 39279 4 VSS
port 42 nsew
rlabel locali s -13260 39279 -13202 39282 4 VSS
port 42 nsew
rlabel locali s -13260 39282 -13000 39316 4 VSS
port 42 nsew
rlabel locali s -10672 40075 -9870 40155 4 VSS
port 42 nsew
rlabel locali s -10131 40155 -9870 40461 4 VSS
port 42 nsew
rlabel locali s -10672 40155 -10576 40351 4 VSS
port 42 nsew
rlabel locali s -12941 40049 -12814 40341 4 VSS
port 42 nsew
rlabel locali s -13007 40341 -12814 40346 4 VSS
port 42 nsew
rlabel locali s -10756 40351 -10576 40356 4 VSS
port 42 nsew
rlabel locali s -10957 40356 -10576 40390 4 VSS
port 42 nsew
rlabel locali s -13208 40346 -12814 40380 4 VSS
port 42 nsew
rlabel locali s -13007 40380 -12814 40384 4 VSS
port 42 nsew
rlabel locali s -10756 40390 -10576 40394 4 VSS
port 42 nsew
rlabel locali s -10672 40394 -10576 40461 4 VSS
port 42 nsew
rlabel locali s -10672 40461 -9870 40658 4 VSS
port 42 nsew
rlabel locali s -10131 40658 -9870 40856 4 VSS
port 42 nsew
rlabel locali s -10672 40658 -10576 40660 4 VSS
port 42 nsew
rlabel locali s -12941 40384 -12814 40650 4 VSS
port 42 nsew
rlabel locali s -13009 40650 -12814 40655 4 VSS
port 42 nsew
rlabel locali s -10758 40660 -10576 40665 4 VSS
port 42 nsew
rlabel locali s -10957 40665 -10576 40699 4 VSS
port 42 nsew
rlabel locali s -13208 40655 -12814 40689 4 VSS
port 42 nsew
rlabel locali s -13009 40689 -12814 40693 4 VSS
port 42 nsew
rlabel locali s -10758 40699 -10576 40703 4 VSS
port 42 nsew
rlabel locali s -10672 40703 -10576 40707 4 VSS
port 42 nsew
rlabel locali s -12941 40693 -12814 40856 4 VSS
port 42 nsew
rlabel locali s -12941 40856 -3747 41117 4 VSS
port 42 nsew
rlabel locali s -4080 41117 -3747 42470 4 VSS
port 42 nsew
rlabel locali s -10819 41117 -10558 41750 4 VSS
port 42 nsew
rlabel locali s -14110 41583 -12539 41637 4 VSS
port 42 nsew
rlabel locali s -15491 10372 -15355 41602 4 VSS
port 42 nsew
rlabel locali s -12579 41637 -12539 41740 4 VSS
port 42 nsew
rlabel locali s -11874 41750 -10558 42011 4 VSS
port 42 nsew
rlabel locali s -12452 41742 -12408 41797 4 VSS
port 42 nsew
rlabel locali s -14110 41698 -12883 41752 4 VSS
port 42 nsew
rlabel locali s -15491 41602 -15353 41738 4 VSS
port 42 nsew
rlabel locali s -12937 41752 -12883 41797 4 VSS
port 42 nsew
rlabel locali s -12937 41797 -12408 41851 4 VSS
port 42 nsew
rlabel locali s -12452 41851 -12408 41865 4 VSS
port 42 nsew
rlabel locali s -14110 41842 -13985 41896 4 VSS
port 42 nsew
rlabel locali s -11874 42011 -11613 42459 4 VSS
port 42 nsew
rlabel locali s -12317 41898 -12269 41940 4 VSS
port 42 nsew
rlabel locali s -14069 41896 -14015 41940 4 VSS
port 42 nsew
rlabel locali s -14069 41940 -12269 41994 4 VSS
port 42 nsew
rlabel locali s -12317 41994 -12269 42046 4 VSS
port 42 nsew
rlabel locali s -4820 42470 -3747 44102 4 VSS
port 42 nsew
rlabel locali s -13915 42459 -11613 42720 4 VSS
port 42 nsew
rlabel locali s -12732 43876 -12664 43885 4 VSS
port 42 nsew
rlabel locali s -12732 43885 -12505 43919 4 VSS
port 42 nsew
rlabel locali s -12732 43919 -12664 44081 4 VSS
port 42 nsew
rlabel locali s -4080 44102 -3747 51579 4 VSS
port 42 nsew
rlabel locali s -12732 44081 -12505 44115 4 VSS
port 42 nsew
rlabel locali s -12732 44115 -12664 44277 4 VSS
port 42 nsew
rlabel locali s -12996 44138 -12957 44139 4 VSS
port 42 nsew
rlabel locali s -12998 44139 -12938 44243 4 VSS
port 42 nsew
rlabel locali s -13915 42720 -13654 44243 4 VSS
port 42 nsew
rlabel locali s -13915 44243 -12938 44271 4 VSS
port 42 nsew
rlabel locali s -12732 44277 -12505 44311 4 VSS
port 42 nsew
rlabel locali s -12732 44311 -12664 44767 4 VSS
port 42 nsew
rlabel locali s -12732 44767 -12505 44801 4 VSS
port 42 nsew
rlabel locali s -12732 44801 -12664 44963 4 VSS
port 42 nsew
rlabel locali s -12732 44963 -12505 44997 4 VSS
port 42 nsew
rlabel locali s -12732 44997 -12664 45159 4 VSS
port 42 nsew
rlabel locali s -12732 45159 -12505 45193 4 VSS
port 42 nsew
rlabel locali s -12732 45193 -12664 45292 4 VSS
port 42 nsew
rlabel locali s -13915 44271 -12957 44504 4 VSS
port 42 nsew
rlabel locali s -12996 44504 -12957 45897 4 VSS
port 42 nsew
rlabel locali s -13112 45672 -13044 45771 4 VSS
port 42 nsew
rlabel locali s -13271 45771 -13044 45805 4 VSS
port 42 nsew
rlabel locali s -13112 45805 -13044 45897 4 VSS
port 42 nsew
rlabel locali s -13112 45897 -12957 45967 4 VSS
port 42 nsew
rlabel locali s -13271 45967 -12957 46001 4 VSS
port 42 nsew
rlabel locali s -13112 46001 -12957 46008 4 VSS
port 42 nsew
rlabel locali s -12732 46501 -12664 46510 4 VSS
port 42 nsew
rlabel locali s -12732 46510 -12505 46544 4 VSS
port 42 nsew
rlabel locali s -12732 46544 -12664 46706 4 VSS
port 42 nsew
rlabel locali s -12732 46706 -12505 46740 4 VSS
port 42 nsew
rlabel locali s -12732 46740 -12664 46902 4 VSS
port 42 nsew
rlabel locali s -12996 46008 -12957 46772 4 VSS
port 42 nsew
rlabel locali s -13112 46008 -13044 46163 4 VSS
port 42 nsew
rlabel locali s -13271 46163 -13044 46183 4 VSS
port 42 nsew
rlabel locali s -13271 46183 -13042 46197 4 VSS
port 42 nsew
rlabel locali s -13112 46197 -13042 46206 4 VSS
port 42 nsew
rlabel locali s -13110 46206 -13042 46509 4 VSS
port 42 nsew
rlabel locali s -13112 46509 -13042 46608 4 VSS
port 42 nsew
rlabel locali s -13271 46608 -13042 46642 4 VSS
port 42 nsew
rlabel locali s -13112 46642 -13042 46703 4 VSS
port 42 nsew
rlabel locali s -12732 46902 -12505 46936 4 VSS
port 42 nsew
rlabel locali s -12998 46772 -12938 46775 4 VSS
port 42 nsew
rlabel locali s -13112 46703 -13044 46775 4 VSS
port 42 nsew
rlabel locali s -13112 46775 -12938 46804 4 VSS
port 42 nsew
rlabel locali s -13271 46804 -12938 46838 4 VSS
port 42 nsew
rlabel locali s -13112 46838 -12938 46886 4 VSS
port 42 nsew
rlabel locali s -12998 46886 -12938 46909 4 VSS
port 42 nsew
rlabel locali s -12732 46936 -12664 47467 4 VSS
port 42 nsew
rlabel locali s -12732 47467 -12505 47501 4 VSS
port 42 nsew
rlabel locali s -12732 47501 -12664 47663 4 VSS
port 42 nsew
rlabel locali s -12732 47663 -12505 47697 4 VSS
port 42 nsew
rlabel locali s -12732 47697 -12664 47859 4 VSS
port 42 nsew
rlabel locali s -12732 47859 -12505 47893 4 VSS
port 42 nsew
rlabel locali s -12732 47893 -12664 47992 4 VSS
port 42 nsew
rlabel locali s -12996 46909 -12957 48573 4 VSS
port 42 nsew
rlabel locali s -13112 46886 -13044 47000 4 VSS
port 42 nsew
rlabel locali s -13271 47000 -13044 47034 4 VSS
port 42 nsew
rlabel locali s -13112 47034 -13044 47043 4 VSS
port 42 nsew
rlabel locali s -13112 48372 -13044 48471 4 VSS
port 42 nsew
rlabel locali s -13271 48471 -13044 48505 4 VSS
port 42 nsew
rlabel locali s -13112 48505 -13044 48573 4 VSS
port 42 nsew
rlabel locali s -13112 48573 -12957 48667 4 VSS
port 42 nsew
rlabel locali s -13271 48667 -12957 48684 4 VSS
port 42 nsew
rlabel locali s -12732 49201 -12664 49210 4 VSS
port 42 nsew
rlabel locali s -12732 49210 -12505 49244 4 VSS
port 42 nsew
rlabel locali s -12732 49244 -12664 49406 4 VSS
port 42 nsew
rlabel locali s -12996 48684 -12957 49369 4 VSS
port 42 nsew
rlabel locali s -13271 48684 -13044 48701 4 VSS
port 42 nsew
rlabel locali s -13112 48701 -13044 48863 4 VSS
port 42 nsew
rlabel locali s -13271 48863 -13044 48897 4 VSS
port 42 nsew
rlabel locali s -13112 48897 -13044 49308 4 VSS
port 42 nsew
rlabel locali s -13271 49308 -13044 49342 4 VSS
port 42 nsew
rlabel locali s -12732 49406 -12505 49440 4 VSS
port 42 nsew
rlabel locali s -12732 49440 -12664 49602 4 VSS
port 42 nsew
rlabel locali s -13004 49369 -12944 49384 4 VSS
port 42 nsew
rlabel locali s -13112 49342 -13044 49384 4 VSS
port 42 nsew
rlabel locali s -13112 49384 -12944 49495 4 VSS
port 42 nsew
rlabel locali s -13004 49495 -12944 49506 4 VSS
port 42 nsew
rlabel locali s -13112 49495 -13044 49504 4 VSS
port 42 nsew
rlabel locali s -12996 49506 -12957 49523 4 VSS
port 42 nsew
rlabel locali s -12732 49602 -12505 49636 4 VSS
port 42 nsew
rlabel locali s -12732 49636 -12664 49735 4 VSS
port 42 nsew
rlabel locali s -13271 49504 -13044 49538 4 VSS
port 42 nsew
rlabel locali s -13112 49538 -13044 49700 4 VSS
port 42 nsew
rlabel locali s -13271 49700 -13044 49734 4 VSS
port 42 nsew
rlabel locali s -13112 49734 -13044 49743 4 VSS
port 42 nsew
rlabel locali s -7694 50681 -7588 50785 4 VSS
port 42 nsew
rlabel locali s -10318 50652 -10229 50781 4 VSS
port 42 nsew
rlabel locali s -10470 50781 -10229 50785 4 VSS
port 42 nsew
rlabel locali s -7840 50785 -7588 50790 4 VSS
port 42 nsew
rlabel locali s -8011 50790 -7588 50824 4 VSS
port 42 nsew
rlabel locali s -10629 50785 -10229 50819 4 VSS
port 42 nsew
rlabel locali s -7840 50824 -7588 50833 4 VSS
port 42 nsew
rlabel locali s -10470 50819 -10229 50825 4 VSS
port 42 nsew
rlabel locali s -7694 50833 -7588 50979 4 VSS
port 42 nsew
rlabel locali s -10318 50825 -10229 50975 4 VSS
port 42 nsew
rlabel locali s -7843 50979 -7588 50986 4 VSS
port 42 nsew
rlabel locali s -10469 50975 -10229 50981 4 VSS
port 42 nsew
rlabel locali s -6124 50996 -5618 51579 4 VSS
port 42 nsew
rlabel locali s -8011 50986 -7588 51020 4 VSS
port 42 nsew
rlabel locali s -10629 50981 -10229 51015 4 VSS
port 42 nsew
rlabel locali s -10469 51015 -10229 51019 4 VSS
port 42 nsew
rlabel locali s -7843 51020 -7588 51027 4 VSS
port 42 nsew
rlabel locali s -7694 51027 -7588 51579 4 VSS
port 42 nsew
rlabel locali s -7694 51579 -3747 51706 4 VSS
port 42 nsew
rlabel locali s -10318 51019 -10229 51706 4 VSS
port 42 nsew
rlabel locali s -10318 51706 -3747 51727 4 VSS
port 42 nsew
rlabel locali s -10470 51727 -3747 51731 4 VSS
port 42 nsew
rlabel locali s -10629 51731 -3747 51765 4 VSS
port 42 nsew
rlabel locali s -10470 51765 -3747 51771 4 VSS
port 42 nsew
rlabel locali s -10318 51771 -3747 51855 4 VSS
port 42 nsew
rlabel locali s -7694 51855 -3747 52124 4 VSS
port 42 nsew
rlabel locali s -10318 51855 -10229 51921 4 VSS
port 42 nsew
rlabel locali s -10469 51921 -10229 51927 4 VSS
port 42 nsew
rlabel locali s -10629 51927 -10229 51961 4 VSS
port 42 nsew
rlabel locali s -10469 51961 -10229 51965 4 VSS
port 42 nsew
rlabel locali s -6124 52124 -5618 61325 4 VSS
port 42 nsew
rlabel locali s -7694 52124 -7588 52267 4 VSS
port 42 nsew
rlabel locali s -8556 52004 -8488 52013 4 VSS
port 42 nsew
rlabel locali s -8715 52013 -8488 52047 4 VSS
port 42 nsew
rlabel locali s -8556 52047 -8488 52209 4 VSS
port 42 nsew
rlabel locali s -8715 52209 -8488 52243 4 VSS
port 42 nsew
rlabel locali s -8263 52266 -8224 52267 4 VSS
port 42 nsew
rlabel locali s -8282 52267 -7588 52399 4 VSS
port 42 nsew
rlabel locali s -8263 52399 -7588 52451 4 VSS
port 42 nsew
rlabel locali s -8176 53800 -8108 53899 4 VSS
port 42 nsew
rlabel locali s -8176 53899 -7949 53933 4 VSS
port 42 nsew
rlabel locali s -8176 53933 -8108 54025 4 VSS
port 42 nsew
rlabel locali s -8263 52451 -8224 54025 4 VSS
port 42 nsew
rlabel locali s -8556 52243 -8488 52405 4 VSS
port 42 nsew
rlabel locali s -8715 52405 -8488 52439 4 VSS
port 42 nsew
rlabel locali s -8556 52439 -8488 52895 4 VSS
port 42 nsew
rlabel locali s -10318 51965 -10229 52501 4 VSS
port 42 nsew
rlabel locali s -10318 52501 -10186 52647 4 VSS
port 42 nsew
rlabel locali s -10748 52647 -10186 52681 4 VSS
port 42 nsew
rlabel locali s -8715 52895 -8488 52929 4 VSS
port 42 nsew
rlabel locali s -8556 52929 -8488 53091 4 VSS
port 42 nsew
rlabel locali s -8715 53091 -8488 53125 4 VSS
port 42 nsew
rlabel locali s -8556 53125 -8488 53287 4 VSS
port 42 nsew
rlabel locali s -8715 53287 -8488 53321 4 VSS
port 42 nsew
rlabel locali s -8556 53321 -8488 53420 4 VSS
port 42 nsew
rlabel locali s -8263 54025 -8108 54095 4 VSS
port 42 nsew
rlabel locali s -8263 54095 -7949 54129 4 VSS
port 42 nsew
rlabel locali s -10251 52681 -10186 53679 4 VSS
port 42 nsew
rlabel locali s -10647 53679 -10186 53713 4 VSS
port 42 nsew
rlabel locali s -10251 53713 -10186 53781 4 VSS
port 42 nsew
rlabel locali s -10302 53781 -10186 54015 4 VSS
port 42 nsew
rlabel locali s -10766 54015 -10186 54096 4 VSS
port 42 nsew
rlabel locali s -10267 54096 -10186 54097 4 VSS
port 42 nsew
rlabel locali s -8263 54129 -8108 54136 4 VSS
port 42 nsew
rlabel locali s -8176 54136 -8108 54291 4 VSS
port 42 nsew
rlabel locali s -8176 54291 -7949 54311 4 VSS
port 42 nsew
rlabel locali s -8178 54311 -7949 54325 4 VSS
port 42 nsew
rlabel locali s -8178 54325 -8108 54334 4 VSS
port 42 nsew
rlabel locali s -8178 54334 -8110 54637 4 VSS
port 42 nsew
rlabel locali s -8178 54637 -8108 54736 4 VSS
port 42 nsew
rlabel locali s -8178 54736 -7949 54770 4 VSS
port 42 nsew
rlabel locali s -8178 54770 -8108 54831 4 VSS
port 42 nsew
rlabel locali s -8176 54831 -8108 54903 4 VSS
port 42 nsew
rlabel locali s -8263 54136 -8224 54900 4 VSS
port 42 nsew
rlabel locali s -10766 54096 -10608 54399 4 VSS
port 42 nsew
rlabel locali s -10809 54399 -10608 54408 4 VSS
port 42 nsew
rlabel locali s -10968 54408 -10608 54425 4 VSS
port 42 nsew
rlabel locali s -10968 54425 -10605 54442 4 VSS
port 42 nsew
rlabel locali s -10809 54442 -10605 54458 4 VSS
port 42 nsew
rlabel locali s -10809 54458 -10293 54492 4 VSS
port 42 nsew
rlabel locali s -10809 54492 -10605 54604 4 VSS
port 42 nsew
rlabel locali s -8556 54629 -8488 54638 4 VSS
port 42 nsew
rlabel locali s -10968 54604 -10605 54638 4 VSS
port 42 nsew
rlabel locali s -8715 54638 -8488 54672 4 VSS
port 42 nsew
rlabel locali s -8556 54672 -8488 54834 4 VSS
port 42 nsew
rlabel locali s -10809 54638 -10605 54800 4 VSS
port 42 nsew
rlabel locali s -10968 54800 -10605 54834 4 VSS
port 42 nsew
rlabel locali s -8715 54834 -8488 54868 4 VSS
port 42 nsew
rlabel locali s -8282 54900 -8222 54903 4 VSS
port 42 nsew
rlabel locali s -8282 54903 -8108 54932 4 VSS
port 42 nsew
rlabel locali s -8282 54932 -7949 54966 4 VSS
port 42 nsew
rlabel locali s -8282 54966 -8108 55014 4 VSS
port 42 nsew
rlabel locali s -8176 55014 -8108 55128 4 VSS
port 42 nsew
rlabel locali s -8282 55014 -8222 55037 4 VSS
port 42 nsew
rlabel locali s -8556 54868 -8488 55030 4 VSS
port 42 nsew
rlabel locali s -10809 54834 -10605 54904 4 VSS
port 42 nsew
rlabel locali s -10809 54904 -10608 54994 4 VSS
port 42 nsew
rlabel locali s -8176 55128 -7949 55162 4 VSS
port 42 nsew
rlabel locali s -8176 55162 -8108 55171 4 VSS
port 42 nsew
rlabel locali s -8176 56500 -8108 56599 4 VSS
port 42 nsew
rlabel locali s -8176 56599 -7949 56633 4 VSS
port 42 nsew
rlabel locali s -8176 56633 -8108 56701 4 VSS
port 42 nsew
rlabel locali s -8263 55037 -8224 56701 4 VSS
port 42 nsew
rlabel locali s -8715 55030 -8488 55064 4 VSS
port 42 nsew
rlabel locali s -10809 54994 -9474 55064 4 VSS
port 42 nsew
rlabel locali s -8556 55064 -8488 55595 4 VSS
port 42 nsew
rlabel locali s -9571 55064 -9474 55288 4 VSS
port 42 nsew
rlabel locali s -10392 55288 -9474 55322 4 VSS
port 42 nsew
rlabel locali s -8715 55595 -8488 55629 4 VSS
port 42 nsew
rlabel locali s -8556 55629 -8488 55791 4 VSS
port 42 nsew
rlabel locali s -9571 55322 -9474 55688 4 VSS
port 42 nsew
rlabel locali s -10392 55688 -9474 55722 4 VSS
port 42 nsew
rlabel locali s -8715 55791 -8488 55825 4 VSS
port 42 nsew
rlabel locali s -8556 55825 -8488 55987 4 VSS
port 42 nsew
rlabel locali s -8715 55987 -8488 56021 4 VSS
port 42 nsew
rlabel locali s -8556 56021 -8488 56120 4 VSS
port 42 nsew
rlabel locali s -8263 56701 -8108 56795 4 VSS
port 42 nsew
rlabel locali s -8263 56795 -7949 56812 4 VSS
port 42 nsew
rlabel locali s -8176 56812 -7949 56829 4 VSS
port 42 nsew
rlabel locali s -8176 56829 -8108 56991 4 VSS
port 42 nsew
rlabel locali s -8176 56991 -7949 57025 4 VSS
port 42 nsew
rlabel locali s -8176 57025 -8108 57436 4 VSS
port 42 nsew
rlabel locali s -8176 57436 -7949 57470 4 VSS
port 42 nsew
rlabel locali s -8176 57470 -8108 57512 4 VSS
port 42 nsew
rlabel locali s -8263 56812 -8224 57497 4 VSS
port 42 nsew
rlabel locali s -9571 55722 -9474 56288 4 VSS
port 42 nsew
rlabel locali s -10392 56288 -9474 56322 4 VSS
port 42 nsew
rlabel locali s -9571 56322 -9474 56688 4 VSS
port 42 nsew
rlabel locali s -10392 56688 -9474 56722 4 VSS
port 42 nsew
rlabel locali s -9571 56722 -9474 57288 4 VSS
port 42 nsew
rlabel locali s -10392 57288 -9474 57322 4 VSS
port 42 nsew
rlabel locali s -8556 57329 -8488 57338 4 VSS
port 42 nsew
rlabel locali s -8715 57338 -8488 57372 4 VSS
port 42 nsew
rlabel locali s -8276 57497 -8216 57512 4 VSS
port 42 nsew
rlabel locali s -8276 57512 -8108 57623 4 VSS
port 42 nsew
rlabel locali s -8176 57623 -8108 57632 4 VSS
port 42 nsew
rlabel locali s -8176 57632 -7949 57666 4 VSS
port 42 nsew
rlabel locali s -8276 57623 -8216 57634 4 VSS
port 42 nsew
rlabel locali s -8556 57372 -8488 57534 4 VSS
port 42 nsew
rlabel locali s -8715 57534 -8488 57568 4 VSS
port 42 nsew
rlabel locali s -8263 57634 -8224 57651 4 VSS
port 42 nsew
rlabel locali s -8176 57666 -8108 57828 4 VSS
port 42 nsew
rlabel locali s -8176 57828 -7949 57862 4 VSS
port 42 nsew
rlabel locali s -8176 57862 -8108 57871 4 VSS
port 42 nsew
rlabel locali s -8556 57568 -8488 57730 4 VSS
port 42 nsew
rlabel locali s -9571 57322 -9474 57688 4 VSS
port 42 nsew
rlabel locali s -10392 57688 -9474 57722 4 VSS
port 42 nsew
rlabel locali s -8715 57730 -8488 57764 4 VSS
port 42 nsew
rlabel locali s -8556 57764 -8488 57863 4 VSS
port 42 nsew
rlabel locali s -9571 57722 -9474 57918 4 VSS
port 42 nsew
rlabel locali s -6838 60229 -6752 60369 4 VSS
port 42 nsew
rlabel locali s -9103 60225 -9042 60342 4 VSS
port 42 nsew
rlabel locali s -9103 60342 -8990 60343 4 VSS
port 42 nsew
rlabel locali s -7094 60369 -6752 60403 4 VSS
port 42 nsew
rlabel locali s -9103 60343 -8682 60377 4 VSS
port 42 nsew
rlabel locali s -6838 60403 -6752 60565 4 VSS
port 42 nsew
rlabel locali s -7094 60565 -6752 60599 4 VSS
port 42 nsew
rlabel locali s -6838 60599 -6752 61081 4 VSS
port 42 nsew
rlabel locali s -9103 60377 -9042 60667 4 VSS
port 42 nsew
rlabel locali s -9103 60667 -9024 60674 4 VSS
port 42 nsew
rlabel locali s -10291 60221 -10205 60361 4 VSS
port 42 nsew
rlabel locali s -12556 60217 -12495 60334 4 VSS
port 42 nsew
rlabel locali s -12556 60334 -12443 60335 4 VSS
port 42 nsew
rlabel locali s -10547 60361 -10205 60395 4 VSS
port 42 nsew
rlabel locali s -12556 60335 -12135 60369 4 VSS
port 42 nsew
rlabel locali s -10291 60395 -10205 60557 4 VSS
port 42 nsew
rlabel locali s -10547 60557 -10205 60591 4 VSS
port 42 nsew
rlabel locali s -8617 60812 -8531 60952 4 VSS
port 42 nsew
rlabel locali s -8617 60952 -8375 60986 4 VSS
port 42 nsew
rlabel locali s -6838 61081 -6585 61167 4 VSS
port 42 nsew
rlabel locali s -8617 60986 -8531 61056 4 VSS
port 42 nsew
rlabel locali s -9085 60674 -9024 61056 4 VSS
port 42 nsew
rlabel locali s -9493 61056 -8531 61117 4 VSS
port 42 nsew
rlabel locali s -10291 60591 -10205 61073 4 VSS
port 42 nsew
rlabel locali s -12556 60369 -12495 60659 4 VSS
port 42 nsew
rlabel locali s -12556 60659 -12477 60666 4 VSS
port 42 nsew
rlabel locali s -12070 60804 -11984 60944 4 VSS
port 42 nsew
rlabel locali s -12070 60944 -11828 60978 4 VSS
port 42 nsew
rlabel locali s -8617 61117 -8531 61148 4 VSS
port 42 nsew
rlabel locali s -6671 61167 -6585 61325 4 VSS
port 42 nsew
rlabel locali s -8617 61148 -8375 61182 4 VSS
port 42 nsew
rlabel locali s -6671 61325 -5618 61341 4 VSS
port 42 nsew
rlabel locali s -6708 61341 -5618 61342 4 VSS
port 42 nsew
rlabel locali s -7016 61342 -5618 61376 4 VSS
port 42 nsew
rlabel locali s -6671 61376 -5618 61608 4 VSS
port 42 nsew
rlabel locali s -8617 61182 -8531 61427 4 VSS
port 42 nsew
rlabel locali s -6124 61608 -5618 69724 4 VSS
port 42 nsew
rlabel locali s -6671 61608 -6585 61666 4 VSS
port 42 nsew
rlabel locali s -6674 61666 -6585 61746 4 VSS
port 42 nsew
rlabel locali s -6674 61746 -6613 62055 4 VSS
port 42 nsew
rlabel locali s -9493 61117 -9380 61783 4 VSS
port 42 nsew
rlabel locali s -10291 61073 -10038 61159 4 VSS
port 42 nsew
rlabel locali s -12070 60978 -11984 61048 4 VSS
port 42 nsew
rlabel locali s -12538 60666 -12477 61048 4 VSS
port 42 nsew
rlabel locali s -12946 61048 -11984 61109 4 VSS
port 42 nsew
rlabel locali s -12070 61109 -11984 61140 4 VSS
port 42 nsew
rlabel locali s -10124 61159 -10038 61333 4 VSS
port 42 nsew
rlabel locali s -12070 61140 -11828 61174 4 VSS
port 42 nsew
rlabel locali s -10161 61333 -10038 61334 4 VSS
port 42 nsew
rlabel locali s -10469 61334 -10038 61368 4 VSS
port 42 nsew
rlabel locali s -10124 61368 -10038 61658 4 VSS
port 42 nsew
rlabel locali s -12070 61174 -11984 61419 4 VSS
port 42 nsew
rlabel locali s -10127 61658 -10038 61738 4 VSS
port 42 nsew
rlabel locali s -9493 61783 -9262 61790 4 VSS
port 42 nsew
rlabel locali s -7167 61811 -7081 61951 4 VSS
port 42 nsew
rlabel locali s -9493 61790 -8968 61824 4 VSS
port 42 nsew
rlabel locali s -9493 61824 -9262 61830 4 VSS
port 42 nsew
rlabel locali s -7323 61951 -7081 61985 4 VSS
port 42 nsew
rlabel locali s -9493 61830 -9380 61979 4 VSS
port 42 nsew
rlabel locali s -7167 61985 -7081 62055 4 VSS
port 42 nsew
rlabel locali s -9493 61979 -9261 61986 4 VSS
port 42 nsew
rlabel locali s -9493 61986 -8968 62020 4 VSS
port 42 nsew
rlabel locali s -9493 62020 -9261 62026 4 VSS
port 42 nsew
rlabel locali s -7167 62055 -6613 62116 4 VSS
port 42 nsew
rlabel locali s -7167 62116 -7081 62147 4 VSS
port 42 nsew
rlabel locali s -7323 62147 -7081 62181 4 VSS
port 42 nsew
rlabel locali s -7167 62181 -7081 62596 4 VSS
port 42 nsew
rlabel locali s -9493 62026 -9380 62221 4 VSS
port 42 nsew
rlabel locali s -10127 61738 -10066 62047 4 VSS
port 42 nsew
rlabel locali s -12946 61109 -12833 61775 4 VSS
port 42 nsew
rlabel locali s -12946 61775 -12715 61782 4 VSS
port 42 nsew
rlabel locali s -10620 61803 -10534 61943 4 VSS
port 42 nsew
rlabel locali s -12946 61782 -12421 61816 4 VSS
port 42 nsew
rlabel locali s -12946 61816 -12715 61822 4 VSS
port 42 nsew
rlabel locali s -10776 61943 -10534 61977 4 VSS
port 42 nsew
rlabel locali s -12946 61822 -12833 61971 4 VSS
port 42 nsew
rlabel locali s -10620 61977 -10534 62047 4 VSS
port 42 nsew
rlabel locali s -12946 61971 -12714 61978 4 VSS
port 42 nsew
rlabel locali s -12946 61978 -12421 62012 4 VSS
port 42 nsew
rlabel locali s -12946 62012 -12714 62018 4 VSS
port 42 nsew
rlabel locali s -10620 62047 -10066 62108 4 VSS
port 42 nsew
rlabel locali s -9493 62221 -9251 62228 4 VSS
port 42 nsew
rlabel locali s -9493 62228 -8968 62262 4 VSS
port 42 nsew
rlabel locali s -9493 62262 -9251 62268 4 VSS
port 42 nsew
rlabel locali s -9493 62268 -9380 63145 4 VSS
port 42 nsew
rlabel locali s -10620 62108 -10534 62139 4 VSS
port 42 nsew
rlabel locali s -10776 62139 -10534 62173 4 VSS
port 42 nsew
rlabel locali s -10620 62173 -10534 62588 4 VSS
port 42 nsew
rlabel locali s -12946 62018 -12833 62213 4 VSS
port 42 nsew
rlabel locali s -12946 62213 -12704 62220 4 VSS
port 42 nsew
rlabel locali s -12946 62220 -12421 62254 4 VSS
port 42 nsew
rlabel locali s -12946 62254 -12704 62260 4 VSS
port 42 nsew
rlabel locali s -12946 62260 -12833 62525 4 VSS
port 42 nsew
rlabel locali s -9493 63145 -9312 63258 4 VSS
port 42 nsew
rlabel locali s -9425 63258 -9312 63606 4 VSS
port 42 nsew
rlabel locali s -9477 63606 -9312 63682 4 VSS
port 42 nsew
rlabel locali s -9477 63682 -9201 63684 4 VSS
port 42 nsew
rlabel locali s -9477 63684 -8910 63718 4 VSS
port 42 nsew
rlabel locali s -9477 63718 -9201 63719 4 VSS
port 42 nsew
rlabel locali s -9477 63719 -9312 63756 4 VSS
port 42 nsew
rlabel locali s -9477 63756 -9316 64474 4 VSS
port 42 nsew
rlabel locali s -9477 64474 -9201 64475 4 VSS
port 42 nsew
rlabel locali s -9477 64475 -8710 64509 4 VSS
port 42 nsew
rlabel locali s -9477 64509 -9201 64511 4 VSS
port 42 nsew
rlabel locali s -9477 64511 -9316 64602 4 VSS
port 42 nsew
rlabel locali s -9477 64602 -9200 64605 4 VSS
port 42 nsew
rlabel locali s -9477 64605 -8710 64639 4 VSS
port 42 nsew
rlabel locali s -9477 64639 -9316 64929 4 VSS
port 42 nsew
rlabel locali s -10322 63889 -10236 64029 4 VSS
port 42 nsew
rlabel locali s -12587 63885 -12526 64002 4 VSS
port 42 nsew
rlabel locali s -12587 64002 -12474 64003 4 VSS
port 42 nsew
rlabel locali s -10578 64029 -10236 64063 4 VSS
port 42 nsew
rlabel locali s -12587 64003 -12166 64037 4 VSS
port 42 nsew
rlabel locali s -10322 64063 -10236 64225 4 VSS
port 42 nsew
rlabel locali s -10578 64225 -10236 64259 4 VSS
port 42 nsew
rlabel locali s -10322 64259 -10236 64741 4 VSS
port 42 nsew
rlabel locali s -12587 64037 -12526 64327 4 VSS
port 42 nsew
rlabel locali s -12587 64327 -12508 64334 4 VSS
port 42 nsew
rlabel locali s -12101 64472 -12015 64612 4 VSS
port 42 nsew
rlabel locali s -12101 64612 -11859 64646 4 VSS
port 42 nsew
rlabel locali s -9477 64929 -9199 64931 4 VSS
port 42 nsew
rlabel locali s -9477 64931 -8910 64965 4 VSS
port 42 nsew
rlabel locali s -9477 64965 -9199 64966 4 VSS
port 42 nsew
rlabel locali s -9477 64966 -9316 65079 4 VSS
port 42 nsew
rlabel locali s -10322 64741 -10069 64827 4 VSS
port 42 nsew
rlabel locali s -12101 64646 -12015 64716 4 VSS
port 42 nsew
rlabel locali s -12569 64334 -12508 64716 4 VSS
port 42 nsew
rlabel locali s -12977 64716 -12015 64777 4 VSS
port 42 nsew
rlabel locali s -12101 64777 -12015 64808 4 VSS
port 42 nsew
rlabel locali s -10155 64827 -10069 65001 4 VSS
port 42 nsew
rlabel locali s -12101 64808 -11859 64842 4 VSS
port 42 nsew
rlabel locali s -10192 65001 -10069 65002 4 VSS
port 42 nsew
rlabel locali s -10500 65002 -10069 65036 4 VSS
port 42 nsew
rlabel locali s -10155 65036 -10069 65326 4 VSS
port 42 nsew
rlabel locali s -12101 64842 -12015 65087 4 VSS
port 42 nsew
rlabel locali s -10158 65326 -10069 65406 4 VSS
port 42 nsew
rlabel locali s -10158 65406 -10097 65715 4 VSS
port 42 nsew
rlabel locali s -12977 64777 -12864 65443 4 VSS
port 42 nsew
rlabel locali s -12977 65443 -12746 65450 4 VSS
port 42 nsew
rlabel locali s -10651 65471 -10565 65611 4 VSS
port 42 nsew
rlabel locali s -12977 65450 -12452 65484 4 VSS
port 42 nsew
rlabel locali s -12977 65484 -12746 65490 4 VSS
port 42 nsew
rlabel locali s -10807 65611 -10565 65645 4 VSS
port 42 nsew
rlabel locali s -12977 65490 -12864 65639 4 VSS
port 42 nsew
rlabel locali s -10651 65645 -10565 65715 4 VSS
port 42 nsew
rlabel locali s -12977 65639 -12745 65646 4 VSS
port 42 nsew
rlabel locali s -12977 65646 -12452 65680 4 VSS
port 42 nsew
rlabel locali s -12977 65680 -12745 65686 4 VSS
port 42 nsew
rlabel locali s -10651 65715 -10097 65776 4 VSS
port 42 nsew
rlabel locali s -10651 65776 -10565 65807 4 VSS
port 42 nsew
rlabel locali s -10807 65807 -10565 65841 4 VSS
port 42 nsew
rlabel locali s -10651 65841 -10565 66256 4 VSS
port 42 nsew
rlabel locali s -12977 65686 -12864 65881 4 VSS
port 42 nsew
rlabel locali s -12977 65881 -12735 65888 4 VSS
port 42 nsew
rlabel locali s -12977 65888 -12452 65922 4 VSS
port 42 nsew
rlabel locali s -12977 65922 -12735 65928 4 VSS
port 42 nsew
rlabel locali s -12977 65928 -12864 66193 4 VSS
port 42 nsew
rlabel locali s -6849 68669 -6763 68809 4 VSS
port 42 nsew
rlabel locali s -9114 68665 -9053 68782 4 VSS
port 42 nsew
rlabel locali s -9114 68782 -9001 68783 4 VSS
port 42 nsew
rlabel locali s -7105 68809 -6763 68843 4 VSS
port 42 nsew
rlabel locali s -9114 68783 -8693 68817 4 VSS
port 42 nsew
rlabel locali s -6849 68843 -6763 69005 4 VSS
port 42 nsew
rlabel locali s -7105 69005 -6763 69039 4 VSS
port 42 nsew
rlabel locali s -6849 69039 -6763 69521 4 VSS
port 42 nsew
rlabel locali s -9114 68817 -9053 69107 4 VSS
port 42 nsew
rlabel locali s -9114 69107 -9035 69114 4 VSS
port 42 nsew
rlabel locali s -10302 68661 -10216 68801 4 VSS
port 42 nsew
rlabel locali s -12567 68657 -12506 68774 4 VSS
port 42 nsew
rlabel locali s -12567 68774 -12454 68775 4 VSS
port 42 nsew
rlabel locali s -10558 68801 -10216 68835 4 VSS
port 42 nsew
rlabel locali s -12567 68775 -12146 68809 4 VSS
port 42 nsew
rlabel locali s -10302 68835 -10216 68997 4 VSS
port 42 nsew
rlabel locali s -10558 68997 -10216 69031 4 VSS
port 42 nsew
rlabel locali s -8628 69252 -8542 69392 4 VSS
port 42 nsew
rlabel locali s -8628 69392 -8386 69426 4 VSS
port 42 nsew
rlabel locali s -6849 69521 -6596 69607 4 VSS
port 42 nsew
rlabel locali s -8628 69426 -8542 69496 4 VSS
port 42 nsew
rlabel locali s -9096 69114 -9035 69496 4 VSS
port 42 nsew
rlabel locali s -9504 69496 -8542 69557 4 VSS
port 42 nsew
rlabel locali s -10302 69031 -10216 69513 4 VSS
port 42 nsew
rlabel locali s -12567 68809 -12506 69099 4 VSS
port 42 nsew
rlabel locali s -12567 69099 -12488 69106 4 VSS
port 42 nsew
rlabel locali s -12081 69244 -11995 69384 4 VSS
port 42 nsew
rlabel locali s -12081 69384 -11839 69418 4 VSS
port 42 nsew
rlabel locali s -8628 69557 -8542 69588 4 VSS
port 42 nsew
rlabel locali s -6682 69607 -6596 69724 4 VSS
port 42 nsew
rlabel locali s -8628 69588 -8386 69622 4 VSS
port 42 nsew
rlabel locali s -6682 69724 -5618 69781 4 VSS
port 42 nsew
rlabel locali s -6719 69781 -5618 69782 4 VSS
port 42 nsew
rlabel locali s -7027 69782 -5618 69816 4 VSS
port 42 nsew
rlabel locali s -6682 69816 -5618 70007 4 VSS
port 42 nsew
rlabel locali s -8628 69622 -8542 69867 4 VSS
port 42 nsew
rlabel locali s -6124 70007 -5618 78636 4 VSS
port 42 nsew
rlabel locali s -6682 70007 -6596 70106 4 VSS
port 42 nsew
rlabel locali s -6685 70106 -6596 70186 4 VSS
port 42 nsew
rlabel locali s -6685 70186 -6624 70495 4 VSS
port 42 nsew
rlabel locali s -9504 69557 -9391 70223 4 VSS
port 42 nsew
rlabel locali s -10302 69513 -10049 69599 4 VSS
port 42 nsew
rlabel locali s -12081 69418 -11995 69488 4 VSS
port 42 nsew
rlabel locali s -12549 69106 -12488 69488 4 VSS
port 42 nsew
rlabel locali s -12957 69488 -11995 69549 4 VSS
port 42 nsew
rlabel locali s -12081 69549 -11995 69580 4 VSS
port 42 nsew
rlabel locali s -10135 69599 -10049 69773 4 VSS
port 42 nsew
rlabel locali s -12081 69580 -11839 69614 4 VSS
port 42 nsew
rlabel locali s -10172 69773 -10049 69774 4 VSS
port 42 nsew
rlabel locali s -10480 69774 -10049 69808 4 VSS
port 42 nsew
rlabel locali s -10135 69808 -10049 70098 4 VSS
port 42 nsew
rlabel locali s -12081 69614 -11995 69859 4 VSS
port 42 nsew
rlabel locali s -10138 70098 -10049 70178 4 VSS
port 42 nsew
rlabel locali s -9504 70223 -9273 70230 4 VSS
port 42 nsew
rlabel locali s -7178 70251 -7092 70391 4 VSS
port 42 nsew
rlabel locali s -9504 70230 -8979 70264 4 VSS
port 42 nsew
rlabel locali s -9504 70264 -9273 70270 4 VSS
port 42 nsew
rlabel locali s -7334 70391 -7092 70425 4 VSS
port 42 nsew
rlabel locali s -9504 70270 -9391 70419 4 VSS
port 42 nsew
rlabel locali s -7178 70425 -7092 70495 4 VSS
port 42 nsew
rlabel locali s -9504 70419 -9272 70426 4 VSS
port 42 nsew
rlabel locali s -9504 70426 -8979 70460 4 VSS
port 42 nsew
rlabel locali s -9504 70460 -9272 70466 4 VSS
port 42 nsew
rlabel locali s -7178 70495 -6624 70556 4 VSS
port 42 nsew
rlabel locali s -7178 70556 -7092 70587 4 VSS
port 42 nsew
rlabel locali s -7334 70587 -7092 70621 4 VSS
port 42 nsew
rlabel locali s -7178 70621 -7092 71036 4 VSS
port 42 nsew
rlabel locali s -9504 70466 -9391 70661 4 VSS
port 42 nsew
rlabel locali s -10138 70178 -10077 70487 4 VSS
port 42 nsew
rlabel locali s -12957 69549 -12844 70215 4 VSS
port 42 nsew
rlabel locali s -12957 70215 -12726 70222 4 VSS
port 42 nsew
rlabel locali s -10631 70243 -10545 70383 4 VSS
port 42 nsew
rlabel locali s -12957 70222 -12432 70256 4 VSS
port 42 nsew
rlabel locali s -12957 70256 -12726 70262 4 VSS
port 42 nsew
rlabel locali s -10787 70383 -10545 70417 4 VSS
port 42 nsew
rlabel locali s -12957 70262 -12844 70411 4 VSS
port 42 nsew
rlabel locali s -10631 70417 -10545 70487 4 VSS
port 42 nsew
rlabel locali s -12957 70411 -12725 70418 4 VSS
port 42 nsew
rlabel locali s -12957 70418 -12432 70452 4 VSS
port 42 nsew
rlabel locali s -12957 70452 -12725 70458 4 VSS
port 42 nsew
rlabel locali s -10631 70487 -10077 70548 4 VSS
port 42 nsew
rlabel locali s -9504 70661 -9262 70668 4 VSS
port 42 nsew
rlabel locali s -9504 70668 -8979 70702 4 VSS
port 42 nsew
rlabel locali s -9504 70702 -9262 70708 4 VSS
port 42 nsew
rlabel locali s -9504 70708 -9391 71585 4 VSS
port 42 nsew
rlabel locali s -10631 70548 -10545 70579 4 VSS
port 42 nsew
rlabel locali s -10787 70579 -10545 70613 4 VSS
port 42 nsew
rlabel locali s -10631 70613 -10545 71028 4 VSS
port 42 nsew
rlabel locali s -12957 70458 -12844 70653 4 VSS
port 42 nsew
rlabel locali s -12957 70653 -12715 70660 4 VSS
port 42 nsew
rlabel locali s -12957 70660 -12432 70694 4 VSS
port 42 nsew
rlabel locali s -12957 70694 -12715 70700 4 VSS
port 42 nsew
rlabel locali s -12957 70700 -12844 70965 4 VSS
port 42 nsew
rlabel locali s -9504 71585 -9323 71698 4 VSS
port 42 nsew
rlabel locali s -9436 71698 -9323 72046 4 VSS
port 42 nsew
rlabel locali s -9488 72046 -9323 72122 4 VSS
port 42 nsew
rlabel locali s -9488 72122 -9212 72124 4 VSS
port 42 nsew
rlabel locali s -9488 72124 -8921 72158 4 VSS
port 42 nsew
rlabel locali s -9488 72158 -9212 72159 4 VSS
port 42 nsew
rlabel locali s -9488 72159 -9323 72196 4 VSS
port 42 nsew
rlabel locali s -9488 72196 -9327 72914 4 VSS
port 42 nsew
rlabel locali s -9488 72914 -9212 72915 4 VSS
port 42 nsew
rlabel locali s -9488 72915 -8721 72949 4 VSS
port 42 nsew
rlabel locali s -9488 72949 -9212 72951 4 VSS
port 42 nsew
rlabel locali s -9488 72951 -9327 73042 4 VSS
port 42 nsew
rlabel locali s -9488 73042 -9211 73045 4 VSS
port 42 nsew
rlabel locali s -9488 73045 -8721 73079 4 VSS
port 42 nsew
rlabel locali s -9488 73079 -9327 73369 4 VSS
port 42 nsew
rlabel locali s -10333 72329 -10247 72469 4 VSS
port 42 nsew
rlabel locali s -12598 72325 -12537 72442 4 VSS
port 42 nsew
rlabel locali s -12598 72442 -12485 72443 4 VSS
port 42 nsew
rlabel locali s -10589 72469 -10247 72503 4 VSS
port 42 nsew
rlabel locali s -12598 72443 -12177 72477 4 VSS
port 42 nsew
rlabel locali s -10333 72503 -10247 72665 4 VSS
port 42 nsew
rlabel locali s -10589 72665 -10247 72699 4 VSS
port 42 nsew
rlabel locali s -10333 72699 -10247 73181 4 VSS
port 42 nsew
rlabel locali s -12598 72477 -12537 72767 4 VSS
port 42 nsew
rlabel locali s -12598 72767 -12519 72774 4 VSS
port 42 nsew
rlabel locali s -12112 72912 -12026 73052 4 VSS
port 42 nsew
rlabel locali s -12112 73052 -11870 73086 4 VSS
port 42 nsew
rlabel locali s -9488 73369 -9210 73371 4 VSS
port 42 nsew
rlabel locali s -9488 73371 -8921 73405 4 VSS
port 42 nsew
rlabel locali s -9488 73405 -9210 73406 4 VSS
port 42 nsew
rlabel locali s -9488 73406 -9327 73519 4 VSS
port 42 nsew
rlabel locali s -10333 73181 -10080 73267 4 VSS
port 42 nsew
rlabel locali s -12112 73086 -12026 73156 4 VSS
port 42 nsew
rlabel locali s -12580 72774 -12519 73156 4 VSS
port 42 nsew
rlabel locali s -12988 73156 -12026 73217 4 VSS
port 42 nsew
rlabel locali s -12112 73217 -12026 73248 4 VSS
port 42 nsew
rlabel locali s -10166 73267 -10080 73441 4 VSS
port 42 nsew
rlabel locali s -12112 73248 -11870 73282 4 VSS
port 42 nsew
rlabel locali s -10203 73441 -10080 73442 4 VSS
port 42 nsew
rlabel locali s -10511 73442 -10080 73476 4 VSS
port 42 nsew
rlabel locali s -10166 73476 -10080 73766 4 VSS
port 42 nsew
rlabel locali s -12112 73282 -12026 73527 4 VSS
port 42 nsew
rlabel locali s -10169 73766 -10080 73846 4 VSS
port 42 nsew
rlabel locali s -10169 73846 -10108 74155 4 VSS
port 42 nsew
rlabel locali s -12988 73217 -12875 73883 4 VSS
port 42 nsew
rlabel locali s -12988 73883 -12757 73890 4 VSS
port 42 nsew
rlabel locali s -10662 73911 -10576 74051 4 VSS
port 42 nsew
rlabel locali s -12988 73890 -12463 73924 4 VSS
port 42 nsew
rlabel locali s -12988 73924 -12757 73930 4 VSS
port 42 nsew
rlabel locali s -10818 74051 -10576 74085 4 VSS
port 42 nsew
rlabel locali s -12988 73930 -12875 74079 4 VSS
port 42 nsew
rlabel locali s -10662 74085 -10576 74155 4 VSS
port 42 nsew
rlabel locali s -12988 74079 -12756 74086 4 VSS
port 42 nsew
rlabel locali s -12988 74086 -12463 74120 4 VSS
port 42 nsew
rlabel locali s -12988 74120 -12756 74126 4 VSS
port 42 nsew
rlabel locali s -10662 74155 -10108 74216 4 VSS
port 42 nsew
rlabel locali s -10662 74216 -10576 74247 4 VSS
port 42 nsew
rlabel locali s -10818 74247 -10576 74281 4 VSS
port 42 nsew
rlabel locali s -10662 74281 -10576 74696 4 VSS
port 42 nsew
rlabel locali s -12988 74126 -12875 74321 4 VSS
port 42 nsew
rlabel locali s -12988 74321 -12746 74328 4 VSS
port 42 nsew
rlabel locali s -12988 74328 -12463 74362 4 VSS
port 42 nsew
rlabel locali s -12988 74362 -12746 74368 4 VSS
port 42 nsew
rlabel locali s -12988 74368 -12875 74633 4 VSS
port 42 nsew
rlabel locali s -6888 77532 -6802 77672 4 VSS
port 42 nsew
rlabel locali s -9153 77528 -9092 77645 4 VSS
port 42 nsew
rlabel locali s -9153 77645 -9040 77646 4 VSS
port 42 nsew
rlabel locali s -7144 77672 -6802 77706 4 VSS
port 42 nsew
rlabel locali s -9153 77646 -8732 77680 4 VSS
port 42 nsew
rlabel locali s -6888 77706 -6802 77868 4 VSS
port 42 nsew
rlabel locali s -7144 77868 -6802 77902 4 VSS
port 42 nsew
rlabel locali s -6888 77902 -6802 78384 4 VSS
port 42 nsew
rlabel locali s -9153 77680 -9092 77970 4 VSS
port 42 nsew
rlabel locali s -9153 77970 -9074 77977 4 VSS
port 42 nsew
rlabel locali s -10341 77524 -10255 77664 4 VSS
port 42 nsew
rlabel locali s -12606 77520 -12545 77637 4 VSS
port 42 nsew
rlabel locali s -12606 77637 -12493 77638 4 VSS
port 42 nsew
rlabel locali s -10597 77664 -10255 77698 4 VSS
port 42 nsew
rlabel locali s -12606 77638 -12185 77672 4 VSS
port 42 nsew
rlabel locali s -10341 77698 -10255 77860 4 VSS
port 42 nsew
rlabel locali s -10597 77860 -10255 77894 4 VSS
port 42 nsew
rlabel locali s -8667 78115 -8581 78255 4 VSS
port 42 nsew
rlabel locali s -8667 78255 -8425 78289 4 VSS
port 42 nsew
rlabel locali s -6888 78384 -6635 78470 4 VSS
port 42 nsew
rlabel locali s -8667 78289 -8581 78359 4 VSS
port 42 nsew
rlabel locali s -9135 77977 -9074 78359 4 VSS
port 42 nsew
rlabel locali s -9543 78359 -8581 78420 4 VSS
port 42 nsew
rlabel locali s -10341 77894 -10255 78376 4 VSS
port 42 nsew
rlabel locali s -12606 77672 -12545 77962 4 VSS
port 42 nsew
rlabel locali s -12606 77962 -12527 77969 4 VSS
port 42 nsew
rlabel locali s -12120 78107 -12034 78247 4 VSS
port 42 nsew
rlabel locali s -12120 78247 -11878 78281 4 VSS
port 42 nsew
rlabel locali s -8667 78420 -8581 78451 4 VSS
port 42 nsew
rlabel locali s -6721 78470 -6635 78636 4 VSS
port 42 nsew
rlabel locali s -8667 78451 -8425 78485 4 VSS
port 42 nsew
rlabel locali s -6721 78636 -5618 78644 4 VSS
port 42 nsew
rlabel locali s -6758 78644 -5618 78645 4 VSS
port 42 nsew
rlabel locali s -7066 78645 -5618 78679 4 VSS
port 42 nsew
rlabel locali s -6721 78679 -5618 78919 4 VSS
port 42 nsew
rlabel locali s -8667 78485 -8581 78730 4 VSS
port 42 nsew
rlabel locali s -6124 78919 -5618 87855 4 VSS
port 42 nsew
rlabel locali s -6721 78919 -6635 78969 4 VSS
port 42 nsew
rlabel locali s -6724 78969 -6635 79049 4 VSS
port 42 nsew
rlabel locali s -6724 79049 -6663 79358 4 VSS
port 42 nsew
rlabel locali s -9543 78420 -9430 79086 4 VSS
port 42 nsew
rlabel locali s -10341 78376 -10088 78462 4 VSS
port 42 nsew
rlabel locali s -12120 78281 -12034 78351 4 VSS
port 42 nsew
rlabel locali s -12588 77969 -12527 78351 4 VSS
port 42 nsew
rlabel locali s -12996 78351 -12034 78412 4 VSS
port 42 nsew
rlabel locali s -12120 78412 -12034 78443 4 VSS
port 42 nsew
rlabel locali s -10174 78462 -10088 78636 4 VSS
port 42 nsew
rlabel locali s -12120 78443 -11878 78477 4 VSS
port 42 nsew
rlabel locali s -10211 78636 -10088 78637 4 VSS
port 42 nsew
rlabel locali s -10519 78637 -10088 78671 4 VSS
port 42 nsew
rlabel locali s -10174 78671 -10088 78961 4 VSS
port 42 nsew
rlabel locali s -12120 78477 -12034 78722 4 VSS
port 42 nsew
rlabel locali s -10177 78961 -10088 79041 4 VSS
port 42 nsew
rlabel locali s -9543 79086 -9312 79093 4 VSS
port 42 nsew
rlabel locali s -7217 79114 -7131 79254 4 VSS
port 42 nsew
rlabel locali s -9543 79093 -9018 79127 4 VSS
port 42 nsew
rlabel locali s -9543 79127 -9312 79133 4 VSS
port 42 nsew
rlabel locali s -7373 79254 -7131 79288 4 VSS
port 42 nsew
rlabel locali s -9543 79133 -9430 79282 4 VSS
port 42 nsew
rlabel locali s -7217 79288 -7131 79358 4 VSS
port 42 nsew
rlabel locali s -9543 79282 -9311 79289 4 VSS
port 42 nsew
rlabel locali s -9543 79289 -9018 79323 4 VSS
port 42 nsew
rlabel locali s -9543 79323 -9311 79329 4 VSS
port 42 nsew
rlabel locali s -7217 79358 -6663 79419 4 VSS
port 42 nsew
rlabel locali s -7217 79419 -7131 79450 4 VSS
port 42 nsew
rlabel locali s -7373 79450 -7131 79484 4 VSS
port 42 nsew
rlabel locali s -7217 79484 -7131 79899 4 VSS
port 42 nsew
rlabel locali s -9543 79329 -9430 79524 4 VSS
port 42 nsew
rlabel locali s -10177 79041 -10116 79350 4 VSS
port 42 nsew
rlabel locali s -12996 78412 -12883 79078 4 VSS
port 42 nsew
rlabel locali s -12996 79078 -12765 79085 4 VSS
port 42 nsew
rlabel locali s -10670 79106 -10584 79246 4 VSS
port 42 nsew
rlabel locali s -12996 79085 -12471 79119 4 VSS
port 42 nsew
rlabel locali s -12996 79119 -12765 79125 4 VSS
port 42 nsew
rlabel locali s -10826 79246 -10584 79280 4 VSS
port 42 nsew
rlabel locali s -12996 79125 -12883 79274 4 VSS
port 42 nsew
rlabel locali s -10670 79280 -10584 79350 4 VSS
port 42 nsew
rlabel locali s -12996 79274 -12764 79281 4 VSS
port 42 nsew
rlabel locali s -12996 79281 -12471 79315 4 VSS
port 42 nsew
rlabel locali s -12996 79315 -12764 79321 4 VSS
port 42 nsew
rlabel locali s -10670 79350 -10116 79411 4 VSS
port 42 nsew
rlabel locali s -9543 79524 -9301 79531 4 VSS
port 42 nsew
rlabel locali s -9543 79531 -9018 79565 4 VSS
port 42 nsew
rlabel locali s -9543 79565 -9301 79571 4 VSS
port 42 nsew
rlabel locali s -9543 79571 -9430 80448 4 VSS
port 42 nsew
rlabel locali s -10670 79411 -10584 79442 4 VSS
port 42 nsew
rlabel locali s -10826 79442 -10584 79476 4 VSS
port 42 nsew
rlabel locali s -10670 79476 -10584 79891 4 VSS
port 42 nsew
rlabel locali s -12996 79321 -12883 79516 4 VSS
port 42 nsew
rlabel locali s -12996 79516 -12754 79523 4 VSS
port 42 nsew
rlabel locali s -12996 79523 -12471 79557 4 VSS
port 42 nsew
rlabel locali s -12996 79557 -12754 79563 4 VSS
port 42 nsew
rlabel locali s -12996 79563 -12883 79828 4 VSS
port 42 nsew
rlabel locali s -9543 80448 -9362 80561 4 VSS
port 42 nsew
rlabel locali s -9475 80561 -9362 80909 4 VSS
port 42 nsew
rlabel locali s -9527 80909 -9362 80985 4 VSS
port 42 nsew
rlabel locali s -9527 80985 -9251 80987 4 VSS
port 42 nsew
rlabel locali s -9527 80987 -8960 81021 4 VSS
port 42 nsew
rlabel locali s -9527 81021 -9251 81022 4 VSS
port 42 nsew
rlabel locali s -9527 81022 -9362 81059 4 VSS
port 42 nsew
rlabel locali s -9527 81059 -9366 81777 4 VSS
port 42 nsew
rlabel locali s -9527 81777 -9251 81778 4 VSS
port 42 nsew
rlabel locali s -9527 81778 -8760 81812 4 VSS
port 42 nsew
rlabel locali s -9527 81812 -9251 81814 4 VSS
port 42 nsew
rlabel locali s -9527 81814 -9366 81905 4 VSS
port 42 nsew
rlabel locali s -9527 81905 -9250 81908 4 VSS
port 42 nsew
rlabel locali s -9527 81908 -8760 81942 4 VSS
port 42 nsew
rlabel locali s -9527 81942 -9366 82232 4 VSS
port 42 nsew
rlabel locali s -10372 81192 -10286 81332 4 VSS
port 42 nsew
rlabel locali s -12637 81188 -12576 81305 4 VSS
port 42 nsew
rlabel locali s -12637 81305 -12524 81306 4 VSS
port 42 nsew
rlabel locali s -10628 81332 -10286 81366 4 VSS
port 42 nsew
rlabel locali s -12637 81306 -12216 81340 4 VSS
port 42 nsew
rlabel locali s -10372 81366 -10286 81528 4 VSS
port 42 nsew
rlabel locali s -10628 81528 -10286 81562 4 VSS
port 42 nsew
rlabel locali s -10372 81562 -10286 82044 4 VSS
port 42 nsew
rlabel locali s -12637 81340 -12576 81630 4 VSS
port 42 nsew
rlabel locali s -12637 81630 -12558 81637 4 VSS
port 42 nsew
rlabel locali s -12151 81775 -12065 81915 4 VSS
port 42 nsew
rlabel locali s -12151 81915 -11909 81949 4 VSS
port 42 nsew
rlabel locali s -9527 82232 -9249 82234 4 VSS
port 42 nsew
rlabel locali s -9527 82234 -8960 82268 4 VSS
port 42 nsew
rlabel locali s -9527 82268 -9249 82269 4 VSS
port 42 nsew
rlabel locali s -9527 82269 -9366 82382 4 VSS
port 42 nsew
rlabel locali s -10372 82044 -10119 82130 4 VSS
port 42 nsew
rlabel locali s -12151 81949 -12065 82019 4 VSS
port 42 nsew
rlabel locali s -12619 81637 -12558 82019 4 VSS
port 42 nsew
rlabel locali s -13027 82019 -12065 82080 4 VSS
port 42 nsew
rlabel locali s -12151 82080 -12065 82111 4 VSS
port 42 nsew
rlabel locali s -10205 82130 -10119 82304 4 VSS
port 42 nsew
rlabel locali s -12151 82111 -11909 82145 4 VSS
port 42 nsew
rlabel locali s -10242 82304 -10119 82305 4 VSS
port 42 nsew
rlabel locali s -10550 82305 -10119 82339 4 VSS
port 42 nsew
rlabel locali s -10205 82339 -10119 82629 4 VSS
port 42 nsew
rlabel locali s -12151 82145 -12065 82390 4 VSS
port 42 nsew
rlabel locali s -10208 82629 -10119 82709 4 VSS
port 42 nsew
rlabel locali s -10208 82709 -10147 83018 4 VSS
port 42 nsew
rlabel locali s -13027 82080 -12914 82746 4 VSS
port 42 nsew
rlabel locali s -13027 82746 -12796 82753 4 VSS
port 42 nsew
rlabel locali s -10701 82774 -10615 82914 4 VSS
port 42 nsew
rlabel locali s -13027 82753 -12502 82787 4 VSS
port 42 nsew
rlabel locali s -13027 82787 -12796 82793 4 VSS
port 42 nsew
rlabel locali s -10857 82914 -10615 82948 4 VSS
port 42 nsew
rlabel locali s -13027 82793 -12914 82942 4 VSS
port 42 nsew
rlabel locali s -10701 82948 -10615 83018 4 VSS
port 42 nsew
rlabel locali s -13027 82942 -12795 82949 4 VSS
port 42 nsew
rlabel locali s -13027 82949 -12502 82983 4 VSS
port 42 nsew
rlabel locali s -13027 82983 -12795 82989 4 VSS
port 42 nsew
rlabel locali s -10701 83018 -10147 83079 4 VSS
port 42 nsew
rlabel locali s -10701 83079 -10615 83110 4 VSS
port 42 nsew
rlabel locali s -10857 83110 -10615 83144 4 VSS
port 42 nsew
rlabel locali s -10701 83144 -10615 83559 4 VSS
port 42 nsew
rlabel locali s -13027 82989 -12914 83184 4 VSS
port 42 nsew
rlabel locali s -13027 83184 -12785 83191 4 VSS
port 42 nsew
rlabel locali s -13027 83191 -12502 83225 4 VSS
port 42 nsew
rlabel locali s -13027 83225 -12785 83231 4 VSS
port 42 nsew
rlabel locali s -13027 83231 -12914 83496 4 VSS
port 42 nsew
rlabel locali s -6854 86730 -6768 86870 4 VSS
port 42 nsew
rlabel locali s -9119 86726 -9058 86843 4 VSS
port 42 nsew
rlabel locali s -9119 86843 -9006 86844 4 VSS
port 42 nsew
rlabel locali s -7110 86870 -6768 86904 4 VSS
port 42 nsew
rlabel locali s -9119 86844 -8698 86878 4 VSS
port 42 nsew
rlabel locali s -6854 86904 -6768 87066 4 VSS
port 42 nsew
rlabel locali s -7110 87066 -6768 87100 4 VSS
port 42 nsew
rlabel locali s -6854 87100 -6768 87582 4 VSS
port 42 nsew
rlabel locali s -9119 86878 -9058 87168 4 VSS
port 42 nsew
rlabel locali s -9119 87168 -9040 87175 4 VSS
port 42 nsew
rlabel locali s -10307 86722 -10221 86862 4 VSS
port 42 nsew
rlabel locali s -12572 86718 -12511 86835 4 VSS
port 42 nsew
rlabel locali s -12572 86835 -12459 86836 4 VSS
port 42 nsew
rlabel locali s -10563 86862 -10221 86896 4 VSS
port 42 nsew
rlabel locali s -12572 86836 -12151 86870 4 VSS
port 42 nsew
rlabel locali s -10307 86896 -10221 87058 4 VSS
port 42 nsew
rlabel locali s -10563 87058 -10221 87092 4 VSS
port 42 nsew
rlabel locali s -8633 87313 -8547 87453 4 VSS
port 42 nsew
rlabel locali s -8633 87453 -8391 87487 4 VSS
port 42 nsew
rlabel locali s -6854 87582 -6601 87668 4 VSS
port 42 nsew
rlabel locali s -8633 87487 -8547 87557 4 VSS
port 42 nsew
rlabel locali s -9101 87175 -9040 87557 4 VSS
port 42 nsew
rlabel locali s -9509 87557 -8547 87618 4 VSS
port 42 nsew
rlabel locali s -10307 87092 -10221 87574 4 VSS
port 42 nsew
rlabel locali s -12572 86870 -12511 87160 4 VSS
port 42 nsew
rlabel locali s -12572 87160 -12493 87167 4 VSS
port 42 nsew
rlabel locali s -12086 87305 -12000 87445 4 VSS
port 42 nsew
rlabel locali s -12086 87445 -11844 87479 4 VSS
port 42 nsew
rlabel locali s -8633 87618 -8547 87649 4 VSS
port 42 nsew
rlabel locali s -6687 87668 -6601 87842 4 VSS
port 42 nsew
rlabel locali s -8633 87649 -8391 87683 4 VSS
port 42 nsew
rlabel locali s -6724 87842 -6601 87843 4 VSS
port 42 nsew
rlabel locali s -7032 87843 -6601 87855 4 VSS
port 42 nsew
rlabel locali s -7032 87855 -5618 87877 4 VSS
port 42 nsew
rlabel locali s -6687 87877 -5618 88138 4 VSS
port 42 nsew
rlabel locali s -8633 87683 -8547 87928 4 VSS
port 42 nsew
rlabel locali s -6124 88138 -5618 96650 4 VSS
port 42 nsew
rlabel locali s -6687 88138 -6601 88167 4 VSS
port 42 nsew
rlabel locali s -6690 88167 -6601 88247 4 VSS
port 42 nsew
rlabel locali s -6690 88247 -6629 88556 4 VSS
port 42 nsew
rlabel locali s -9509 87618 -9396 88284 4 VSS
port 42 nsew
rlabel locali s -10307 87574 -10054 87660 4 VSS
port 42 nsew
rlabel locali s -12086 87479 -12000 87549 4 VSS
port 42 nsew
rlabel locali s -12554 87167 -12493 87549 4 VSS
port 42 nsew
rlabel locali s -12962 87549 -12000 87610 4 VSS
port 42 nsew
rlabel locali s -12086 87610 -12000 87641 4 VSS
port 42 nsew
rlabel locali s -10140 87660 -10054 87834 4 VSS
port 42 nsew
rlabel locali s -12086 87641 -11844 87675 4 VSS
port 42 nsew
rlabel locali s -10177 87834 -10054 87835 4 VSS
port 42 nsew
rlabel locali s -10485 87835 -10054 87869 4 VSS
port 42 nsew
rlabel locali s -10140 87869 -10054 88159 4 VSS
port 42 nsew
rlabel locali s -12086 87675 -12000 87920 4 VSS
port 42 nsew
rlabel locali s -10143 88159 -10054 88239 4 VSS
port 42 nsew
rlabel locali s -9509 88284 -9278 88291 4 VSS
port 42 nsew
rlabel locali s -7183 88312 -7097 88452 4 VSS
port 42 nsew
rlabel locali s -9509 88291 -8984 88325 4 VSS
port 42 nsew
rlabel locali s -9509 88325 -9278 88331 4 VSS
port 42 nsew
rlabel locali s -7339 88452 -7097 88486 4 VSS
port 42 nsew
rlabel locali s -9509 88331 -9396 88480 4 VSS
port 42 nsew
rlabel locali s -7183 88486 -7097 88556 4 VSS
port 42 nsew
rlabel locali s -9509 88480 -9277 88487 4 VSS
port 42 nsew
rlabel locali s -9509 88487 -8984 88521 4 VSS
port 42 nsew
rlabel locali s -9509 88521 -9277 88527 4 VSS
port 42 nsew
rlabel locali s -7183 88556 -6629 88617 4 VSS
port 42 nsew
rlabel locali s -7183 88617 -7097 88648 4 VSS
port 42 nsew
rlabel locali s -7339 88648 -7097 88682 4 VSS
port 42 nsew
rlabel locali s -7183 88682 -7097 89097 4 VSS
port 42 nsew
rlabel locali s -9509 88527 -9396 88722 4 VSS
port 42 nsew
rlabel locali s -10143 88239 -10082 88548 4 VSS
port 42 nsew
rlabel locali s -12962 87610 -12849 88276 4 VSS
port 42 nsew
rlabel locali s -12962 88276 -12731 88283 4 VSS
port 42 nsew
rlabel locali s -10636 88304 -10550 88444 4 VSS
port 42 nsew
rlabel locali s -12962 88283 -12437 88317 4 VSS
port 42 nsew
rlabel locali s -12962 88317 -12731 88323 4 VSS
port 42 nsew
rlabel locali s -10792 88444 -10550 88478 4 VSS
port 42 nsew
rlabel locali s -12962 88323 -12849 88472 4 VSS
port 42 nsew
rlabel locali s -10636 88478 -10550 88548 4 VSS
port 42 nsew
rlabel locali s -12962 88472 -12730 88479 4 VSS
port 42 nsew
rlabel locali s -12962 88479 -12437 88513 4 VSS
port 42 nsew
rlabel locali s -12962 88513 -12730 88519 4 VSS
port 42 nsew
rlabel locali s -10636 88548 -10082 88609 4 VSS
port 42 nsew
rlabel locali s -9509 88722 -9267 88729 4 VSS
port 42 nsew
rlabel locali s -9509 88729 -8984 88763 4 VSS
port 42 nsew
rlabel locali s -9509 88763 -9267 88769 4 VSS
port 42 nsew
rlabel locali s -9509 88769 -9396 89646 4 VSS
port 42 nsew
rlabel locali s -10636 88609 -10550 88640 4 VSS
port 42 nsew
rlabel locali s -10792 88640 -10550 88674 4 VSS
port 42 nsew
rlabel locali s -10636 88674 -10550 89089 4 VSS
port 42 nsew
rlabel locali s -12962 88519 -12849 88714 4 VSS
port 42 nsew
rlabel locali s -12962 88714 -12720 88721 4 VSS
port 42 nsew
rlabel locali s -12962 88721 -12437 88755 4 VSS
port 42 nsew
rlabel locali s -12962 88755 -12720 88761 4 VSS
port 42 nsew
rlabel locali s -12962 88761 -12849 89026 4 VSS
port 42 nsew
rlabel locali s -9509 89646 -9328 89759 4 VSS
port 42 nsew
rlabel locali s -9441 89759 -9328 90107 4 VSS
port 42 nsew
rlabel locali s -9493 90107 -9328 90183 4 VSS
port 42 nsew
rlabel locali s -9493 90183 -9217 90185 4 VSS
port 42 nsew
rlabel locali s -9493 90185 -8926 90219 4 VSS
port 42 nsew
rlabel locali s -9493 90219 -9217 90220 4 VSS
port 42 nsew
rlabel locali s -9493 90220 -9328 90257 4 VSS
port 42 nsew
rlabel locali s -9493 90257 -9332 90975 4 VSS
port 42 nsew
rlabel locali s -9493 90975 -9217 90976 4 VSS
port 42 nsew
rlabel locali s -9493 90976 -8726 91010 4 VSS
port 42 nsew
rlabel locali s -9493 91010 -9217 91012 4 VSS
port 42 nsew
rlabel locali s -9493 91012 -9332 91103 4 VSS
port 42 nsew
rlabel locali s -9493 91103 -9216 91106 4 VSS
port 42 nsew
rlabel locali s -9493 91106 -8726 91140 4 VSS
port 42 nsew
rlabel locali s -9493 91140 -9332 91430 4 VSS
port 42 nsew
rlabel locali s -10338 90390 -10252 90530 4 VSS
port 42 nsew
rlabel locali s -12603 90386 -12542 90503 4 VSS
port 42 nsew
rlabel locali s -12603 90503 -12490 90504 4 VSS
port 42 nsew
rlabel locali s -10594 90530 -10252 90564 4 VSS
port 42 nsew
rlabel locali s -12603 90504 -12182 90538 4 VSS
port 42 nsew
rlabel locali s -10338 90564 -10252 90726 4 VSS
port 42 nsew
rlabel locali s -10594 90726 -10252 90760 4 VSS
port 42 nsew
rlabel locali s -10338 90760 -10252 91242 4 VSS
port 42 nsew
rlabel locali s -12603 90538 -12542 90828 4 VSS
port 42 nsew
rlabel locali s -12603 90828 -12524 90835 4 VSS
port 42 nsew
rlabel locali s -12117 90973 -12031 91113 4 VSS
port 42 nsew
rlabel locali s -12117 91113 -11875 91147 4 VSS
port 42 nsew
rlabel locali s -9493 91430 -9215 91432 4 VSS
port 42 nsew
rlabel locali s -9493 91432 -8926 91466 4 VSS
port 42 nsew
rlabel locali s -9493 91466 -9215 91467 4 VSS
port 42 nsew
rlabel locali s -9493 91467 -9332 91580 4 VSS
port 42 nsew
rlabel locali s -10338 91242 -10085 91328 4 VSS
port 42 nsew
rlabel locali s -12117 91147 -12031 91217 4 VSS
port 42 nsew
rlabel locali s -12585 90835 -12524 91217 4 VSS
port 42 nsew
rlabel locali s -12993 91217 -12031 91278 4 VSS
port 42 nsew
rlabel locali s -12117 91278 -12031 91309 4 VSS
port 42 nsew
rlabel locali s -10171 91328 -10085 91502 4 VSS
port 42 nsew
rlabel locali s -12117 91309 -11875 91343 4 VSS
port 42 nsew
rlabel locali s -10208 91502 -10085 91503 4 VSS
port 42 nsew
rlabel locali s -10516 91503 -10085 91537 4 VSS
port 42 nsew
rlabel locali s -10171 91537 -10085 91827 4 VSS
port 42 nsew
rlabel locali s -12117 91343 -12031 91588 4 VSS
port 42 nsew
rlabel locali s -10174 91827 -10085 91907 4 VSS
port 42 nsew
rlabel locali s -10174 91907 -10113 92216 4 VSS
port 42 nsew
rlabel locali s -12993 91278 -12880 91944 4 VSS
port 42 nsew
rlabel locali s -12993 91944 -12762 91951 4 VSS
port 42 nsew
rlabel locali s -10667 91972 -10581 92112 4 VSS
port 42 nsew
rlabel locali s -12993 91951 -12468 91985 4 VSS
port 42 nsew
rlabel locali s -12993 91985 -12762 91991 4 VSS
port 42 nsew
rlabel locali s -10823 92112 -10581 92146 4 VSS
port 42 nsew
rlabel locali s -12993 91991 -12880 92140 4 VSS
port 42 nsew
rlabel locali s -10667 92146 -10581 92216 4 VSS
port 42 nsew
rlabel locali s -12993 92140 -12761 92147 4 VSS
port 42 nsew
rlabel locali s -12993 92147 -12468 92181 4 VSS
port 42 nsew
rlabel locali s -12993 92181 -12761 92187 4 VSS
port 42 nsew
rlabel locali s -10667 92216 -10113 92277 4 VSS
port 42 nsew
rlabel locali s -10667 92277 -10581 92308 4 VSS
port 42 nsew
rlabel locali s -10823 92308 -10581 92342 4 VSS
port 42 nsew
rlabel locali s -10667 92342 -10581 92757 4 VSS
port 42 nsew
rlabel locali s -12993 92187 -12880 92382 4 VSS
port 42 nsew
rlabel locali s -12993 92382 -12751 92389 4 VSS
port 42 nsew
rlabel locali s -12993 92389 -12468 92423 4 VSS
port 42 nsew
rlabel locali s -12993 92423 -12751 92429 4 VSS
port 42 nsew
rlabel locali s -12993 92429 -12880 92694 4 VSS
port 42 nsew
rlabel locali s -11943 94859 -11907 95042 4 VSS
port 42 nsew
rlabel locali s -15491 41738 -15355 95042 4 VSS
port 42 nsew
rlabel locali s -15491 95042 -11907 95178 4 VSS
port 42 nsew
rlabel locali s -11943 95178 -11907 95387 4 VSS
port 42 nsew
rlabel locali s -11945 95387 -11905 95407 4 VSS
port 42 nsew
rlabel locali s -6788 95484 -6702 95624 4 VSS
port 42 nsew
rlabel locali s -9053 95480 -8992 95597 4 VSS
port 42 nsew
rlabel locali s -9053 95597 -8940 95598 4 VSS
port 42 nsew
rlabel locali s -7044 95624 -6702 95658 4 VSS
port 42 nsew
rlabel locali s -9053 95598 -8632 95632 4 VSS
port 42 nsew
rlabel locali s -6788 95658 -6702 95820 4 VSS
port 42 nsew
rlabel locali s -7044 95820 -6702 95854 4 VSS
port 42 nsew
rlabel locali s -6788 95854 -6702 96336 4 VSS
port 42 nsew
rlabel locali s -9053 95632 -8992 95922 4 VSS
port 42 nsew
rlabel locali s -9053 95922 -8974 95929 4 VSS
port 42 nsew
rlabel locali s -10241 95476 -10155 95616 4 VSS
port 42 nsew
rlabel locali s -11953 95407 -11899 95542 4 VSS
port 42 nsew
rlabel locali s -12506 95472 -12445 95589 4 VSS
port 42 nsew
rlabel locali s -12506 95589 -12393 95590 4 VSS
port 42 nsew
rlabel locali s -10497 95616 -10155 95650 4 VSS
port 42 nsew
rlabel locali s -12506 95590 -12085 95624 4 VSS
port 42 nsew
rlabel locali s -10241 95650 -10155 95812 4 VSS
port 42 nsew
rlabel locali s -10497 95812 -10155 95846 4 VSS
port 42 nsew
rlabel locali s -8567 96067 -8481 96207 4 VSS
port 42 nsew
rlabel locali s -8567 96207 -8325 96241 4 VSS
port 42 nsew
rlabel locali s -6788 96336 -6535 96422 4 VSS
port 42 nsew
rlabel locali s -8567 96241 -8481 96311 4 VSS
port 42 nsew
rlabel locali s -9035 95929 -8974 96311 4 VSS
port 42 nsew
rlabel locali s -9443 96311 -8481 96372 4 VSS
port 42 nsew
rlabel locali s -10241 95846 -10155 96328 4 VSS
port 42 nsew
rlabel locali s -12506 95624 -12445 95914 4 VSS
port 42 nsew
rlabel locali s -12506 95914 -12427 95921 4 VSS
port 42 nsew
rlabel locali s -12020 96059 -11934 96199 4 VSS
port 42 nsew
rlabel locali s -12020 96199 -11778 96233 4 VSS
port 42 nsew
rlabel locali s -8567 96372 -8481 96403 4 VSS
port 42 nsew
rlabel locali s -6621 96422 -6535 96596 4 VSS
port 42 nsew
rlabel locali s -8567 96403 -8325 96437 4 VSS
port 42 nsew
rlabel locali s -6658 96596 -6535 96597 4 VSS
port 42 nsew
rlabel locali s -6966 96597 -6535 96631 4 VSS
port 42 nsew
rlabel locali s -6621 96631 -6535 96650 4 VSS
port 42 nsew
rlabel locali s -6621 96650 -5618 96921 4 VSS
port 42 nsew
rlabel locali s -8567 96437 -8481 96682 4 VSS
port 42 nsew
rlabel locali s -6624 96921 -5618 96957 4 VSS
port 42 nsew
rlabel locali s -6124 96957 -5618 105756 4 VSS
port 42 nsew
rlabel locali s -6624 96957 -6535 97001 4 VSS
port 42 nsew
rlabel locali s -6624 97001 -6563 97310 4 VSS
port 42 nsew
rlabel locali s -9443 96372 -9330 97038 4 VSS
port 42 nsew
rlabel locali s -10241 96328 -9988 96414 4 VSS
port 42 nsew
rlabel locali s -12020 96233 -11934 96303 4 VSS
port 42 nsew
rlabel locali s -12488 95921 -12427 96303 4 VSS
port 42 nsew
rlabel locali s -12896 96303 -11934 96364 4 VSS
port 42 nsew
rlabel locali s -12020 96364 -11934 96395 4 VSS
port 42 nsew
rlabel locali s -10074 96414 -9988 96588 4 VSS
port 42 nsew
rlabel locali s -12020 96395 -11778 96429 4 VSS
port 42 nsew
rlabel locali s -10111 96588 -9988 96589 4 VSS
port 42 nsew
rlabel locali s -10419 96589 -9988 96623 4 VSS
port 42 nsew
rlabel locali s -10074 96623 -9988 96913 4 VSS
port 42 nsew
rlabel locali s -12020 96429 -11934 96674 4 VSS
port 42 nsew
rlabel locali s -10077 96913 -9988 96993 4 VSS
port 42 nsew
rlabel locali s -9443 97038 -9212 97045 4 VSS
port 42 nsew
rlabel locali s -7117 97066 -7031 97206 4 VSS
port 42 nsew
rlabel locali s -9443 97045 -8918 97079 4 VSS
port 42 nsew
rlabel locali s -9443 97079 -9212 97085 4 VSS
port 42 nsew
rlabel locali s -7273 97206 -7031 97240 4 VSS
port 42 nsew
rlabel locali s -9443 97085 -9330 97234 4 VSS
port 42 nsew
rlabel locali s -7117 97240 -7031 97310 4 VSS
port 42 nsew
rlabel locali s -9443 97234 -9211 97241 4 VSS
port 42 nsew
rlabel locali s -9443 97241 -8918 97275 4 VSS
port 42 nsew
rlabel locali s -9443 97275 -9211 97281 4 VSS
port 42 nsew
rlabel locali s -7117 97310 -6563 97371 4 VSS
port 42 nsew
rlabel locali s -7117 97371 -7031 97402 4 VSS
port 42 nsew
rlabel locali s -7273 97402 -7031 97436 4 VSS
port 42 nsew
rlabel locali s -7117 97436 -7031 97851 4 VSS
port 42 nsew
rlabel locali s -9443 97281 -9330 97476 4 VSS
port 42 nsew
rlabel locali s -10077 96993 -10016 97302 4 VSS
port 42 nsew
rlabel locali s -12896 96364 -12783 97030 4 VSS
port 42 nsew
rlabel locali s -12896 97030 -12665 97037 4 VSS
port 42 nsew
rlabel locali s -10570 97058 -10484 97198 4 VSS
port 42 nsew
rlabel locali s -12896 97037 -12371 97071 4 VSS
port 42 nsew
rlabel locali s -12896 97071 -12665 97077 4 VSS
port 42 nsew
rlabel locali s -10726 97198 -10484 97232 4 VSS
port 42 nsew
rlabel locali s -12896 97077 -12783 97226 4 VSS
port 42 nsew
rlabel locali s -10570 97232 -10484 97302 4 VSS
port 42 nsew
rlabel locali s -12896 97226 -12664 97233 4 VSS
port 42 nsew
rlabel locali s -12896 97233 -12371 97267 4 VSS
port 42 nsew
rlabel locali s -12896 97267 -12664 97273 4 VSS
port 42 nsew
rlabel locali s -10570 97302 -10016 97363 4 VSS
port 42 nsew
rlabel locali s -9443 97476 -9201 97483 4 VSS
port 42 nsew
rlabel locali s -9443 97483 -8918 97517 4 VSS
port 42 nsew
rlabel locali s -9443 97517 -9201 97523 4 VSS
port 42 nsew
rlabel locali s -9443 97523 -9330 98400 4 VSS
port 42 nsew
rlabel locali s -10570 97363 -10484 97394 4 VSS
port 42 nsew
rlabel locali s -10726 97394 -10484 97428 4 VSS
port 42 nsew
rlabel locali s -10570 97428 -10484 97843 4 VSS
port 42 nsew
rlabel locali s -12896 97273 -12783 97468 4 VSS
port 42 nsew
rlabel locali s -12896 97468 -12654 97475 4 VSS
port 42 nsew
rlabel locali s -12896 97475 -12371 97509 4 VSS
port 42 nsew
rlabel locali s -12896 97509 -12654 97515 4 VSS
port 42 nsew
rlabel locali s -12896 97515 -12783 97780 4 VSS
port 42 nsew
rlabel locali s -9443 98400 -9262 98513 4 VSS
port 42 nsew
rlabel locali s -9375 98513 -9262 98861 4 VSS
port 42 nsew
rlabel locali s -13106 95178 -12970 98641 4 VSS
port 42 nsew
rlabel locali s -13106 98641 -11938 98777 4 VSS
port 42 nsew
rlabel locali s -9427 98861 -9262 98937 4 VSS
port 42 nsew
rlabel locali s -9427 98937 -9151 98939 4 VSS
port 42 nsew
rlabel locali s -9427 98939 -8860 98973 4 VSS
port 42 nsew
rlabel locali s -9427 98973 -9151 98974 4 VSS
port 42 nsew
rlabel locali s -9427 98974 -9262 99011 4 VSS
port 42 nsew
rlabel locali s -9427 99011 -9266 99729 4 VSS
port 42 nsew
rlabel locali s -11974 98777 -11938 99055 4 VSS
port 42 nsew
rlabel locali s -11976 99055 -11936 99075 4 VSS
port 42 nsew
rlabel locali s -9427 99729 -9151 99730 4 VSS
port 42 nsew
rlabel locali s -9427 99730 -8660 99764 4 VSS
port 42 nsew
rlabel locali s -9427 99764 -9151 99766 4 VSS
port 42 nsew
rlabel locali s -9427 99766 -9266 99857 4 VSS
port 42 nsew
rlabel locali s -9427 99857 -9150 99860 4 VSS
port 42 nsew
rlabel locali s -9427 99860 -8660 99894 4 VSS
port 42 nsew
rlabel locali s -9427 99894 -9266 100184 4 VSS
port 42 nsew
rlabel locali s -10272 99144 -10186 99284 4 VSS
port 42 nsew
rlabel locali s -11984 99075 -11930 99210 4 VSS
port 42 nsew
rlabel locali s -12537 99140 -12476 99257 4 VSS
port 42 nsew
rlabel locali s -12537 99257 -12424 99258 4 VSS
port 42 nsew
rlabel locali s -10528 99284 -10186 99318 4 VSS
port 42 nsew
rlabel locali s -12537 99258 -12116 99292 4 VSS
port 42 nsew
rlabel locali s -10272 99318 -10186 99480 4 VSS
port 42 nsew
rlabel locali s -10528 99480 -10186 99514 4 VSS
port 42 nsew
rlabel locali s -10272 99514 -10186 99996 4 VSS
port 42 nsew
rlabel locali s -12537 99292 -12476 99582 4 VSS
port 42 nsew
rlabel locali s -12537 99582 -12458 99589 4 VSS
port 42 nsew
rlabel locali s -12051 99727 -11965 99867 4 VSS
port 42 nsew
rlabel locali s -12051 99867 -11809 99901 4 VSS
port 42 nsew
rlabel locali s -9427 100184 -9149 100186 4 VSS
port 42 nsew
rlabel locali s -9427 100186 -8860 100220 4 VSS
port 42 nsew
rlabel locali s -9427 100220 -9149 100221 4 VSS
port 42 nsew
rlabel locali s -9427 100221 -9266 100334 4 VSS
port 42 nsew
rlabel locali s -10272 99996 -10019 100082 4 VSS
port 42 nsew
rlabel locali s -12051 99901 -11965 99971 4 VSS
port 42 nsew
rlabel locali s -12519 99589 -12458 99971 4 VSS
port 42 nsew
rlabel locali s -12927 99971 -11965 100032 4 VSS
port 42 nsew
rlabel locali s -12051 100032 -11965 100063 4 VSS
port 42 nsew
rlabel locali s -10105 100082 -10019 100256 4 VSS
port 42 nsew
rlabel locali s -12051 100063 -11809 100097 4 VSS
port 42 nsew
rlabel locali s -10142 100256 -10019 100257 4 VSS
port 42 nsew
rlabel locali s -10450 100257 -10019 100291 4 VSS
port 42 nsew
rlabel locali s -10105 100291 -10019 100581 4 VSS
port 42 nsew
rlabel locali s -12051 100097 -11965 100342 4 VSS
port 42 nsew
rlabel locali s -10108 100581 -10019 100661 4 VSS
port 42 nsew
rlabel locali s -10108 100661 -10047 100970 4 VSS
port 42 nsew
rlabel locali s -12927 100032 -12814 100698 4 VSS
port 42 nsew
rlabel locali s -12927 100698 -12696 100705 4 VSS
port 42 nsew
rlabel locali s -10601 100726 -10515 100866 4 VSS
port 42 nsew
rlabel locali s -12927 100705 -12402 100739 4 VSS
port 42 nsew
rlabel locali s -12927 100739 -12696 100745 4 VSS
port 42 nsew
rlabel locali s -10757 100866 -10515 100900 4 VSS
port 42 nsew
rlabel locali s -12927 100745 -12814 100894 4 VSS
port 42 nsew
rlabel locali s -10601 100900 -10515 100970 4 VSS
port 42 nsew
rlabel locali s -12927 100894 -12695 100901 4 VSS
port 42 nsew
rlabel locali s -12927 100901 -12402 100935 4 VSS
port 42 nsew
rlabel locali s -12927 100935 -12695 100941 4 VSS
port 42 nsew
rlabel locali s -10601 100970 -10047 101031 4 VSS
port 42 nsew
rlabel locali s -10601 101031 -10515 101062 4 VSS
port 42 nsew
rlabel locali s -10757 101062 -10515 101096 4 VSS
port 42 nsew
rlabel locali s -10601 101096 -10515 101511 4 VSS
port 42 nsew
rlabel locali s -12927 100941 -12814 101136 4 VSS
port 42 nsew
rlabel locali s -12927 101136 -12685 101143 4 VSS
port 42 nsew
rlabel locali s -12927 101143 -12402 101177 4 VSS
port 42 nsew
rlabel locali s -12927 101177 -12685 101183 4 VSS
port 42 nsew
rlabel locali s -12927 101183 -12814 101448 4 VSS
port 42 nsew
rlabel locali s -11926 104012 -11890 104195 4 VSS
port 42 nsew
rlabel locali s -15790 8555 -15654 104195 4 VSS
port 42 nsew
rlabel locali s -15790 104195 -11890 104331 4 VSS
port 42 nsew
rlabel locali s -11926 104331 -11890 104540 4 VSS
port 42 nsew
rlabel locali s -11928 104540 -11888 104560 4 VSS
port 42 nsew
rlabel locali s -6771 104637 -6685 104777 4 VSS
port 42 nsew
rlabel locali s -9036 104633 -8975 104750 4 VSS
port 42 nsew
rlabel locali s -9036 104750 -8923 104751 4 VSS
port 42 nsew
rlabel locali s -7027 104777 -6685 104811 4 VSS
port 42 nsew
rlabel locali s -9036 104751 -8615 104785 4 VSS
port 42 nsew
rlabel locali s -6771 104811 -6685 104973 4 VSS
port 42 nsew
rlabel locali s -7027 104973 -6685 105007 4 VSS
port 42 nsew
rlabel locali s -6771 105007 -6685 105489 4 VSS
port 42 nsew
rlabel locali s -9036 104785 -8975 105075 4 VSS
port 42 nsew
rlabel locali s -9036 105075 -8957 105082 4 VSS
port 42 nsew
rlabel locali s -10224 104629 -10138 104769 4 VSS
port 42 nsew
rlabel locali s -11936 104560 -11882 104695 4 VSS
port 42 nsew
rlabel locali s -12489 104625 -12428 104742 4 VSS
port 42 nsew
rlabel locali s -12489 104742 -12376 104743 4 VSS
port 42 nsew
rlabel locali s -10480 104769 -10138 104803 4 VSS
port 42 nsew
rlabel locali s -12489 104743 -12068 104777 4 VSS
port 42 nsew
rlabel locali s -10224 104803 -10138 104965 4 VSS
port 42 nsew
rlabel locali s -10480 104965 -10138 104999 4 VSS
port 42 nsew
rlabel locali s -8550 105220 -8464 105360 4 VSS
port 42 nsew
rlabel locali s -8550 105360 -8308 105394 4 VSS
port 42 nsew
rlabel locali s -6771 105489 -6518 105575 4 VSS
port 42 nsew
rlabel locali s -8550 105394 -8464 105464 4 VSS
port 42 nsew
rlabel locali s -9018 105082 -8957 105464 4 VSS
port 42 nsew
rlabel locali s -9426 105464 -8464 105525 4 VSS
port 42 nsew
rlabel locali s -10224 104999 -10138 105481 4 VSS
port 42 nsew
rlabel locali s -12489 104777 -12428 105067 4 VSS
port 42 nsew
rlabel locali s -12489 105067 -12410 105074 4 VSS
port 42 nsew
rlabel locali s -12003 105212 -11917 105352 4 VSS
port 42 nsew
rlabel locali s -12003 105352 -11761 105386 4 VSS
port 42 nsew
rlabel locali s -8550 105525 -8464 105556 4 VSS
port 42 nsew
rlabel locali s -6604 105575 -6518 105749 4 VSS
port 42 nsew
rlabel locali s -8550 105556 -8308 105590 4 VSS
port 42 nsew
rlabel locali s -6641 105749 -6518 105750 4 VSS
port 42 nsew
rlabel locali s -6949 105750 -6518 105756 4 VSS
port 42 nsew
rlabel locali s -6949 105756 -5618 105784 4 VSS
port 42 nsew
rlabel locali s -6604 105784 -5618 106074 4 VSS
port 42 nsew
rlabel locali s -8550 105590 -8464 105835 4 VSS
port 42 nsew
rlabel locali s -6607 106074 -5618 106096 4 VSS
port 42 nsew
rlabel locali s -6124 106096 -5618 115092 4 VSS
port 42 nsew
rlabel locali s -6607 106096 -6518 106154 4 VSS
port 42 nsew
rlabel locali s -6607 106154 -6546 106463 4 VSS
port 42 nsew
rlabel locali s -9426 105525 -9313 106191 4 VSS
port 42 nsew
rlabel locali s -10224 105481 -9971 105567 4 VSS
port 42 nsew
rlabel locali s -12003 105386 -11917 105456 4 VSS
port 42 nsew
rlabel locali s -12471 105074 -12410 105456 4 VSS
port 42 nsew
rlabel locali s -12879 105456 -11917 105517 4 VSS
port 42 nsew
rlabel locali s -12003 105517 -11917 105548 4 VSS
port 42 nsew
rlabel locali s -10057 105567 -9971 105741 4 VSS
port 42 nsew
rlabel locali s -12003 105548 -11761 105582 4 VSS
port 42 nsew
rlabel locali s -10094 105741 -9971 105742 4 VSS
port 42 nsew
rlabel locali s -10402 105742 -9971 105776 4 VSS
port 42 nsew
rlabel locali s -10057 105776 -9971 106066 4 VSS
port 42 nsew
rlabel locali s -12003 105582 -11917 105827 4 VSS
port 42 nsew
rlabel locali s -10060 106066 -9971 106146 4 VSS
port 42 nsew
rlabel locali s -9426 106191 -9195 106198 4 VSS
port 42 nsew
rlabel locali s -7100 106219 -7014 106359 4 VSS
port 42 nsew
rlabel locali s -9426 106198 -8901 106232 4 VSS
port 42 nsew
rlabel locali s -9426 106232 -9195 106238 4 VSS
port 42 nsew
rlabel locali s -7256 106359 -7014 106393 4 VSS
port 42 nsew
rlabel locali s -9426 106238 -9313 106387 4 VSS
port 42 nsew
rlabel locali s -7100 106393 -7014 106463 4 VSS
port 42 nsew
rlabel locali s -9426 106387 -9194 106394 4 VSS
port 42 nsew
rlabel locali s -9426 106394 -8901 106428 4 VSS
port 42 nsew
rlabel locali s -9426 106428 -9194 106434 4 VSS
port 42 nsew
rlabel locali s -7100 106463 -6546 106524 4 VSS
port 42 nsew
rlabel locali s -7100 106524 -7014 106555 4 VSS
port 42 nsew
rlabel locali s -7256 106555 -7014 106589 4 VSS
port 42 nsew
rlabel locali s -7100 106589 -7014 107004 4 VSS
port 42 nsew
rlabel locali s -9426 106434 -9313 106629 4 VSS
port 42 nsew
rlabel locali s -10060 106146 -9999 106455 4 VSS
port 42 nsew
rlabel locali s -12879 105517 -12766 106183 4 VSS
port 42 nsew
rlabel locali s -12879 106183 -12648 106190 4 VSS
port 42 nsew
rlabel locali s -10553 106211 -10467 106351 4 VSS
port 42 nsew
rlabel locali s -12879 106190 -12354 106224 4 VSS
port 42 nsew
rlabel locali s -12879 106224 -12648 106230 4 VSS
port 42 nsew
rlabel locali s -10709 106351 -10467 106385 4 VSS
port 42 nsew
rlabel locali s -12879 106230 -12766 106379 4 VSS
port 42 nsew
rlabel locali s -10553 106385 -10467 106455 4 VSS
port 42 nsew
rlabel locali s -12879 106379 -12647 106386 4 VSS
port 42 nsew
rlabel locali s -12879 106386 -12354 106420 4 VSS
port 42 nsew
rlabel locali s -12879 106420 -12647 106426 4 VSS
port 42 nsew
rlabel locali s -10553 106455 -9999 106516 4 VSS
port 42 nsew
rlabel locali s -9426 106629 -9184 106636 4 VSS
port 42 nsew
rlabel locali s -9426 106636 -8901 106670 4 VSS
port 42 nsew
rlabel locali s -9426 106670 -9184 106676 4 VSS
port 42 nsew
rlabel locali s -9426 106676 -9313 107553 4 VSS
port 42 nsew
rlabel locali s -10553 106516 -10467 106547 4 VSS
port 42 nsew
rlabel locali s -10709 106547 -10467 106581 4 VSS
port 42 nsew
rlabel locali s -10553 106581 -10467 106996 4 VSS
port 42 nsew
rlabel locali s -12879 106426 -12766 106621 4 VSS
port 42 nsew
rlabel locali s -12879 106621 -12637 106628 4 VSS
port 42 nsew
rlabel locali s -12879 106628 -12354 106662 4 VSS
port 42 nsew
rlabel locali s -12879 106662 -12637 106668 4 VSS
port 42 nsew
rlabel locali s -12879 106668 -12766 106933 4 VSS
port 42 nsew
rlabel locali s -9426 107553 -9245 107666 4 VSS
port 42 nsew
rlabel locali s -9358 107666 -9245 108014 4 VSS
port 42 nsew
rlabel locali s -13089 104331 -12953 107794 4 VSS
port 42 nsew
rlabel locali s -13089 107794 -11921 107930 4 VSS
port 42 nsew
rlabel locali s -9410 108014 -9245 108090 4 VSS
port 42 nsew
rlabel locali s -9410 108090 -9134 108092 4 VSS
port 42 nsew
rlabel locali s -9410 108092 -8843 108126 4 VSS
port 42 nsew
rlabel locali s -9410 108126 -9134 108127 4 VSS
port 42 nsew
rlabel locali s -9410 108127 -9245 108164 4 VSS
port 42 nsew
rlabel locali s -9410 108164 -9249 108882 4 VSS
port 42 nsew
rlabel locali s -11957 107930 -11921 108208 4 VSS
port 42 nsew
rlabel locali s -11959 108208 -11919 108228 4 VSS
port 42 nsew
rlabel locali s -9410 108882 -9134 108883 4 VSS
port 42 nsew
rlabel locali s -9410 108883 -8643 108917 4 VSS
port 42 nsew
rlabel locali s -9410 108917 -9134 108919 4 VSS
port 42 nsew
rlabel locali s -9410 108919 -9249 109010 4 VSS
port 42 nsew
rlabel locali s -9410 109010 -9133 109013 4 VSS
port 42 nsew
rlabel locali s -9410 109013 -8643 109047 4 VSS
port 42 nsew
rlabel locali s -9410 109047 -9249 109337 4 VSS
port 42 nsew
rlabel locali s -10255 108297 -10169 108437 4 VSS
port 42 nsew
rlabel locali s -11967 108228 -11913 108363 4 VSS
port 42 nsew
rlabel locali s -12520 108293 -12459 108410 4 VSS
port 42 nsew
rlabel locali s -12520 108410 -12407 108411 4 VSS
port 42 nsew
rlabel locali s -10511 108437 -10169 108471 4 VSS
port 42 nsew
rlabel locali s -12520 108411 -12099 108445 4 VSS
port 42 nsew
rlabel locali s -10255 108471 -10169 108633 4 VSS
port 42 nsew
rlabel locali s -10511 108633 -10169 108667 4 VSS
port 42 nsew
rlabel locali s -10255 108667 -10169 109149 4 VSS
port 42 nsew
rlabel locali s -12520 108445 -12459 108735 4 VSS
port 42 nsew
rlabel locali s -12520 108735 -12441 108742 4 VSS
port 42 nsew
rlabel locali s -12034 108880 -11948 109020 4 VSS
port 42 nsew
rlabel locali s -12034 109020 -11792 109054 4 VSS
port 42 nsew
rlabel locali s -9410 109337 -9132 109339 4 VSS
port 42 nsew
rlabel locali s -9410 109339 -8843 109373 4 VSS
port 42 nsew
rlabel locali s -9410 109373 -9132 109374 4 VSS
port 42 nsew
rlabel locali s -9410 109374 -9249 109487 4 VSS
port 42 nsew
rlabel locali s -10255 109149 -10002 109235 4 VSS
port 42 nsew
rlabel locali s -12034 109054 -11948 109124 4 VSS
port 42 nsew
rlabel locali s -12502 108742 -12441 109124 4 VSS
port 42 nsew
rlabel locali s -12910 109124 -11948 109185 4 VSS
port 42 nsew
rlabel locali s -12034 109185 -11948 109216 4 VSS
port 42 nsew
rlabel locali s -10088 109235 -10002 109409 4 VSS
port 42 nsew
rlabel locali s -12034 109216 -11792 109250 4 VSS
port 42 nsew
rlabel locali s -10125 109409 -10002 109410 4 VSS
port 42 nsew
rlabel locali s -10433 109410 -10002 109444 4 VSS
port 42 nsew
rlabel locali s -10088 109444 -10002 109734 4 VSS
port 42 nsew
rlabel locali s -12034 109250 -11948 109495 4 VSS
port 42 nsew
rlabel locali s -10091 109734 -10002 109814 4 VSS
port 42 nsew
rlabel locali s -10091 109814 -10030 110123 4 VSS
port 42 nsew
rlabel locali s -12910 109185 -12797 109851 4 VSS
port 42 nsew
rlabel locali s -12910 109851 -12679 109858 4 VSS
port 42 nsew
rlabel locali s -10584 109879 -10498 110019 4 VSS
port 42 nsew
rlabel locali s -12910 109858 -12385 109892 4 VSS
port 42 nsew
rlabel locali s -12910 109892 -12679 109898 4 VSS
port 42 nsew
rlabel locali s -10740 110019 -10498 110053 4 VSS
port 42 nsew
rlabel locali s -12910 109898 -12797 110047 4 VSS
port 42 nsew
rlabel locali s -10584 110053 -10498 110123 4 VSS
port 42 nsew
rlabel locali s -12910 110047 -12678 110054 4 VSS
port 42 nsew
rlabel locali s -12910 110054 -12385 110088 4 VSS
port 42 nsew
rlabel locali s -12910 110088 -12678 110094 4 VSS
port 42 nsew
rlabel locali s -10584 110123 -10030 110184 4 VSS
port 42 nsew
rlabel locali s -10584 110184 -10498 110215 4 VSS
port 42 nsew
rlabel locali s -10740 110215 -10498 110249 4 VSS
port 42 nsew
rlabel locali s -10584 110249 -10498 110664 4 VSS
port 42 nsew
rlabel locali s -12910 110094 -12797 110289 4 VSS
port 42 nsew
rlabel locali s -12910 110289 -12668 110296 4 VSS
port 42 nsew
rlabel locali s -12910 110296 -12385 110330 4 VSS
port 42 nsew
rlabel locali s -12910 110330 -12668 110336 4 VSS
port 42 nsew
rlabel locali s -12910 110336 -12797 110601 4 VSS
port 42 nsew
rlabel locali s -11888 113376 -11852 113559 4 VSS
port 42 nsew
rlabel locali s -13051 113559 -11852 113583 4 VSS
port 42 nsew
rlabel locali s -16160 8555 -16024 113583 4 VSS
port 42 nsew
rlabel locali s -16160 113583 -11852 113695 4 VSS
port 42 nsew
rlabel locali s -11888 113695 -11852 113904 4 VSS
port 42 nsew
rlabel locali s -16160 113695 -12915 113719 4 VSS
port 42 nsew
rlabel locali s -11890 113904 -11850 113924 4 VSS
port 42 nsew
rlabel locali s -6733 114001 -6647 114141 4 VSS
port 42 nsew
rlabel locali s -8998 113997 -8937 114114 4 VSS
port 42 nsew
rlabel locali s -8998 114114 -8885 114115 4 VSS
port 42 nsew
rlabel locali s -6989 114141 -6647 114175 4 VSS
port 42 nsew
rlabel locali s -8998 114115 -8577 114149 4 VSS
port 42 nsew
rlabel locali s -6733 114175 -6647 114337 4 VSS
port 42 nsew
rlabel locali s -6989 114337 -6647 114371 4 VSS
port 42 nsew
rlabel locali s -6733 114371 -6647 114853 4 VSS
port 42 nsew
rlabel locali s -8998 114149 -8937 114439 4 VSS
port 42 nsew
rlabel locali s -8998 114439 -8919 114446 4 VSS
port 42 nsew
rlabel locali s -10186 113993 -10100 114133 4 VSS
port 42 nsew
rlabel locali s -11898 113924 -11844 114059 4 VSS
port 42 nsew
rlabel locali s -12451 113989 -12390 114106 4 VSS
port 42 nsew
rlabel locali s -12451 114106 -12338 114107 4 VSS
port 42 nsew
rlabel locali s -10442 114133 -10100 114167 4 VSS
port 42 nsew
rlabel locali s -12451 114107 -12030 114141 4 VSS
port 42 nsew
rlabel locali s -10186 114167 -10100 114329 4 VSS
port 42 nsew
rlabel locali s -10442 114329 -10100 114363 4 VSS
port 42 nsew
rlabel locali s -8512 114584 -8426 114724 4 VSS
port 42 nsew
rlabel locali s -8512 114724 -8270 114758 4 VSS
port 42 nsew
rlabel locali s -6733 114853 -6480 114939 4 VSS
port 42 nsew
rlabel locali s -8512 114758 -8426 114828 4 VSS
port 42 nsew
rlabel locali s -8980 114446 -8919 114828 4 VSS
port 42 nsew
rlabel locali s -9388 114828 -8426 114889 4 VSS
port 42 nsew
rlabel locali s -10186 114363 -10100 114845 4 VSS
port 42 nsew
rlabel locali s -12451 114141 -12390 114431 4 VSS
port 42 nsew
rlabel locali s -12451 114431 -12372 114438 4 VSS
port 42 nsew
rlabel locali s -11965 114576 -11879 114716 4 VSS
port 42 nsew
rlabel locali s -11965 114716 -11723 114750 4 VSS
port 42 nsew
rlabel locali s -8512 114889 -8426 114920 4 VSS
port 42 nsew
rlabel locali s -6566 114939 -6480 115092 4 VSS
port 42 nsew
rlabel locali s -8512 114920 -8270 114954 4 VSS
port 42 nsew
rlabel locali s -6566 115092 -5618 115113 4 VSS
port 42 nsew
rlabel locali s -6603 115113 -5618 115114 4 VSS
port 42 nsew
rlabel locali s -6911 115114 -5618 115148 4 VSS
port 42 nsew
rlabel locali s -6566 115148 -5618 115303 4 VSS
port 42 nsew
rlabel locali s -8512 114954 -8426 115199 4 VSS
port 42 nsew
rlabel locali s -6124 115303 -5618 116969 4 VSS
port 42 nsew
rlabel locali s -6566 115303 -6480 115438 4 VSS
port 42 nsew
rlabel locali s -6569 115438 -6480 115518 4 VSS
port 42 nsew
rlabel locali s -6569 115518 -6508 115827 4 VSS
port 42 nsew
rlabel locali s -9388 114889 -9275 115555 4 VSS
port 42 nsew
rlabel locali s -10186 114845 -9933 114931 4 VSS
port 42 nsew
rlabel locali s -11965 114750 -11879 114820 4 VSS
port 42 nsew
rlabel locali s -12433 114438 -12372 114820 4 VSS
port 42 nsew
rlabel locali s -12841 114820 -11879 114881 4 VSS
port 42 nsew
rlabel locali s -11965 114881 -11879 114912 4 VSS
port 42 nsew
rlabel locali s -10019 114931 -9933 115105 4 VSS
port 42 nsew
rlabel locali s -11965 114912 -11723 114946 4 VSS
port 42 nsew
rlabel locali s -10056 115105 -9933 115106 4 VSS
port 42 nsew
rlabel locali s -10364 115106 -9933 115140 4 VSS
port 42 nsew
rlabel locali s -10019 115140 -9933 115430 4 VSS
port 42 nsew
rlabel locali s -11965 114946 -11879 115191 4 VSS
port 42 nsew
rlabel locali s -10022 115430 -9933 115510 4 VSS
port 42 nsew
rlabel locali s -9388 115555 -9157 115562 4 VSS
port 42 nsew
rlabel locali s -7062 115583 -6976 115723 4 VSS
port 42 nsew
rlabel locali s -9388 115562 -8863 115596 4 VSS
port 42 nsew
rlabel locali s -9388 115596 -9157 115602 4 VSS
port 42 nsew
rlabel locali s -7218 115723 -6976 115757 4 VSS
port 42 nsew
rlabel locali s -9388 115602 -9275 115751 4 VSS
port 42 nsew
rlabel locali s -7062 115757 -6976 115827 4 VSS
port 42 nsew
rlabel locali s -9388 115751 -9156 115758 4 VSS
port 42 nsew
rlabel locali s -9388 115758 -8863 115792 4 VSS
port 42 nsew
rlabel locali s -9388 115792 -9156 115798 4 VSS
port 42 nsew
rlabel locali s -7062 115827 -6508 115888 4 VSS
port 42 nsew
rlabel locali s -7062 115888 -6976 115919 4 VSS
port 42 nsew
rlabel locali s -7218 115919 -6976 115953 4 VSS
port 42 nsew
rlabel locali s -7062 115953 -6976 116368 4 VSS
port 42 nsew
rlabel locali s -9388 115798 -9275 115993 4 VSS
port 42 nsew
rlabel locali s -10022 115510 -9961 115819 4 VSS
port 42 nsew
rlabel locali s -12841 114881 -12728 115547 4 VSS
port 42 nsew
rlabel locali s -12841 115547 -12610 115554 4 VSS
port 42 nsew
rlabel locali s -10515 115575 -10429 115715 4 VSS
port 42 nsew
rlabel locali s -12841 115554 -12316 115588 4 VSS
port 42 nsew
rlabel locali s -12841 115588 -12610 115594 4 VSS
port 42 nsew
rlabel locali s -10671 115715 -10429 115749 4 VSS
port 42 nsew
rlabel locali s -12841 115594 -12728 115743 4 VSS
port 42 nsew
rlabel locali s -10515 115749 -10429 115819 4 VSS
port 42 nsew
rlabel locali s -12841 115743 -12609 115750 4 VSS
port 42 nsew
rlabel locali s -12841 115750 -12316 115784 4 VSS
port 42 nsew
rlabel locali s -12841 115784 -12609 115790 4 VSS
port 42 nsew
rlabel locali s -10515 115819 -9961 115880 4 VSS
port 42 nsew
rlabel locali s -9388 115993 -9146 116000 4 VSS
port 42 nsew
rlabel locali s -9388 116000 -8863 116034 4 VSS
port 42 nsew
rlabel locali s -9388 116034 -9146 116040 4 VSS
port 42 nsew
rlabel locali s -9388 116040 -9275 116917 4 VSS
port 42 nsew
rlabel locali s -10515 115880 -10429 115911 4 VSS
port 42 nsew
rlabel locali s -10671 115911 -10429 115945 4 VSS
port 42 nsew
rlabel locali s -10515 115945 -10429 116360 4 VSS
port 42 nsew
rlabel locali s -12841 115790 -12728 115985 4 VSS
port 42 nsew
rlabel locali s -12841 115985 -12599 115992 4 VSS
port 42 nsew
rlabel locali s -12841 115992 -12316 116026 4 VSS
port 42 nsew
rlabel locali s -12841 116026 -12599 116032 4 VSS
port 42 nsew
rlabel locali s -12841 116032 -12728 116297 4 VSS
port 42 nsew
rlabel locali s -9388 116917 -9207 117030 4 VSS
port 42 nsew
rlabel locali s -9320 117030 -9207 117378 4 VSS
port 42 nsew
rlabel locali s -13051 113719 -12915 117158 4 VSS
port 42 nsew
rlabel locali s -13051 117158 -11883 117294 4 VSS
port 42 nsew
rlabel locali s -9372 117378 -9207 117454 4 VSS
port 42 nsew
rlabel locali s -9372 117454 -9096 117456 4 VSS
port 42 nsew
rlabel locali s -9372 117456 -8805 117490 4 VSS
port 42 nsew
rlabel locali s -9372 117490 -9096 117491 4 VSS
port 42 nsew
rlabel locali s -9372 117491 -9207 117528 4 VSS
port 42 nsew
rlabel locali s -9372 117528 -9211 118246 4 VSS
port 42 nsew
rlabel locali s -11919 117294 -11883 117572 4 VSS
port 42 nsew
rlabel locali s -11921 117572 -11881 117592 4 VSS
port 42 nsew
rlabel locali s -9372 118246 -9096 118247 4 VSS
port 42 nsew
rlabel locali s -9372 118247 -8605 118281 4 VSS
port 42 nsew
rlabel locali s -9372 118281 -9096 118283 4 VSS
port 42 nsew
rlabel locali s -9372 118283 -9211 118374 4 VSS
port 42 nsew
rlabel locali s -9372 118374 -9095 118377 4 VSS
port 42 nsew
rlabel locali s -9372 118377 -8605 118411 4 VSS
port 42 nsew
rlabel locali s -9372 118411 -9211 118701 4 VSS
port 42 nsew
rlabel locali s -10217 117661 -10131 117801 4 VSS
port 42 nsew
rlabel locali s -11929 117592 -11875 117727 4 VSS
port 42 nsew
rlabel locali s -12482 117657 -12421 117774 4 VSS
port 42 nsew
rlabel locali s -12482 117774 -12369 117775 4 VSS
port 42 nsew
rlabel locali s -10473 117801 -10131 117835 4 VSS
port 42 nsew
rlabel locali s -12482 117775 -12061 117809 4 VSS
port 42 nsew
rlabel locali s -10217 117835 -10131 117997 4 VSS
port 42 nsew
rlabel locali s -10473 117997 -10131 118031 4 VSS
port 42 nsew
rlabel locali s -10217 118031 -10131 118513 4 VSS
port 42 nsew
rlabel locali s -12482 117809 -12421 118099 4 VSS
port 42 nsew
rlabel locali s -12482 118099 -12403 118106 4 VSS
port 42 nsew
rlabel locali s -11996 118244 -11910 118384 4 VSS
port 42 nsew
rlabel locali s -11996 118384 -11754 118418 4 VSS
port 42 nsew
rlabel locali s -9372 118701 -9094 118703 4 VSS
port 42 nsew
rlabel locali s -9372 118703 -8805 118737 4 VSS
port 42 nsew
rlabel locali s -9372 118737 -9094 118738 4 VSS
port 42 nsew
rlabel locali s -9372 118738 -9211 118851 4 VSS
port 42 nsew
rlabel locali s -10217 118513 -9964 118599 4 VSS
port 42 nsew
rlabel locali s -11996 118418 -11910 118488 4 VSS
port 42 nsew
rlabel locali s -12464 118106 -12403 118488 4 VSS
port 42 nsew
rlabel locali s -12872 118488 -11910 118549 4 VSS
port 42 nsew
rlabel locali s -11996 118549 -11910 118580 4 VSS
port 42 nsew
rlabel locali s -10050 118599 -9964 118773 4 VSS
port 42 nsew
rlabel locali s -11996 118580 -11754 118614 4 VSS
port 42 nsew
rlabel locali s -10087 118773 -9964 118774 4 VSS
port 42 nsew
rlabel locali s -10395 118774 -9964 118808 4 VSS
port 42 nsew
rlabel locali s -10050 118808 -9964 119098 4 VSS
port 42 nsew
rlabel locali s -11996 118614 -11910 118859 4 VSS
port 42 nsew
rlabel locali s -10053 119098 -9964 119178 4 VSS
port 42 nsew
rlabel locali s -10053 119178 -9992 119487 4 VSS
port 42 nsew
rlabel locali s -12872 118549 -12759 119215 4 VSS
port 42 nsew
rlabel locali s -12872 119215 -12641 119222 4 VSS
port 42 nsew
rlabel locali s -10546 119243 -10460 119383 4 VSS
port 42 nsew
rlabel locali s -12872 119222 -12347 119256 4 VSS
port 42 nsew
rlabel locali s -12872 119256 -12641 119262 4 VSS
port 42 nsew
rlabel locali s -10702 119383 -10460 119417 4 VSS
port 42 nsew
rlabel locali s -12872 119262 -12759 119411 4 VSS
port 42 nsew
rlabel locali s -10546 119417 -10460 119487 4 VSS
port 42 nsew
rlabel locali s -12872 119411 -12640 119418 4 VSS
port 42 nsew
rlabel locali s -12872 119418 -12347 119452 4 VSS
port 42 nsew
rlabel locali s -12872 119452 -12640 119458 4 VSS
port 42 nsew
rlabel locali s -10546 119487 -9992 119548 4 VSS
port 42 nsew
rlabel locali s -10546 119548 -10460 119579 4 VSS
port 42 nsew
rlabel locali s -10702 119579 -10460 119613 4 VSS
port 42 nsew
rlabel locali s -10546 119613 -10460 120028 4 VSS
port 42 nsew
rlabel locali s -12872 119458 -12759 119653 4 VSS
port 42 nsew
rlabel locali s -12872 119653 -12630 119660 4 VSS
port 42 nsew
rlabel locali s -12872 119660 -12347 119694 4 VSS
port 42 nsew
rlabel locali s -12872 119694 -12630 119700 4 VSS
port 42 nsew
rlabel locali s -12872 119700 -12759 119965 4 VSS
port 42 nsew
rlabel pwell s 50911 -4368 58164 -4190 8 VSS
port 42 nsew
rlabel pwell s 63208 -3604 63794 -3484 8 VSS
port 42 nsew
rlabel pwell s 63208 -3467 63794 -3347 8 VSS
port 42 nsew
rlabel pwell s 62358 -3467 62944 -3347 8 VSS
port 42 nsew
rlabel pwell s 7795 -1943 15048 -1765 8 VSS
port 42 nsew
rlabel pwell s 50911 -1321 58164 -1143 8 VSS
port 42 nsew
rlabel pwell s 25581 -1450 47660 -1203 8 VSS
port 42 nsew
rlabel pwell s 51114 1590 58367 1768 6 VSS
port 42 nsew
rlabel pwell s 47413 -1203 47660 3506 6 VSS
port 42 nsew
rlabel pwell s 36735 -459 38123 -282 8 VSS
port 42 nsew
rlabel pwell s 35014 -502 36402 -325 8 VSS
port 42 nsew
rlabel pwell s 30279 -525 31667 -348 8 VSS
port 42 nsew
rlabel pwell s 32593 -291 34344 -148 8 VSS
port 42 nsew
rlabel pwell s 27738 -284 29489 -141 8 VSS
port 42 nsew
rlabel pwell s 45544 2016 46130 2136 6 VSS
port 42 nsew
rlabel pwell s 44484 1926 45070 2046 6 VSS
port 42 nsew
rlabel pwell s 43647 1926 44233 2046 6 VSS
port 42 nsew
rlabel pwell s 41784 1926 42370 2046 6 VSS
port 42 nsew
rlabel pwell s 40947 1926 41533 2046 6 VSS
port 42 nsew
rlabel pwell s 44476 2306 45062 2426 6 VSS
port 42 nsew
rlabel pwell s 42733 2306 43319 2426 6 VSS
port 42 nsew
rlabel pwell s 41776 2306 42362 2426 6 VSS
port 42 nsew
rlabel pwell s 40033 2306 40619 2426 6 VSS
port 42 nsew
rlabel pwell s 39151 2306 39737 2426 6 VSS
port 42 nsew
rlabel pwell s 36735 2607 38123 2784 6 VSS
port 42 nsew
rlabel pwell s 35014 2650 36402 2827 6 VSS
port 42 nsew
rlabel pwell s 30279 2628 31667 2805 6 VSS
port 42 nsew
rlabel pwell s 25581 -1203 25828 3506 6 VSS
port 42 nsew
rlabel pwell s 5345 -1243 5931 -1123 8 VSS
port 42 nsew
rlabel pwell s 5345 -1106 5931 -986 8 VSS
port 42 nsew
rlabel pwell s 4495 -1106 5081 -986 8 VSS
port 42 nsew
rlabel pwell s 20781 -738 21367 -618 8 VSS
port 42 nsew
rlabel pwell s 20781 -601 21367 -481 8 VSS
port 42 nsew
rlabel pwell s 19931 -601 20517 -481 8 VSS
port 42 nsew
rlabel pwell s 539 469 2991 602 6 VSS
port 42 nsew
rlabel pwell s 1535 602 2991 616 6 VSS
port 42 nsew
rlabel pwell s 539 602 1153 616 6 VSS
port 42 nsew
rlabel pwell s 2429 616 2991 716 6 VSS
port 42 nsew
rlabel pwell s 565 616 818 716 6 VSS
port 42 nsew
rlabel pwell s 7836 813 15089 991 6 VSS
port 42 nsew
rlabel pwell s 5330 1447 5916 1567 6 VSS
port 42 nsew
rlabel pwell s 5330 1584 5916 1704 6 VSS
port 42 nsew
rlabel pwell s 4480 1584 5066 1704 6 VSS
port 42 nsew
rlabel pwell s 2429 2146 2991 2246 6 VSS
port 42 nsew
rlabel pwell s 565 2146 818 2246 6 VSS
port 42 nsew
rlabel pwell s 1535 2246 2991 2248 6 VSS
port 42 nsew
rlabel pwell s 1535 2248 3125 2260 6 VSS
port 42 nsew
rlabel pwell s 539 2246 1153 2260 6 VSS
port 42 nsew
rlabel pwell s 539 2260 3125 2393 6 VSS
port 42 nsew
rlabel pwell s 2794 2393 3125 2534 6 VSS
port 42 nsew
rlabel pwell s 20609 2612 21195 2732 6 VSS
port 42 nsew
rlabel pwell s 20609 2749 21195 2869 6 VSS
port 42 nsew
rlabel pwell s 19759 2749 20345 2869 6 VSS
port 42 nsew
rlabel pwell s 25581 3506 47660 3753 6 VSS
port 42 nsew
rlabel pwell s 8082 4332 12576 4530 6 VSS
port 42 nsew
rlabel pwell s 69208 9612 92372 10082 6 VSS
port 42 nsew
rlabel pwell s 17109 8966 17341 10210 6 VSS
port 42 nsew
rlabel pwell s -6844 10549 -6727 11875 4 VSS
port 42 nsew
rlabel pwell s -8664 10586 -8551 11087 4 VSS
port 42 nsew
rlabel pwell s -8173 11229 -8042 11810 4 VSS
port 42 nsew
rlabel pwell s -12287 10660 -12129 11569 4 VSS
port 42 nsew
rlabel pwell s -12822 10420 -12705 11746 4 VSS
port 42 nsew
rlabel pwell s -6755 12528 -6642 13029 4 VSS
port 42 nsew
rlabel pwell s -6264 13171 -6133 13752 4 VSS
port 42 nsew
rlabel pwell s -8780 12379 -8663 13705 4 VSS
port 42 nsew
rlabel pwell s -11921 11842 -11780 12491 4 VSS
port 42 nsew
rlabel pwell s -11922 12747 -11781 13396 4 VSS
port 42 nsew
rlabel pwell s -6170 14164 -6057 14665 4 VSS
port 42 nsew
rlabel pwell s -8455 14224 -8324 14805 4 VSS
port 42 nsew
rlabel pwell s -11170 14164 -11057 14665 4 VSS
port 42 nsew
rlabel pwell s -13455 14224 -13324 14805 4 VSS
port 42 nsew
rlabel pwell s -6679 14807 -6548 15388 4 VSS
port 42 nsew
rlabel pwell s -5831 15640 -5697 16439 4 VSS
port 42 nsew
rlabel pwell s -8617 15163 -8504 15664 4 VSS
port 42 nsew
rlabel pwell s -11679 14807 -11548 15388 4 VSS
port 42 nsew
rlabel pwell s -8126 15806 -7995 16387 4 VSS
port 42 nsew
rlabel pwell s -10831 15640 -10697 16439 4 VSS
port 42 nsew
rlabel pwell s -13617 15163 -13504 15664 4 VSS
port 42 nsew
rlabel pwell s -13126 15806 -12995 16387 4 VSS
port 42 nsew
rlabel pwell s -5495 18139 -5375 18725 4 VSS
port 42 nsew
rlabel pwell s -5875 18147 -5755 18733 4 VSS
port 42 nsew
rlabel pwell s -10422 18139 -10302 18725 4 VSS
port 42 nsew
rlabel pwell s -10802 18147 -10682 18733 4 VSS
port 42 nsew
rlabel pwell s -5495 18976 -5375 19562 4 VSS
port 42 nsew
rlabel pwell s -7146 19153 -7033 19654 4 VSS
port 42 nsew
rlabel pwell s -9431 19213 -9300 19794 4 VSS
port 42 nsew
rlabel pwell s -10422 18976 -10302 19562 4 VSS
port 42 nsew
rlabel pwell s -5875 19890 -5755 20476 4 VSS
port 42 nsew
rlabel pwell s -7655 19796 -7524 20377 4 VSS
port 42 nsew
rlabel pwell s -5495 20839 -5375 21425 4 VSS
port 42 nsew
rlabel pwell s -5875 20847 -5755 21433 4 VSS
port 42 nsew
rlabel pwell s -6807 20629 -6673 21428 4 VSS
port 42 nsew
rlabel pwell s -9593 20152 -9480 20653 4 VSS
port 42 nsew
rlabel pwell s -10802 19890 -10682 20476 4 VSS
port 42 nsew
rlabel pwell s -9102 20795 -8971 21376 4 VSS
port 42 nsew
rlabel pwell s -10422 20839 -10302 21425 4 VSS
port 42 nsew
rlabel pwell s -10802 20847 -10682 21433 4 VSS
port 42 nsew
rlabel pwell s -5495 21676 -5375 22262 4 VSS
port 42 nsew
rlabel pwell s -10422 21676 -10302 22262 4 VSS
port 42 nsew
rlabel pwell s -5875 22590 -5755 23176 4 VSS
port 42 nsew
rlabel pwell s -10802 22590 -10682 23176 4 VSS
port 42 nsew
rlabel pwell s -5875 23472 -5755 24058 4 VSS
port 42 nsew
rlabel pwell s -10802 23472 -10682 24058 4 VSS
port 42 nsew
rlabel pwell s -6305 24407 -6171 25206 4 VSS
port 42 nsew
rlabel pwell s -11239 24434 -11105 25233 4 VSS
port 42 nsew
rlabel pwell s -6092 26270 -5972 26856 4 VSS
port 42 nsew
rlabel pwell s -7933 26021 -7813 26607 4 VSS
port 42 nsew
rlabel pwell s -8313 26013 -8193 26599 4 VSS
port 42 nsew
rlabel pwell s -10689 26013 -10569 26599 4 VSS
port 42 nsew
rlabel pwell s -11069 26021 -10949 26607 4 VSS
port 42 nsew
rlabel pwell s -6081 27039 -5933 27723 4 VSS
port 42 nsew
rlabel pwell s -8313 26850 -8193 27436 4 VSS
port 42 nsew
rlabel pwell s -10689 26850 -10569 27436 4 VSS
port 42 nsew
rlabel pwell s -12949 27039 -12801 27723 4 VSS
port 42 nsew
rlabel pwell s -7933 27764 -7813 28350 4 VSS
port 42 nsew
rlabel pwell s -11069 27764 -10949 28350 4 VSS
port 42 nsew
rlabel pwell s -7933 28721 -7813 29307 4 VSS
port 42 nsew
rlabel pwell s -8313 28713 -8193 29299 4 VSS
port 42 nsew
rlabel pwell s -10689 28713 -10569 29299 4 VSS
port 42 nsew
rlabel pwell s -11069 28721 -10949 29307 4 VSS
port 42 nsew
rlabel pwell s -6081 29539 -5933 30223 4 VSS
port 42 nsew
rlabel pwell s -8313 29550 -8193 30136 4 VSS
port 42 nsew
rlabel pwell s -10689 29550 -10569 30136 4 VSS
port 42 nsew
rlabel pwell s -12949 29539 -12801 30223 4 VSS
port 42 nsew
rlabel pwell s -7933 30464 -7813 31050 4 VSS
port 42 nsew
rlabel pwell s -11069 30464 -10949 31050 4 VSS
port 42 nsew
rlabel pwell s -7933 31346 -7813 31932 4 VSS
port 42 nsew
rlabel pwell s -11069 31346 -10949 31932 4 VSS
port 42 nsew
rlabel pwell s -6081 32039 -5933 32723 4 VSS
port 42 nsew
rlabel pwell s -8512 32265 -8395 33591 4 VSS
port 42 nsew
rlabel pwell s -10487 32265 -10370 33591 4 VSS
port 42 nsew
rlabel pwell s -12949 32039 -12801 32723 4 VSS
port 42 nsew
rlabel pwell s -6081 34539 -5933 35223 4 VSS
port 42 nsew
rlabel pwell s -7824 33991 -7693 34572 4 VSS
port 42 nsew
rlabel pwell s -11189 33991 -11058 34572 4 VSS
port 42 nsew
rlabel pwell s -8315 34714 -8202 35215 4 VSS
port 42 nsew
rlabel pwell s -10680 34714 -10567 35215 4 VSS
port 42 nsew
rlabel pwell s -12949 34539 -12801 35223 4 VSS
port 42 nsew
rlabel pwell s -7826 35596 -7695 36177 4 VSS
port 42 nsew
rlabel pwell s -11187 35596 -11056 36177 4 VSS
port 42 nsew
rlabel pwell s -8317 36319 -8204 36820 4 VSS
port 42 nsew
rlabel pwell s -10678 36319 -10565 36820 4 VSS
port 42 nsew
rlabel pwell s -6081 37039 -5933 37723 4 VSS
port 42 nsew
rlabel pwell s -8503 37227 -8386 38553 4 VSS
port 42 nsew
rlabel pwell s -10496 37227 -10379 38553 4 VSS
port 42 nsew
rlabel pwell s -12949 37039 -12801 37723 4 VSS
port 42 nsew
rlabel pwell s -6081 40039 -5933 40723 4 VSS
port 42 nsew
rlabel pwell s -8332 40049 -8184 40733 4 VSS
port 42 nsew
rlabel pwell s -10698 40049 -10550 40733 4 VSS
port 42 nsew
rlabel pwell s -12949 40039 -12801 40723 4 VSS
port 42 nsew
rlabel pwell s -12758 43850 -12638 44436 4 VSS
port 42 nsew
rlabel pwell s -12758 44732 -12638 45318 4 VSS
port 42 nsew
rlabel pwell s -13138 45646 -13018 46232 4 VSS
port 42 nsew
rlabel pwell s -12758 46475 -12638 47061 4 VSS
port 42 nsew
rlabel pwell s -13138 46483 -13018 47069 4 VSS
port 42 nsew
rlabel pwell s -12758 47432 -12638 48018 4 VSS
port 42 nsew
rlabel pwell s -13138 48346 -13018 48932 4 VSS
port 42 nsew
rlabel pwell s -12758 49175 -12638 49761 4 VSS
port 42 nsew
rlabel pwell s -13138 49183 -13018 49769 4 VSS
port 42 nsew
rlabel pwell s -7720 50655 -7562 51564 4 VSS
port 42 nsew
rlabel pwell s -10344 50626 -10203 51275 4 VSS
port 42 nsew
rlabel pwell s -8582 51978 -8462 52564 4 VSS
port 42 nsew
rlabel pwell s -10344 51572 -10203 52221 4 VSS
port 42 nsew
rlabel pwell s -8582 52860 -8462 53446 4 VSS
port 42 nsew
rlabel pwell s -8202 53774 -8082 54360 4 VSS
port 42 nsew
rlabel pwell s -10277 52523 -10160 53849 4 VSS
port 42 nsew
rlabel pwell s -8202 54611 -8082 55197 4 VSS
port 42 nsew
rlabel pwell s -8582 54603 -8462 55189 4 VSS
port 42 nsew
rlabel pwell s -10712 54399 -10579 54930 4 VSS
port 42 nsew
rlabel pwell s -10835 54373 -10715 54959 4 VSS
port 42 nsew
rlabel pwell s -8582 55560 -8462 56146 4 VSS
port 42 nsew
rlabel pwell s -8202 56474 -8082 57060 4 VSS
port 42 nsew
rlabel pwell s -8202 57311 -8082 57897 4 VSS
port 42 nsew
rlabel pwell s -8582 57303 -8462 57889 4 VSS
port 42 nsew
rlabel pwell s -9597 55165 -9448 57944 4 VSS
port 42 nsew
rlabel pwell s -6862 60259 -6731 60840 4 VSS
port 42 nsew
rlabel pwell s -9129 60199 -9016 60700 4 VSS
port 42 nsew
rlabel pwell s -10315 60251 -10184 60832 4 VSS
port 42 nsew
rlabel pwell s -12582 60191 -12469 60692 4 VSS
port 42 nsew
rlabel pwell s -6682 61198 -6569 61699 4 VSS
port 42 nsew
rlabel pwell s -8638 60842 -8507 61423 4 VSS
port 42 nsew
rlabel pwell s -7191 61841 -7060 62422 4 VSS
port 42 nsew
rlabel pwell s -9489 61675 -9355 62474 4 VSS
port 42 nsew
rlabel pwell s -10135 61190 -10022 61691 4 VSS
port 42 nsew
rlabel pwell s -12091 60834 -11960 61415 4 VSS
port 42 nsew
rlabel pwell s -10644 61833 -10513 62414 4 VSS
port 42 nsew
rlabel pwell s -12942 61667 -12808 62466 4 VSS
port 42 nsew
rlabel pwell s -9503 63580 -9290 65105 4 VSS
port 42 nsew
rlabel pwell s -10346 63919 -10215 64500 4 VSS
port 42 nsew
rlabel pwell s -12613 63859 -12500 64360 4 VSS
port 42 nsew
rlabel pwell s -10166 64858 -10053 65359 4 VSS
port 42 nsew
rlabel pwell s -12122 64502 -11991 65083 4 VSS
port 42 nsew
rlabel pwell s -10675 65501 -10544 66082 4 VSS
port 42 nsew
rlabel pwell s -12973 65335 -12839 66134 4 VSS
port 42 nsew
rlabel pwell s -6873 68699 -6742 69280 4 VSS
port 42 nsew
rlabel pwell s -9140 68639 -9027 69140 4 VSS
port 42 nsew
rlabel pwell s -10326 68691 -10195 69272 4 VSS
port 42 nsew
rlabel pwell s -12593 68631 -12480 69132 4 VSS
port 42 nsew
rlabel pwell s -6693 69638 -6580 70139 4 VSS
port 42 nsew
rlabel pwell s -8649 69282 -8518 69863 4 VSS
port 42 nsew
rlabel pwell s -7202 70281 -7071 70862 4 VSS
port 42 nsew
rlabel pwell s -9500 70115 -9366 70914 4 VSS
port 42 nsew
rlabel pwell s -10146 69630 -10033 70131 4 VSS
port 42 nsew
rlabel pwell s -12102 69274 -11971 69855 4 VSS
port 42 nsew
rlabel pwell s -10655 70273 -10524 70854 4 VSS
port 42 nsew
rlabel pwell s -12953 70107 -12819 70906 4 VSS
port 42 nsew
rlabel pwell s -9514 72020 -9301 73545 4 VSS
port 42 nsew
rlabel pwell s -10357 72359 -10226 72940 4 VSS
port 42 nsew
rlabel pwell s -12624 72299 -12511 72800 4 VSS
port 42 nsew
rlabel pwell s -10177 73298 -10064 73799 4 VSS
port 42 nsew
rlabel pwell s -12133 72942 -12002 73523 4 VSS
port 42 nsew
rlabel pwell s -10686 73941 -10555 74522 4 VSS
port 42 nsew
rlabel pwell s -12984 73775 -12850 74574 4 VSS
port 42 nsew
rlabel pwell s -6912 77562 -6781 78143 4 VSS
port 42 nsew
rlabel pwell s -9179 77502 -9066 78003 4 VSS
port 42 nsew
rlabel pwell s -10365 77554 -10234 78135 4 VSS
port 42 nsew
rlabel pwell s -12632 77494 -12519 77995 4 VSS
port 42 nsew
rlabel pwell s -6732 78501 -6619 79002 4 VSS
port 42 nsew
rlabel pwell s -8688 78145 -8557 78726 4 VSS
port 42 nsew
rlabel pwell s -7241 79144 -7110 79725 4 VSS
port 42 nsew
rlabel pwell s -9539 78978 -9405 79777 4 VSS
port 42 nsew
rlabel pwell s -10185 78493 -10072 78994 4 VSS
port 42 nsew
rlabel pwell s -12141 78137 -12010 78718 4 VSS
port 42 nsew
rlabel pwell s -10694 79136 -10563 79717 4 VSS
port 42 nsew
rlabel pwell s -12992 78970 -12858 79769 4 VSS
port 42 nsew
rlabel pwell s -9553 80883 -9340 82408 4 VSS
port 42 nsew
rlabel pwell s -10396 81222 -10265 81803 4 VSS
port 42 nsew
rlabel pwell s -12663 81162 -12550 81663 4 VSS
port 42 nsew
rlabel pwell s -10216 82161 -10103 82662 4 VSS
port 42 nsew
rlabel pwell s -12172 81805 -12041 82386 4 VSS
port 42 nsew
rlabel pwell s -10725 82804 -10594 83385 4 VSS
port 42 nsew
rlabel pwell s -13023 82638 -12889 83437 4 VSS
port 42 nsew
rlabel pwell s -6878 86760 -6747 87341 4 VSS
port 42 nsew
rlabel pwell s -9145 86700 -9032 87201 4 VSS
port 42 nsew
rlabel pwell s -10331 86752 -10200 87333 4 VSS
port 42 nsew
rlabel pwell s -12598 86692 -12485 87193 4 VSS
port 42 nsew
rlabel pwell s -6698 87699 -6585 88200 4 VSS
port 42 nsew
rlabel pwell s -8654 87343 -8523 87924 4 VSS
port 42 nsew
rlabel pwell s -7207 88342 -7076 88923 4 VSS
port 42 nsew
rlabel pwell s -9505 88176 -9371 88975 4 VSS
port 42 nsew
rlabel pwell s -10151 87691 -10038 88192 4 VSS
port 42 nsew
rlabel pwell s -12107 87335 -11976 87916 4 VSS
port 42 nsew
rlabel pwell s -10660 88334 -10529 88915 4 VSS
port 42 nsew
rlabel pwell s -12958 88168 -12824 88967 4 VSS
port 42 nsew
rlabel pwell s -9519 90081 -9306 91606 4 VSS
port 42 nsew
rlabel pwell s -10362 90420 -10231 91001 4 VSS
port 42 nsew
rlabel pwell s -12629 90360 -12516 90861 4 VSS
port 42 nsew
rlabel pwell s -10182 91359 -10069 91860 4 VSS
port 42 nsew
rlabel pwell s -12138 91003 -12007 91584 4 VSS
port 42 nsew
rlabel pwell s -10691 92002 -10560 92583 4 VSS
port 42 nsew
rlabel pwell s -12989 91836 -12855 92635 4 VSS
port 42 nsew
rlabel pwell s -6812 95514 -6681 96095 4 VSS
port 42 nsew
rlabel pwell s -9079 95454 -8966 95955 4 VSS
port 42 nsew
rlabel pwell s -10265 95506 -10134 96087 4 VSS
port 42 nsew
rlabel pwell s -12532 95446 -12419 95947 4 VSS
port 42 nsew
rlabel pwell s -6632 96453 -6519 96954 4 VSS
port 42 nsew
rlabel pwell s -8588 96097 -8457 96678 4 VSS
port 42 nsew
rlabel pwell s -7141 97096 -7010 97677 4 VSS
port 42 nsew
rlabel pwell s -9439 96930 -9305 97729 4 VSS
port 42 nsew
rlabel pwell s -10085 96445 -9972 96946 4 VSS
port 42 nsew
rlabel pwell s -12041 96089 -11910 96670 4 VSS
port 42 nsew
rlabel pwell s -10594 97088 -10463 97669 4 VSS
port 42 nsew
rlabel pwell s -12892 96922 -12758 97721 4 VSS
port 42 nsew
rlabel pwell s -9453 98835 -9240 100360 4 VSS
port 42 nsew
rlabel pwell s -10296 99174 -10165 99755 4 VSS
port 42 nsew
rlabel pwell s -12563 99114 -12450 99615 4 VSS
port 42 nsew
rlabel pwell s -10116 100113 -10003 100614 4 VSS
port 42 nsew
rlabel pwell s -12072 99757 -11941 100338 4 VSS
port 42 nsew
rlabel pwell s -10625 100756 -10494 101337 4 VSS
port 42 nsew
rlabel pwell s -12923 100590 -12789 101389 4 VSS
port 42 nsew
rlabel pwell s -6795 104667 -6664 105248 4 VSS
port 42 nsew
rlabel pwell s -9062 104607 -8949 105108 4 VSS
port 42 nsew
rlabel pwell s -10248 104659 -10117 105240 4 VSS
port 42 nsew
rlabel pwell s -12515 104599 -12402 105100 4 VSS
port 42 nsew
rlabel pwell s -6615 105606 -6502 106107 4 VSS
port 42 nsew
rlabel pwell s -8571 105250 -8440 105831 4 VSS
port 42 nsew
rlabel pwell s -7124 106249 -6993 106830 4 VSS
port 42 nsew
rlabel pwell s -9422 106083 -9288 106882 4 VSS
port 42 nsew
rlabel pwell s -10068 105598 -9955 106099 4 VSS
port 42 nsew
rlabel pwell s -12024 105242 -11893 105823 4 VSS
port 42 nsew
rlabel pwell s -10577 106241 -10446 106822 4 VSS
port 42 nsew
rlabel pwell s -12875 106075 -12741 106874 4 VSS
port 42 nsew
rlabel pwell s -9436 107988 -9223 109513 4 VSS
port 42 nsew
rlabel pwell s -10279 108327 -10148 108908 4 VSS
port 42 nsew
rlabel pwell s -12546 108267 -12433 108768 4 VSS
port 42 nsew
rlabel pwell s -10099 109266 -9986 109767 4 VSS
port 42 nsew
rlabel pwell s -12055 108910 -11924 109491 4 VSS
port 42 nsew
rlabel pwell s -10608 109909 -10477 110490 4 VSS
port 42 nsew
rlabel pwell s -12906 109743 -12772 110542 4 VSS
port 42 nsew
rlabel pwell s -6757 114031 -6626 114612 4 VSS
port 42 nsew
rlabel pwell s -9024 113971 -8911 114472 4 VSS
port 42 nsew
rlabel pwell s -10210 114023 -10079 114604 4 VSS
port 42 nsew
rlabel pwell s -12477 113963 -12364 114464 4 VSS
port 42 nsew
rlabel pwell s -6577 114970 -6464 115471 4 VSS
port 42 nsew
rlabel pwell s -8533 114614 -8402 115195 4 VSS
port 42 nsew
rlabel pwell s -7086 115613 -6955 116194 4 VSS
port 42 nsew
rlabel pwell s -9384 115447 -9250 116246 4 VSS
port 42 nsew
rlabel pwell s -10030 114962 -9917 115463 4 VSS
port 42 nsew
rlabel pwell s -11986 114606 -11855 115187 4 VSS
port 42 nsew
rlabel pwell s -10539 115605 -10408 116186 4 VSS
port 42 nsew
rlabel pwell s -12837 115439 -12703 116238 4 VSS
port 42 nsew
rlabel pwell s -9398 117352 -9185 118877 4 VSS
port 42 nsew
rlabel pwell s -10241 117691 -10110 118272 4 VSS
port 42 nsew
rlabel pwell s -12508 117631 -12395 118132 4 VSS
port 42 nsew
rlabel pwell s -10061 118630 -9948 119131 4 VSS
port 42 nsew
rlabel pwell s -12017 118274 -11886 118855 4 VSS
port 42 nsew
rlabel pwell s -10570 119273 -10439 119854 4 VSS
port 42 nsew
rlabel pwell s -12868 119107 -12734 119906 4 VSS
port 42 nsew
<< properties >>
string FIXED_BBOX -34505 -65703 98798 121313
string LEFclass BLOCK
string LEFview TRUE
string GDS_FILE ../gds/sky130_aa_ip__programmable_pll.gds.gz
string GDS_START 0
<< end >>
