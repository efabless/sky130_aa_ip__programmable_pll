magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect 1193 1383 1220 1391
<< pwell >>
rect 2254 1774 2585 2060
<< psubdiff >>
rect 2280 1800 2559 2034
<< locali >>
rect -278 2068 571 2121
rect -278 504 -225 2068
rect 494 2027 571 2068
rect 507 1971 546 2027
rect 2280 1993 2559 2034
rect 2280 1991 2471 1993
rect 2280 1957 2328 1991
rect 2362 1959 2471 1991
rect 2505 1959 2559 1993
rect 2362 1957 2559 1959
rect 2280 1878 2559 1957
rect 2280 1867 2477 1878
rect 2280 1833 2327 1867
rect 2361 1844 2477 1867
rect 2511 1844 2559 1878
rect 2361 1833 2559 1844
rect 2280 1800 2559 1833
rect 978 1436 1038 1449
rect 978 1402 991 1436
rect 1025 1402 1038 1436
rect 2463 1410 2721 1449
rect 978 1390 1038 1402
rect 407 849 895 1065
rect -278 465 6 504
rect 2476 465 2730 504
rect -278 451 -54 465
rect 2245 119 2415 121
rect 2224 89 2559 119
rect 2224 76 2476 89
rect 2224 42 2311 76
rect 2345 55 2476 76
rect 2510 55 2559 89
rect 2345 42 2559 55
rect 2224 -46 2559 42
rect 2224 -53 2444 -46
rect 2224 -87 2300 -53
rect 2334 -80 2444 -53
rect 2478 -80 2559 -46
rect 2334 -87 2559 -80
rect 2224 -138 2559 -87
<< viali >>
rect 2328 1957 2362 1991
rect 2471 1959 2505 1993
rect 2327 1833 2361 1867
rect 2477 1844 2511 1878
rect 991 1402 1025 1436
rect 2311 42 2345 76
rect 2476 55 2510 89
rect 2300 -87 2334 -53
rect 2444 -80 2478 -46
<< metal1 >>
rect -539 2236 917 2342
rect 811 1961 917 2236
rect 2269 1993 2695 2034
rect 2269 1991 2471 1993
rect 2269 1957 2328 1991
rect 2362 1959 2471 1991
rect 2505 1959 2695 1993
rect 2362 1957 2695 1959
rect 2269 1878 2695 1957
rect 2269 1867 2477 1878
rect 2269 1833 2327 1867
rect 2361 1844 2477 1867
rect 2511 1844 2695 1878
rect 2361 1833 2695 1844
rect 2269 1798 2695 1833
rect 959 1445 1050 1459
rect 959 1393 982 1445
rect 1034 1393 1050 1445
rect 959 1380 1050 1393
rect 1159 1391 1254 1425
rect 1193 1383 1254 1391
rect -129 1218 89 1295
rect -129 -166 -52 1218
rect 1220 979 1254 1383
rect 968 933 1254 979
rect 968 738 1014 933
rect 1098 522 1178 526
rect 1098 470 1112 522
rect 1164 470 1178 522
rect 1098 467 1178 470
rect 2521 115 2695 1798
rect 2254 89 2695 115
rect 2254 76 2476 89
rect 480 -166 572 -112
rect -129 -243 572 -166
rect 811 -368 917 44
rect 2254 42 2311 76
rect 2345 55 2476 76
rect 2510 55 2695 89
rect 2345 42 2695 55
rect 2254 -35 2695 42
rect 2254 -46 2559 -35
rect 2254 -53 2444 -46
rect 2254 -87 2300 -53
rect 2334 -80 2444 -53
rect 2478 -80 2559 -46
rect 2334 -87 2559 -80
rect 2254 -119 2559 -87
rect -539 -474 917 -368
<< via1 >>
rect 982 1436 1034 1445
rect 982 1402 991 1436
rect 991 1402 1025 1436
rect 1025 1402 1034 1436
rect 982 1393 1034 1402
rect 1112 470 1164 522
<< metal2 >>
rect 959 1445 1178 1459
rect 959 1393 982 1445
rect 1034 1393 1178 1445
rect 959 1380 1178 1393
rect 1095 522 1178 1380
rect 1095 470 1112 522
rect 1164 470 1178 522
rect 1095 457 1178 470
use PFD_UP  PFD_UP_0
timestamp 1726359333
transform 1 0 373 0 1 457
box -506 -610 2335 500
use PFD_UP  PFD_UP_1
timestamp 1726359333
transform 1 0 373 0 -1 1457
box -506 -610 2335 500
<< labels >>
flabel metal1 s -450 2298 -450 2298 0 FreeSans 1000 0 0 0 FIN
flabel metal1 s -450 -421 -450 -421 0 FreeSans 1000 0 0 0 FDIV
flabel locali s 2605 1430 2605 1430 0 FreeSans 1000 0 0 0 UP
flabel locali s 2668 482 2668 482 0 FreeSans 1000 0 0 0 DOWN
flabel metal1 s 2539 -101 2539 -101 0 FreeSans 1000 0 0 0 VSS
flabel locali s 702 931 702 931 0 FreeSans 1000 0 0 0 VDD
<< end >>
