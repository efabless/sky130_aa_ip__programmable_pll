magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect -114 -412 114 412
<< pmos >>
rect -20 -350 20 350
<< pdiff >>
rect -78 323 -20 350
rect -78 289 -66 323
rect -32 289 -20 323
rect -78 255 -20 289
rect -78 221 -66 255
rect -32 221 -20 255
rect -78 187 -20 221
rect -78 153 -66 187
rect -32 153 -20 187
rect -78 119 -20 153
rect -78 85 -66 119
rect -32 85 -20 119
rect -78 51 -20 85
rect -78 17 -66 51
rect -32 17 -20 51
rect -78 -17 -20 17
rect -78 -51 -66 -17
rect -32 -51 -20 -17
rect -78 -85 -20 -51
rect -78 -119 -66 -85
rect -32 -119 -20 -85
rect -78 -153 -20 -119
rect -78 -187 -66 -153
rect -32 -187 -20 -153
rect -78 -221 -20 -187
rect -78 -255 -66 -221
rect -32 -255 -20 -221
rect -78 -289 -20 -255
rect -78 -323 -66 -289
rect -32 -323 -20 -289
rect -78 -350 -20 -323
rect 20 323 78 350
rect 20 289 32 323
rect 66 289 78 323
rect 20 255 78 289
rect 20 221 32 255
rect 66 221 78 255
rect 20 187 78 221
rect 20 153 32 187
rect 66 153 78 187
rect 20 119 78 153
rect 20 85 32 119
rect 66 85 78 119
rect 20 51 78 85
rect 20 17 32 51
rect 66 17 78 51
rect 20 -17 78 17
rect 20 -51 32 -17
rect 66 -51 78 -17
rect 20 -85 78 -51
rect 20 -119 32 -85
rect 66 -119 78 -85
rect 20 -153 78 -119
rect 20 -187 32 -153
rect 66 -187 78 -153
rect 20 -221 78 -187
rect 20 -255 32 -221
rect 66 -255 78 -221
rect 20 -289 78 -255
rect 20 -323 32 -289
rect 66 -323 78 -289
rect 20 -350 78 -323
<< pdiffc >>
rect -66 289 -32 323
rect -66 221 -32 255
rect -66 153 -32 187
rect -66 85 -32 119
rect -66 17 -32 51
rect -66 -51 -32 -17
rect -66 -119 -32 -85
rect -66 -187 -32 -153
rect -66 -255 -32 -221
rect -66 -323 -32 -289
rect 32 289 66 323
rect 32 221 66 255
rect 32 153 66 187
rect 32 85 66 119
rect 32 17 66 51
rect 32 -51 66 -17
rect 32 -119 66 -85
rect 32 -187 66 -153
rect 32 -255 66 -221
rect 32 -323 66 -289
<< poly >>
rect -20 350 20 376
rect -20 -376 20 -350
<< locali >>
rect -66 323 -32 354
rect -66 255 -32 271
rect -66 187 -32 199
rect -66 119 -32 127
rect -66 51 -32 55
rect -66 -55 -32 -51
rect -66 -127 -32 -119
rect -66 -199 -32 -187
rect -66 -271 -32 -255
rect -66 -354 -32 -323
rect 32 323 66 354
rect 32 255 66 271
rect 32 187 66 199
rect 32 119 66 127
rect 32 51 66 55
rect 32 -55 66 -51
rect 32 -127 66 -119
rect 32 -199 66 -187
rect 32 -271 66 -255
rect 32 -354 66 -323
<< viali >>
rect -66 289 -32 305
rect -66 271 -32 289
rect -66 221 -32 233
rect -66 199 -32 221
rect -66 153 -32 161
rect -66 127 -32 153
rect -66 85 -32 89
rect -66 55 -32 85
rect -66 -17 -32 17
rect -66 -85 -32 -55
rect -66 -89 -32 -85
rect -66 -153 -32 -127
rect -66 -161 -32 -153
rect -66 -221 -32 -199
rect -66 -233 -32 -221
rect -66 -289 -32 -271
rect -66 -305 -32 -289
rect 32 289 66 305
rect 32 271 66 289
rect 32 221 66 233
rect 32 199 66 221
rect 32 153 66 161
rect 32 127 66 153
rect 32 85 66 89
rect 32 55 66 85
rect 32 -17 66 17
rect 32 -85 66 -55
rect 32 -89 66 -85
rect 32 -153 66 -127
rect 32 -161 66 -153
rect 32 -221 66 -199
rect 32 -233 66 -221
rect 32 -289 66 -271
rect 32 -305 66 -289
<< metal1 >>
rect -72 305 -26 350
rect -72 271 -66 305
rect -32 271 -26 305
rect -72 233 -26 271
rect -72 199 -66 233
rect -32 199 -26 233
rect -72 161 -26 199
rect -72 127 -66 161
rect -32 127 -26 161
rect -72 89 -26 127
rect -72 55 -66 89
rect -32 55 -26 89
rect -72 17 -26 55
rect -72 -17 -66 17
rect -32 -17 -26 17
rect -72 -55 -26 -17
rect -72 -89 -66 -55
rect -32 -89 -26 -55
rect -72 -127 -26 -89
rect -72 -161 -66 -127
rect -32 -161 -26 -127
rect -72 -199 -26 -161
rect -72 -233 -66 -199
rect -32 -233 -26 -199
rect -72 -271 -26 -233
rect -72 -305 -66 -271
rect -32 -305 -26 -271
rect -72 -350 -26 -305
rect 26 305 72 350
rect 26 271 32 305
rect 66 271 72 305
rect 26 233 72 271
rect 26 199 32 233
rect 66 199 72 233
rect 26 161 72 199
rect 26 127 32 161
rect 66 127 72 161
rect 26 89 72 127
rect 26 55 32 89
rect 66 55 72 89
rect 26 17 72 55
rect 26 -17 32 17
rect 66 -17 72 17
rect 26 -55 72 -17
rect 26 -89 32 -55
rect 66 -89 72 -55
rect 26 -127 72 -89
rect 26 -161 32 -127
rect 66 -161 72 -127
rect 26 -199 72 -161
rect 26 -233 32 -199
rect 66 -233 72 -199
rect 26 -271 72 -233
rect 26 -305 32 -271
rect 66 -305 72 -271
rect 26 -350 72 -305
<< end >>
