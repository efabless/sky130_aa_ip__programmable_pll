magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect 2439 4146 2529 4215
rect 2702 4128 2765 4226
rect 2839 4142 2977 4209
rect 4518 4038 7244 4246
rect 4566 3976 4600 4038
rect 4762 3976 4796 4038
rect 4839 3214 5543 4038
rect 5566 3976 5600 4038
rect 5762 3976 5796 4038
rect 5823 3214 5933 4038
rect 5966 3976 6000 4038
rect 6162 3976 6196 4038
rect 6229 3214 6537 4038
rect 6566 3976 6600 4038
rect 6762 3976 7199 4038
rect 6794 3214 7199 3976
rect 3677 2133 4209 2254
rect -79 1532 2237 1985
rect 3677 1981 4210 2133
rect 3677 1980 4209 1981
rect 3743 1968 3988 1980
<< pwell >>
rect 4443 2151 7222 2300
<< psubdiff >>
rect 4469 2242 7196 2274
rect 4469 2208 4509 2242
rect 4543 2208 4577 2242
rect 4611 2208 4645 2242
rect 4679 2208 4713 2242
rect 4747 2208 4781 2242
rect 4815 2208 4849 2242
rect 4883 2208 4917 2242
rect 4951 2208 4985 2242
rect 5019 2208 5053 2242
rect 5087 2208 5121 2242
rect 5155 2208 5459 2242
rect 5493 2208 5527 2242
rect 5561 2208 5595 2242
rect 5629 2208 5663 2242
rect 5697 2208 5731 2242
rect 5765 2208 5799 2242
rect 5833 2208 5867 2242
rect 5901 2208 5935 2242
rect 5969 2208 6003 2242
rect 6037 2208 6071 2242
rect 6105 2208 6409 2242
rect 6443 2208 6477 2242
rect 6511 2208 6545 2242
rect 6579 2208 6613 2242
rect 6647 2208 6681 2242
rect 6715 2208 6749 2242
rect 6783 2208 6817 2242
rect 6851 2208 6885 2242
rect 6919 2208 6953 2242
rect 6987 2208 7021 2242
rect 7055 2208 7196 2242
rect 4469 2177 7196 2208
<< nsubdiff >>
rect 4556 4173 7208 4210
rect 4556 4139 4614 4173
rect 4648 4139 4682 4173
rect 4716 4139 4750 4173
rect 4784 4139 4818 4173
rect 4852 4139 4886 4173
rect 4920 4139 4954 4173
rect 4988 4139 5022 4173
rect 5056 4139 5090 4173
rect 5124 4139 5158 4173
rect 5192 4139 5226 4173
rect 5260 4139 5514 4173
rect 5548 4139 5582 4173
rect 5616 4139 5650 4173
rect 5684 4139 5718 4173
rect 5752 4139 5786 4173
rect 5820 4139 5854 4173
rect 5888 4139 5922 4173
rect 5956 4139 5990 4173
rect 6024 4139 6058 4173
rect 6092 4139 6126 4173
rect 6160 4139 6414 4173
rect 6448 4139 6482 4173
rect 6516 4139 6550 4173
rect 6584 4139 6618 4173
rect 6652 4139 6686 4173
rect 6720 4139 6754 4173
rect 6788 4139 6822 4173
rect 6856 4139 6890 4173
rect 6924 4139 6958 4173
rect 6992 4139 7026 4173
rect 7060 4139 7208 4173
rect 4556 4107 7208 4139
<< psubdiffcont >>
rect 4509 2208 4543 2242
rect 4577 2208 4611 2242
rect 4645 2208 4679 2242
rect 4713 2208 4747 2242
rect 4781 2208 4815 2242
rect 4849 2208 4883 2242
rect 4917 2208 4951 2242
rect 4985 2208 5019 2242
rect 5053 2208 5087 2242
rect 5121 2208 5155 2242
rect 5459 2208 5493 2242
rect 5527 2208 5561 2242
rect 5595 2208 5629 2242
rect 5663 2208 5697 2242
rect 5731 2208 5765 2242
rect 5799 2208 5833 2242
rect 5867 2208 5901 2242
rect 5935 2208 5969 2242
rect 6003 2208 6037 2242
rect 6071 2208 6105 2242
rect 6409 2208 6443 2242
rect 6477 2208 6511 2242
rect 6545 2208 6579 2242
rect 6613 2208 6647 2242
rect 6681 2208 6715 2242
rect 6749 2208 6783 2242
rect 6817 2208 6851 2242
rect 6885 2208 6919 2242
rect 6953 2208 6987 2242
rect 7021 2208 7055 2242
<< nsubdiffcont >>
rect 4614 4139 4648 4173
rect 4682 4139 4716 4173
rect 4750 4139 4784 4173
rect 4818 4139 4852 4173
rect 4886 4139 4920 4173
rect 4954 4139 4988 4173
rect 5022 4139 5056 4173
rect 5090 4139 5124 4173
rect 5158 4139 5192 4173
rect 5226 4139 5260 4173
rect 5514 4139 5548 4173
rect 5582 4139 5616 4173
rect 5650 4139 5684 4173
rect 5718 4139 5752 4173
rect 5786 4139 5820 4173
rect 5854 4139 5888 4173
rect 5922 4139 5956 4173
rect 5990 4139 6024 4173
rect 6058 4139 6092 4173
rect 6126 4139 6160 4173
rect 6414 4139 6448 4173
rect 6482 4139 6516 4173
rect 6550 4139 6584 4173
rect 6618 4139 6652 4173
rect 6686 4139 6720 4173
rect 6754 4139 6788 4173
rect 6822 4139 6856 4173
rect 6890 4139 6924 4173
rect 6958 4139 6992 4173
rect 7026 4139 7060 4173
<< poly >>
rect 4612 3259 4638 3262
rect 4612 3250 4652 3259
rect 5012 3250 5052 3276
rect 5110 3250 5150 3276
rect 4612 3214 4750 3250
rect 5012 3214 5150 3250
rect 5612 3252 5638 3262
rect 5612 3250 5652 3252
rect 6012 3250 6052 3276
rect 6110 3250 6150 3276
rect 5612 3214 5750 3250
rect 6012 3214 6150 3250
rect 6612 3250 6652 3276
rect 6710 3250 6750 3276
rect 6612 3214 6750 3250
rect 7012 3250 7052 3276
rect 7110 3250 7150 3276
rect 7012 3214 7150 3250
rect 4612 3207 4652 3214
rect 4494 3197 4652 3207
rect 4494 3163 4510 3197
rect 4544 3163 4578 3197
rect 4612 3163 4652 3197
rect 5012 3192 5052 3214
rect 5612 3205 5652 3214
rect 6012 3207 6052 3214
rect 6612 3212 6652 3214
rect 4494 3153 4652 3163
rect 4612 3091 4652 3153
rect 4896 3182 5052 3192
rect 4896 3148 4912 3182
rect 4946 3148 4980 3182
rect 5014 3148 5052 3182
rect 5483 3195 5652 3205
rect 5483 3161 5499 3195
rect 5533 3161 5567 3195
rect 5601 3161 5652 3195
rect 5483 3151 5652 3161
rect 5896 3197 6052 3207
rect 5896 3163 5912 3197
rect 5946 3163 5980 3197
rect 6014 3163 6052 3197
rect 5896 3153 6052 3163
rect 6483 3202 6652 3212
rect 7012 3209 7052 3214
rect 6483 3168 6499 3202
rect 6533 3168 6567 3202
rect 6601 3168 6652 3202
rect 6483 3158 6652 3168
rect 4896 3138 5052 3148
rect 5012 3091 5052 3138
rect 5612 3091 5652 3151
rect 6012 3091 6052 3153
rect 6612 3091 6652 3158
rect 6889 3199 7052 3209
rect 6889 3165 6905 3199
rect 6939 3165 6973 3199
rect 7007 3165 7052 3199
rect 6889 3155 7052 3165
rect 7012 3091 7052 3155
<< polycont >>
rect 4510 3163 4544 3197
rect 4578 3163 4612 3197
rect 4912 3148 4946 3182
rect 4980 3148 5014 3182
rect 5499 3161 5533 3195
rect 5567 3161 5601 3195
rect 5912 3163 5946 3197
rect 5980 3163 6014 3197
rect 6499 3168 6533 3202
rect 6567 3168 6601 3202
rect 6905 3165 6939 3199
rect 6973 3165 7007 3199
<< locali >>
rect 1582 4215 1668 4219
rect 2702 4215 2765 4226
rect 1582 4203 1970 4215
rect 491 4134 938 4203
rect 1407 4146 1970 4203
rect 2439 4209 2765 4215
rect 3383 4209 3457 4215
rect 2439 4146 2977 4209
rect 1407 4134 1668 4146
rect 1582 4126 1668 4134
rect 2702 4142 2977 4146
rect 3178 4202 3457 4209
rect 3178 4142 3700 4202
rect 2702 4128 2765 4142
rect 3383 4134 3700 4142
rect 4100 4173 7389 4210
rect 4100 4139 4614 4173
rect 4648 4139 4682 4173
rect 4716 4139 4750 4173
rect 4784 4139 4818 4173
rect 4852 4139 4886 4173
rect 4920 4139 4954 4173
rect 4988 4139 5022 4173
rect 5056 4139 5090 4173
rect 5124 4139 5158 4173
rect 5192 4139 5226 4173
rect 5260 4139 5514 4173
rect 5548 4139 5582 4173
rect 5616 4139 5650 4173
rect 5684 4139 5718 4173
rect 5752 4139 5786 4173
rect 5820 4139 5854 4173
rect 5888 4139 5922 4173
rect 5956 4139 5990 4173
rect 6024 4139 6058 4173
rect 6092 4139 6126 4173
rect 6160 4139 6414 4173
rect 6448 4139 6482 4173
rect 6516 4139 6550 4173
rect 6584 4139 6618 4173
rect 6652 4139 6686 4173
rect 6720 4139 6754 4173
rect 6788 4139 6822 4173
rect 6856 4139 6890 4173
rect 6924 4139 6958 4173
rect 6992 4139 7026 4173
rect 7060 4139 7389 4173
rect 3383 4128 3457 4134
rect 4100 4107 7389 4139
rect 4566 3976 4600 4107
rect 4762 3976 4796 4107
rect 4966 3976 5000 4107
rect 5162 3976 5196 4107
rect 5566 3976 5600 4107
rect 5762 3976 5796 4107
rect 5966 3976 6000 4107
rect 6162 3976 6196 4107
rect 6566 3976 6600 4107
rect 6762 3976 6796 4107
rect 6966 3976 7000 4107
rect 7162 3976 7196 4107
rect 1618 3891 1678 3898
rect 1618 3857 1631 3891
rect 1665 3857 1678 3891
rect 1618 3813 1678 3857
rect 1618 3779 1631 3813
rect 1665 3801 1678 3813
rect 1665 3779 1766 3801
rect 1618 3766 1766 3779
rect 3574 3752 3706 3765
rect 1503 3682 1777 3720
rect 3574 3718 3581 3752
rect 3615 3718 3659 3752
rect 3693 3718 3706 3752
rect 3574 3705 3706 3718
rect 4176 3716 4469 3786
rect 1503 3641 1563 3682
rect 1503 3607 1516 3641
rect 1550 3607 1563 3641
rect 1503 3563 1563 3607
rect 1503 3529 1516 3563
rect 1550 3529 1563 3563
rect 1503 3516 1563 3529
rect -140 3464 -37 3500
rect 1138 3494 1270 3507
rect 1138 3460 1145 3494
rect 1179 3460 1223 3494
rect 1257 3460 1270 3494
rect 1138 3447 1270 3460
rect 467 3420 599 3433
rect -140 3375 -54 3411
rect 467 3386 474 3420
rect 508 3386 552 3420
rect 586 3386 599 3420
rect 467 3373 599 3386
rect 915 3414 1047 3427
rect 1738 3417 1772 3638
rect 3201 3582 3332 3595
rect 3201 3571 3208 3582
rect 3055 3548 3208 3571
rect 3242 3548 3286 3582
rect 3320 3548 3332 3582
rect 3055 3535 3332 3548
rect 3677 3469 4342 3512
rect 915 3380 922 3414
rect 956 3380 1000 3414
rect 1034 3380 1047 3414
rect 1483 3413 1772 3417
rect 915 3367 1047 3380
rect 1479 3379 1772 3413
rect 1483 3372 1772 3379
rect 3293 3311 4342 3469
rect 521 2932 904 3021
rect -242 922 -100 963
rect -251 833 -103 874
rect 816 795 948 808
rect -245 741 -109 782
rect 816 761 823 795
rect 857 761 901 795
rect 935 761 948 795
rect 816 748 948 761
rect 984 397 1133 2979
rect 1448 2932 1953 3021
rect 3293 3005 3374 3311
rect 1779 2889 1953 2932
rect 3059 2970 3374 3005
rect 3059 2889 3375 2970
rect 3561 2950 3720 2951
rect 3561 2939 3721 2950
rect 3561 2905 3574 2939
rect 3608 2905 3674 2939
rect 3708 2905 3721 2939
rect 3561 2892 3721 2905
rect 4174 2925 4234 2933
rect 3561 2891 3720 2892
rect 4174 2891 4187 2925
rect 4221 2891 4234 2925
rect 3208 2837 3340 2850
rect 3208 2803 3215 2837
rect 3249 2803 3293 2837
rect 3327 2836 3340 2837
rect 4174 2847 4234 2891
rect 3327 2803 3667 2836
rect 3208 2800 3667 2803
rect 4174 2813 4187 2847
rect 4221 2813 4234 2847
rect 3208 2790 3340 2800
rect 4174 2799 4234 2813
rect 3311 2460 3471 2467
rect 3311 2426 3324 2460
rect 3358 2426 3424 2460
rect 3458 2426 3471 2460
rect 3311 2382 3471 2426
rect 3311 2348 3324 2382
rect 3358 2348 3424 2382
rect 3458 2348 3471 2382
rect 3311 2335 3471 2348
rect 3321 2152 3456 2335
rect 4272 2274 4342 3311
rect 4399 3207 4469 3716
rect 4399 3197 4628 3207
rect 4399 3163 4510 3197
rect 4544 3163 4578 3197
rect 4612 3163 4628 3197
rect 4399 3153 4628 3163
rect 4664 3185 4698 3279
rect 4896 3185 5030 3192
rect 4664 3182 5030 3185
rect 4399 2531 4469 3153
rect 4664 3151 4912 3182
rect 4664 3093 4698 3151
rect 4896 3148 4912 3151
rect 4946 3148 4980 3182
rect 5014 3148 5030 3182
rect 4896 3138 5030 3148
rect 5064 3175 5098 3277
rect 5443 3195 5617 3205
rect 5172 3175 5290 3187
rect 5064 3141 5178 3175
rect 5212 3141 5250 3175
rect 5284 3141 5290 3175
rect 5064 3091 5098 3141
rect 5172 3129 5290 3141
rect 5443 3161 5499 3195
rect 5533 3161 5567 3195
rect 5601 3161 5617 3195
rect 5443 3151 5617 3161
rect 5664 3200 5698 3300
rect 5896 3200 6030 3207
rect 5664 3197 6030 3200
rect 5664 3163 5912 3197
rect 5946 3163 5980 3197
rect 6014 3163 6030 3197
rect 5664 3161 6030 3163
rect 5443 3082 5513 3151
rect 5664 3091 5698 3161
rect 5896 3153 6030 3161
rect 6064 3202 6098 3300
rect 6249 3202 6367 3214
rect 6064 3168 6255 3202
rect 6289 3168 6327 3202
rect 6361 3168 6367 3202
rect 6064 3091 6098 3168
rect 6249 3156 6367 3168
rect 6434 3202 6617 3212
rect 6434 3168 6499 3202
rect 6533 3168 6567 3202
rect 6601 3168 6617 3202
rect 6434 3158 6617 3168
rect 6664 3201 6698 3300
rect 6889 3201 7023 3209
rect 6664 3199 7023 3201
rect 6664 3165 6905 3199
rect 6939 3165 6973 3199
rect 7007 3165 7023 3199
rect 6664 3162 7023 3165
rect 5443 3048 5463 3082
rect 5497 3048 5513 3082
rect 5443 3010 5513 3048
rect 5443 2976 5463 3010
rect 5497 2976 5513 3010
rect 5443 2970 5513 2976
rect 6434 3083 6504 3158
rect 6664 3091 6698 3162
rect 6889 3155 7023 3162
rect 7064 3186 7098 3300
rect 7145 3190 7263 3202
rect 7145 3186 7151 3190
rect 7064 3156 7151 3186
rect 7185 3156 7223 3190
rect 7257 3186 7263 3190
rect 7257 3156 7266 3186
rect 7064 3152 7266 3156
rect 7064 3091 7098 3152
rect 7145 3144 7263 3152
rect 6434 3049 6450 3083
rect 6484 3049 6504 3083
rect 6434 3011 6504 3049
rect 6434 2977 6450 3011
rect 6484 2977 6504 3011
rect 6434 2971 6504 2977
rect 4399 2497 4418 2531
rect 4452 2497 4469 2531
rect 4399 2459 4469 2497
rect 4399 2425 4418 2459
rect 4452 2425 4469 2459
rect 4399 2419 4469 2425
rect 4566 2274 4600 2389
rect 4966 2274 5000 2387
rect 5566 2274 5600 2387
rect 5966 2274 6000 2387
rect 6566 2274 6600 2387
rect 6966 2274 7000 2388
rect 4272 2242 7196 2274
rect 4272 2208 4509 2242
rect 4543 2208 4577 2242
rect 4611 2208 4645 2242
rect 4679 2208 4713 2242
rect 4747 2208 4781 2242
rect 4815 2208 4849 2242
rect 4883 2208 4917 2242
rect 4951 2208 4985 2242
rect 5019 2208 5053 2242
rect 5087 2208 5121 2242
rect 5155 2208 5459 2242
rect 5493 2208 5527 2242
rect 5561 2208 5595 2242
rect 5629 2208 5663 2242
rect 5697 2208 5731 2242
rect 5765 2208 5799 2242
rect 5833 2208 5867 2242
rect 5901 2208 5935 2242
rect 5969 2208 6003 2242
rect 6037 2208 6071 2242
rect 6105 2208 6409 2242
rect 6443 2208 6477 2242
rect 6511 2208 6545 2242
rect 6579 2208 6613 2242
rect 6647 2208 6681 2242
rect 6715 2208 6749 2242
rect 6783 2208 6817 2242
rect 6851 2208 6885 2242
rect 6919 2208 6953 2242
rect 6987 2208 7021 2242
rect 7055 2208 7196 2242
rect 3314 2145 3474 2152
rect 3314 2111 3327 2145
rect 3361 2111 3427 2145
rect 3461 2111 3474 2145
rect 3314 2067 3474 2111
rect 3314 2033 3327 2067
rect 3361 2033 3427 2067
rect 3461 2033 3474 2067
rect 3314 2020 3474 2033
rect 3784 1905 4016 2199
rect 4272 2177 7196 2208
rect 7300 1733 7389 4107
rect 1199 1058 1238 1349
rect 1199 684 1305 1058
rect 1199 671 1331 684
rect 1199 637 1206 671
rect 1240 637 1284 671
rect 1318 637 1331 671
rect 1199 596 1331 637
rect 1199 562 1206 596
rect 1240 562 1284 596
rect 1318 562 1331 596
rect 1199 549 1331 562
rect 1545 397 1729 964
rect 798 291 1729 397
<< viali >>
rect 1631 3857 1665 3891
rect 1631 3779 1665 3813
rect 3581 3718 3615 3752
rect 3659 3718 3693 3752
rect 1516 3607 1550 3641
rect 1516 3529 1550 3563
rect 1145 3460 1179 3494
rect 1223 3460 1257 3494
rect 474 3386 508 3420
rect 552 3386 586 3420
rect 3208 3548 3242 3582
rect 3286 3548 3320 3582
rect 922 3380 956 3414
rect 1000 3380 1034 3414
rect 823 761 857 795
rect 901 761 935 795
rect 3574 2905 3608 2939
rect 3674 2905 3708 2939
rect 4187 2891 4221 2925
rect 3215 2803 3249 2837
rect 3293 2803 3327 2837
rect 4187 2813 4221 2847
rect 3324 2426 3358 2460
rect 3424 2426 3458 2460
rect 3324 2348 3358 2382
rect 3424 2348 3458 2382
rect 5178 3141 5212 3175
rect 5250 3141 5284 3175
rect 6255 3168 6289 3202
rect 6327 3168 6361 3202
rect 5463 3048 5497 3082
rect 5463 2976 5497 3010
rect 7151 3156 7185 3190
rect 7223 3156 7257 3190
rect 6450 3049 6484 3083
rect 6450 2977 6484 3011
rect 4418 2497 4452 2531
rect 4418 2425 4452 2459
rect 3327 2111 3361 2145
rect 3427 2111 3461 2145
rect 3327 2033 3361 2067
rect 3427 2033 3461 2067
rect 1206 637 1240 671
rect 1284 637 1318 671
rect 1206 562 1240 596
rect 1284 562 1318 596
<< metal1 >>
rect 5345 4076 7475 4110
rect 1618 3891 1678 3898
rect 1618 3857 1631 3891
rect 1665 3857 1678 3891
rect 1618 3813 1678 3857
rect 1618 3779 1631 3813
rect 1665 3779 1678 3813
rect 1618 3766 1678 3779
rect 1503 3641 1563 3648
rect 1503 3607 1516 3641
rect 1550 3607 1563 3641
rect 1503 3588 1563 3607
rect 554 3563 1563 3588
rect 554 3546 1516 3563
rect 554 3433 596 3546
rect 1503 3529 1516 3546
rect 1550 3529 1563 3563
rect 1503 3516 1563 3529
rect 1138 3500 1270 3507
rect 709 3494 1270 3500
rect 709 3460 1145 3494
rect 1179 3460 1223 3494
rect 1257 3460 1270 3494
rect 709 3458 1270 3460
rect 467 3420 599 3433
rect 467 3386 474 3420
rect 508 3386 552 3420
rect 586 3386 599 3420
rect 467 3373 599 3386
rect 709 2887 751 3458
rect 1138 3447 1270 3458
rect 915 3416 1047 3427
rect -201 2845 751 2887
rect 799 3414 1047 3416
rect 799 3380 922 3414
rect 956 3380 1000 3414
rect 1034 3380 1047 3414
rect 799 3374 1047 3380
rect 799 2813 841 3374
rect 915 3367 1047 3374
rect 1626 2884 1668 3766
rect 3379 3752 3706 3765
rect 3379 3718 3581 3752
rect 3615 3718 3659 3752
rect 3693 3718 3706 3752
rect 3379 3705 3706 3718
rect 3201 3582 3332 3595
rect 3201 3548 3208 3582
rect 3242 3548 3286 3582
rect 3320 3548 3332 3582
rect 3201 3535 3332 3548
rect -196 2771 841 2813
rect 898 2842 1668 2884
rect 3240 2850 3300 3535
rect 3379 2951 3439 3705
rect 5172 3175 5290 3187
rect 5345 3175 5379 4076
rect 6255 4011 7479 4045
rect 6255 3214 6289 4011
rect 5172 3141 5178 3175
rect 5212 3141 5250 3175
rect 5284 3141 5379 3175
rect 6249 3202 6367 3214
rect 6249 3168 6255 3202
rect 6289 3168 6327 3202
rect 6361 3168 6367 3202
rect 6249 3156 6367 3168
rect 7145 3193 7263 3202
rect 7145 3190 7480 3193
rect 7145 3156 7151 3190
rect 7185 3156 7223 3190
rect 7257 3156 7480 3190
rect 7145 3148 7480 3156
rect 7145 3144 7263 3148
rect 5172 3129 5290 3141
rect 5443 3082 5513 3088
rect 5443 3048 5463 3082
rect 5497 3048 5513 3082
rect 5443 3010 5513 3048
rect 5443 2976 5463 3010
rect 5497 2976 5513 3010
rect 3379 2950 3720 2951
rect 3379 2939 3721 2950
rect 3379 2905 3574 2939
rect 3608 2905 3674 2939
rect 3708 2905 3721 2939
rect 3379 2892 3721 2905
rect 4174 2925 4260 2933
rect 3379 2891 3720 2892
rect 4174 2891 4187 2925
rect 4221 2891 4260 2925
rect 898 808 940 2842
rect 3208 2837 3340 2850
rect 3208 2803 3215 2837
rect 3249 2803 3293 2837
rect 3327 2803 3340 2837
rect 3208 2790 3340 2803
rect 3379 2467 3439 2891
rect 4174 2847 4260 2891
rect 4174 2813 4187 2847
rect 4221 2813 4260 2847
rect 4174 2799 4260 2813
rect 3311 2460 3471 2467
rect 3311 2426 3324 2460
rect 3358 2426 3424 2460
rect 3458 2426 3471 2460
rect 3311 2382 3471 2426
rect 3311 2348 3324 2382
rect 3358 2348 3424 2382
rect 3458 2348 3471 2382
rect 3311 2335 3471 2348
rect 4203 2277 4260 2799
rect 4399 2531 4469 2537
rect 4399 2497 4418 2531
rect 4452 2497 4469 2531
rect 4399 2459 4469 2497
rect 4399 2425 4418 2459
rect 4452 2425 4469 2459
rect 4399 2358 4469 2425
rect 5443 2358 5513 2976
rect 6434 3083 6504 3089
rect 6434 3049 6450 3083
rect 6484 3049 6504 3083
rect 6434 3011 6504 3049
rect 6434 2977 6450 3011
rect 6484 2977 6504 3011
rect 6434 2358 6504 2977
rect 4399 2288 7549 2358
rect 988 2220 4260 2277
rect 988 869 1045 2220
rect 3314 2145 3474 2152
rect 3314 2111 3327 2145
rect 3361 2111 3427 2145
rect 3461 2111 3474 2145
rect 3314 2067 3474 2111
rect 3314 2033 3327 2067
rect 3361 2033 3427 2067
rect 3461 2061 3474 2067
rect 3461 2033 7346 2061
rect 3314 1971 7346 2033
rect 7256 1037 7346 1971
rect 988 812 1255 869
rect 816 795 948 808
rect 816 761 823 795
rect 857 761 901 795
rect 935 761 948 795
rect 816 748 948 761
rect 898 744 940 748
rect 1199 671 1331 684
rect 1199 637 1206 671
rect 1240 637 1284 671
rect 1318 637 1331 671
rect 1199 596 1331 637
rect 1199 562 1206 596
rect 1240 562 1284 596
rect 1318 562 1331 596
rect 1199 549 1331 562
rect 1226 474 1301 549
rect -266 399 1301 474
use 3_INPUT_NOR_MAG  3_INPUT_NOR_MAG_0
timestamp 1726359333
transform 1 0 -74 0 1 1001
box -80 -736 945 956
use 3AND_MAGIC  3AND_MAGIC_0
timestamp 1726359333
transform 1 0 1779 0 1 3792
box -48 -929 1456 459
use DFF_MAG  DFF_MAG_0
timestamp 1726359333
transform 1 0 3809 0 1 1189
box -2665 -1137 3660 829
use inverter  inverter_0
timestamp 1726359333
transform 1 0 3354 0 1 3871
box 220 -453 904 367
use NAND_MAGIC  NAND_MAGIC_0
timestamp 1726359333
transform 1 0 3676 0 -1 2800
box -48 -615 534 667
use NOR_MAGIC  NOR_MAGIC_0
timestamp 1726359333
transform 1 0 863 0 1 3558
box -13 -652 636 681
use NOR_MAGIC  NOR_MAGIC_1
timestamp 1726359333
transform 1 0 -83 0 1 3558
box -13 -652 636 681
use sky130_fd_pr__nfet_01v8_T7BQPS  sky130_fd_pr__nfet_01v8_T7BQPS_0 paramcells
timestamp 1726359333
transform 1 0 7032 0 1 2741
box -104 -376 104 376
use sky130_fd_pr__nfet_01v8_T7BQPS  sky130_fd_pr__nfet_01v8_T7BQPS_1
timestamp 1726359333
transform 1 0 4632 0 1 2741
box -104 -376 104 376
use sky130_fd_pr__nfet_01v8_T7BQPS  sky130_fd_pr__nfet_01v8_T7BQPS_2
timestamp 1726359333
transform 1 0 5032 0 1 2741
box -104 -376 104 376
use sky130_fd_pr__nfet_01v8_T7BQPS  sky130_fd_pr__nfet_01v8_T7BQPS_3
timestamp 1726359333
transform 1 0 6632 0 1 2741
box -104 -376 104 376
use sky130_fd_pr__nfet_01v8_T7BQPS  sky130_fd_pr__nfet_01v8_T7BQPS_4
timestamp 1726359333
transform 1 0 5632 0 1 2741
box -104 -376 104 376
use sky130_fd_pr__nfet_01v8_T7BQPS  sky130_fd_pr__nfet_01v8_T7BQPS_5
timestamp 1726359333
transform 1 0 6032 0 1 2741
box -104 -376 104 376
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_0 paramcells
timestamp 1726359333
transform 1 0 7130 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_1
timestamp 1726359333
transform 1 0 7032 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_2
timestamp 1726359333
transform 1 0 4730 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_3
timestamp 1726359333
transform 1 0 4632 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_4
timestamp 1726359333
transform 1 0 5130 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_5
timestamp 1726359333
transform 1 0 5032 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_6
timestamp 1726359333
transform 1 0 6730 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_7
timestamp 1726359333
transform 1 0 6632 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_8
timestamp 1726359333
transform 1 0 5730 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_9
timestamp 1726359333
transform 1 0 5632 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_10
timestamp 1726359333
transform 1 0 6032 0 1 3626
box -114 -412 114 412
use sky130_fd_pr__pfet_01v8_WNVYTC  sky130_fd_pr__pfet_01v8_WNVYTC_11
timestamp 1726359333
transform 1 0 6130 0 1 3626
box -114 -412 114 412
<< labels >>
flabel locali s -215 847 -215 847 0 FreeSans 1563 0 0 0 Q2
flabel locali s -228 759 -228 759 0 FreeSans 1563 0 0 0 Q3
flabel metal1 s -177 2868 -177 2868 0 FreeSans 1563 0 0 0 Q4
flabel metal1 s -183 2787 -183 2787 0 FreeSans 1563 0 0 0 Q5
flabel locali s -129 3477 -129 3477 0 FreeSans 1563 0 0 0 Q6
flabel locali s -125 3395 -125 3395 0 FreeSans 1563 0 0 0 Q7
flabel metal1 s -245 435 -245 435 0 FreeSans 1563 0 0 0 G_CLK
flabel locali s 4380 4169 4380 4169 0 FreeSans 3125 0 0 0 VDD
flabel locali s 1602 362 1602 362 0 FreeSans 3125 0 0 0 VSS
flabel metal1 s 7488 2319 7488 2319 0 FreeSans 3125 0 0 0 LD
flabel metal1 s 7440 3171 7440 3171 0 FreeSans 3125 0 0 0 LD1
flabel metal1 s 7443 4033 7443 4033 0 FreeSans 3125 0 0 0 LD2
flabel metal1 s 7416 4101 7416 4101 0 FreeSans 3125 0 0 0 LD3
flabel locali s -219 936 -219 936 0 FreeSans 1563 0 0 0 Q1
<< end >>
