magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect -114 -162 114 162
<< pmos >>
rect -20 -100 20 100
<< pdiff >>
rect -78 85 -20 100
rect -78 51 -66 85
rect -32 51 -20 85
rect -78 17 -20 51
rect -78 -17 -66 17
rect -32 -17 -20 17
rect -78 -51 -20 -17
rect -78 -85 -66 -51
rect -32 -85 -20 -51
rect -78 -100 -20 -85
rect 20 85 78 100
rect 20 51 32 85
rect 66 51 78 85
rect 20 17 78 51
rect 20 -17 32 17
rect 66 -17 78 17
rect 20 -51 78 -17
rect 20 -85 32 -51
rect 66 -85 78 -51
rect 20 -100 78 -85
<< pdiffc >>
rect -66 51 -32 85
rect -66 -17 -32 17
rect -66 -85 -32 -51
rect 32 51 66 85
rect 32 -17 66 17
rect 32 -85 66 -51
<< poly >>
rect -20 100 20 126
rect -20 -126 20 -100
<< locali >>
rect -66 85 -32 104
rect -66 17 -32 19
rect -66 -19 -32 -17
rect -66 -104 -32 -85
rect 32 85 66 104
rect 32 17 66 19
rect 32 -19 66 -17
rect 32 -104 66 -85
<< viali >>
rect -66 51 -32 53
rect -66 19 -32 51
rect -66 -51 -32 -19
rect -66 -53 -32 -51
rect 32 51 66 53
rect 32 19 66 51
rect 32 -51 66 -19
rect 32 -53 66 -51
<< metal1 >>
rect -72 53 -26 100
rect -72 19 -66 53
rect -32 19 -26 53
rect -72 -19 -26 19
rect -72 -53 -66 -19
rect -32 -53 -26 -19
rect -72 -100 -26 -53
rect 26 53 72 100
rect 26 19 32 53
rect 66 19 72 53
rect 26 -19 72 19
rect 26 -53 32 -19
rect 66 -53 72 -19
rect 26 -100 72 -53
<< end >>
