magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect 12 416 534 567
rect 12 415 338 416
<< pwell >>
rect 14 -626 515 -513
<< psubdiff >>
rect 40 -553 489 -539
rect 40 -587 77 -553
rect 111 -587 145 -553
rect 179 -587 213 -553
rect 247 -587 281 -553
rect 315 -587 349 -553
rect 383 -587 417 -553
rect 451 -587 489 -553
rect 40 -600 489 -587
<< nsubdiff >>
rect 50 516 492 531
rect 50 482 114 516
rect 148 482 182 516
rect 216 482 250 516
rect 284 482 318 516
rect 352 482 386 516
rect 420 482 492 516
rect 50 467 492 482
<< psubdiffcont >>
rect 77 -587 111 -553
rect 145 -587 179 -553
rect 213 -587 247 -553
rect 281 -587 315 -553
rect 349 -587 383 -553
rect 417 -587 451 -553
<< nsubdiffcont >>
rect 114 482 148 516
rect 182 482 216 516
rect 250 482 284 516
rect 318 482 352 516
rect 386 482 420 516
<< poly >>
rect 106 7 146 28
rect -25 -3 146 7
rect -25 -37 -9 -3
rect 25 -37 60 -3
rect 94 -13 146 -3
rect 204 -13 244 28
rect 94 -37 244 -13
rect -25 -43 244 -37
rect -25 -47 146 -43
rect 106 -174 146 -47
rect 204 -157 244 -43
rect 302 -6 342 28
rect 400 -6 440 28
rect 302 -38 440 -6
rect 302 -157 342 -38
rect 400 -71 440 -38
rect 400 -88 514 -71
rect 400 -122 459 -88
rect 493 -122 514 -88
rect 400 -142 514 -122
rect 400 -157 440 -142
<< polycont >>
rect -9 -37 25 -3
rect 60 -37 94 -3
rect 459 -122 493 -88
<< locali >>
rect 50 516 492 531
rect 50 482 114 516
rect 148 482 182 516
rect 216 482 250 516
rect 284 482 318 516
rect 352 482 386 516
rect 420 482 492 516
rect 50 467 492 482
rect 60 354 94 467
rect 256 354 290 467
rect 452 354 486 467
rect 158 14 192 57
rect 354 14 388 51
rect -25 1 110 7
rect -45 -3 110 1
rect -45 -37 -9 -3
rect 25 -37 60 -3
rect 94 -37 110 -3
rect 158 -24 577 14
rect -45 -39 110 -37
rect -25 -47 110 -39
rect 440 -88 514 -71
rect 440 -97 459 -88
rect 28 -122 459 -97
rect 493 -122 514 -88
rect 28 -136 514 -122
rect 28 -137 99 -136
rect 440 -142 514 -136
rect 157 -539 192 -487
rect 40 -553 489 -539
rect 40 -587 77 -553
rect 111 -587 145 -553
rect 179 -587 213 -553
rect 247 -587 281 -553
rect 315 -587 349 -553
rect 383 -587 417 -553
rect 451 -587 489 -553
rect 40 -600 489 -587
<< metal1 >>
rect 348 -183 394 55
rect 53 -519 100 -482
rect 250 -519 296 -482
rect 446 -519 492 -483
rect 53 -566 492 -519
use sky130_fd_pr__nfet_01v8_FQGQPXv0  sky130_fd_pr__nfet_01v8_FQGQPX_0 paramcells
timestamp 1726359333
transform 1 0 224 0 1 -333
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPXv0  sky130_fd_pr__nfet_01v8_FQGQPX_1
timestamp 1726359333
transform 1 0 126 0 1 -333
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPXv0  sky130_fd_pr__nfet_01v8_FQGQPX_2
timestamp 1726359333
transform 1 0 420 0 1 -333
box -104 -176 104 176
use sky130_fd_pr__nfet_01v8_FQGQPXv0  sky130_fd_pr__nfet_01v8_FQGQPX_3
timestamp 1726359333
transform 1 0 322 0 1 -333
box -104 -176 104 176
use sky130_fd_pr__pfet_01v8_WNFSTCv0  sky130_fd_pr__pfet_01v8_WNFSTC_0 paramcells
timestamp 1726359333
transform 1 0 126 0 1 204
box -114 -212 114 212
use sky130_fd_pr__pfet_01v8_WNFSTCv0  sky130_fd_pr__pfet_01v8_WNFSTC_1
timestamp 1726359333
transform 1 0 322 0 1 204
box -114 -212 114 212
use sky130_fd_pr__pfet_01v8_WNFSTCv0  sky130_fd_pr__pfet_01v8_WNFSTC_2
timestamp 1726359333
transform 1 0 224 0 1 204
box -114 -212 114 212
use sky130_fd_pr__pfet_01v8_WNFSTCv0  sky130_fd_pr__pfet_01v8_WNFSTC_3
timestamp 1726359333
transform 1 0 420 0 1 204
box -114 -212 114 212
<< labels >>
flabel locali s 253 522 253 522 0 FreeSans 750 0 0 0 VDD
flabel locali s -38 -19 -38 -19 0 FreeSans 750 0 0 0 B
flabel locali s 276 -570 276 -570 0 FreeSans 2500 0 0 0 VSS
flabel locali s 571 -13 571 -13 0 FreeSans 1250 0 0 0 VOUT
<< end >>
