magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect -301 -262 301 262
<< pmos >>
rect -207 -200 -147 200
rect -89 -200 -29 200
rect 29 -200 89 200
rect 147 -200 207 200
<< pdiff >>
rect -265 187 -207 200
rect -265 153 -253 187
rect -219 153 -207 187
rect -265 119 -207 153
rect -265 85 -253 119
rect -219 85 -207 119
rect -265 51 -207 85
rect -265 17 -253 51
rect -219 17 -207 51
rect -265 -17 -207 17
rect -265 -51 -253 -17
rect -219 -51 -207 -17
rect -265 -85 -207 -51
rect -265 -119 -253 -85
rect -219 -119 -207 -85
rect -265 -153 -207 -119
rect -265 -187 -253 -153
rect -219 -187 -207 -153
rect -265 -200 -207 -187
rect -147 187 -89 200
rect -147 153 -135 187
rect -101 153 -89 187
rect -147 119 -89 153
rect -147 85 -135 119
rect -101 85 -89 119
rect -147 51 -89 85
rect -147 17 -135 51
rect -101 17 -89 51
rect -147 -17 -89 17
rect -147 -51 -135 -17
rect -101 -51 -89 -17
rect -147 -85 -89 -51
rect -147 -119 -135 -85
rect -101 -119 -89 -85
rect -147 -153 -89 -119
rect -147 -187 -135 -153
rect -101 -187 -89 -153
rect -147 -200 -89 -187
rect -29 187 29 200
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -200 29 -187
rect 89 187 147 200
rect 89 153 101 187
rect 135 153 147 187
rect 89 119 147 153
rect 89 85 101 119
rect 135 85 147 119
rect 89 51 147 85
rect 89 17 101 51
rect 135 17 147 51
rect 89 -17 147 17
rect 89 -51 101 -17
rect 135 -51 147 -17
rect 89 -85 147 -51
rect 89 -119 101 -85
rect 135 -119 147 -85
rect 89 -153 147 -119
rect 89 -187 101 -153
rect 135 -187 147 -153
rect 89 -200 147 -187
rect 207 187 265 200
rect 207 153 219 187
rect 253 153 265 187
rect 207 119 265 153
rect 207 85 219 119
rect 253 85 265 119
rect 207 51 265 85
rect 207 17 219 51
rect 253 17 265 51
rect 207 -17 265 17
rect 207 -51 219 -17
rect 253 -51 265 -17
rect 207 -85 265 -51
rect 207 -119 219 -85
rect 253 -119 265 -85
rect 207 -153 265 -119
rect 207 -187 219 -153
rect 253 -187 265 -153
rect 207 -200 265 -187
<< pdiffc >>
rect -253 153 -219 187
rect -253 85 -219 119
rect -253 17 -219 51
rect -253 -51 -219 -17
rect -253 -119 -219 -85
rect -253 -187 -219 -153
rect -135 153 -101 187
rect -135 85 -101 119
rect -135 17 -101 51
rect -135 -51 -101 -17
rect -135 -119 -101 -85
rect -135 -187 -101 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 101 153 135 187
rect 101 85 135 119
rect 101 17 135 51
rect 101 -51 135 -17
rect 101 -119 135 -85
rect 101 -187 135 -153
rect 219 153 253 187
rect 219 85 253 119
rect 219 17 253 51
rect 219 -51 253 -17
rect 219 -119 253 -85
rect 219 -187 253 -153
<< poly >>
rect -207 200 -147 226
rect -89 200 -29 226
rect 29 200 89 226
rect 147 200 207 226
rect -207 -226 -147 -200
rect -89 -226 -29 -200
rect 29 -226 89 -200
rect 147 -226 207 -200
<< locali >>
rect -253 187 -219 204
rect -253 119 -219 127
rect -253 51 -219 55
rect -253 -55 -219 -51
rect -253 -127 -219 -119
rect -253 -204 -219 -187
rect -135 187 -101 204
rect -135 119 -101 127
rect -135 51 -101 55
rect -135 -55 -101 -51
rect -135 -127 -101 -119
rect -135 -204 -101 -187
rect -17 187 17 204
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -204 17 -187
rect 101 187 135 204
rect 101 119 135 127
rect 101 51 135 55
rect 101 -55 135 -51
rect 101 -127 135 -119
rect 101 -204 135 -187
rect 219 187 253 204
rect 219 119 253 127
rect 219 51 253 55
rect 219 -55 253 -51
rect 219 -127 253 -119
rect 219 -204 253 -187
<< viali >>
rect -253 153 -219 161
rect -253 127 -219 153
rect -253 85 -219 89
rect -253 55 -219 85
rect -253 -17 -219 17
rect -253 -85 -219 -55
rect -253 -89 -219 -85
rect -253 -153 -219 -127
rect -253 -161 -219 -153
rect -135 153 -101 161
rect -135 127 -101 153
rect -135 85 -101 89
rect -135 55 -101 85
rect -135 -17 -101 17
rect -135 -85 -101 -55
rect -135 -89 -101 -85
rect -135 -153 -101 -127
rect -135 -161 -101 -153
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect 101 153 135 161
rect 101 127 135 153
rect 101 85 135 89
rect 101 55 135 85
rect 101 -17 135 17
rect 101 -85 135 -55
rect 101 -89 135 -85
rect 101 -153 135 -127
rect 101 -161 135 -153
rect 219 153 253 161
rect 219 127 253 153
rect 219 85 253 89
rect 219 55 253 85
rect 219 -17 253 17
rect 219 -85 253 -55
rect 219 -89 253 -85
rect 219 -153 253 -127
rect 219 -161 253 -153
<< metal1 >>
rect -259 161 -213 200
rect -259 127 -253 161
rect -219 127 -213 161
rect -259 89 -213 127
rect -259 55 -253 89
rect -219 55 -213 89
rect -259 17 -213 55
rect -259 -17 -253 17
rect -219 -17 -213 17
rect -259 -55 -213 -17
rect -259 -89 -253 -55
rect -219 -89 -213 -55
rect -259 -127 -213 -89
rect -259 -161 -253 -127
rect -219 -161 -213 -127
rect -259 -200 -213 -161
rect -141 161 -95 200
rect -141 127 -135 161
rect -101 127 -95 161
rect -141 89 -95 127
rect -141 55 -135 89
rect -101 55 -95 89
rect -141 17 -95 55
rect -141 -17 -135 17
rect -101 -17 -95 17
rect -141 -55 -95 -17
rect -141 -89 -135 -55
rect -101 -89 -95 -55
rect -141 -127 -95 -89
rect -141 -161 -135 -127
rect -101 -161 -95 -127
rect -141 -200 -95 -161
rect -23 161 23 200
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -200 23 -161
rect 95 161 141 200
rect 95 127 101 161
rect 135 127 141 161
rect 95 89 141 127
rect 95 55 101 89
rect 135 55 141 89
rect 95 17 141 55
rect 95 -17 101 17
rect 135 -17 141 17
rect 95 -55 141 -17
rect 95 -89 101 -55
rect 135 -89 141 -55
rect 95 -127 141 -89
rect 95 -161 101 -127
rect 135 -161 141 -127
rect 95 -200 141 -161
rect 213 161 259 200
rect 213 127 219 161
rect 253 127 259 161
rect 213 89 259 127
rect 213 55 219 89
rect 253 55 259 89
rect 213 17 259 55
rect 213 -17 219 17
rect 253 -17 259 17
rect 213 -55 259 -17
rect 213 -89 219 -55
rect 253 -89 259 -55
rect 213 -127 259 -89
rect 213 -161 219 -127
rect 253 -161 259 -127
rect 213 -200 259 -161
<< end >>
