magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect 1529 2669 6198 3030
rect 1529 1781 1621 2669
rect 1638 2606 1672 2669
rect 2554 1803 2718 2669
rect 4400 2607 4434 2669
rect 6115 2607 6149 2669
rect 5258 1781 5292 1807
rect 1529 1745 6104 1781
rect 1580 1700 6104 1745
<< pwell >>
rect 1718 -557 6212 -359
<< psubdiff >>
rect 1744 -443 6186 -385
rect 1744 -477 1816 -443
rect 1850 -477 1884 -443
rect 1918 -477 1952 -443
rect 1986 -477 2020 -443
rect 2054 -477 2088 -443
rect 2122 -477 2156 -443
rect 2190 -477 2224 -443
rect 2258 -477 2292 -443
rect 2326 -477 2360 -443
rect 2394 -477 2428 -443
rect 2462 -477 2496 -443
rect 2530 -477 2564 -443
rect 2598 -477 2632 -443
rect 2666 -477 2700 -443
rect 2734 -477 2768 -443
rect 2802 -477 2836 -443
rect 2870 -477 2904 -443
rect 2938 -477 2972 -443
rect 3006 -477 3040 -443
rect 3074 -477 3108 -443
rect 3142 -477 3176 -443
rect 3210 -477 3244 -443
rect 3278 -477 3312 -443
rect 3346 -477 3380 -443
rect 3414 -477 3448 -443
rect 3482 -477 3516 -443
rect 3550 -477 3584 -443
rect 3618 -477 3652 -443
rect 3686 -477 3720 -443
rect 3754 -477 3788 -443
rect 3822 -477 3856 -443
rect 3890 -477 3924 -443
rect 3958 -477 3992 -443
rect 4026 -477 4060 -443
rect 4094 -477 4128 -443
rect 4162 -477 4196 -443
rect 4230 -477 4264 -443
rect 4298 -477 4332 -443
rect 4366 -477 4400 -443
rect 4434 -477 4468 -443
rect 4502 -477 4536 -443
rect 4570 -477 4604 -443
rect 4638 -477 4672 -443
rect 4706 -477 4740 -443
rect 4774 -477 4808 -443
rect 4842 -477 4876 -443
rect 4910 -477 4944 -443
rect 4978 -477 5012 -443
rect 5046 -477 5080 -443
rect 5114 -477 5148 -443
rect 5182 -477 5216 -443
rect 5250 -477 5284 -443
rect 5318 -477 5352 -443
rect 5386 -477 5420 -443
rect 5454 -477 5488 -443
rect 5522 -477 5556 -443
rect 5590 -477 5624 -443
rect 5658 -477 5692 -443
rect 5726 -477 5760 -443
rect 5794 -477 5828 -443
rect 5862 -477 5896 -443
rect 5930 -477 5964 -443
rect 5998 -477 6032 -443
rect 6066 -477 6100 -443
rect 6134 -477 6186 -443
rect 1744 -531 6186 -477
<< nsubdiff >>
rect 1580 2905 6150 2951
rect 1580 2803 1695 2905
rect 6013 2803 6150 2905
rect 1580 2769 6150 2803
<< psubdiffcont >>
rect 1816 -477 1850 -443
rect 1884 -477 1918 -443
rect 1952 -477 1986 -443
rect 2020 -477 2054 -443
rect 2088 -477 2122 -443
rect 2156 -477 2190 -443
rect 2224 -477 2258 -443
rect 2292 -477 2326 -443
rect 2360 -477 2394 -443
rect 2428 -477 2462 -443
rect 2496 -477 2530 -443
rect 2564 -477 2598 -443
rect 2632 -477 2666 -443
rect 2700 -477 2734 -443
rect 2768 -477 2802 -443
rect 2836 -477 2870 -443
rect 2904 -477 2938 -443
rect 2972 -477 3006 -443
rect 3040 -477 3074 -443
rect 3108 -477 3142 -443
rect 3176 -477 3210 -443
rect 3244 -477 3278 -443
rect 3312 -477 3346 -443
rect 3380 -477 3414 -443
rect 3448 -477 3482 -443
rect 3516 -477 3550 -443
rect 3584 -477 3618 -443
rect 3652 -477 3686 -443
rect 3720 -477 3754 -443
rect 3788 -477 3822 -443
rect 3856 -477 3890 -443
rect 3924 -477 3958 -443
rect 3992 -477 4026 -443
rect 4060 -477 4094 -443
rect 4128 -477 4162 -443
rect 4196 -477 4230 -443
rect 4264 -477 4298 -443
rect 4332 -477 4366 -443
rect 4400 -477 4434 -443
rect 4468 -477 4502 -443
rect 4536 -477 4570 -443
rect 4604 -477 4638 -443
rect 4672 -477 4706 -443
rect 4740 -477 4774 -443
rect 4808 -477 4842 -443
rect 4876 -477 4910 -443
rect 4944 -477 4978 -443
rect 5012 -477 5046 -443
rect 5080 -477 5114 -443
rect 5148 -477 5182 -443
rect 5216 -477 5250 -443
rect 5284 -477 5318 -443
rect 5352 -477 5386 -443
rect 5420 -477 5454 -443
rect 5488 -477 5522 -443
rect 5556 -477 5590 -443
rect 5624 -477 5658 -443
rect 5692 -477 5726 -443
rect 5760 -477 5794 -443
rect 5828 -477 5862 -443
rect 5896 -477 5930 -443
rect 5964 -477 5998 -443
rect 6032 -477 6066 -443
rect 6100 -477 6134 -443
<< nsubdiffcont >>
rect 1695 2803 6013 2905
<< poly >>
rect 1580 1700 6104 1781
rect 3744 1666 3785 1700
rect 3819 1666 3860 1700
rect 3744 1642 3860 1666
rect 4044 1666 4085 1700
rect 4119 1666 4160 1700
rect 4044 1642 4160 1666
rect 4344 1666 4385 1700
rect 4419 1666 4460 1700
rect 4344 1642 4460 1666
rect 4644 1666 4685 1700
rect 4719 1666 4760 1700
rect 4644 1642 4760 1666
rect 4944 1666 4985 1700
rect 5019 1666 5060 1700
rect 4944 1642 5060 1666
rect 1999 765 2479 821
rect 1999 731 2053 765
rect 2087 731 2121 765
rect 2155 731 2189 765
rect 2223 731 2257 765
rect 2291 731 2325 765
rect 2359 731 2393 765
rect 2427 731 2479 765
rect 1999 728 2479 731
rect 1836 675 6068 728
rect 1836 641 3504 675
rect 3538 667 6068 675
rect 3538 641 5222 667
rect 1836 633 5222 641
rect 5256 633 6068 667
rect 1836 580 6068 633
<< polycont >>
rect 3785 1666 3819 1700
rect 4085 1666 4119 1700
rect 4385 1666 4419 1700
rect 4685 1666 4719 1700
rect 4985 1666 5019 1700
rect 2053 731 2087 765
rect 2121 731 2155 765
rect 2189 731 2223 765
rect 2257 731 2291 765
rect 2325 731 2359 765
rect 2393 731 2427 765
rect 3504 641 3538 675
rect 5222 633 5256 667
<< locali >>
rect 1580 2905 6150 2951
rect 1580 2803 1695 2905
rect 6013 2803 6150 2905
rect 1580 2769 6150 2803
rect 1638 2606 1672 2769
rect 2096 1639 2130 1806
rect 2554 1803 2718 2769
rect 4400 2607 4434 2769
rect 6116 2607 6150 2769
rect 3542 1669 3576 1807
rect 3744 1700 3860 1725
rect 3744 1669 3785 1700
rect 3506 1666 3785 1669
rect 3819 1669 3860 1700
rect 4044 1700 4160 1725
rect 4044 1669 4085 1700
rect 3819 1666 4085 1669
rect 4119 1669 4160 1700
rect 4344 1700 4460 1725
rect 4344 1669 4385 1700
rect 4119 1666 4385 1669
rect 4419 1669 4460 1700
rect 4644 1700 4760 1725
rect 4644 1669 4685 1700
rect 4419 1666 4685 1669
rect 4719 1669 4760 1700
rect 4944 1700 5060 1725
rect 4944 1669 4985 1700
rect 4719 1666 4985 1669
rect 5019 1669 5060 1700
rect 5258 1669 5292 1807
rect 5019 1666 5292 1669
rect 3506 1635 5292 1666
rect 3506 1556 3540 1635
rect 5222 1554 5256 1635
rect 2158 821 2271 934
rect 1999 765 2479 821
rect 1999 731 2053 765
rect 2087 731 2121 765
rect 2155 731 2189 765
rect 2223 731 2257 765
rect 2291 731 2325 765
rect 2359 731 2393 765
rect 2427 731 2479 765
rect 1790 554 1824 731
rect 1999 676 2479 731
rect 2648 554 2682 752
rect 3457 675 3583 703
rect 3457 641 3504 675
rect 3538 641 3583 675
rect 3457 612 3583 641
rect 3506 555 3540 612
rect 4364 554 4398 752
rect 5196 667 5282 693
rect 5196 633 5222 667
rect 5256 633 5282 667
rect 5196 607 5282 633
rect 5222 554 5256 607
rect 6080 554 6114 752
rect 2647 -385 2682 -246
rect 4364 -385 4398 -248
rect 6080 -385 6114 -249
rect 1744 -443 6186 -385
rect 1744 -477 1816 -443
rect 1850 -477 1884 -443
rect 1918 -477 1952 -443
rect 1986 -477 2020 -443
rect 2054 -477 2088 -443
rect 2122 -477 2156 -443
rect 2190 -477 2224 -443
rect 2258 -477 2292 -443
rect 2326 -477 2360 -443
rect 2394 -477 2428 -443
rect 2462 -477 2496 -443
rect 2530 -477 2564 -443
rect 2598 -477 2632 -443
rect 2666 -477 2700 -443
rect 2734 -477 2768 -443
rect 2802 -477 2836 -443
rect 2870 -477 2904 -443
rect 2938 -477 2972 -443
rect 3006 -477 3040 -443
rect 3074 -477 3108 -443
rect 3142 -477 3176 -443
rect 3210 -477 3244 -443
rect 3278 -477 3312 -443
rect 3346 -477 3380 -443
rect 3414 -477 3448 -443
rect 3482 -477 3516 -443
rect 3550 -477 3584 -443
rect 3618 -477 3652 -443
rect 3686 -477 3720 -443
rect 3754 -477 3788 -443
rect 3822 -477 3856 -443
rect 3890 -477 3924 -443
rect 3958 -477 3992 -443
rect 4026 -477 4060 -443
rect 4094 -477 4128 -443
rect 4162 -477 4196 -443
rect 4230 -477 4264 -443
rect 4298 -477 4332 -443
rect 4366 -477 4400 -443
rect 4434 -477 4468 -443
rect 4502 -477 4536 -443
rect 4570 -477 4604 -443
rect 4638 -477 4672 -443
rect 4706 -477 4740 -443
rect 4774 -477 4808 -443
rect 4842 -477 4876 -443
rect 4910 -477 4944 -443
rect 4978 -477 5012 -443
rect 5046 -477 5080 -443
rect 5114 -477 5148 -443
rect 5182 -477 5216 -443
rect 5250 -477 5284 -443
rect 5318 -477 5352 -443
rect 5386 -477 5420 -443
rect 5454 -477 5488 -443
rect 5522 -477 5556 -443
rect 5590 -477 5624 -443
rect 5658 -477 5692 -443
rect 5726 -477 5760 -443
rect 5794 -477 5828 -443
rect 5862 -477 5896 -443
rect 5930 -477 5964 -443
rect 5998 -477 6032 -443
rect 6066 -477 6100 -443
rect 6134 -477 6186 -443
rect 1744 -531 6186 -477
use sky130_fd_pr__nfet_01v8_lvt_QAGZKG  sky130_fd_pr__nfet_01v8_lvt_QAGZKG_0
timestamp 1717691374
transform 1 0 4381 0 1 1154
box -1771 -426 1771 426
use sky130_fd_pr__nfet_01v8_lvt_QAGZKG  sky130_fd_pr__nfet_01v8_lvt_QAGZKG_1
timestamp 1717691374
transform 1 0 4381 0 1 154
box -1771 -426 1771 426
use sky130_fd_pr__nfet_01v8_lvt_X7SJAL  sky130_fd_pr__nfet_01v8_lvt_X7SJAL_0
timestamp 1717691374
transform 1 0 2236 0 1 154
box -484 -426 484 426
use sky130_fd_pr__pfet_01v8_lvt_VFL754  sky130_fd_pr__pfet_01v8_lvt_VFL754_0
timestamp 1717691374
transform 1 0 4417 0 1 2207
box -1781 -462 1781 462
use sky130_fd_pr__pfet_01v8_YFYKQQ  sky130_fd_pr__pfet_01v8_YFYKQQ_0
timestamp 1717691374
transform 1 0 2113 0 1 2207
box -523 -462 523 462
<< labels >>
flabel locali s 3524 1650 3524 1650 0 FreeSans 2000 0 0 0 G_source_up
flabel locali s 2845 2923 2845 2923 0 FreeSans 2000 0 0 0 VDD
flabel locali s 3159 -514 3159 -514 0 FreeSans 2000 0 0 0 VSS
flabel locali s 1800 667 1800 667 0 FreeSans 2000 0 0 0 ITAIL_SINK
flabel locali s 2207 921 2207 921 0 FreeSans 2000 0 0 0 ITAIL
flabel locali s 2112 1662 2112 1662 0 FreeSans 2000 0 0 0 ITAIL_SRC
<< end >>
