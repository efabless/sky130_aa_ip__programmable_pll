magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect 0 524 7600 769
rect 886 464 920 524
rect 1122 465 1156 524
rect 1358 465 1392 524
rect 1594 465 1628 524
rect 1724 464 1758 524
rect 1960 464 1994 524
rect 2196 465 2230 524
rect 2432 465 2466 524
rect 2668 465 2702 524
rect 2904 465 2938 524
rect 3140 465 3174 524
rect 3376 465 3410 524
rect 3612 464 3646 524
rect 3860 464 3894 524
rect 4096 465 4130 524
rect 4332 465 4366 524
rect 4568 465 4602 524
rect 4804 465 4838 524
rect 5040 465 5074 524
rect 5276 465 5310 524
rect 5512 465 5546 524
rect 5748 465 5782 524
rect 5984 465 6018 524
rect 6220 464 6254 524
rect 6456 465 6490 524
rect 6692 464 6726 524
rect 6928 464 6962 524
rect 7164 464 7198 524
rect 7400 464 7434 524
<< pwell >>
rect 266 -982 7519 -804
<< psubdiff >>
rect 292 -878 7493 -830
rect 292 -912 339 -878
rect 373 -912 407 -878
rect 441 -912 475 -878
rect 509 -912 543 -878
rect 577 -912 611 -878
rect 645 -912 679 -878
rect 713 -912 747 -878
rect 781 -912 815 -878
rect 849 -912 883 -878
rect 917 -912 951 -878
rect 985 -912 1019 -878
rect 1053 -912 1087 -878
rect 1121 -912 1155 -878
rect 1189 -912 1223 -878
rect 1257 -912 1291 -878
rect 1325 -912 1359 -878
rect 1393 -912 1427 -878
rect 1461 -912 1495 -878
rect 1529 -912 1563 -878
rect 1597 -912 1631 -878
rect 1665 -912 1699 -878
rect 1733 -912 1767 -878
rect 1801 -912 1835 -878
rect 1869 -912 1903 -878
rect 1937 -912 1971 -878
rect 2005 -912 2039 -878
rect 2073 -912 2107 -878
rect 2141 -912 2175 -878
rect 2209 -912 2243 -878
rect 2277 -912 2311 -878
rect 2345 -912 2379 -878
rect 2413 -912 2447 -878
rect 2481 -912 2515 -878
rect 2549 -912 2583 -878
rect 2617 -912 2651 -878
rect 2685 -912 2719 -878
rect 2753 -912 2787 -878
rect 2821 -912 2855 -878
rect 2889 -912 2923 -878
rect 2957 -912 2991 -878
rect 3025 -912 3059 -878
rect 3093 -912 3127 -878
rect 3161 -912 3195 -878
rect 3229 -912 3263 -878
rect 3297 -912 3331 -878
rect 3365 -912 3399 -878
rect 3433 -912 3467 -878
rect 3501 -912 3535 -878
rect 3569 -912 3603 -878
rect 3637 -912 3671 -878
rect 3705 -912 3739 -878
rect 3773 -912 3807 -878
rect 3841 -912 3875 -878
rect 3909 -912 3943 -878
rect 3977 -912 4011 -878
rect 4045 -912 4079 -878
rect 4113 -912 4147 -878
rect 4181 -912 4215 -878
rect 4249 -912 4283 -878
rect 4317 -912 4351 -878
rect 4385 -912 4419 -878
rect 4453 -912 4487 -878
rect 4521 -912 4555 -878
rect 4589 -912 4623 -878
rect 4657 -912 4691 -878
rect 4725 -912 4759 -878
rect 4793 -912 4827 -878
rect 4861 -912 4895 -878
rect 4929 -912 4963 -878
rect 4997 -912 5031 -878
rect 5065 -912 5099 -878
rect 5133 -912 5167 -878
rect 5201 -912 5235 -878
rect 5269 -912 5303 -878
rect 5337 -912 5371 -878
rect 5405 -912 5439 -878
rect 5473 -912 5507 -878
rect 5541 -912 5575 -878
rect 5609 -912 5643 -878
rect 5677 -912 5711 -878
rect 5745 -912 5779 -878
rect 5813 -912 5847 -878
rect 5881 -912 5915 -878
rect 5949 -912 5983 -878
rect 6017 -912 6051 -878
rect 6085 -912 6119 -878
rect 6153 -912 6187 -878
rect 6221 -912 6255 -878
rect 6289 -912 6323 -878
rect 6357 -912 6391 -878
rect 6425 -912 6459 -878
rect 6493 -912 6527 -878
rect 6561 -912 6595 -878
rect 6629 -912 6663 -878
rect 6697 -912 6731 -878
rect 6765 -912 6799 -878
rect 6833 -912 6867 -878
rect 6901 -912 6935 -878
rect 6969 -912 7003 -878
rect 7037 -912 7071 -878
rect 7105 -912 7139 -878
rect 7173 -912 7207 -878
rect 7241 -912 7275 -878
rect 7309 -912 7343 -878
rect 7377 -912 7411 -878
rect 7445 -912 7493 -878
rect 292 -956 7493 -912
<< nsubdiff >>
rect 47 675 7515 706
rect 47 641 129 675
rect 163 641 197 675
rect 231 641 265 675
rect 299 641 333 675
rect 367 641 401 675
rect 435 641 469 675
rect 503 641 537 675
rect 571 641 605 675
rect 639 641 673 675
rect 707 641 741 675
rect 775 641 809 675
rect 843 641 877 675
rect 911 641 945 675
rect 979 641 1013 675
rect 1047 641 1081 675
rect 1115 641 1149 675
rect 1183 641 1217 675
rect 1251 641 1285 675
rect 1319 641 1353 675
rect 1387 641 1421 675
rect 1455 641 1489 675
rect 1523 641 1557 675
rect 1591 641 1625 675
rect 1659 641 1693 675
rect 1727 641 1761 675
rect 1795 641 1829 675
rect 1863 641 1897 675
rect 1931 641 1965 675
rect 1999 641 2033 675
rect 2067 641 2101 675
rect 2135 641 2169 675
rect 2203 641 2237 675
rect 2271 641 2305 675
rect 2339 641 2373 675
rect 2407 641 2441 675
rect 2475 641 2509 675
rect 2543 641 2577 675
rect 2611 641 2645 675
rect 2679 641 2713 675
rect 2747 641 2781 675
rect 2815 641 2849 675
rect 2883 641 2917 675
rect 2951 641 2985 675
rect 3019 641 3053 675
rect 3087 641 3121 675
rect 3155 641 3189 675
rect 3223 641 3257 675
rect 3291 641 3325 675
rect 3359 641 3393 675
rect 3427 641 3461 675
rect 3495 641 3529 675
rect 3563 641 3597 675
rect 3631 641 3665 675
rect 3699 641 3733 675
rect 3767 641 3801 675
rect 3835 641 3869 675
rect 3903 641 3937 675
rect 3971 641 4005 675
rect 4039 641 4073 675
rect 4107 641 4141 675
rect 4175 641 4209 675
rect 4243 641 4277 675
rect 4311 641 4345 675
rect 4379 641 4413 675
rect 4447 641 4481 675
rect 4515 641 4549 675
rect 4583 641 4617 675
rect 4651 641 4685 675
rect 4719 641 4753 675
rect 4787 641 4821 675
rect 4855 641 4889 675
rect 4923 641 4957 675
rect 4991 641 5025 675
rect 5059 641 5093 675
rect 5127 641 5161 675
rect 5195 641 5229 675
rect 5263 641 5297 675
rect 5331 641 5365 675
rect 5399 641 5433 675
rect 5467 641 5501 675
rect 5535 641 5569 675
rect 5603 641 5637 675
rect 5671 641 5705 675
rect 5739 641 5773 675
rect 5807 641 5841 675
rect 5875 641 5909 675
rect 5943 641 5977 675
rect 6011 641 6045 675
rect 6079 641 6113 675
rect 6147 641 6181 675
rect 6215 641 6249 675
rect 6283 641 6317 675
rect 6351 641 6385 675
rect 6419 641 6453 675
rect 6487 641 6521 675
rect 6555 641 6589 675
rect 6623 641 6657 675
rect 6691 641 6725 675
rect 6759 641 6793 675
rect 6827 641 6861 675
rect 6895 641 6929 675
rect 6963 641 6997 675
rect 7031 641 7065 675
rect 7099 641 7133 675
rect 7167 641 7201 675
rect 7235 641 7269 675
rect 7303 641 7337 675
rect 7371 641 7405 675
rect 7439 641 7515 675
rect 47 615 7515 641
<< psubdiffcont >>
rect 339 -912 373 -878
rect 407 -912 441 -878
rect 475 -912 509 -878
rect 543 -912 577 -878
rect 611 -912 645 -878
rect 679 -912 713 -878
rect 747 -912 781 -878
rect 815 -912 849 -878
rect 883 -912 917 -878
rect 951 -912 985 -878
rect 1019 -912 1053 -878
rect 1087 -912 1121 -878
rect 1155 -912 1189 -878
rect 1223 -912 1257 -878
rect 1291 -912 1325 -878
rect 1359 -912 1393 -878
rect 1427 -912 1461 -878
rect 1495 -912 1529 -878
rect 1563 -912 1597 -878
rect 1631 -912 1665 -878
rect 1699 -912 1733 -878
rect 1767 -912 1801 -878
rect 1835 -912 1869 -878
rect 1903 -912 1937 -878
rect 1971 -912 2005 -878
rect 2039 -912 2073 -878
rect 2107 -912 2141 -878
rect 2175 -912 2209 -878
rect 2243 -912 2277 -878
rect 2311 -912 2345 -878
rect 2379 -912 2413 -878
rect 2447 -912 2481 -878
rect 2515 -912 2549 -878
rect 2583 -912 2617 -878
rect 2651 -912 2685 -878
rect 2719 -912 2753 -878
rect 2787 -912 2821 -878
rect 2855 -912 2889 -878
rect 2923 -912 2957 -878
rect 2991 -912 3025 -878
rect 3059 -912 3093 -878
rect 3127 -912 3161 -878
rect 3195 -912 3229 -878
rect 3263 -912 3297 -878
rect 3331 -912 3365 -878
rect 3399 -912 3433 -878
rect 3467 -912 3501 -878
rect 3535 -912 3569 -878
rect 3603 -912 3637 -878
rect 3671 -912 3705 -878
rect 3739 -912 3773 -878
rect 3807 -912 3841 -878
rect 3875 -912 3909 -878
rect 3943 -912 3977 -878
rect 4011 -912 4045 -878
rect 4079 -912 4113 -878
rect 4147 -912 4181 -878
rect 4215 -912 4249 -878
rect 4283 -912 4317 -878
rect 4351 -912 4385 -878
rect 4419 -912 4453 -878
rect 4487 -912 4521 -878
rect 4555 -912 4589 -878
rect 4623 -912 4657 -878
rect 4691 -912 4725 -878
rect 4759 -912 4793 -878
rect 4827 -912 4861 -878
rect 4895 -912 4929 -878
rect 4963 -912 4997 -878
rect 5031 -912 5065 -878
rect 5099 -912 5133 -878
rect 5167 -912 5201 -878
rect 5235 -912 5269 -878
rect 5303 -912 5337 -878
rect 5371 -912 5405 -878
rect 5439 -912 5473 -878
rect 5507 -912 5541 -878
rect 5575 -912 5609 -878
rect 5643 -912 5677 -878
rect 5711 -912 5745 -878
rect 5779 -912 5813 -878
rect 5847 -912 5881 -878
rect 5915 -912 5949 -878
rect 5983 -912 6017 -878
rect 6051 -912 6085 -878
rect 6119 -912 6153 -878
rect 6187 -912 6221 -878
rect 6255 -912 6289 -878
rect 6323 -912 6357 -878
rect 6391 -912 6425 -878
rect 6459 -912 6493 -878
rect 6527 -912 6561 -878
rect 6595 -912 6629 -878
rect 6663 -912 6697 -878
rect 6731 -912 6765 -878
rect 6799 -912 6833 -878
rect 6867 -912 6901 -878
rect 6935 -912 6969 -878
rect 7003 -912 7037 -878
rect 7071 -912 7105 -878
rect 7139 -912 7173 -878
rect 7207 -912 7241 -878
rect 7275 -912 7309 -878
rect 7343 -912 7377 -878
rect 7411 -912 7445 -878
<< nsubdiffcont >>
rect 129 641 163 675
rect 197 641 231 675
rect 265 641 299 675
rect 333 641 367 675
rect 401 641 435 675
rect 469 641 503 675
rect 537 641 571 675
rect 605 641 639 675
rect 673 641 707 675
rect 741 641 775 675
rect 809 641 843 675
rect 877 641 911 675
rect 945 641 979 675
rect 1013 641 1047 675
rect 1081 641 1115 675
rect 1149 641 1183 675
rect 1217 641 1251 675
rect 1285 641 1319 675
rect 1353 641 1387 675
rect 1421 641 1455 675
rect 1489 641 1523 675
rect 1557 641 1591 675
rect 1625 641 1659 675
rect 1693 641 1727 675
rect 1761 641 1795 675
rect 1829 641 1863 675
rect 1897 641 1931 675
rect 1965 641 1999 675
rect 2033 641 2067 675
rect 2101 641 2135 675
rect 2169 641 2203 675
rect 2237 641 2271 675
rect 2305 641 2339 675
rect 2373 641 2407 675
rect 2441 641 2475 675
rect 2509 641 2543 675
rect 2577 641 2611 675
rect 2645 641 2679 675
rect 2713 641 2747 675
rect 2781 641 2815 675
rect 2849 641 2883 675
rect 2917 641 2951 675
rect 2985 641 3019 675
rect 3053 641 3087 675
rect 3121 641 3155 675
rect 3189 641 3223 675
rect 3257 641 3291 675
rect 3325 641 3359 675
rect 3393 641 3427 675
rect 3461 641 3495 675
rect 3529 641 3563 675
rect 3597 641 3631 675
rect 3665 641 3699 675
rect 3733 641 3767 675
rect 3801 641 3835 675
rect 3869 641 3903 675
rect 3937 641 3971 675
rect 4005 641 4039 675
rect 4073 641 4107 675
rect 4141 641 4175 675
rect 4209 641 4243 675
rect 4277 641 4311 675
rect 4345 641 4379 675
rect 4413 641 4447 675
rect 4481 641 4515 675
rect 4549 641 4583 675
rect 4617 641 4651 675
rect 4685 641 4719 675
rect 4753 641 4787 675
rect 4821 641 4855 675
rect 4889 641 4923 675
rect 4957 641 4991 675
rect 5025 641 5059 675
rect 5093 641 5127 675
rect 5161 641 5195 675
rect 5229 641 5263 675
rect 5297 641 5331 675
rect 5365 641 5399 675
rect 5433 641 5467 675
rect 5501 641 5535 675
rect 5569 641 5603 675
rect 5637 641 5671 675
rect 5705 641 5739 675
rect 5773 641 5807 675
rect 5841 641 5875 675
rect 5909 641 5943 675
rect 5977 641 6011 675
rect 6045 641 6079 675
rect 6113 641 6147 675
rect 6181 641 6215 675
rect 6249 641 6283 675
rect 6317 641 6351 675
rect 6385 641 6419 675
rect 6453 641 6487 675
rect 6521 641 6555 675
rect 6589 641 6623 675
rect 6657 641 6691 675
rect 6725 641 6759 675
rect 6793 641 6827 675
rect 6861 641 6895 675
rect 6929 641 6963 675
rect 6997 641 7031 675
rect 7065 641 7099 675
rect 7133 641 7167 675
rect 7201 641 7235 675
rect 7269 641 7303 675
rect 7337 641 7371 675
rect 7405 641 7439 675
<< poly >>
rect 94 487 508 524
rect 696 488 1582 525
rect 1770 488 3600 525
rect 3788 488 7506 525
rect 94 -24 508 37
rect 386 -125 446 -24
rect 696 -25 1582 36
rect 1770 -24 3600 36
rect 3788 -24 7506 37
rect 386 -159 398 -125
rect 432 -159 446 -125
rect 386 -225 446 -159
rect 386 -259 398 -225
rect 432 -259 446 -225
rect 386 -278 446 -259
rect 976 -95 1036 -25
rect 976 -129 988 -95
rect 1022 -129 1036 -95
rect 976 -170 1036 -129
rect 976 -204 988 -170
rect 1022 -204 1036 -170
rect 976 -278 1036 -204
rect 1920 -73 1980 -24
rect 1920 -107 1933 -73
rect 1967 -107 1980 -73
rect 1920 -157 1980 -107
rect 1920 -191 1933 -157
rect 1967 -191 1980 -157
rect 1920 -278 1980 -191
rect 3808 -112 3868 -24
rect 3808 -146 3820 -112
rect 3854 -146 3868 -112
rect 3808 -191 3868 -146
rect 3808 -225 3821 -191
rect 3855 -225 3868 -191
rect 3808 -278 3868 -225
rect 386 -320 564 -278
rect 622 -320 1036 -278
rect 1094 -320 1980 -278
rect 2038 -320 3868 -278
rect 3926 -272 7408 -259
rect 3926 -306 4064 -272
rect 4098 -306 4164 -272
rect 4198 -306 4264 -272
rect 4298 -306 4364 -272
rect 4398 -306 4464 -272
rect 4498 -306 4564 -272
rect 4598 -306 4664 -272
rect 4698 -306 7408 -272
rect 3926 -320 7408 -306
rect 386 -338 446 -320
rect 976 -338 1036 -320
rect 1920 -338 1980 -320
rect 3808 -338 3868 -320
<< polycont >>
rect 398 -159 432 -125
rect 398 -259 432 -225
rect 988 -129 1022 -95
rect 988 -204 1022 -170
rect 1933 -107 1967 -73
rect 1933 -191 1967 -157
rect 3820 -146 3854 -112
rect 3821 -225 3855 -191
rect 4064 -306 4098 -272
rect 4164 -306 4198 -272
rect 4264 -306 4298 -272
rect 4364 -306 4398 -272
rect 4464 -306 4498 -272
rect 4564 -306 4598 -272
rect 4664 -306 4698 -272
<< locali >>
rect 52 675 7490 691
rect 52 641 129 675
rect 163 641 197 675
rect 231 641 265 675
rect 299 641 333 675
rect 367 641 401 675
rect 435 641 469 675
rect 503 641 537 675
rect 571 641 605 675
rect 639 641 673 675
rect 707 641 741 675
rect 775 641 809 675
rect 843 641 877 675
rect 911 641 945 675
rect 979 641 1013 675
rect 1047 641 1081 675
rect 1115 641 1149 675
rect 1183 641 1217 675
rect 1251 641 1285 675
rect 1319 641 1353 675
rect 1387 641 1421 675
rect 1455 641 1489 675
rect 1523 641 1557 675
rect 1591 641 1625 675
rect 1659 641 1693 675
rect 1727 641 1761 675
rect 1795 641 1829 675
rect 1863 641 1897 675
rect 1931 641 1965 675
rect 1999 641 2033 675
rect 2067 641 2101 675
rect 2135 641 2169 675
rect 2203 641 2237 675
rect 2271 641 2305 675
rect 2339 641 2373 675
rect 2407 641 2441 675
rect 2475 641 2509 675
rect 2543 641 2577 675
rect 2611 641 2645 675
rect 2679 641 2713 675
rect 2747 641 2781 675
rect 2815 641 2849 675
rect 2883 641 2917 675
rect 2951 641 2985 675
rect 3019 641 3053 675
rect 3087 641 3121 675
rect 3155 641 3189 675
rect 3223 641 3257 675
rect 3291 641 3325 675
rect 3359 641 3393 675
rect 3427 641 3461 675
rect 3495 641 3529 675
rect 3563 641 3597 675
rect 3631 641 3665 675
rect 3699 641 3733 675
rect 3767 641 3801 675
rect 3835 641 3869 675
rect 3903 641 3937 675
rect 3971 641 4005 675
rect 4039 641 4073 675
rect 4107 641 4141 675
rect 4175 641 4209 675
rect 4243 641 4277 675
rect 4311 641 4345 675
rect 4379 641 4413 675
rect 4447 641 4481 675
rect 4515 641 4549 675
rect 4583 641 4617 675
rect 4651 641 4685 675
rect 4719 641 4753 675
rect 4787 641 4821 675
rect 4855 641 4889 675
rect 4923 641 4957 675
rect 4991 641 5025 675
rect 5059 641 5093 675
rect 5127 641 5161 675
rect 5195 641 5229 675
rect 5263 641 5297 675
rect 5331 641 5365 675
rect 5399 641 5433 675
rect 5467 641 5501 675
rect 5535 641 5569 675
rect 5603 641 5637 675
rect 5671 641 5705 675
rect 5739 641 5773 675
rect 5807 641 5841 675
rect 5875 641 5909 675
rect 5943 641 5977 675
rect 6011 641 6045 675
rect 6079 641 6113 675
rect 6147 641 6181 675
rect 6215 641 6249 675
rect 6283 641 6317 675
rect 6351 641 6385 675
rect 6419 641 6453 675
rect 6487 641 6521 675
rect 6555 641 6589 675
rect 6623 641 6657 675
rect 6691 641 6725 675
rect 6759 641 6793 675
rect 6827 641 6861 675
rect 6895 641 6929 675
rect 6963 641 6997 675
rect 7031 641 7065 675
rect 7099 641 7133 675
rect 7167 641 7201 675
rect 7235 641 7269 675
rect 7303 641 7337 675
rect 7371 641 7405 675
rect 7439 641 7490 675
rect 52 625 7490 641
rect 253 553 312 625
rect 841 553 900 625
rect 1112 553 1171 625
rect 1353 553 1412 625
rect 1585 553 1644 625
rect 2191 553 2250 625
rect 2420 553 2479 625
rect 2659 553 2718 625
rect 2894 553 2953 625
rect 3130 553 3189 625
rect 3361 553 3420 625
rect 4086 553 4145 625
rect 4320 553 4379 625
rect 4554 553 4613 625
rect 4791 553 4850 625
rect 5021 553 5080 625
rect 5261 553 5320 625
rect 5499 553 5558 625
rect 5735 553 5794 625
rect 5966 553 6025 625
rect 6443 553 6502 625
rect 48 505 7600 553
rect 48 465 82 505
rect 284 466 318 505
rect 520 445 554 505
rect 650 463 684 505
rect 886 464 920 505
rect 1122 465 1156 505
rect 1358 465 1392 505
rect 1594 465 1628 505
rect 1724 464 1758 505
rect 1960 464 1994 505
rect 2196 465 2230 505
rect 2432 465 2466 505
rect 2668 465 2702 505
rect 2904 465 2938 505
rect 3140 465 3174 505
rect 3376 465 3410 505
rect 3612 464 3646 505
rect 3860 464 3894 505
rect 4096 465 4130 505
rect 4332 465 4366 505
rect 4568 465 4602 505
rect 4804 465 4838 505
rect 5040 465 5074 505
rect 5276 465 5310 505
rect 5512 465 5546 505
rect 5748 465 5782 505
rect 5984 465 6018 505
rect 6220 464 6254 505
rect 6456 465 6490 505
rect 6692 464 6726 505
rect 6928 464 6962 505
rect 7164 464 7198 505
rect 7400 464 7434 505
rect 402 -8 436 62
rect 402 -42 610 -8
rect 377 -125 453 -101
rect 377 -159 398 -125
rect 432 -159 453 -125
rect 377 -161 453 -159
rect -156 -222 453 -161
rect 576 -131 610 -42
rect 953 -95 1055 -83
rect 953 -129 988 -95
rect 1022 -129 1055 -95
rect 953 -131 1055 -129
rect 576 -165 1055 -131
rect 1476 -128 1510 59
rect 1914 -73 1986 -54
rect 1914 -107 1933 -73
rect 1967 -107 1986 -73
rect 1914 -128 1986 -107
rect 1476 -157 1986 -128
rect 1476 -162 1933 -157
rect 377 -225 453 -222
rect 953 -170 1055 -165
rect 953 -204 988 -170
rect 1022 -204 1055 -170
rect 953 -223 1055 -204
rect 1914 -191 1933 -162
rect 1967 -191 1986 -157
rect 3494 -142 3528 60
rect 7518 -88 7552 66
rect 3802 -112 3874 -88
rect 3802 -142 3820 -112
rect 3494 -146 3820 -142
rect 3854 -146 3874 -112
rect 7518 -122 7721 -88
rect 3494 -176 3874 -146
rect 1914 -210 1986 -191
rect 3802 -191 3874 -176
rect 377 -259 398 -225
rect 432 -259 453 -225
rect 3802 -225 3821 -191
rect 3855 -225 3874 -191
rect 3802 -244 3874 -225
rect 377 -278 453 -259
rect 3998 -272 7480 -250
rect 3998 -278 4064 -272
rect 3850 -306 4064 -278
rect 4098 -306 4164 -272
rect 4198 -306 4264 -272
rect 4298 -306 4364 -272
rect 4398 -306 4464 -272
rect 4498 -306 4564 -272
rect 4598 -306 4664 -272
rect 4698 -306 7480 -272
rect 3850 -342 7480 -306
rect 340 -835 374 -749
rect 576 -835 610 -749
rect 812 -835 846 -748
rect 1048 -835 1082 -749
rect 1284 -835 1318 -748
rect 1520 -835 1554 -747
rect 1756 -835 1790 -747
rect 1992 -835 2026 -748
rect 2228 -835 2262 -749
rect 2464 -835 2498 -749
rect 2700 -835 2734 -748
rect 2936 -835 2970 -749
rect 3172 -835 3206 -747
rect 3408 -835 3442 -749
rect 3644 -835 3678 -748
rect 3880 -835 3914 -749
rect 298 -878 7485 -835
rect 298 -912 339 -878
rect 373 -912 407 -878
rect 441 -912 475 -878
rect 509 -912 543 -878
rect 577 -912 611 -878
rect 645 -912 679 -878
rect 713 -912 747 -878
rect 781 -912 815 -878
rect 849 -912 883 -878
rect 917 -912 951 -878
rect 985 -912 1019 -878
rect 1053 -912 1087 -878
rect 1121 -912 1155 -878
rect 1189 -912 1223 -878
rect 1257 -912 1291 -878
rect 1325 -912 1359 -878
rect 1393 -912 1427 -878
rect 1461 -912 1495 -878
rect 1529 -912 1563 -878
rect 1597 -912 1631 -878
rect 1665 -912 1699 -878
rect 1733 -912 1767 -878
rect 1801 -912 1835 -878
rect 1869 -912 1903 -878
rect 1937 -912 1971 -878
rect 2005 -912 2039 -878
rect 2073 -912 2107 -878
rect 2141 -912 2175 -878
rect 2209 -912 2243 -878
rect 2277 -912 2311 -878
rect 2345 -912 2379 -878
rect 2413 -912 2447 -878
rect 2481 -912 2515 -878
rect 2549 -912 2583 -878
rect 2617 -912 2651 -878
rect 2685 -912 2719 -878
rect 2753 -912 2787 -878
rect 2821 -912 2855 -878
rect 2889 -912 2923 -878
rect 2957 -912 2991 -878
rect 3025 -912 3059 -878
rect 3093 -912 3127 -878
rect 3161 -912 3195 -878
rect 3229 -912 3263 -878
rect 3297 -912 3331 -878
rect 3365 -912 3399 -878
rect 3433 -912 3467 -878
rect 3501 -912 3535 -878
rect 3569 -912 3603 -878
rect 3637 -912 3671 -878
rect 3705 -912 3739 -878
rect 3773 -912 3807 -878
rect 3841 -912 3875 -878
rect 3909 -912 3943 -878
rect 3977 -912 4011 -878
rect 4045 -912 4079 -878
rect 4113 -912 4147 -878
rect 4181 -912 4215 -878
rect 4249 -912 4283 -878
rect 4317 -912 4351 -878
rect 4385 -912 4419 -878
rect 4453 -912 4487 -878
rect 4521 -912 4555 -878
rect 4589 -912 4623 -878
rect 4657 -912 4691 -878
rect 4725 -912 4759 -878
rect 4793 -912 4827 -878
rect 4861 -912 4895 -878
rect 4929 -912 4963 -878
rect 4997 -912 5031 -878
rect 5065 -912 5099 -878
rect 5133 -912 5167 -878
rect 5201 -912 5235 -878
rect 5269 -912 5303 -878
rect 5337 -912 5371 -878
rect 5405 -912 5439 -878
rect 5473 -912 5507 -878
rect 5541 -912 5575 -878
rect 5609 -912 5643 -878
rect 5677 -912 5711 -878
rect 5745 -912 5779 -878
rect 5813 -912 5847 -878
rect 5881 -912 5915 -878
rect 5949 -912 5983 -878
rect 6017 -912 6051 -878
rect 6085 -912 6119 -878
rect 6153 -912 6187 -878
rect 6221 -912 6255 -878
rect 6289 -912 6323 -878
rect 6357 -912 6391 -878
rect 6425 -912 6459 -878
rect 6493 -912 6527 -878
rect 6561 -912 6595 -878
rect 6629 -912 6663 -878
rect 6697 -912 6731 -878
rect 6765 -912 6799 -878
rect 6833 -912 6867 -878
rect 6901 -912 6935 -878
rect 6969 -912 7003 -878
rect 7037 -912 7071 -878
rect 7105 -912 7139 -878
rect 7173 -912 7207 -878
rect 7241 -912 7275 -878
rect 7309 -912 7343 -878
rect 7377 -912 7411 -878
rect 7445 -912 7485 -878
rect 298 -955 7485 -912
<< metal1 >>
rect 160 -9 206 67
rect 396 -9 442 68
rect 762 -9 808 63
rect 998 -9 1044 65
rect 1234 -9 1280 63
rect 1470 -9 1516 65
rect 1836 -9 1882 64
rect 2072 -9 2118 63
rect 2308 -9 2354 64
rect 2544 -9 2590 64
rect 2780 -9 2826 65
rect 3016 -9 3062 65
rect 3252 -9 3298 65
rect 3488 -9 3534 66
rect 3736 -9 3782 66
rect 3972 -9 4018 65
rect 4208 -9 4254 66
rect 4444 -9 4490 65
rect 4680 -9 4726 65
rect 4916 -9 4962 66
rect 5152 -9 5198 66
rect 5388 -9 5434 66
rect 5624 -9 5670 66
rect 5860 -9 5906 63
rect 6096 -9 6142 64
rect 6332 -9 6378 65
rect 6568 -9 6614 65
rect 6804 -9 6850 65
rect 7040 -9 7086 64
rect 7276 -9 7322 66
rect 7512 -9 7558 64
rect 155 -83 572 -9
rect 633 -83 1643 -9
rect 1704 -83 3649 -9
rect 3710 -83 7587 -9
rect 452 -348 498 -83
rect 847 -223 893 -83
rect 1829 -211 1875 -83
rect 3756 -199 3802 -83
rect 688 -269 970 -223
rect 688 -346 734 -269
rect 924 -346 970 -269
rect 1160 -257 1914 -211
rect 1160 -346 1206 -257
rect 1396 -346 1442 -257
rect 1632 -346 1678 -257
rect 1868 -346 1914 -257
rect 2104 -245 3802 -199
rect 2104 -346 2150 -245
rect 2340 -346 2386 -245
rect 2576 -346 2622 -245
rect 2812 -346 2858 -245
rect 3048 -346 3094 -245
rect 3284 -346 3330 -245
rect 3520 -346 3566 -245
rect 3756 -346 3802 -245
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_15 paramcells
timestamp 1726359333
transform 1 0 475 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_16
timestamp 1726359333
transform 1 0 711 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_17
timestamp 1726359333
transform 1 0 947 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_18
timestamp 1726359333
transform 1 0 1183 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_19
timestamp 1726359333
transform 1 0 1419 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_20
timestamp 1726359333
transform 1 0 1891 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_21
timestamp 1726359333
transform 1 0 1655 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_22
timestamp 1726359333
transform 1 0 2127 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_23
timestamp 1726359333
transform 1 0 2363 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_24
timestamp 1726359333
transform 1 0 2599 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_25
timestamp 1726359333
transform 1 0 2835 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_26
timestamp 1726359333
transform 1 0 3071 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_27
timestamp 1726359333
transform 1 0 3307 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_28
timestamp 1726359333
transform 1 0 3543 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_29
timestamp 1726359333
transform 1 0 3779 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_30
timestamp 1726359333
transform 1 0 5195 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_31
timestamp 1726359333
transform 1 0 4959 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_32
timestamp 1726359333
transform 1 0 4251 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_33
timestamp 1726359333
transform 1 0 4487 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_34
timestamp 1726359333
transform 1 0 4723 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_35
timestamp 1726359333
transform 1 0 4015 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_36
timestamp 1726359333
transform 1 0 6611 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_37
timestamp 1726359333
transform 1 0 6375 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_38
timestamp 1726359333
transform 1 0 6139 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_39
timestamp 1726359333
transform 1 0 5903 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_40
timestamp 1726359333
transform 1 0 5667 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_41
timestamp 1726359333
transform 1 0 5431 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_42
timestamp 1726359333
transform 1 0 7319 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_43
timestamp 1726359333
transform 1 0 6847 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__nfet_01v8_4LH2UU  sky130_fd_pr__nfet_01v8_4LH2UU_44
timestamp 1726359333
transform 1 0 7083 0 1 -546
box -173 -226 173 226
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_0 paramcells
timestamp 1726359333
transform 1 0 1977 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_1
timestamp 1726359333
transform 1 0 301 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_2
timestamp 1726359333
transform 1 0 2449 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_3
timestamp 1726359333
transform 1 0 1375 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_4
timestamp 1726359333
transform 1 0 903 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_5
timestamp 1726359333
transform 1 0 2921 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_6
timestamp 1726359333
transform 1 0 3393 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_7
timestamp 1726359333
transform 1 0 3995 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_8
timestamp 1726359333
transform 1 0 4467 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_9
timestamp 1726359333
transform 1 0 4939 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_10
timestamp 1726359333
transform 1 0 5411 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_11
timestamp 1726359333
transform 1 0 5883 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_12
timestamp 1726359333
transform 1 0 6355 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_13
timestamp 1726359333
transform 1 0 6827 0 1 262
box -301 -262 301 262
use sky130_fd_pr__pfet_01v8_2PR8SB  sky130_fd_pr__pfet_01v8_2PR8SB_14
timestamp 1726359333
transform 1 0 7299 0 1 262
box -301 -262 301 262
<< labels >>
flabel locali s -124 -196 -124 -196 0 FreeSans 1250 0 0 0 IN
flabel locali s 7699 -107 7699 -107 0 FreeSans 1250 0 0 0 OUT
flabel locali s 2857 673 2857 673 0 FreeSans 1250 0 0 0 VDD
flabel locali s 2625 -896 2625 -896 0 FreeSans 1250 0 0 0 VSS
<< end >>
