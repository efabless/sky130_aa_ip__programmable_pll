magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect -697 -262 697 262
<< pmos >>
rect -603 -200 -503 200
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
rect 503 -200 603 200
<< pdiff >>
rect -661 187 -603 200
rect -661 153 -649 187
rect -615 153 -603 187
rect -661 119 -603 153
rect -661 85 -649 119
rect -615 85 -603 119
rect -661 51 -603 85
rect -661 17 -649 51
rect -615 17 -603 51
rect -661 -17 -603 17
rect -661 -51 -649 -17
rect -615 -51 -603 -17
rect -661 -85 -603 -51
rect -661 -119 -649 -85
rect -615 -119 -603 -85
rect -661 -153 -603 -119
rect -661 -187 -649 -153
rect -615 -187 -603 -153
rect -661 -200 -603 -187
rect -503 187 -445 200
rect -503 153 -491 187
rect -457 153 -445 187
rect -503 119 -445 153
rect -503 85 -491 119
rect -457 85 -445 119
rect -503 51 -445 85
rect -503 17 -491 51
rect -457 17 -445 51
rect -503 -17 -445 17
rect -503 -51 -491 -17
rect -457 -51 -445 -17
rect -503 -85 -445 -51
rect -503 -119 -491 -85
rect -457 -119 -445 -85
rect -503 -153 -445 -119
rect -503 -187 -491 -153
rect -457 -187 -445 -153
rect -503 -200 -445 -187
rect -345 187 -287 200
rect -345 153 -333 187
rect -299 153 -287 187
rect -345 119 -287 153
rect -345 85 -333 119
rect -299 85 -287 119
rect -345 51 -287 85
rect -345 17 -333 51
rect -299 17 -287 51
rect -345 -17 -287 17
rect -345 -51 -333 -17
rect -299 -51 -287 -17
rect -345 -85 -287 -51
rect -345 -119 -333 -85
rect -299 -119 -287 -85
rect -345 -153 -287 -119
rect -345 -187 -333 -153
rect -299 -187 -287 -153
rect -345 -200 -287 -187
rect -187 187 -129 200
rect -187 153 -175 187
rect -141 153 -129 187
rect -187 119 -129 153
rect -187 85 -175 119
rect -141 85 -129 119
rect -187 51 -129 85
rect -187 17 -175 51
rect -141 17 -129 51
rect -187 -17 -129 17
rect -187 -51 -175 -17
rect -141 -51 -129 -17
rect -187 -85 -129 -51
rect -187 -119 -175 -85
rect -141 -119 -129 -85
rect -187 -153 -129 -119
rect -187 -187 -175 -153
rect -141 -187 -129 -153
rect -187 -200 -129 -187
rect -29 187 29 200
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -200 29 -187
rect 129 187 187 200
rect 129 153 141 187
rect 175 153 187 187
rect 129 119 187 153
rect 129 85 141 119
rect 175 85 187 119
rect 129 51 187 85
rect 129 17 141 51
rect 175 17 187 51
rect 129 -17 187 17
rect 129 -51 141 -17
rect 175 -51 187 -17
rect 129 -85 187 -51
rect 129 -119 141 -85
rect 175 -119 187 -85
rect 129 -153 187 -119
rect 129 -187 141 -153
rect 175 -187 187 -153
rect 129 -200 187 -187
rect 287 187 345 200
rect 287 153 299 187
rect 333 153 345 187
rect 287 119 345 153
rect 287 85 299 119
rect 333 85 345 119
rect 287 51 345 85
rect 287 17 299 51
rect 333 17 345 51
rect 287 -17 345 17
rect 287 -51 299 -17
rect 333 -51 345 -17
rect 287 -85 345 -51
rect 287 -119 299 -85
rect 333 -119 345 -85
rect 287 -153 345 -119
rect 287 -187 299 -153
rect 333 -187 345 -153
rect 287 -200 345 -187
rect 445 187 503 200
rect 445 153 457 187
rect 491 153 503 187
rect 445 119 503 153
rect 445 85 457 119
rect 491 85 503 119
rect 445 51 503 85
rect 445 17 457 51
rect 491 17 503 51
rect 445 -17 503 17
rect 445 -51 457 -17
rect 491 -51 503 -17
rect 445 -85 503 -51
rect 445 -119 457 -85
rect 491 -119 503 -85
rect 445 -153 503 -119
rect 445 -187 457 -153
rect 491 -187 503 -153
rect 445 -200 503 -187
rect 603 187 661 200
rect 603 153 615 187
rect 649 153 661 187
rect 603 119 661 153
rect 603 85 615 119
rect 649 85 661 119
rect 603 51 661 85
rect 603 17 615 51
rect 649 17 661 51
rect 603 -17 661 17
rect 603 -51 615 -17
rect 649 -51 661 -17
rect 603 -85 661 -51
rect 603 -119 615 -85
rect 649 -119 661 -85
rect 603 -153 661 -119
rect 603 -187 615 -153
rect 649 -187 661 -153
rect 603 -200 661 -187
<< pdiffc >>
rect -649 153 -615 187
rect -649 85 -615 119
rect -649 17 -615 51
rect -649 -51 -615 -17
rect -649 -119 -615 -85
rect -649 -187 -615 -153
rect -491 153 -457 187
rect -491 85 -457 119
rect -491 17 -457 51
rect -491 -51 -457 -17
rect -491 -119 -457 -85
rect -491 -187 -457 -153
rect -333 153 -299 187
rect -333 85 -299 119
rect -333 17 -299 51
rect -333 -51 -299 -17
rect -333 -119 -299 -85
rect -333 -187 -299 -153
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 299 153 333 187
rect 299 85 333 119
rect 299 17 333 51
rect 299 -51 333 -17
rect 299 -119 333 -85
rect 299 -187 333 -153
rect 457 153 491 187
rect 457 85 491 119
rect 457 17 491 51
rect 457 -51 491 -17
rect 457 -119 491 -85
rect 457 -187 491 -153
rect 615 153 649 187
rect 615 85 649 119
rect 615 17 649 51
rect 615 -51 649 -17
rect 615 -119 649 -85
rect 615 -187 649 -153
<< poly >>
rect -603 200 -503 226
rect -445 200 -345 226
rect -287 200 -187 226
rect -129 200 -29 226
rect 29 200 129 226
rect 187 200 287 226
rect 345 200 445 226
rect 503 200 603 226
rect -603 -226 -503 -200
rect -445 -226 -345 -200
rect -287 -226 -187 -200
rect -129 -226 -29 -200
rect 29 -226 129 -200
rect 187 -226 287 -200
rect 345 -226 445 -200
rect 503 -226 603 -200
<< locali >>
rect -649 187 -615 204
rect -649 119 -615 127
rect -649 51 -615 55
rect -649 -55 -615 -51
rect -649 -127 -615 -119
rect -649 -204 -615 -187
rect -491 187 -457 204
rect -491 119 -457 127
rect -491 51 -457 55
rect -491 -55 -457 -51
rect -491 -127 -457 -119
rect -491 -204 -457 -187
rect -333 187 -299 204
rect -333 119 -299 127
rect -333 51 -299 55
rect -333 -55 -299 -51
rect -333 -127 -299 -119
rect -333 -204 -299 -187
rect -175 187 -141 204
rect -175 119 -141 127
rect -175 51 -141 55
rect -175 -55 -141 -51
rect -175 -127 -141 -119
rect -175 -204 -141 -187
rect -17 187 17 204
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -204 17 -187
rect 141 187 175 204
rect 141 119 175 127
rect 141 51 175 55
rect 141 -55 175 -51
rect 141 -127 175 -119
rect 141 -204 175 -187
rect 299 187 333 204
rect 299 119 333 127
rect 299 51 333 55
rect 299 -55 333 -51
rect 299 -127 333 -119
rect 299 -204 333 -187
rect 457 187 491 204
rect 457 119 491 127
rect 457 51 491 55
rect 457 -55 491 -51
rect 457 -127 491 -119
rect 457 -204 491 -187
rect 615 187 649 204
rect 615 119 649 127
rect 615 51 649 55
rect 615 -55 649 -51
rect 615 -127 649 -119
rect 615 -204 649 -187
<< viali >>
rect -649 153 -615 161
rect -649 127 -615 153
rect -649 85 -615 89
rect -649 55 -615 85
rect -649 -17 -615 17
rect -649 -85 -615 -55
rect -649 -89 -615 -85
rect -649 -153 -615 -127
rect -649 -161 -615 -153
rect -491 153 -457 161
rect -491 127 -457 153
rect -491 85 -457 89
rect -491 55 -457 85
rect -491 -17 -457 17
rect -491 -85 -457 -55
rect -491 -89 -457 -85
rect -491 -153 -457 -127
rect -491 -161 -457 -153
rect -333 153 -299 161
rect -333 127 -299 153
rect -333 85 -299 89
rect -333 55 -299 85
rect -333 -17 -299 17
rect -333 -85 -299 -55
rect -333 -89 -299 -85
rect -333 -153 -299 -127
rect -333 -161 -299 -153
rect -175 153 -141 161
rect -175 127 -141 153
rect -175 85 -141 89
rect -175 55 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -55
rect -175 -89 -141 -85
rect -175 -153 -141 -127
rect -175 -161 -141 -153
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect 141 153 175 161
rect 141 127 175 153
rect 141 85 175 89
rect 141 55 175 85
rect 141 -17 175 17
rect 141 -85 175 -55
rect 141 -89 175 -85
rect 141 -153 175 -127
rect 141 -161 175 -153
rect 299 153 333 161
rect 299 127 333 153
rect 299 85 333 89
rect 299 55 333 85
rect 299 -17 333 17
rect 299 -85 333 -55
rect 299 -89 333 -85
rect 299 -153 333 -127
rect 299 -161 333 -153
rect 457 153 491 161
rect 457 127 491 153
rect 457 85 491 89
rect 457 55 491 85
rect 457 -17 491 17
rect 457 -85 491 -55
rect 457 -89 491 -85
rect 457 -153 491 -127
rect 457 -161 491 -153
rect 615 153 649 161
rect 615 127 649 153
rect 615 85 649 89
rect 615 55 649 85
rect 615 -17 649 17
rect 615 -85 649 -55
rect 615 -89 649 -85
rect 615 -153 649 -127
rect 615 -161 649 -153
<< metal1 >>
rect -655 161 -609 200
rect -655 127 -649 161
rect -615 127 -609 161
rect -655 89 -609 127
rect -655 55 -649 89
rect -615 55 -609 89
rect -655 17 -609 55
rect -655 -17 -649 17
rect -615 -17 -609 17
rect -655 -55 -609 -17
rect -655 -89 -649 -55
rect -615 -89 -609 -55
rect -655 -127 -609 -89
rect -655 -161 -649 -127
rect -615 -161 -609 -127
rect -655 -200 -609 -161
rect -497 161 -451 200
rect -497 127 -491 161
rect -457 127 -451 161
rect -497 89 -451 127
rect -497 55 -491 89
rect -457 55 -451 89
rect -497 17 -451 55
rect -497 -17 -491 17
rect -457 -17 -451 17
rect -497 -55 -451 -17
rect -497 -89 -491 -55
rect -457 -89 -451 -55
rect -497 -127 -451 -89
rect -497 -161 -491 -127
rect -457 -161 -451 -127
rect -497 -200 -451 -161
rect -339 161 -293 200
rect -339 127 -333 161
rect -299 127 -293 161
rect -339 89 -293 127
rect -339 55 -333 89
rect -299 55 -293 89
rect -339 17 -293 55
rect -339 -17 -333 17
rect -299 -17 -293 17
rect -339 -55 -293 -17
rect -339 -89 -333 -55
rect -299 -89 -293 -55
rect -339 -127 -293 -89
rect -339 -161 -333 -127
rect -299 -161 -293 -127
rect -339 -200 -293 -161
rect -181 161 -135 200
rect -181 127 -175 161
rect -141 127 -135 161
rect -181 89 -135 127
rect -181 55 -175 89
rect -141 55 -135 89
rect -181 17 -135 55
rect -181 -17 -175 17
rect -141 -17 -135 17
rect -181 -55 -135 -17
rect -181 -89 -175 -55
rect -141 -89 -135 -55
rect -181 -127 -135 -89
rect -181 -161 -175 -127
rect -141 -161 -135 -127
rect -181 -200 -135 -161
rect -23 161 23 200
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -200 23 -161
rect 135 161 181 200
rect 135 127 141 161
rect 175 127 181 161
rect 135 89 181 127
rect 135 55 141 89
rect 175 55 181 89
rect 135 17 181 55
rect 135 -17 141 17
rect 175 -17 181 17
rect 135 -55 181 -17
rect 135 -89 141 -55
rect 175 -89 181 -55
rect 135 -127 181 -89
rect 135 -161 141 -127
rect 175 -161 181 -127
rect 135 -200 181 -161
rect 293 161 339 200
rect 293 127 299 161
rect 333 127 339 161
rect 293 89 339 127
rect 293 55 299 89
rect 333 55 339 89
rect 293 17 339 55
rect 293 -17 299 17
rect 333 -17 339 17
rect 293 -55 339 -17
rect 293 -89 299 -55
rect 333 -89 339 -55
rect 293 -127 339 -89
rect 293 -161 299 -127
rect 333 -161 339 -127
rect 293 -200 339 -161
rect 451 161 497 200
rect 451 127 457 161
rect 491 127 497 161
rect 451 89 497 127
rect 451 55 457 89
rect 491 55 497 89
rect 451 17 497 55
rect 451 -17 457 17
rect 491 -17 497 17
rect 451 -55 497 -17
rect 451 -89 457 -55
rect 491 -89 497 -55
rect 451 -127 497 -89
rect 451 -161 457 -127
rect 491 -161 497 -127
rect 451 -200 497 -161
rect 609 161 655 200
rect 609 127 615 161
rect 649 127 655 161
rect 609 89 655 127
rect 609 55 615 89
rect 649 55 655 89
rect 609 17 655 55
rect 609 -17 615 17
rect 649 -17 655 17
rect 609 -55 655 -17
rect 609 -89 615 -55
rect 649 -89 655 -55
rect 609 -127 655 -89
rect 609 -161 615 -127
rect 649 -161 655 -127
rect 609 -200 655 -161
<< end >>
