magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect -581 -162 581 162
<< pmoslvt >>
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
<< pdiff >>
rect -545 85 -487 100
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -100 -487 -85
rect -287 85 -229 100
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -100 -229 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 229 85 287 100
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -100 287 -85
rect 487 85 545 100
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -100 545 -85
<< pdiffc >>
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
<< poly >>
rect -487 100 -287 126
rect -229 100 -29 126
rect 29 100 229 126
rect 287 100 487 126
rect -487 -126 -287 -100
rect -229 -126 -29 -100
rect 29 -126 229 -100
rect 287 -126 487 -100
<< locali >>
rect -533 85 -499 104
rect -533 17 -499 19
rect -533 -19 -499 -17
rect -533 -104 -499 -85
rect -275 85 -241 104
rect -275 17 -241 19
rect -275 -19 -241 -17
rect -275 -104 -241 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 241 85 275 104
rect 241 17 275 19
rect 241 -19 275 -17
rect 241 -104 275 -85
rect 499 85 533 104
rect 499 17 533 19
rect 499 -19 533 -17
rect 499 -104 533 -85
<< viali >>
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
<< metal1 >>
rect -539 53 -493 100
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -100 -493 -53
rect -281 53 -235 100
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -100 -235 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 235 53 281 100
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -100 281 -53
rect 493 53 539 100
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -100 539 -53
<< end >>
