magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< nwell >>
rect -381 -162 381 162
<< pmos >>
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
<< pdiff >>
rect -345 85 -287 100
rect -345 51 -333 85
rect -299 51 -287 85
rect -345 17 -287 51
rect -345 -17 -333 17
rect -299 -17 -287 17
rect -345 -51 -287 -17
rect -345 -85 -333 -51
rect -299 -85 -287 -51
rect -345 -100 -287 -85
rect -187 85 -129 100
rect -187 51 -175 85
rect -141 51 -129 85
rect -187 17 -129 51
rect -187 -17 -175 17
rect -141 -17 -129 17
rect -187 -51 -129 -17
rect -187 -85 -175 -51
rect -141 -85 -129 -51
rect -187 -100 -129 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 129 85 187 100
rect 129 51 141 85
rect 175 51 187 85
rect 129 17 187 51
rect 129 -17 141 17
rect 175 -17 187 17
rect 129 -51 187 -17
rect 129 -85 141 -51
rect 175 -85 187 -51
rect 129 -100 187 -85
rect 287 85 345 100
rect 287 51 299 85
rect 333 51 345 85
rect 287 17 345 51
rect 287 -17 299 17
rect 333 -17 345 17
rect 287 -51 345 -17
rect 287 -85 299 -51
rect 333 -85 345 -51
rect 287 -100 345 -85
<< pdiffc >>
rect -333 51 -299 85
rect -333 -17 -299 17
rect -333 -85 -299 -51
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 299 51 333 85
rect 299 -17 333 17
rect 299 -85 333 -51
<< poly >>
rect -287 100 -187 126
rect -129 100 -29 126
rect 29 100 129 126
rect 187 100 287 126
rect -287 -126 -187 -100
rect -129 -126 -29 -100
rect 29 -126 129 -100
rect 187 -126 287 -100
<< locali >>
rect -333 85 -299 104
rect -333 17 -299 19
rect -333 -19 -299 -17
rect -333 -104 -299 -85
rect -175 85 -141 104
rect -175 17 -141 19
rect -175 -19 -141 -17
rect -175 -104 -141 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 141 85 175 104
rect 141 17 175 19
rect 141 -19 175 -17
rect 141 -104 175 -85
rect 299 85 333 104
rect 299 17 333 19
rect 299 -19 333 -17
rect 299 -104 333 -85
<< viali >>
rect -333 51 -299 53
rect -333 19 -299 51
rect -333 -51 -299 -19
rect -333 -53 -299 -51
rect -175 51 -141 53
rect -175 19 -141 51
rect -175 -51 -141 -19
rect -175 -53 -141 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 141 51 175 53
rect 141 19 175 51
rect 141 -51 175 -19
rect 141 -53 175 -51
rect 299 51 333 53
rect 299 19 333 51
rect 299 -51 333 -19
rect 299 -53 333 -51
<< metal1 >>
rect -339 53 -293 100
rect -339 19 -333 53
rect -299 19 -293 53
rect -339 -19 -293 19
rect -339 -53 -333 -19
rect -299 -53 -293 -19
rect -339 -100 -293 -53
rect -181 53 -135 100
rect -181 19 -175 53
rect -141 19 -135 53
rect -181 -19 -135 19
rect -181 -53 -175 -19
rect -141 -53 -135 -19
rect -181 -100 -135 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 135 53 181 100
rect 135 19 141 53
rect 175 19 181 53
rect 135 -19 181 19
rect 135 -53 141 -19
rect 175 -53 181 -19
rect 135 -100 181 -53
rect 293 53 339 100
rect 293 19 299 53
rect 333 19 339 53
rect 293 -19 339 19
rect 293 -53 299 -19
rect 333 -53 339 -19
rect 293 -100 339 -53
<< end >>
