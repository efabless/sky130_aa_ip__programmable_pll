magic
tech sky130A
magscale 1 2
timestamp 1717691374
<< nwell >>
rect 568 1540 740 1632
rect 997 1540 1359 1906
rect 360 1404 1359 1540
rect 360 1394 1373 1404
rect 360 1347 2124 1394
rect 360 1258 2654 1347
rect 360 1243 2588 1258
rect 360 1230 2124 1243
rect 360 1172 1817 1230
rect 947 1157 1817 1172
rect 1589 791 1817 1157
<< poly >>
rect 1322 1907 1450 1955
<< locali >>
rect 1244 2437 1909 2523
rect 1244 2356 1330 2437
rect 1006 2270 1330 2356
rect 240 2050 370 2072
rect 240 2016 288 2050
rect 322 2016 370 2050
rect 240 1978 370 2016
rect 827 2008 1290 2048
rect 240 1944 288 1978
rect 322 1944 370 1978
rect 2495 1997 2759 2027
rect 2495 1996 2671 1997
rect 2495 1995 2589 1996
rect 2495 1961 2511 1995
rect 2545 1962 2589 1995
rect 2623 1963 2671 1996
rect 2705 1963 2759 1997
rect 2623 1962 2759 1963
rect 2545 1961 2759 1962
rect 1322 1950 1450 1955
rect 240 1922 370 1944
rect 1117 1949 1450 1950
rect 1117 1948 1412 1949
rect 1117 1914 1332 1948
rect 1366 1915 1412 1948
rect 1446 1915 1450 1949
rect 2495 1941 2759 1961
rect 1366 1914 1450 1915
rect 1322 1906 1450 1914
rect 2714 1726 2878 1796
rect 568 1337 740 1547
rect 1396 1354 1839 1383
rect 1396 1337 2014 1354
rect 398 1184 2509 1337
rect 800 1177 1026 1184
rect 837 1170 1026 1177
rect -88 568 107 604
rect 112 568 204 604
rect 150 506 374 510
rect 150 472 175 506
rect 209 472 249 506
rect 283 472 374 506
rect 150 470 374 472
rect 1709 327 1779 792
rect 2808 389 2878 1726
rect 2797 372 2902 389
rect 2797 338 2833 372
rect 2867 338 2902 372
rect 1709 291 1956 327
rect 2797 317 2902 338
rect 1709 289 1779 291
rect 1849 218 1907 228
rect 1849 184 1861 218
rect 1895 184 1907 218
rect 1849 174 1907 184
rect 1945 217 1987 221
rect 1945 183 1949 217
rect 1983 183 1987 217
rect 1945 180 1987 183
rect 2609 171 3361 214
rect 1219 -272 1280 99
rect 1219 -337 2696 -272
rect 1219 -371 2549 -337
rect 2583 -338 2696 -337
rect 2583 -371 2624 -338
rect 1219 -372 2624 -371
rect 2658 -372 2696 -338
rect 1219 -385 2696 -372
<< viali >>
rect 288 2016 322 2050
rect 288 1944 322 1978
rect 2511 1961 2545 1995
rect 2589 1962 2623 1996
rect 2671 1963 2705 1997
rect 1332 1914 1366 1948
rect 1412 1915 1446 1949
rect 175 472 209 506
rect 249 472 283 506
rect 2833 338 2867 372
rect 1861 184 1895 218
rect 1949 183 1983 217
rect 2549 -371 2583 -337
rect 2624 -372 2658 -338
<< metal1 >>
rect 14 2362 1111 2416
rect 1057 2072 1111 2362
rect 240 2050 370 2072
rect 240 2016 288 2050
rect 322 2016 370 2050
rect 1057 2018 1385 2072
rect 240 1978 370 2016
rect 240 1944 288 1978
rect 322 1944 370 1978
rect 1331 1963 1385 2018
rect 2495 1997 3203 2037
rect 2495 1996 2671 1997
rect 2495 1995 2589 1996
rect 240 1922 370 1944
rect 1305 1949 1464 1963
rect 1305 1948 1412 1949
rect 290 518 344 1922
rect 1305 1914 1332 1948
rect 1366 1915 1412 1948
rect 1446 1915 1464 1949
rect 2495 1961 2511 1995
rect 2545 1962 2589 1995
rect 2623 1963 2671 1996
rect 2705 1963 3203 1997
rect 2623 1962 3203 1963
rect 2545 1961 3203 1962
rect 2495 1924 3203 1961
rect 1366 1914 1464 1915
rect 1305 1905 1464 1914
rect 147 506 344 518
rect 147 472 175 506
rect 209 472 249 506
rect 283 472 344 506
rect 147 464 344 472
rect 2797 372 2902 389
rect 2797 338 2833 372
rect 2867 338 2902 372
rect 2797 317 2902 338
rect 2803 234 2868 317
rect 1848 218 2868 234
rect 1848 184 1861 218
rect 1895 217 2868 218
rect 1895 184 1949 217
rect 1848 183 1949 184
rect 1983 183 2868 217
rect 1848 169 2868 183
rect 3090 -272 3203 1924
rect 2526 -337 3203 -272
rect 2526 -371 2549 -337
rect 2583 -338 3203 -337
rect 2583 -371 2624 -338
rect 2526 -372 2624 -371
rect 2658 -372 3203 -338
rect 2526 -385 3203 -372
use AND_1  AND_1_0
timestamp 1717691374
transform 1 0 300 0 1 0
box -204 -132 1711 1174
use AND_1  AND_1_1
timestamp 1717691374
transform 1 0 1299 0 -1 2518
box -204 -132 1711 1174
use inverter_1  inverter_1_0
timestamp 1717691374
transform 1 0 386 0 -1 1950
box -72 -427 777 423
use OR_MAGIC  OR_MAGIC_0
timestamp 1717691374
transform 1 0 3843 0 1 -1096
box -2036 715 -1189 2359
<< labels >>
flabel locali s 2846 934 2846 934 0 FreeSans 2500 0 0 0 a4
flabel locali s 1744 450 1744 450 0 FreeSans 2500 0 0 0 a3
flabel locali s 1242 2028 1242 2028 0 FreeSans 2500 0 0 0 a1
flabel metal1 s 270 2038 270 2038 0 FreeSans 2500 0 0 0 SEL
flabel locali s 1352 1228 1352 1228 0 FreeSans 2500 0 0 0 VDD
flabel locali s 3317 189 3317 189 0 FreeSans 2500 0 0 0 VOUT
flabel locali s -18 580 -18 580 0 FreeSans 750 0 0 0 IN2
flabel metal1 s 84 2392 84 2392 0 FreeSans 750 0 0 0 IN1
flabel locali s 1222 2302 1222 2302 0 FreeSans 750 0 0 0 VSS
<< end >>
