magic
tech sky130A
magscale 1 2
timestamp 1726361494
<< pwell >>
rect -4222 1453 -4082 1548
rect -3591 1428 -3506 1523
<< psubdiff >>
rect -4196 1479 -4108 1522
rect -3565 1454 -3532 1497
<< locali >>
rect -4820 43955 -3786 44102
rect -4820 42553 -4688 43955
rect -3934 42553 -3786 43955
rect -4820 42470 -3786 42553
rect -2105 43971 -746 44258
rect -2105 42569 -1796 43971
rect -1042 42569 -746 43971
rect -3742 40390 -2527 40571
rect -3742 39564 -3582 40390
rect -2684 39564 -2527 40390
rect -3742 39356 -2527 39564
rect -16160 8555 -16024 8692
rect -15790 8555 -15654 8720
rect -15496 8555 -15355 8722
rect -16182 8439 -15355 8555
rect -16182 8117 -16054 8439
rect -15588 8210 -15355 8439
rect -15588 8117 -15367 8210
rect -16182 8044 -15367 8117
rect -15205 7856 -15069 8692
rect -19000 7720 -15069 7856
rect -14950 7153 -14814 8692
rect -19851 7017 -14814 7153
rect -14717 5489 -14581 8724
rect -19980 5353 -14581 5489
rect -14717 5310 -14581 5353
rect -14518 4472 -14382 8692
rect -9654 7738 -9468 9038
rect -2105 8544 -746 42569
rect 3428 9172 14566 9807
rect -20516 4336 -14382 4472
rect -13709 7552 -9468 7738
rect -6647 8380 -745 8544
rect -13709 2685 -13523 7552
rect -6647 7410 -6465 8380
rect -5567 7410 -745 8380
rect 3428 8200 4063 9172
rect 14586 8869 14773 8899
rect 14586 8763 14616 8869
rect 14722 8817 14773 8869
rect 14722 8764 15071 8817
rect 14722 8763 14773 8764
rect 6966 8709 7312 8756
rect 14586 8746 14773 8763
rect 6966 8531 7017 8709
rect 7267 8691 7312 8709
rect 15942 8691 15978 8805
rect 7267 8531 16005 8691
rect 16226 8688 16396 8743
rect 16226 8654 16266 8688
rect 16300 8654 16338 8688
rect 16372 8654 16396 8688
rect 16226 8605 16396 8654
rect 6966 8530 16005 8531
rect 6966 8466 7312 8530
rect 7289 8261 7635 8307
rect 16722 8261 16775 8824
rect 26753 8619 38073 8844
rect 7289 8250 16799 8261
rect 3375 8050 4103 8200
rect 3375 7656 3512 8050
rect 3906 7918 4103 8050
rect 7289 8072 7357 8250
rect 7535 8079 16799 8250
rect 7535 8072 7635 8079
rect 7289 8017 7635 8072
rect 3906 7659 8854 7918
rect 16664 7877 16961 7884
rect 14552 7821 14795 7846
rect 16664 7821 16687 7877
rect 14552 7793 16687 7821
rect 14552 7687 14612 7793
rect 14718 7687 16687 7793
rect 14552 7685 16687 7687
rect 3906 7656 4103 7659
rect 3375 7565 4103 7656
rect 14552 7642 14795 7685
rect 16664 7627 16687 7685
rect 16937 7627 16961 7877
rect 16664 7621 16961 7627
rect 26753 7793 27007 8619
rect 37625 7793 38073 8619
rect 26753 7623 38073 7793
rect -6647 7185 -745 7410
rect -12975 6803 -11404 6943
rect -12975 6735 -2388 6803
rect -12975 5693 -12793 6735
rect -11679 6667 -2388 6735
rect -11679 5769 -3460 6667
rect -2562 5769 -2388 6667
rect -11679 5693 -2388 5769
rect -12975 5558 -2388 5693
rect -12975 5372 -11404 5558
rect -2105 4551 -746 7185
rect 19201 6977 19643 7085
rect 14997 6931 15211 6970
rect 19201 6931 19319 6977
rect 14997 6910 19319 6931
rect 14997 6804 15045 6910
rect 15151 6807 19319 6910
rect 15151 6804 15211 6807
rect 14997 6756 15211 6804
rect 19201 6727 19319 6807
rect 19569 6931 19643 6977
rect 22939 6990 23303 7116
rect 22939 6931 23024 6990
rect 19569 6807 23024 6931
rect 19569 6727 19643 6807
rect 16227 6562 16406 6623
rect 19201 6620 19643 6727
rect 22939 6740 23024 6807
rect 23202 6740 23303 6990
rect 22939 6666 23303 6740
rect 12164 6549 16406 6562
rect 12164 6515 16262 6549
rect 16296 6515 16334 6549
rect 16368 6515 16406 6549
rect 12164 6480 16406 6515
rect 16227 6444 16406 6480
rect 14443 6172 14691 6213
rect 14443 6151 14508 6172
rect 12023 6066 14508 6151
rect 14614 6066 14691 6172
rect 12023 6038 14691 6066
rect 12023 5692 12136 6038
rect 14443 6016 14691 6038
rect 13866 5924 14130 5964
rect 13866 5898 13910 5924
rect 12465 5746 13910 5898
rect 14088 5746 14130 5924
rect 12465 5641 14130 5746
rect 12470 5556 12504 5641
rect 18791 5522 19168 5573
rect 18791 5272 18862 5522
rect 19112 5272 19168 5522
rect 18791 5216 19168 5272
rect 23929 4724 61121 4741
rect 2866 4551 3250 4560
rect -2197 4458 12654 4551
rect -2197 4208 2928 4458
rect 3178 4208 12654 4458
rect -2197 4085 12654 4208
rect 23929 4330 41740 4724
rect 44510 4367 61121 4724
rect 44510 4330 98798 4367
rect 23929 4290 98798 4330
rect 15817 4168 16331 4171
rect 23929 4168 24380 4290
rect 14819 4098 24380 4168
rect 14819 3776 15899 4098
rect 16221 3776 24380 4098
rect 14819 3717 24380 3776
rect 26583 3803 38866 3886
rect 14819 3692 15270 3717
rect -13207 3541 15270 3692
rect 21388 3567 21612 3717
rect -13207 3497 3593 3541
rect -13207 3391 -13067 3497
rect -9289 3391 3593 3497
rect -13207 3363 3593 3391
rect 3771 3363 15270 3541
rect 26583 3553 26677 3803
rect 38663 3553 38866 3803
rect 26583 3483 38866 3553
rect -13207 3241 15270 3363
rect -5845 2711 -5539 2764
rect -5845 2685 -5790 2711
rect -13709 2548 -5790 2685
rect -5845 2533 -5790 2548
rect -5612 2533 -5539 2711
rect -5845 2483 -5539 2533
rect -13326 2292 -9322 2305
rect -13326 2186 -13321 2292
rect -9327 2186 -9322 2292
rect -2198 2241 -1747 3241
rect 6011 2400 6354 3241
rect 11748 2486 12550 3241
rect 41815 3199 44205 3238
rect 51135 3226 51730 4290
rect 53312 3230 53907 4290
rect 55261 3230 55856 4290
rect 57618 3209 58213 4290
rect 18156 3138 18330 3181
rect 18156 3032 18185 3138
rect 18291 3110 18330 3138
rect 41815 3165 41866 3199
rect 41900 3165 41938 3199
rect 41972 3165 42010 3199
rect 42044 3165 42082 3199
rect 42116 3165 42154 3199
rect 42188 3165 42226 3199
rect 42260 3165 42298 3199
rect 42332 3165 42370 3199
rect 42404 3165 42442 3199
rect 42476 3165 42514 3199
rect 42548 3165 42586 3199
rect 42620 3165 42658 3199
rect 42692 3165 42730 3199
rect 42764 3165 42802 3199
rect 42836 3165 42874 3199
rect 42908 3165 42946 3199
rect 42980 3165 43018 3199
rect 43052 3165 43090 3199
rect 43124 3165 43162 3199
rect 43196 3165 43234 3199
rect 43268 3165 43306 3199
rect 43340 3165 43378 3199
rect 43412 3165 43450 3199
rect 43484 3165 43522 3199
rect 43556 3165 43594 3199
rect 43628 3165 43666 3199
rect 43700 3165 43738 3199
rect 43772 3165 43810 3199
rect 43844 3165 43882 3199
rect 43916 3165 43954 3199
rect 43988 3165 44026 3199
rect 44060 3165 44098 3199
rect 44132 3165 44205 3199
rect 18291 3036 19662 3110
rect 41815 3072 44205 3165
rect 18291 3032 18330 3036
rect 18156 2985 18330 3032
rect 19567 2877 19632 2878
rect 19563 2855 19636 2877
rect 19563 2821 19582 2855
rect 19616 2821 19636 2855
rect 22316 2856 22554 2900
rect 19563 2800 19636 2821
rect 19826 2837 20301 2844
rect 19826 2803 19830 2837
rect 19864 2803 19902 2837
rect 19936 2803 19974 2837
rect 20008 2803 20046 2837
rect 20080 2803 20118 2837
rect 20152 2803 20190 2837
rect 20224 2803 20262 2837
rect 20296 2803 20301 2837
rect 19341 2564 19481 2579
rect 18629 2540 18739 2549
rect 19341 2540 19401 2564
rect 18629 2530 19401 2540
rect 19435 2530 19481 2564
rect 18629 2511 19481 2530
rect 18629 2477 18667 2511
rect 18701 2492 19481 2511
rect 18701 2477 19401 2492
rect 18629 2458 19401 2477
rect 19435 2458 19481 2492
rect 18629 2447 19481 2458
rect 18629 2441 18739 2447
rect 19341 2444 19481 2447
rect -13326 2173 -9322 2186
rect 7054 2043 7303 2079
rect 3222 1884 4073 1923
rect 3500 1595 3875 1654
rect 4034 1638 4073 1884
rect 7054 1865 7089 2043
rect 7267 1865 7303 2043
rect 7054 1845 7303 1865
rect 3500 1574 3553 1595
rect -5642 1514 -5574 1521
rect -5779 1492 -5574 1514
rect -22664 1391 -13491 1425
rect -5779 1386 -5730 1492
rect -5624 1386 -5574 1492
rect -4212 1517 -4099 1535
rect -4212 1483 -4169 1517
rect -4135 1483 -4099 1517
rect -4212 1461 -4099 1483
rect -3565 1493 -3532 1497
rect -3565 1492 -3098 1493
rect -5779 1352 -5574 1386
rect -5779 1299 -5642 1352
rect -13321 689 -6175 692
rect -13321 583 -13293 689
rect -6203 680 -6175 689
rect -4187 680 -4102 1461
rect -3565 1458 -3512 1492
rect -3478 1458 -3440 1492
rect -3406 1458 -3368 1492
rect -3334 1458 -3296 1492
rect -3262 1458 -3224 1492
rect -3190 1458 -3152 1492
rect -3118 1458 -3098 1492
rect -3565 1454 -3532 1458
rect 2935 1345 3553 1574
rect 3803 1345 3875 1595
rect 3990 1624 4106 1638
rect 3990 1590 4029 1624
rect 4063 1590 4106 1624
rect 3990 1552 4106 1590
rect 3990 1518 4029 1552
rect 4063 1518 4106 1552
rect 3990 1499 4106 1518
rect 4626 1517 4768 1644
rect 7096 1568 7234 1845
rect 15522 1770 15742 1833
rect 15522 1707 15576 1770
rect 7337 1640 7470 1680
rect 15184 1673 15576 1707
rect 7337 1606 7381 1640
rect 7415 1606 7470 1640
rect 2935 1319 3875 1345
rect 3500 1279 3875 1319
rect 4196 1465 4326 1504
rect 4196 1431 4245 1465
rect 4279 1431 4326 1465
rect -6203 595 -4102 680
rect -6203 583 -6175 595
rect -13321 581 -6175 583
rect -18039 534 -17604 565
rect -18039 457 -17981 534
rect -22512 356 -17981 457
rect -17659 457 -17604 534
rect -6543 457 -5591 465
rect -17659 431 -5591 457
rect -17659 356 -6478 431
rect -22512 325 -6478 356
rect -5652 325 -5591 431
rect -22512 320 -5591 325
rect -6543 299 -5591 320
rect -3695 212 -3643 1090
rect 3563 1017 3725 1039
rect 3563 978 3591 1017
rect 3231 939 3591 978
rect 3563 911 3591 939
rect 3697 911 3725 1017
rect 3563 885 3725 911
rect -2404 576 -2375 608
rect 4196 595 4326 1431
rect 4600 1468 4817 1517
rect 4600 1434 4649 1468
rect 4683 1434 4721 1468
rect 4755 1434 4817 1468
rect 4600 1392 4817 1434
rect 7029 1506 7278 1568
rect 7337 1562 7470 1606
rect 15522 1664 15576 1673
rect 15682 1664 15742 1770
rect 15522 1597 15742 1664
rect 7029 1400 7121 1506
rect 7227 1400 7278 1506
rect 7029 1334 7278 1400
rect 4415 1243 4467 1266
rect 4388 1205 4549 1243
rect 19567 1242 19632 2800
rect 19826 2796 20301 2803
rect 22316 2750 22385 2856
rect 22491 2750 22554 2856
rect 22316 2711 22554 2750
rect 26688 2858 26963 2876
rect 26688 2820 28014 2858
rect 26688 2714 26734 2820
rect 26912 2714 28014 2820
rect 22376 2297 22532 2711
rect 26688 2669 28014 2714
rect 26688 2653 26963 2669
rect 58711 2522 58930 2597
rect 58711 2484 58776 2522
rect 50510 2421 50749 2467
rect 58493 2450 58776 2484
rect 25061 2314 25333 2372
rect 25061 2297 25092 2314
rect 22376 2141 25092 2297
rect 25061 2136 25092 2141
rect 25270 2136 25333 2314
rect 25061 2085 25333 2136
rect 25955 2313 26111 2333
rect 25955 2135 25980 2313
rect 26086 2273 26111 2313
rect 26086 2145 27166 2273
rect 50510 2243 50542 2421
rect 50720 2243 50749 2421
rect 58711 2416 58776 2450
rect 58882 2416 58930 2522
rect 58711 2334 58930 2416
rect 50510 2215 50749 2243
rect 26086 2135 26111 2145
rect 25955 2116 26111 2135
rect 4388 1099 4417 1205
rect 4523 1099 4549 1205
rect 4388 1066 4549 1099
rect 19404 1241 19736 1242
rect 19404 1164 19770 1241
rect 19404 986 19522 1164
rect 19700 986 19770 1164
rect 5730 747 6208 775
rect 5730 713 5767 747
rect 5801 713 5839 747
rect 5873 713 5911 747
rect 5945 713 5983 747
rect 6017 713 6055 747
rect 6089 713 6127 747
rect 6161 713 6208 747
rect 8203 744 8571 936
rect 9394 744 9762 971
rect 10640 744 11008 885
rect 12204 744 12572 911
rect 13329 744 13697 920
rect 14498 744 14866 947
rect 19404 943 19770 986
rect 19404 744 19742 943
rect 5730 686 6208 713
rect 8089 595 19742 744
rect -2404 364 -2075 576
rect 3030 382 19742 595
rect -22962 160 -3643 212
rect -3192 35 -2075 364
rect 15818 275 16268 345
rect 5857 270 16268 275
rect 3985 219 4186 265
rect 3985 213 4030 219
rect -1806 113 4030 213
rect 4136 113 4186 219
rect -1806 100 4186 113
rect -13197 -205 -7163 -135
rect -3192 -153 -2863 35
rect -13197 -383 -13046 -205
rect -7324 -274 -7163 -205
rect -7324 -304 -5720 -274
rect -7324 -338 -6020 -304
rect -5986 -338 -5948 -304
rect -5914 -338 -5876 -304
rect -5842 -338 -5804 -304
rect -5770 -338 -5720 -304
rect -7324 -378 -5720 -338
rect -7324 -383 -7163 -378
rect -13197 -453 -7163 -383
rect -25553 -704 -25165 -654
rect -22114 -677 -5221 -603
rect -25553 -954 -25480 -704
rect -25230 -806 -25165 -704
rect -5976 -806 -5800 -784
rect -25230 -807 -5800 -806
rect -25230 -943 -5939 -807
rect -25230 -954 -25165 -943
rect -25553 -1050 -25165 -954
rect -5976 -985 -5939 -943
rect -5833 -985 -5800 -807
rect -5038 -876 -4568 -869
rect -5038 -910 -5036 -876
rect -5002 -910 -4964 -876
rect -4930 -910 -4892 -876
rect -4858 -910 -4820 -876
rect -4786 -910 -4748 -876
rect -4714 -910 -4676 -876
rect -4642 -910 -4604 -876
rect -4570 -910 -4568 -876
rect -5038 -916 -4568 -910
rect -5976 -1005 -5800 -985
rect -4169 -1022 -4077 -1007
rect -4169 -1056 -4140 -1022
rect -4106 -1056 -4077 -1022
rect -4169 -1070 -4077 -1056
rect -1806 -1962 -1693 100
rect 3985 76 4186 100
rect 5857 162 15880 270
rect 4383 -36 4585 -15
rect -1577 -62 4585 -36
rect -1577 -85 4424 -62
rect -1581 -117 4424 -85
rect -1581 -295 -1548 -117
rect -1370 -168 4424 -117
rect 4530 -168 4585 -62
rect -1370 -175 4585 -168
rect -1370 -295 -1323 -175
rect 4383 -213 4585 -175
rect 5857 -88 5919 162
rect 6169 -88 15880 162
rect 5857 -124 15880 -88
rect 16202 -124 16268 270
rect 21288 224 21541 1919
rect 21915 199 22067 1925
rect 46637 1919 46961 1997
rect 46637 1741 46686 1919
rect 46864 1741 46961 1919
rect 46637 1686 46961 1741
rect 47896 1953 48216 1992
rect 47896 1703 47959 1953
rect 48137 1900 48216 1953
rect 50541 1900 50720 2215
rect 48137 1721 50720 1900
rect 48137 1703 48216 1721
rect 47896 1636 48216 1703
rect 22419 1248 25673 1356
rect 22419 926 22486 1248
rect 22808 926 25673 1248
rect 22419 876 25673 926
rect 51870 824 52157 1672
rect 60670 1398 98798 4290
rect 60670 1310 61121 1398
rect 47592 537 52157 824
rect 53362 859 64533 1310
rect 53362 326 54000 859
rect 54759 326 55397 859
rect 56173 343 56811 859
rect 57259 326 57897 859
rect 5857 -176 16268 -124
rect 5877 -291 6211 -176
rect -1581 -342 -1323 -295
rect 8303 -302 8754 -176
rect 9891 -302 10342 -176
rect 11432 -321 11883 -176
rect 12650 -283 13101 -176
rect 13848 -283 14299 -176
rect 15818 -209 16268 -176
rect 60613 -382 61078 -338
rect 60613 -427 60645 -382
rect 58332 -445 60645 -427
rect 19992 -518 20496 -512
rect 19992 -552 20011 -518
rect 20045 -552 20083 -518
rect 20117 -552 20155 -518
rect 20189 -552 20227 -518
rect 20261 -552 20299 -518
rect 20333 -552 20371 -518
rect 20405 -552 20443 -518
rect 20477 -552 20496 -518
rect 19992 -557 20496 -552
rect 50434 -572 50725 -478
rect 47758 -600 50725 -572
rect 3281 -699 3574 -645
rect 3281 -877 3355 -699
rect 3533 -745 3574 -699
rect 47758 -706 47797 -600
rect 47903 -632 50725 -600
rect 58324 -618 60645 -445
rect 60613 -632 60645 -618
rect 61039 -632 61078 -382
rect 47903 -706 50588 -632
rect 60613 -669 61078 -632
rect 47758 -726 50588 -706
rect 3533 -819 4361 -745
rect 47758 -752 47953 -726
rect 3533 -877 3574 -819
rect 3281 -911 3574 -877
rect 16101 -928 16445 -871
rect 4545 -1022 4984 -1020
rect 16101 -1021 16129 -928
rect 4545 -1056 4567 -1022
rect 4601 -1056 4639 -1022
rect 4673 -1056 4711 -1022
rect 4745 -1056 4783 -1022
rect 4817 -1056 4855 -1022
rect 4889 -1056 4927 -1022
rect 4961 -1056 4984 -1022
rect 4545 -1058 4984 -1056
rect 7334 -1131 7443 -1093
rect 15047 -1127 16129 -1021
rect 7334 -1165 7372 -1131
rect 7406 -1165 7443 -1131
rect 7334 -1207 7443 -1165
rect 16101 -1178 16129 -1127
rect 16379 -1178 16445 -928
rect 16101 -1228 16445 -1178
rect 19836 -1048 20098 -916
rect 19836 -1226 19870 -1048
rect 20048 -1129 20098 -1048
rect 20048 -1226 20093 -1129
rect 19836 -1279 20093 -1226
rect -26391 -2075 -1693 -1962
rect 8336 -1966 8557 -1837
rect 9274 -1966 9547 -1837
rect 10255 -1966 10528 -1871
rect 11457 -1966 11730 -1845
rect 12412 -1966 12685 -1879
rect 13206 -1966 13479 -1845
rect 13931 -1966 14204 -1845
rect 26281 -1966 26638 -1361
rect 4310 -2187 4465 -2171
rect 4310 -2204 4333 -2187
rect -26307 -2293 4333 -2204
rect 4439 -2293 4465 -2187
rect -26307 -2300 4465 -2293
rect 4310 -2309 4465 -2300
rect 8168 -2323 26638 -1966
rect 46864 -1737 47369 -1268
rect 52463 -1737 52968 -1175
rect 55332 -1517 55783 -1516
rect 56669 -1517 57120 -1516
rect 57856 -1517 58307 -1516
rect 64082 -1517 64533 859
rect 46864 -2109 52968 -1737
rect -1585 -2393 -1283 -2369
rect -26253 -2419 -1283 -2393
rect -26253 -2525 -1533 -2419
rect -1355 -2525 -1283 -2419
rect 46864 -2431 46934 -2109
rect 47256 -2242 52968 -2109
rect 53892 -1968 64533 -1517
rect 47256 -2431 47369 -2242
rect 46864 -2515 47369 -2431
rect -26253 -2533 -1283 -2525
rect -1585 -2584 -1283 -2533
rect 3196 -2596 3624 -2539
rect 3196 -2628 3300 -2596
rect -26211 -2846 3300 -2628
rect 3550 -2846 3624 -2596
rect 53892 -2712 54343 -1968
rect 55332 -2712 55783 -1968
rect 56669 -2731 57120 -1968
rect 57856 -2731 58307 -1968
rect 64082 -2655 64533 -1968
rect -26211 -2873 3624 -2846
rect 3196 -2900 3624 -2873
rect 15440 -2934 15853 -2842
rect -26114 -2967 15853 -2934
rect -26114 -3145 15515 -2967
rect 15765 -3145 15853 -2967
rect -26114 -3188 15853 -3145
rect 15440 -3211 15853 -3188
rect 87785 -3285 88210 -3189
rect 87785 -3288 87949 -3285
rect 16088 -3296 16483 -3292
rect -26140 -3356 16483 -3296
rect -26140 -3534 16158 -3356
rect 16408 -3534 16483 -3356
rect -26140 -3586 16483 -3534
rect 16088 -3623 16483 -3586
rect 48966 -3402 49277 -3371
rect 48966 -3652 49025 -3402
rect 49203 -3547 49277 -3402
rect 62387 -3378 62911 -3375
rect 62387 -3385 62884 -3378
rect 61873 -3432 62067 -3407
rect 58166 -3442 62067 -3432
rect 62387 -3419 62412 -3385
rect 62446 -3419 62484 -3385
rect 62518 -3419 62556 -3385
rect 62590 -3419 62628 -3385
rect 62662 -3419 62700 -3385
rect 62734 -3419 62772 -3385
rect 62806 -3419 62844 -3385
rect 62878 -3419 62884 -3385
rect 62387 -3428 62884 -3419
rect 62908 -3428 62911 -3378
rect 62387 -3436 62911 -3428
rect 65127 -3386 87949 -3288
rect 65127 -3420 65205 -3386
rect 65239 -3420 65277 -3386
rect 65311 -3420 87949 -3386
rect 58166 -3456 61914 -3442
rect 58163 -3476 61914 -3456
rect 61948 -3476 61986 -3442
rect 62020 -3474 62067 -3442
rect 65127 -3463 87949 -3420
rect 88127 -3463 88210 -3285
rect 62020 -3476 62096 -3474
rect 58163 -3490 62096 -3476
rect 58332 -3508 62096 -3490
rect 65127 -3507 88210 -3463
rect 61873 -3516 62067 -3508
rect 49203 -3608 50651 -3547
rect 87785 -3581 88210 -3507
rect 49203 -3652 49277 -3608
rect 48966 -3697 49277 -3652
rect 62432 -3844 62779 -3786
rect 62432 -4094 62474 -3844
rect 62724 -4094 62779 -3844
rect 62432 -4139 62779 -4094
rect 17293 -4336 17906 -4235
rect 16975 -4345 17906 -4336
rect 16975 -4354 17422 -4345
rect -26205 -4739 17422 -4354
rect 17816 -4739 17906 -4345
rect -26205 -4766 17906 -4739
rect 17293 -4848 17906 -4766
rect 46778 -4698 47398 -4670
rect 52571 -4698 53148 -4252
rect 95829 -4698 98798 1398
rect 46778 -4775 92959 -4698
rect 17978 -5013 18468 -4849
rect -26311 -5014 18468 -5013
rect -26311 -5336 18053 -5014
rect 18375 -5336 18468 -5014
rect 46778 -5169 46926 -4775
rect 47248 -4841 92959 -4775
rect 47248 -4947 61332 -4841
rect 61438 -4947 92959 -4841
rect 47248 -5063 92959 -4947
rect 47248 -5169 90388 -5063
rect 46778 -5275 90388 -5169
rect 46778 -5304 47412 -5275
rect -26311 -5399 18468 -5336
rect 17978 -5437 18468 -5399
rect 18534 -5592 18990 -5587
rect 18534 -5664 18565 -5592
rect -26321 -6058 18565 -5664
rect 18959 -6058 18990 -5592
rect -26321 -6062 18990 -6058
rect -26321 -6098 18704 -6062
rect 18949 -6346 19611 -6293
rect -26653 -6417 19611 -6346
rect -26653 -6739 19129 -6417
rect 19451 -6739 19611 -6417
rect -26653 -6787 19611 -6739
rect 18949 -6850 19611 -6787
rect 19665 -7100 20295 -7025
rect -26746 -7122 20295 -7100
rect -26746 -7516 19786 -7122
rect 20180 -7516 20295 -7122
rect -26746 -7593 20295 -7516
rect 19665 -7634 20295 -7593
rect 70077 -7257 90388 -5275
rect 92654 -7257 92959 -5063
rect 70077 -7667 92959 -7257
rect 95743 -7667 98798 -4698
rect 70077 -7803 73046 -7667
rect 81551 -7803 84520 -7667
rect -31467 -8993 -30570 -8797
rect -31467 -9060 -31392 -8993
rect -34283 -9713 -31392 -9060
rect -31467 -9819 -31392 -9713
rect -30710 -9060 -30570 -8993
rect 58913 -9030 59860 -8831
rect 58913 -9060 59146 -9030
rect -30710 -9712 59146 -9060
rect 59756 -9712 59860 -9030
rect -30710 -9713 59860 -9712
rect -30710 -9819 -30570 -9713
rect -31467 -10014 -30570 -9819
rect 58913 -9909 59860 -9713
rect 60423 -9806 61454 -9617
rect -29173 -9983 -28472 -9982
rect 60423 -9983 60630 -9806
rect -29347 -10522 60630 -9983
rect -29564 -10560 60630 -10522
rect 61312 -10560 61454 -9806
rect -29564 -10681 61454 -10560
rect -29564 -10704 -28286 -10681
rect -29564 -11602 -29366 -10704
rect -28468 -11602 -28286 -10704
rect 60423 -10731 61454 -10681
rect -29564 -11751 -28286 -11602
rect -26907 -11088 -25983 -10980
rect -24373 -11062 -23278 -10959
rect -24373 -11088 -24141 -11062
rect -26907 -11091 -24141 -11088
rect -29173 -12595 -28472 -11751
rect -26907 -11773 -26776 -11091
rect -26094 -11672 -24141 -11091
rect -23459 -11672 -23278 -11062
rect -26094 -11732 -23278 -11672
rect -26094 -11773 -25983 -11732
rect -26907 -11904 -25983 -11773
rect -24373 -11840 -23278 -11732
rect -6611 -11268 -5937 -11153
rect -6611 -11806 -6514 -11268
rect -6048 -11274 -5937 -11268
rect 61366 -11264 62272 -11116
rect 61366 -11274 61636 -11264
rect -6048 -11730 61636 -11274
rect 62174 -11730 62272 -11264
rect -6048 -11806 62272 -11730
rect -6611 -11839 62272 -11806
rect -6611 -11894 -5937 -11839
rect 61366 -11971 62272 -11839
rect 62246 -12546 63072 -12441
rect -34369 -13296 -28472 -12595
rect -26996 -12584 63072 -12546
rect -26996 -13050 62412 -12584
rect 62950 -13050 63072 -12584
rect 95829 -12668 98798 -7667
rect -26996 -13121 63072 -13050
rect -26996 -13991 -26421 -13121
rect 62246 -13180 63072 -13121
rect -34505 -14566 -26421 -13991
rect -25931 -14188 -24870 -14108
rect -25931 -14352 -7185 -14188
rect -25931 -14746 -25638 -14352
rect -25028 -14746 -7185 -14352
rect -25931 -14808 -7185 -14746
rect -25931 -14876 -24870 -14808
rect -12874 -15051 -7870 -14969
rect -12874 -15157 -12791 -15051
rect -8005 -15157 -7870 -15051
rect -12874 -15238 -7870 -15157
rect -34293 -15952 -15114 -15892
rect -7536 -15913 -7185 -14808
rect 81378 -15816 98798 -12668
rect -34293 -15986 -15075 -15952
rect -34293 -16022 -15114 -15986
rect -14106 -18273 -13756 -16708
rect -11883 -18273 -11533 -16708
rect -9810 -18248 -9410 -16724
rect 81378 -16770 84526 -15816
rect 90329 -17748 91702 -17504
rect 90329 -18041 90552 -17748
rect 88428 -18574 90552 -18041
rect 91450 -18574 91702 -17748
rect 88428 -18579 91702 -18574
rect 90329 -18877 91702 -18579
rect -25664 -22895 -25039 -22779
rect -25664 -23289 -25536 -22895
rect -25142 -22999 -25039 -22895
rect -25142 -23185 -24246 -22999
rect -25142 -23289 -25039 -23185
rect -25664 -23404 -25039 -23289
rect -32565 -28049 -24427 -27913
rect -32538 -28248 -24481 -28112
rect 95829 -28339 98798 -15816
rect -32538 -28481 -24400 -28345
rect -32592 -28736 -24400 -28600
rect -33001 -29027 -24533 -28886
rect -32755 -29321 -24481 -29185
rect -32917 -29691 -24454 -29555
rect 83333 -31308 98798 -28339
rect -32225 -33190 -26140 -32972
rect -26347 -33893 -26140 -33190
rect 83333 -33215 86302 -31308
rect 90604 -34284 92221 -33888
rect 90604 -34632 90887 -34284
rect 88763 -35110 90887 -34632
rect 91785 -35110 92221 -34284
rect 88763 -35170 92221 -35110
rect 90604 -35414 92221 -35170
rect -25408 -35732 -23381 -35460
rect -25408 -36532 -23381 -36260
rect -27604 -37050 -27464 -37004
rect -27604 -37084 -27563 -37050
rect -27529 -37084 -27464 -37050
rect -27604 -37122 -27464 -37084
rect -27604 -37156 -27563 -37122
rect -27529 -37156 -27464 -37122
rect -27604 -37174 -27464 -37156
rect -27604 -37194 -26938 -37174
rect -27604 -37228 -27563 -37194
rect -27529 -37228 -26938 -37194
rect -27604 -37266 -26938 -37228
rect -27604 -37300 -27563 -37266
rect -27529 -37300 -26938 -37266
rect -27604 -37338 -26938 -37300
rect -27604 -37372 -27563 -37338
rect -27529 -37351 -26938 -37338
rect -27529 -37372 -27464 -37351
rect -27604 -37410 -27464 -37372
rect -27604 -37444 -27563 -37410
rect -27529 -37444 -27464 -37410
rect -27604 -37482 -27464 -37444
rect -27604 -37516 -27563 -37482
rect -27529 -37516 -27464 -37482
rect -27604 -37554 -27464 -37516
rect -27604 -37588 -27563 -37554
rect -27529 -37588 -27464 -37554
rect -27604 -37626 -27464 -37588
rect -25408 -37593 -23381 -37321
rect -27604 -37660 -27563 -37626
rect -27529 -37660 -27464 -37626
rect -27604 -37685 -27464 -37660
rect -27604 -37698 -26953 -37685
rect -27604 -37732 -27563 -37698
rect -27529 -37732 -26953 -37698
rect -27604 -37770 -26953 -37732
rect -27604 -37804 -27563 -37770
rect -27529 -37804 -26953 -37770
rect -27604 -37842 -26953 -37804
rect -27604 -37876 -27563 -37842
rect -27529 -37862 -26953 -37842
rect -27529 -37876 -27464 -37862
rect -27604 -37914 -27464 -37876
rect -27604 -37948 -27563 -37914
rect -27529 -37948 -27464 -37914
rect -27604 -37986 -27464 -37948
rect -27604 -38020 -27563 -37986
rect -27529 -38020 -27464 -37986
rect -27604 -38058 -27464 -38020
rect -27604 -38092 -27563 -38058
rect -27529 -38092 -27464 -38058
rect -27604 -38130 -27464 -38092
rect -27604 -38164 -27563 -38130
rect -27529 -38164 -27464 -38130
rect -27604 -38202 -27464 -38164
rect -27604 -38236 -27563 -38202
rect -27529 -38236 -27464 -38202
rect -27604 -38274 -27464 -38236
rect -27604 -38308 -27563 -38274
rect -27529 -38300 -27464 -38274
rect -27529 -38308 -26975 -38300
rect -27604 -38346 -26975 -38308
rect -27604 -38380 -27563 -38346
rect -27529 -38380 -26975 -38346
rect -27604 -38418 -26975 -38380
rect -27604 -38452 -27563 -38418
rect -27529 -38452 -26975 -38418
rect -27604 -38477 -26975 -38452
rect -27604 -38490 -27464 -38477
rect -27604 -38524 -27563 -38490
rect -27529 -38524 -27464 -38490
rect -27604 -38562 -27464 -38524
rect -27604 -38596 -27563 -38562
rect -27529 -38596 -27464 -38562
rect -27604 -38634 -27464 -38596
rect -27604 -38668 -27563 -38634
rect -27529 -38668 -27464 -38634
rect -27604 -38706 -27464 -38668
rect -27604 -38740 -27563 -38706
rect -27529 -38740 -27464 -38706
rect -27604 -38778 -27464 -38740
rect -27604 -38812 -27563 -38778
rect -27529 -38812 -27464 -38778
rect -27604 -38850 -27464 -38812
rect -27604 -38884 -27563 -38850
rect -27529 -38884 -27464 -38850
rect -27604 -38922 -27464 -38884
rect -20537 -38893 -20422 -38680
rect -27604 -38956 -27563 -38922
rect -27529 -38956 -27464 -38922
rect -27604 -38994 -27464 -38956
rect -27604 -39028 -27563 -38994
rect -27529 -39028 -27464 -38994
rect -27604 -39066 -27464 -39028
rect -27604 -39100 -27563 -39066
rect -27529 -39092 -27464 -39066
rect -24450 -39008 -20422 -38893
rect -27529 -39100 -26953 -39092
rect -27604 -39138 -26953 -39100
rect -27604 -39172 -27563 -39138
rect -27529 -39172 -26953 -39138
rect -27604 -39210 -26953 -39172
rect -27604 -39244 -27563 -39210
rect -27529 -39244 -26953 -39210
rect -27604 -39269 -26953 -39244
rect -27604 -39282 -27464 -39269
rect -27604 -39316 -27563 -39282
rect -27529 -39316 -27464 -39282
rect -27604 -39354 -27464 -39316
rect -27604 -39388 -27563 -39354
rect -27529 -39388 -27464 -39354
rect -27604 -39426 -27464 -39388
rect -27604 -39460 -27563 -39426
rect -27529 -39460 -27464 -39426
rect -27604 -39498 -27464 -39460
rect -27604 -39532 -27563 -39498
rect -27529 -39532 -27464 -39498
rect -27604 -39570 -27464 -39532
rect -27604 -39604 -27563 -39570
rect -27529 -39604 -27464 -39570
rect -27604 -39642 -27464 -39604
rect -27604 -39676 -27563 -39642
rect -27529 -39676 -27464 -39642
rect -27604 -39714 -27464 -39676
rect -27604 -39748 -27563 -39714
rect -27529 -39748 -27464 -39714
rect -27604 -39786 -27464 -39748
rect -27604 -39820 -27563 -39786
rect -27529 -39820 -27464 -39786
rect -27604 -39858 -27464 -39820
rect -27604 -39892 -27563 -39858
rect -27529 -39892 -27464 -39858
rect -27604 -39930 -27464 -39892
rect -27604 -39964 -27563 -39930
rect -27529 -39964 -27464 -39930
rect -27604 -39973 -27464 -39964
rect -27604 -40002 -26953 -39973
rect -27604 -40036 -27563 -40002
rect -27529 -40036 -26953 -40002
rect -27604 -40074 -26953 -40036
rect -27604 -40108 -27563 -40074
rect -27529 -40108 -26953 -40074
rect -27604 -40146 -26953 -40108
rect -27604 -40180 -27563 -40146
rect -27529 -40150 -26953 -40146
rect -27529 -40180 -27464 -40150
rect -27604 -40218 -27464 -40180
rect -27604 -40252 -27563 -40218
rect -27529 -40252 -27464 -40218
rect -27604 -40290 -27464 -40252
rect -27604 -40324 -27563 -40290
rect -27529 -40324 -27464 -40290
rect -27604 -40362 -27464 -40324
rect -27604 -40396 -27563 -40362
rect -27529 -40396 -27464 -40362
rect -27604 -40434 -27464 -40396
rect -27604 -40468 -27563 -40434
rect -27529 -40468 -27464 -40434
rect -27604 -40506 -27464 -40468
rect -27604 -40540 -27563 -40506
rect -27529 -40540 -27464 -40506
rect -27604 -40578 -27464 -40540
rect -27604 -40612 -27563 -40578
rect -27529 -40612 -27464 -40578
rect -27604 -40650 -27464 -40612
rect -27604 -40684 -27563 -40650
rect -27529 -40684 -27464 -40650
rect -27604 -40722 -27464 -40684
rect -27604 -40756 -27563 -40722
rect -27529 -40756 -27464 -40722
rect -27604 -40794 -27464 -40756
rect -27604 -40828 -27563 -40794
rect -27529 -40795 -27464 -40794
rect -27529 -40828 -26953 -40795
rect -27604 -40866 -26953 -40828
rect -27604 -40900 -27563 -40866
rect -27529 -40900 -26953 -40866
rect -27604 -40938 -26953 -40900
rect -27604 -40972 -27563 -40938
rect -27529 -40972 -26953 -40938
rect -27604 -41010 -27464 -40972
rect -27604 -41044 -27563 -41010
rect -27529 -41044 -27464 -41010
rect -27604 -41082 -27464 -41044
rect -27604 -41116 -27563 -41082
rect -27529 -41116 -27464 -41082
rect -27604 -41184 -27464 -41116
rect -26388 -41420 -26202 -41401
rect -26388 -44174 -26195 -41420
rect -25977 -42849 -25639 -42789
rect -25977 -43027 -25880 -42849
rect -25702 -42872 -25639 -42849
rect -24450 -42872 -24335 -39008
rect -25702 -42987 -24335 -42872
rect -25702 -43027 -25639 -42987
rect -25977 -43127 -25639 -43027
rect -23728 -44174 -23542 -39590
rect -26388 -44360 -23542 -44174
rect -32434 -44640 -16322 -44504
rect -32450 -44839 -16322 -44703
rect -32458 -45072 -15025 -44936
rect -32482 -45327 -16322 -45191
rect -29580 -45439 -28157 -45411
rect -29580 -46337 -29421 -45439
rect -28307 -46337 -28157 -45439
rect -24214 -45613 -14730 -45477
rect -24214 -45618 -24059 -45613
rect -24214 -45776 -24078 -45618
rect -24214 -45912 -16322 -45776
rect -24214 -46146 -24078 -45912
rect 95829 -46113 98798 -31308
rect -24214 -46282 -16322 -46146
rect -29580 -46390 -28157 -46337
rect -29580 -46526 -16322 -46390
rect 83333 -49082 98798 -46113
rect -32776 -50847 -27886 -50668
rect -28065 -52016 -27886 -50847
rect 83333 -51532 86302 -49082
rect 91309 -52499 92592 -52202
rect 91309 -52743 91497 -52499
rect 89400 -53281 91497 -52743
rect 91309 -53325 91497 -53281
rect 92395 -53325 92592 -52499
rect 91309 -53546 92592 -53325
rect -27203 -54080 -22678 -53808
rect -29448 -54844 -29178 -54761
rect -29448 -58982 -29370 -54844
rect -29264 -54911 -29178 -54844
rect -27217 -54866 -22678 -54594
rect -29264 -55189 -28800 -54911
rect -29264 -56093 -29178 -55189
rect -27203 -55600 -22678 -55328
rect -29264 -56371 -28814 -56093
rect -29264 -57168 -29178 -56371
rect -19804 -57056 -19689 -56823
rect -29264 -57446 -28793 -57168
rect -26527 -57171 -19689 -57056
rect -29264 -58329 -29178 -57446
rect -29264 -58607 -28821 -58329
rect -29264 -58982 -29178 -58607
rect -29448 -59163 -29178 -58982
rect -28147 -62311 -28010 -59815
rect -27236 -60583 -26896 -60567
rect -27236 -60977 -27227 -60583
rect -26905 -60736 -26896 -60583
rect -26527 -60736 -26412 -57171
rect -26905 -60851 -26412 -60736
rect -26905 -60977 -26896 -60851
rect -27236 -60993 -26896 -60977
rect -23096 -62272 -22910 -57701
rect -23449 -62311 -22910 -62272
rect -28147 -62448 -22910 -62311
rect -23449 -62458 -22910 -62448
rect -33062 -62751 -16322 -62615
rect -33463 -62950 -16322 -62814
rect -32991 -63183 -16322 -63047
rect -32976 -63438 -16322 -63302
rect -31679 -63836 -30520 -63625
rect -23846 -63729 -23123 -63588
rect -31679 -63855 -30522 -63836
rect -31679 -64753 -31520 -63855
rect -30694 -64501 -30522 -63855
rect -23846 -63887 -23710 -63729
rect -23846 -64023 -22771 -63887
rect -23846 -64257 -23710 -64023
rect -23846 -64393 -23184 -64257
rect -30694 -64637 -22352 -64501
rect -30694 -64753 -30522 -64637
rect -31679 -64865 -30522 -64753
<< viali >>
rect -4688 42553 -3934 43955
rect -1796 42569 -1042 43971
rect -3582 39564 -2684 40390
rect -16054 8117 -15588 8439
rect -6465 7410 -5567 8380
rect 14616 8763 14722 8869
rect 7017 8531 7267 8709
rect 16266 8654 16300 8688
rect 16338 8654 16372 8688
rect 3512 7656 3906 8050
rect 7357 8072 7535 8250
rect 14612 7687 14718 7793
rect 16687 7627 16937 7877
rect 27007 7793 37625 8619
rect -12793 5693 -11679 6735
rect -3460 5769 -2562 6667
rect 15045 6804 15151 6910
rect 19319 6727 19569 6977
rect 23024 6740 23202 6990
rect 16262 6515 16296 6549
rect 16334 6515 16368 6549
rect 14508 6066 14614 6172
rect 13910 5746 14088 5924
rect 18862 5272 19112 5522
rect 2928 4208 3178 4458
rect 41740 4330 44510 4724
rect 15899 3776 16221 4098
rect -13067 3391 -9289 3497
rect 3593 3363 3771 3541
rect 26677 3553 38663 3803
rect -5790 2533 -5612 2711
rect -13321 2186 -9327 2292
rect 18185 3032 18291 3138
rect 41866 3165 41900 3199
rect 41938 3165 41972 3199
rect 42010 3165 42044 3199
rect 42082 3165 42116 3199
rect 42154 3165 42188 3199
rect 42226 3165 42260 3199
rect 42298 3165 42332 3199
rect 42370 3165 42404 3199
rect 42442 3165 42476 3199
rect 42514 3165 42548 3199
rect 42586 3165 42620 3199
rect 42658 3165 42692 3199
rect 42730 3165 42764 3199
rect 42802 3165 42836 3199
rect 42874 3165 42908 3199
rect 42946 3165 42980 3199
rect 43018 3165 43052 3199
rect 43090 3165 43124 3199
rect 43162 3165 43196 3199
rect 43234 3165 43268 3199
rect 43306 3165 43340 3199
rect 43378 3165 43412 3199
rect 43450 3165 43484 3199
rect 43522 3165 43556 3199
rect 43594 3165 43628 3199
rect 43666 3165 43700 3199
rect 43738 3165 43772 3199
rect 43810 3165 43844 3199
rect 43882 3165 43916 3199
rect 43954 3165 43988 3199
rect 44026 3165 44060 3199
rect 44098 3165 44132 3199
rect 19582 2821 19616 2855
rect 19830 2803 19864 2837
rect 19902 2803 19936 2837
rect 19974 2803 20008 2837
rect 20046 2803 20080 2837
rect 20118 2803 20152 2837
rect 20190 2803 20224 2837
rect 20262 2803 20296 2837
rect 19401 2530 19435 2564
rect 18667 2477 18701 2511
rect 19401 2458 19435 2492
rect 7089 1865 7267 2043
rect -5730 1386 -5624 1492
rect -4169 1483 -4135 1517
rect -13293 583 -6203 689
rect -3512 1458 -3478 1492
rect -3440 1458 -3406 1492
rect -3368 1458 -3334 1492
rect -3296 1458 -3262 1492
rect -3224 1458 -3190 1492
rect -3152 1458 -3118 1492
rect 3553 1345 3803 1595
rect 4029 1590 4063 1624
rect 4029 1518 4063 1552
rect 7381 1606 7415 1640
rect 4245 1431 4279 1465
rect -17981 356 -17659 534
rect -6478 325 -5652 431
rect 3591 911 3697 1017
rect 4649 1434 4683 1468
rect 4721 1434 4755 1468
rect 15576 1664 15682 1770
rect 7121 1400 7227 1506
rect 22385 2750 22491 2856
rect 26734 2714 26912 2820
rect 25092 2136 25270 2314
rect 25980 2135 26086 2313
rect 50542 2243 50720 2421
rect 58776 2416 58882 2522
rect 4417 1099 4523 1205
rect 19522 986 19700 1164
rect 5767 713 5801 747
rect 5839 713 5873 747
rect 5911 713 5945 747
rect 5983 713 6017 747
rect 6055 713 6089 747
rect 6127 713 6161 747
rect 4030 113 4136 219
rect -13046 -383 -7324 -205
rect -6020 -338 -5986 -304
rect -5948 -338 -5914 -304
rect -5876 -338 -5842 -304
rect -5804 -338 -5770 -304
rect -25480 -954 -25230 -704
rect -5939 -985 -5833 -807
rect -5036 -910 -5002 -876
rect -4964 -910 -4930 -876
rect -4892 -910 -4858 -876
rect -4820 -910 -4786 -876
rect -4748 -910 -4714 -876
rect -4676 -910 -4642 -876
rect -4604 -910 -4570 -876
rect -4140 -1056 -4106 -1022
rect -1548 -295 -1370 -117
rect 4424 -168 4530 -62
rect 5919 -88 6169 162
rect 15880 -124 16202 270
rect 46686 1741 46864 1919
rect 47959 1703 48137 1953
rect 22486 926 22808 1248
rect 20011 -552 20045 -518
rect 20083 -552 20117 -518
rect 20155 -552 20189 -518
rect 20227 -552 20261 -518
rect 20299 -552 20333 -518
rect 20371 -552 20405 -518
rect 20443 -552 20477 -518
rect 3355 -877 3533 -699
rect 47797 -706 47903 -600
rect 60645 -632 61039 -382
rect 4567 -1056 4601 -1022
rect 4639 -1056 4673 -1022
rect 4711 -1056 4745 -1022
rect 4783 -1056 4817 -1022
rect 4855 -1056 4889 -1022
rect 4927 -1056 4961 -1022
rect 7372 -1165 7406 -1131
rect 16129 -1178 16379 -928
rect 19870 -1226 20048 -1048
rect 4333 -2293 4439 -2187
rect -1533 -2525 -1355 -2419
rect 46934 -2431 47256 -2109
rect 3300 -2846 3550 -2596
rect 15515 -3145 15765 -2967
rect 16158 -3534 16408 -3356
rect 49025 -3652 49203 -3402
rect 62412 -3419 62446 -3385
rect 62484 -3419 62518 -3385
rect 62556 -3419 62590 -3385
rect 62628 -3419 62662 -3385
rect 62700 -3419 62734 -3385
rect 62772 -3419 62806 -3385
rect 62844 -3419 62878 -3385
rect 65205 -3420 65239 -3386
rect 65277 -3420 65311 -3386
rect 61914 -3476 61948 -3442
rect 61986 -3476 62020 -3442
rect 87949 -3463 88127 -3285
rect 62474 -4094 62724 -3844
rect 17422 -4739 17816 -4345
rect 18053 -5336 18375 -5014
rect 46926 -5169 47248 -4775
rect 61332 -4947 61438 -4841
rect 18565 -6058 18959 -5592
rect 19129 -6739 19451 -6417
rect 19786 -7516 20180 -7122
rect 90388 -7257 92654 -5063
rect -31392 -9819 -30710 -8993
rect 59146 -9712 59756 -9030
rect 60630 -10560 61312 -9806
rect -29366 -11602 -28468 -10704
rect -26776 -11773 -26094 -11091
rect -24141 -11672 -23459 -11062
rect -6514 -11806 -6048 -11268
rect 61636 -11730 62174 -11264
rect 62412 -13050 62950 -12584
rect -25638 -14746 -25028 -14352
rect -12791 -15157 -8005 -15051
rect 90552 -18574 91450 -17748
rect -25536 -23289 -25142 -22895
rect 90887 -35110 91785 -34284
rect -27563 -37084 -27529 -37050
rect -27563 -37156 -27529 -37122
rect -27563 -37228 -27529 -37194
rect -27563 -37300 -27529 -37266
rect -27563 -37372 -27529 -37338
rect -27563 -37444 -27529 -37410
rect -27563 -37516 -27529 -37482
rect -27563 -37588 -27529 -37554
rect -27563 -37660 -27529 -37626
rect -27563 -37732 -27529 -37698
rect -27563 -37804 -27529 -37770
rect -27563 -37876 -27529 -37842
rect -27563 -37948 -27529 -37914
rect -27563 -38020 -27529 -37986
rect -27563 -38092 -27529 -38058
rect -27563 -38164 -27529 -38130
rect -27563 -38236 -27529 -38202
rect -27563 -38308 -27529 -38274
rect -27563 -38380 -27529 -38346
rect -27563 -38452 -27529 -38418
rect -27563 -38524 -27529 -38490
rect -27563 -38596 -27529 -38562
rect -27563 -38668 -27529 -38634
rect -27563 -38740 -27529 -38706
rect -27563 -38812 -27529 -38778
rect -27563 -38884 -27529 -38850
rect -27563 -38956 -27529 -38922
rect -27563 -39028 -27529 -38994
rect -27563 -39100 -27529 -39066
rect -27563 -39172 -27529 -39138
rect -27563 -39244 -27529 -39210
rect -27563 -39316 -27529 -39282
rect -27563 -39388 -27529 -39354
rect -27563 -39460 -27529 -39426
rect -27563 -39532 -27529 -39498
rect -27563 -39604 -27529 -39570
rect -27563 -39676 -27529 -39642
rect -27563 -39748 -27529 -39714
rect -27563 -39820 -27529 -39786
rect -27563 -39892 -27529 -39858
rect -27563 -39964 -27529 -39930
rect -27563 -40036 -27529 -40002
rect -27563 -40108 -27529 -40074
rect -27563 -40180 -27529 -40146
rect -27563 -40252 -27529 -40218
rect -27563 -40324 -27529 -40290
rect -27563 -40396 -27529 -40362
rect -27563 -40468 -27529 -40434
rect -27563 -40540 -27529 -40506
rect -27563 -40612 -27529 -40578
rect -27563 -40684 -27529 -40650
rect -27563 -40756 -27529 -40722
rect -27563 -40828 -27529 -40794
rect -27563 -40900 -27529 -40866
rect -27563 -40972 -27529 -40938
rect -27563 -41044 -27529 -41010
rect -27563 -41116 -27529 -41082
rect -25880 -43027 -25702 -42849
rect -29421 -46337 -28307 -45439
rect 91497 -53325 92395 -52499
rect -29370 -58982 -29264 -54844
rect -27227 -60977 -26905 -60583
rect -31520 -64753 -30694 -63855
<< metal1 >>
rect -4820 44054 -3786 44102
rect -1993 44054 -862 44070
rect -4820 43971 -797 44054
rect -4820 43955 -1796 43971
rect -4820 42553 -4688 43955
rect -3934 42569 -1796 43955
rect -1042 42569 -797 43971
rect -3934 42553 -797 42569
rect -4820 42503 -797 42553
rect -4820 42470 -3786 42503
rect -1993 42470 -862 42503
rect -3742 40390 -2527 40571
rect -3742 39564 -3582 40390
rect -2684 40236 -2527 40390
rect -2684 39564 -2367 40236
rect -3742 39356 -2367 39564
rect -17836 9129 -15919 9265
rect -17836 565 -17700 9129
rect -16277 8494 -5438 8555
rect -16277 8439 -5433 8494
rect -16277 8117 -16054 8439
rect -15588 8380 -5433 8439
rect -15588 8117 -6465 8380
rect -16277 8032 -6465 8117
rect -6540 7410 -6465 8032
rect -5567 7410 -5433 8380
rect -6540 7273 -5433 7410
rect -12975 6735 -11404 6943
rect -12975 5693 -12793 6735
rect -11679 5693 -11404 6735
rect -12975 3566 -11404 5693
rect -3582 6667 -2367 39356
rect 13898 8915 14773 8919
rect 13898 8869 14775 8915
rect 13898 8763 14616 8869
rect 14722 8763 14775 8869
rect 6966 8709 7312 8756
rect 6966 8531 7017 8709
rect 7267 8531 7312 8709
rect 6966 8466 7312 8531
rect 13898 8737 14775 8763
rect 3375 8050 4103 8200
rect 3375 7656 3512 8050
rect 3906 7656 4103 8050
rect 3375 7565 4103 7656
rect -3582 5769 -3460 6667
rect -2562 5769 -2367 6667
rect -3582 5554 -2367 5769
rect 2866 4458 3250 4560
rect 2866 4208 2928 4458
rect 3178 4208 3250 4458
rect 2866 4116 3250 4208
rect -13122 3497 -8953 3566
rect -13122 3391 -13067 3497
rect -9289 3391 -8953 3497
rect -13122 3329 -8953 3391
rect -13011 2361 -12663 3329
rect -11909 2361 -11561 3329
rect -11015 2361 -10667 3329
rect -10239 2361 -9891 3329
rect -9633 2361 -9285 3329
rect -5845 2711 -5539 2764
rect -5845 2533 -5790 2711
rect -5612 2533 -5539 2711
rect -5845 2483 -5539 2533
rect -613 2710 538 2816
rect -13395 2292 -9226 2361
rect -13395 2186 -13321 2292
rect -9327 2186 -9226 2292
rect -13395 2124 -9226 2186
rect -5742 1521 -5581 2483
rect -613 1575 -456 2710
rect 3061 2090 3235 4116
rect 3500 3541 3875 7565
rect 3500 3363 3593 3541
rect 3771 3363 3875 3541
rect -5774 1492 -5574 1521
rect -5774 1386 -5730 1492
rect -5624 1415 -5574 1492
rect -4212 1517 -4099 1535
rect -4212 1483 -4169 1517
rect -4135 1498 -4099 1517
rect -3572 1498 -3060 1502
rect -4135 1492 -3060 1498
rect -4135 1483 -3512 1492
rect -4212 1461 -3512 1483
rect -3572 1458 -3512 1461
rect -3478 1458 -3440 1492
rect -3406 1458 -3368 1492
rect -3334 1458 -3296 1492
rect -3262 1458 -3224 1492
rect -3190 1458 -3152 1492
rect -3118 1458 -3060 1492
rect -3572 1449 -3060 1458
rect -1188 1423 -456 1575
rect 3500 1595 3875 3363
rect 7080 2079 7229 8466
rect 7289 8250 7635 8307
rect 7289 8072 7357 8250
rect 7535 8072 7635 8250
rect 7289 8017 7635 8072
rect 7054 2043 7303 2079
rect 7054 1865 7089 2043
rect 7267 1865 7303 2043
rect 7054 1845 7303 1865
rect 7341 1680 7460 8017
rect 13898 5964 14080 8737
rect 14547 8736 14775 8737
rect 14484 7856 14591 7858
rect 14484 7793 14796 7856
rect 14484 7687 14612 7793
rect 14718 7749 14796 7793
rect 14718 7687 14795 7749
rect 14484 7642 14795 7687
rect 14484 6213 14653 7642
rect 15079 6970 15125 8735
rect 16226 8688 16396 8743
rect 16226 8654 16266 8688
rect 16300 8654 16338 8688
rect 16372 8654 16396 8688
rect 16226 8605 16396 8654
rect 26753 8619 38073 8844
rect 14997 6910 15211 6970
rect 14997 6804 15045 6910
rect 15151 6804 15211 6910
rect 14997 6756 15211 6804
rect 16250 6623 16388 8605
rect 16519 7877 17132 8006
rect 16519 7627 16687 7877
rect 16937 7627 17132 7877
rect 16227 6549 16406 6623
rect 16227 6515 16262 6549
rect 16296 6515 16334 6549
rect 16368 6515 16406 6549
rect 16227 6444 16406 6515
rect 14443 6172 14691 6213
rect 14443 6066 14508 6172
rect 14614 6066 14691 6172
rect 14443 6016 14691 6066
rect 13866 5924 14130 5964
rect 13866 5746 13910 5924
rect 14088 5746 14130 5924
rect 13866 5703 14130 5746
rect 15814 4098 16331 4171
rect 15814 3776 15899 4098
rect 16221 3776 16331 4098
rect 15814 3722 16331 3776
rect 15522 1770 15742 1833
rect 7337 1670 7470 1680
rect 6982 1640 7470 1670
rect -5624 1386 -3699 1415
rect -5774 1371 -3699 1386
rect -5774 1352 -5574 1371
rect 3500 1345 3553 1595
rect 3803 1345 3875 1595
rect 3990 1624 4106 1638
rect 6982 1624 7381 1640
rect 3990 1590 4029 1624
rect 4063 1591 4106 1624
rect 7337 1606 7381 1624
rect 7415 1606 7470 1640
rect 4063 1590 4392 1591
rect 3990 1552 4392 1590
rect 7337 1562 7470 1606
rect 15522 1664 15576 1770
rect 15682 1664 15742 1770
rect 15522 1597 15742 1664
rect 3990 1518 4029 1552
rect 4063 1547 4392 1552
rect 4063 1518 4106 1547
rect 3990 1499 4106 1518
rect 4186 1468 4963 1519
rect 4186 1465 4649 1468
rect 4186 1431 4245 1465
rect 4279 1434 4649 1465
rect 4683 1434 4721 1468
rect 4755 1434 4963 1468
rect 4279 1431 4963 1434
rect 4186 1385 4963 1431
rect 7061 1506 7270 1554
rect 7061 1400 7121 1506
rect 7227 1400 7270 1506
rect 4580 1384 4827 1385
rect 7061 1355 7270 1400
rect 3500 1279 3875 1345
rect 4064 1310 4362 1354
rect -5243 1073 -3681 1219
rect 3161 1101 3899 1159
rect -13350 689 -6080 721
rect -13350 583 -13293 689
rect -6203 583 -6080 689
rect -18039 534 -17604 565
rect -13350 548 -6080 583
rect -18039 356 -17981 534
rect -17659 356 -17604 534
rect -18039 321 -17604 356
rect -12759 -135 -12272 548
rect -11199 -135 -10712 548
rect -10006 -135 -9519 548
rect -8823 -135 -8336 548
rect -7809 -135 -7322 548
rect -5243 473 -5078 1073
rect 3563 1017 3725 1039
rect 3563 911 3591 1017
rect 3697 973 3725 1017
rect 3697 929 3812 973
rect 3697 911 3725 929
rect 3563 885 3725 911
rect -6599 431 -5077 473
rect -6599 389 -6478 431
rect -6600 325 -6478 389
rect -5652 325 -5077 431
rect -6600 308 -5077 325
rect -6600 257 -5078 308
rect -6601 224 -5078 257
rect -13197 -205 -7163 -135
rect -13197 -383 -13046 -205
rect -7324 -383 -7163 -205
rect -13197 -453 -7163 -383
rect -25553 -704 -25165 -654
rect -25553 -954 -25480 -704
rect -25230 -954 -25165 -704
rect -25553 -1050 -25165 -954
rect -31679 -8993 -30522 -8679
rect -31679 -9819 -31392 -8993
rect -30710 -9819 -30522 -8993
rect -31679 -62597 -30522 -9819
rect -29580 -10704 -28157 -10506
rect -29580 -11602 -29366 -10704
rect -28468 -11602 -28157 -10704
rect -26907 -11091 -25983 -10980
rect -26907 -11153 -26776 -11091
rect -29580 -45439 -28157 -11602
rect -27809 -11705 -26776 -11153
rect -27809 -37050 -27257 -11705
rect -26907 -11773 -26776 -11705
rect -26094 -11773 -25983 -11091
rect -26907 -11904 -25983 -11773
rect -25501 -14108 -25219 -1050
rect -12865 -10939 -11924 -453
rect -24248 -11062 -11923 -10939
rect -24248 -11672 -24141 -11062
rect -23459 -11672 -11923 -11062
rect -24248 -11880 -11923 -11672
rect -25931 -14352 -24870 -14108
rect -25931 -14746 -25638 -14352
rect -25028 -14746 -24870 -14352
rect -25931 -14876 -24870 -14746
rect -25501 -22779 -25219 -14876
rect -12865 -14969 -11924 -11880
rect -10614 -14969 -9673 -453
rect -8935 -14969 -7994 -453
rect -6601 -11153 -6294 224
rect -2521 0 182 106
rect -6059 -304 -5507 -276
rect -6059 -338 -6020 -304
rect -5986 -338 -5948 -304
rect -5914 -338 -5876 -304
rect -5842 -338 -5804 -304
rect -5770 -338 -5507 -304
rect -6059 -378 -5507 -338
rect -5976 -807 -5800 -784
rect -5976 -985 -5939 -807
rect -5833 -957 -5800 -807
rect -5544 -873 -5507 -378
rect -2521 -665 -2415 0
rect -1581 -117 -1323 -85
rect -1581 -295 -1548 -117
rect -1370 -295 -1323 -117
rect -1581 -342 -1323 -295
rect -2521 -779 -2422 -665
rect -5056 -873 -4533 -861
rect -5544 -876 -4533 -873
rect -5544 -910 -5036 -876
rect -5002 -910 -4964 -876
rect -4930 -910 -4892 -876
rect -4858 -910 -4820 -876
rect -4786 -910 -4748 -876
rect -4714 -910 -4676 -876
rect -4642 -910 -4604 -876
rect -4570 -910 -4533 -876
rect -2650 -887 -2422 -779
rect -5056 -922 -4533 -910
rect -2598 -924 -2422 -887
rect -5833 -985 -5194 -957
rect -5976 -1001 -5194 -985
rect -5976 -1005 -5800 -1001
rect -4185 -1022 -4062 -989
rect -4185 -1056 -4140 -1022
rect -4106 -1056 -4062 -1022
rect -4185 -1079 -4062 -1056
rect -4182 -1094 -4138 -1079
rect -1517 -2369 -1361 -342
rect 3281 -699 3574 -645
rect 3281 -877 3355 -699
rect 3533 -877 3574 -699
rect 3281 -911 3574 -877
rect -1585 -2419 -1283 -2369
rect -1585 -2525 -1533 -2419
rect -1355 -2525 -1283 -2419
rect -1585 -2584 -1283 -2525
rect 3313 -2539 3558 -911
rect 3768 -1099 3812 929
rect 3841 -1011 3899 1101
rect 4064 265 4108 1310
rect 4388 1205 4549 1243
rect 4388 1099 4417 1205
rect 4523 1099 4549 1205
rect 4388 1066 4549 1099
rect 3985 219 4186 265
rect 3985 113 4030 219
rect 4136 113 4186 219
rect 3985 76 4186 113
rect 4408 -15 4507 1066
rect 5730 747 6208 775
rect 5730 713 5767 747
rect 5801 713 5839 747
rect 5873 713 5911 747
rect 5945 713 5983 747
rect 6017 713 6055 747
rect 6089 713 6127 747
rect 6161 713 6208 747
rect 5730 686 6208 713
rect 5943 223 6135 686
rect 5891 162 6236 223
rect 4383 -62 4585 -15
rect 4383 -168 4424 -62
rect 4530 -168 4585 -62
rect 5891 -88 5919 162
rect 6169 -88 6236 162
rect 5891 -122 6236 -88
rect 4383 -213 4585 -168
rect 3841 -1022 4999 -1011
rect 7131 -1020 7230 1355
rect 3841 -1056 4567 -1022
rect 4601 -1056 4639 -1022
rect 4673 -1056 4711 -1022
rect 4745 -1056 4783 -1022
rect 4817 -1056 4855 -1022
rect 4889 -1056 4927 -1022
rect 4961 -1056 4999 -1022
rect 3841 -1066 4999 -1056
rect 6997 -1066 7412 -1020
rect 3841 -1069 4601 -1066
rect 7334 -1093 7412 -1066
rect 3768 -1143 4387 -1099
rect 7334 -1131 7443 -1093
rect 7334 -1165 7372 -1131
rect 7406 -1165 7443 -1131
rect 7334 -1207 7443 -1165
rect 4353 -2171 4397 -1336
rect 4310 -2187 4465 -2171
rect 4310 -2293 4333 -2187
rect 4439 -2293 4465 -2187
rect 4310 -2309 4465 -2293
rect 3196 -2596 3624 -2539
rect 3196 -2846 3300 -2596
rect 3550 -2846 3624 -2596
rect 15547 -2842 15703 1597
rect 15814 270 16329 3722
rect 16519 909 17132 7627
rect 26753 7793 27007 8619
rect 37625 7793 38073 8619
rect 26753 7623 38073 7793
rect 19201 6977 19643 7085
rect 19201 6727 19319 6977
rect 19569 6727 19643 6977
rect 19201 6620 19643 6727
rect 22939 6990 23303 7116
rect 22939 6740 23024 6990
rect 23202 6740 23303 6990
rect 22939 6666 23303 6740
rect 18791 5522 19168 5573
rect 18791 5272 18862 5522
rect 19112 5272 19168 5522
rect 18791 5216 19168 5272
rect 18137 3181 18324 3184
rect 18137 3138 18330 3181
rect 18137 3032 18185 3138
rect 18291 3032 18330 3138
rect 18137 2985 18330 3032
rect 16519 296 17906 909
rect 15814 -124 15880 270
rect 16202 -124 16329 270
rect 15814 -255 16329 -124
rect 16101 -928 16445 -871
rect 16101 -1178 16129 -928
rect 16379 -1178 16445 -928
rect 16101 -1228 16445 -1178
rect 3196 -2900 3624 -2846
rect 15440 -2967 15853 -2842
rect 15440 -3145 15515 -2967
rect 15765 -3145 15853 -2967
rect 15440 -3211 15853 -3145
rect 16133 -3292 16375 -1228
rect 16088 -3356 16483 -3292
rect 16088 -3534 16158 -3356
rect 16408 -3534 16483 -3356
rect 16088 -3623 16483 -3534
rect 17293 -4345 17906 296
rect 17293 -4739 17422 -4345
rect 17816 -4739 17906 -4345
rect 17293 -4848 17906 -4739
rect 18137 -4849 18324 2985
rect 18621 2511 18758 2557
rect 18621 2477 18667 2511
rect 18701 2477 18758 2511
rect 17978 -5014 18468 -4849
rect 17978 -5336 18053 -5014
rect 18375 -5336 18468 -5014
rect 17978 -5437 18468 -5336
rect 18621 -5532 18758 2477
rect 18861 -594 19153 5216
rect 19341 2756 19470 6620
rect 19552 2862 19650 2892
rect 22316 2875 22554 2900
rect 19552 2858 19659 2862
rect 19552 2855 20314 2858
rect 19552 2821 19582 2855
rect 19616 2837 20314 2855
rect 19616 2821 19830 2837
rect 19552 2803 19830 2821
rect 19864 2803 19902 2837
rect 19936 2803 19974 2837
rect 20008 2803 20046 2837
rect 20080 2803 20118 2837
rect 20152 2803 20190 2837
rect 20224 2803 20262 2837
rect 20296 2803 20314 2837
rect 19552 2787 20314 2803
rect 22188 2856 22554 2875
rect 19341 2712 19648 2756
rect 22188 2750 22385 2856
rect 22491 2750 22554 2856
rect 22188 2745 22554 2750
rect 19341 2700 19470 2712
rect 22316 2711 22554 2745
rect 19341 2564 19481 2579
rect 19341 2530 19401 2564
rect 19435 2530 19481 2564
rect 19341 2519 19481 2530
rect 19341 2492 19671 2519
rect 19341 2458 19401 2492
rect 19435 2475 19671 2492
rect 19435 2458 19481 2475
rect 19341 2444 19481 2458
rect 22436 1248 22925 1317
rect 22436 1241 22486 1248
rect 19472 1164 22486 1241
rect 19472 986 19522 1164
rect 19700 986 22486 1164
rect 19472 943 22486 986
rect 19472 -496 19542 943
rect 22436 926 22486 943
rect 22808 926 22925 1248
rect 22436 895 22925 926
rect 22358 -353 22513 -345
rect 23046 -353 23217 6666
rect 26836 3886 28029 7623
rect 29111 3886 30304 7623
rect 31275 3886 32468 7623
rect 33884 3886 35077 7623
rect 36381 3886 37574 7623
rect 41672 4724 44640 4844
rect 41672 4330 41740 4724
rect 44510 4330 44640 4724
rect 41672 4185 44640 4330
rect 26583 3803 38866 3886
rect 26583 3553 26677 3803
rect 38663 3553 38866 3803
rect 26583 3483 38866 3553
rect 41865 3233 42195 4185
rect 42554 3233 42884 4185
rect 43243 3233 43573 4185
rect 43752 3233 44082 4185
rect 41827 3199 44196 3233
rect 41827 3165 41866 3199
rect 41900 3165 41938 3199
rect 41972 3165 42010 3199
rect 42044 3165 42082 3199
rect 42116 3165 42154 3199
rect 42188 3165 42226 3199
rect 42260 3165 42298 3199
rect 42332 3165 42370 3199
rect 42404 3165 42442 3199
rect 42476 3165 42514 3199
rect 42548 3165 42586 3199
rect 42620 3165 42658 3199
rect 42692 3165 42730 3199
rect 42764 3165 42802 3199
rect 42836 3165 42874 3199
rect 42908 3165 42946 3199
rect 42980 3165 43018 3199
rect 43052 3165 43090 3199
rect 43124 3165 43162 3199
rect 43196 3165 43234 3199
rect 43268 3165 43306 3199
rect 43340 3165 43378 3199
rect 43412 3165 43450 3199
rect 43484 3165 43522 3199
rect 43556 3165 43594 3199
rect 43628 3165 43666 3199
rect 43700 3165 43738 3199
rect 43772 3165 43810 3199
rect 43844 3165 43882 3199
rect 43916 3165 43954 3199
rect 43988 3165 44026 3199
rect 44060 3165 44098 3199
rect 44132 3165 44196 3199
rect 41827 3129 44196 3165
rect 26688 2820 26963 2876
rect 26688 2714 26734 2820
rect 26912 2714 26963 2820
rect 26688 2653 26963 2714
rect 25061 2314 25333 2372
rect 25061 2136 25092 2314
rect 25270 2295 25333 2314
rect 25947 2313 26150 2357
rect 25947 2295 25980 2313
rect 25270 2136 25980 2295
rect 25061 2135 25980 2136
rect 26086 2135 26150 2313
rect 25061 2124 26150 2135
rect 25061 2085 25333 2124
rect 25947 2092 26150 2124
rect 26762 646 26890 2653
rect 58706 2522 59616 2704
rect 50510 2421 50749 2467
rect 50510 2243 50542 2421
rect 50720 2243 50749 2421
rect 58706 2416 58776 2522
rect 58882 2416 59616 2522
rect 58706 2260 59616 2416
rect 50510 2215 50749 2243
rect 46637 1919 46961 1997
rect 46637 1741 46686 1919
rect 46864 1917 46961 1919
rect 47896 1953 48216 1992
rect 47896 1917 47959 1953
rect 46864 1741 47959 1917
rect 46637 1738 47959 1741
rect 46637 1686 46961 1738
rect 47896 1703 47959 1738
rect 48137 1884 48216 1953
rect 50542 1917 50721 2215
rect 48137 1705 49256 1884
rect 48137 1703 48216 1705
rect 47896 1636 48216 1703
rect 26762 518 27180 646
rect 27052 -166 27180 518
rect 19472 -518 20517 -496
rect 19472 -552 20011 -518
rect 20045 -552 20083 -518
rect 20117 -552 20155 -518
rect 20189 -552 20227 -518
rect 20261 -552 20299 -518
rect 20333 -552 20371 -518
rect 20405 -552 20443 -518
rect 20477 -552 20517 -518
rect 22342 -524 23217 -353
rect 22358 -525 22513 -524
rect 19472 -566 20517 -552
rect 22433 -561 22513 -525
rect 18861 -638 19820 -594
rect 46227 -632 46301 1314
rect 47758 -600 47953 -572
rect 47758 -632 47797 -600
rect 46227 -706 47797 -632
rect 47903 -706 47953 -600
rect 47758 -752 47953 -706
rect 19212 -831 19359 -829
rect 19212 -875 20074 -831
rect 18424 -5592 19081 -5532
rect 18424 -6058 18565 -5592
rect 18959 -6058 19081 -5592
rect 18424 -6171 19081 -6058
rect 19212 -6293 19542 -875
rect 19836 -1048 20093 -990
rect 19836 -1226 19870 -1048
rect 20048 -1226 20093 -1048
rect 19836 -1279 20093 -1226
rect 18949 -6417 19611 -6293
rect 18949 -6739 19129 -6417
rect 19451 -6739 19611 -6417
rect 18949 -6850 19611 -6739
rect 19868 -7025 20066 -1279
rect 46850 -2109 47412 -1960
rect 46850 -2431 46934 -2109
rect 47256 -2431 47412 -2109
rect 46850 -4670 47412 -2431
rect 49077 -3371 49256 1705
rect 48966 -3402 49277 -3371
rect 48966 -3652 49025 -3402
rect 49203 -3652 49277 -3402
rect 48966 -3697 49277 -3652
rect 46778 -4775 47412 -4670
rect 46778 -5169 46926 -4775
rect 47248 -5169 47412 -4775
rect 46778 -5304 47412 -5169
rect 19665 -7122 20295 -7025
rect 19665 -7516 19786 -7122
rect 20180 -7516 20295 -7122
rect 19665 -7634 20295 -7516
rect 59172 -8831 59616 2260
rect 60549 -382 61159 -228
rect 60549 -632 60645 -382
rect 61039 -632 61159 -382
rect 58913 -9030 59860 -8831
rect 58913 -9712 59146 -9030
rect 59756 -9712 59860 -9030
rect 60549 -9617 61159 -632
rect 61353 -3293 62176 -3228
rect 61353 -4779 61418 -3293
rect 62111 -3360 62176 -3293
rect 87785 -3285 88210 -3189
rect 62111 -3385 62910 -3360
rect 65187 -3381 65330 -3337
rect 61873 -3442 62067 -3407
rect 62111 -3419 62412 -3385
rect 62446 -3419 62484 -3385
rect 62518 -3419 62556 -3385
rect 62590 -3419 62628 -3385
rect 62662 -3419 62700 -3385
rect 62734 -3419 62772 -3385
rect 62806 -3419 62844 -3385
rect 62878 -3419 62910 -3385
rect 62111 -3425 62910 -3419
rect 62387 -3431 62910 -3425
rect 64860 -3386 65330 -3381
rect 64860 -3420 65205 -3386
rect 65239 -3420 65277 -3386
rect 65311 -3420 65330 -3386
rect 64860 -3427 65330 -3420
rect 61873 -3476 61914 -3442
rect 61948 -3476 61986 -3442
rect 62020 -3460 62067 -3442
rect 62020 -3476 62250 -3460
rect 65187 -3468 65330 -3427
rect 87785 -3463 87949 -3285
rect 88127 -3463 88210 -3285
rect 61873 -3504 62250 -3476
rect 61873 -3516 62067 -3504
rect 87785 -3581 88210 -3463
rect 61655 -3741 62267 -3697
rect 61261 -4841 61482 -4779
rect 61261 -4947 61332 -4841
rect 61438 -4947 61482 -4841
rect 61261 -5041 61482 -4947
rect 58913 -9909 59860 -9712
rect 60423 -9806 61454 -9617
rect 60423 -10560 60630 -9806
rect 61312 -10560 61454 -9806
rect 60423 -10731 61454 -10560
rect 61655 -11116 62108 -3741
rect 62432 -3844 62779 -3786
rect 62432 -4094 62474 -3844
rect 62724 -4094 62779 -3844
rect 62432 -4139 62779 -4094
rect -6611 -11268 -5937 -11153
rect -6611 -11806 -6514 -11268
rect -6048 -11806 -5937 -11268
rect -6611 -11894 -5937 -11806
rect 61366 -11264 62272 -11116
rect 61366 -11730 61636 -11264
rect 62174 -11730 62272 -11264
rect 61366 -11971 62272 -11730
rect 62465 -12441 62732 -4139
rect 62246 -12584 63072 -12441
rect 62246 -13050 62412 -12584
rect 62950 -13050 63072 -12584
rect 62246 -13180 63072 -13050
rect -12874 -15051 -7870 -14969
rect -12874 -15157 -12791 -15051
rect -8005 -15157 -7870 -15051
rect -12874 -15238 -7870 -15157
rect -12865 -15240 -11924 -15238
rect -25664 -22895 -25039 -22779
rect -25664 -23289 -25536 -22895
rect -25142 -23289 -25039 -22895
rect -25664 -23404 -25039 -23289
rect 87916 -26943 88161 -3581
rect 89990 -5063 92959 -4698
rect 89990 -7257 90388 -5063
rect 92654 -7257 92959 -5063
rect 89990 -7667 92959 -7257
rect 84040 -27188 88161 -26943
rect 90119 -17748 92731 -7667
rect 90119 -18574 90552 -17748
rect 91450 -18574 92731 -17748
rect 84612 -27482 84857 -27188
rect 80867 -27727 84857 -27482
rect -27809 -37084 -27563 -37050
rect -27529 -37084 -27257 -37050
rect -27809 -37122 -27257 -37084
rect -27809 -37156 -27563 -37122
rect -27529 -37156 -27257 -37122
rect -27809 -37194 -27257 -37156
rect -27809 -37228 -27563 -37194
rect -27529 -37228 -27257 -37194
rect -27809 -37266 -27257 -37228
rect -27809 -37300 -27563 -37266
rect -27529 -37300 -27257 -37266
rect -27809 -37338 -27257 -37300
rect -27809 -37372 -27563 -37338
rect -27529 -37372 -27257 -37338
rect -27809 -37410 -27257 -37372
rect -27809 -37444 -27563 -37410
rect -27529 -37444 -27257 -37410
rect -27809 -37482 -27257 -37444
rect -27809 -37516 -27563 -37482
rect -27529 -37516 -27257 -37482
rect -27809 -37554 -27257 -37516
rect -27809 -37588 -27563 -37554
rect -27529 -37588 -27257 -37554
rect -27809 -37626 -27257 -37588
rect -27809 -37660 -27563 -37626
rect -27529 -37660 -27257 -37626
rect -27809 -37698 -27257 -37660
rect -27809 -37732 -27563 -37698
rect -27529 -37732 -27257 -37698
rect -27809 -37770 -27257 -37732
rect -27809 -37804 -27563 -37770
rect -27529 -37804 -27257 -37770
rect -27809 -37842 -27257 -37804
rect -27809 -37876 -27563 -37842
rect -27529 -37876 -27257 -37842
rect -27809 -37914 -27257 -37876
rect -27809 -37948 -27563 -37914
rect -27529 -37948 -27257 -37914
rect -27809 -37986 -27257 -37948
rect -27809 -38020 -27563 -37986
rect -27529 -38020 -27257 -37986
rect -27809 -38058 -27257 -38020
rect -27809 -38092 -27563 -38058
rect -27529 -38092 -27257 -38058
rect -27809 -38130 -27257 -38092
rect -27809 -38164 -27563 -38130
rect -27529 -38164 -27257 -38130
rect -27809 -38202 -27257 -38164
rect -27809 -38236 -27563 -38202
rect -27529 -38236 -27257 -38202
rect -27809 -38274 -27257 -38236
rect -27809 -38308 -27563 -38274
rect -27529 -38308 -27257 -38274
rect -27809 -38346 -27257 -38308
rect -27809 -38380 -27563 -38346
rect -27529 -38380 -27257 -38346
rect -27809 -38418 -27257 -38380
rect -27809 -38452 -27563 -38418
rect -27529 -38452 -27257 -38418
rect -27809 -38490 -27257 -38452
rect -27809 -38524 -27563 -38490
rect -27529 -38524 -27257 -38490
rect -27809 -38562 -27257 -38524
rect -27809 -38596 -27563 -38562
rect -27529 -38596 -27257 -38562
rect -27809 -38634 -27257 -38596
rect -27809 -38668 -27563 -38634
rect -27529 -38668 -27257 -38634
rect -27809 -38706 -27257 -38668
rect -27809 -38740 -27563 -38706
rect -27529 -38740 -27257 -38706
rect -27809 -38778 -27257 -38740
rect -27809 -38812 -27563 -38778
rect -27529 -38812 -27257 -38778
rect -27809 -38850 -27257 -38812
rect -27809 -38884 -27563 -38850
rect -27529 -38884 -27257 -38850
rect -27809 -38922 -27257 -38884
rect -27809 -38956 -27563 -38922
rect -27529 -38956 -27257 -38922
rect -27809 -38994 -27257 -38956
rect -27809 -39028 -27563 -38994
rect -27529 -39028 -27257 -38994
rect -27809 -39066 -27257 -39028
rect -27809 -39100 -27563 -39066
rect -27529 -39100 -27257 -39066
rect -27809 -39138 -27257 -39100
rect -27809 -39172 -27563 -39138
rect -27529 -39172 -27257 -39138
rect -27809 -39210 -27257 -39172
rect -27809 -39244 -27563 -39210
rect -27529 -39244 -27257 -39210
rect -27809 -39282 -27257 -39244
rect -27809 -39316 -27563 -39282
rect -27529 -39316 -27257 -39282
rect -27809 -39354 -27257 -39316
rect -27809 -39388 -27563 -39354
rect -27529 -39388 -27257 -39354
rect -27809 -39426 -27257 -39388
rect -27809 -39460 -27563 -39426
rect -27529 -39460 -27257 -39426
rect -27809 -39498 -27257 -39460
rect -27809 -39532 -27563 -39498
rect -27529 -39532 -27257 -39498
rect -27809 -39570 -27257 -39532
rect -27809 -39604 -27563 -39570
rect -27529 -39604 -27257 -39570
rect -27809 -39642 -27257 -39604
rect -27809 -39676 -27563 -39642
rect -27529 -39676 -27257 -39642
rect -27809 -39714 -27257 -39676
rect -27809 -39748 -27563 -39714
rect -27529 -39748 -27257 -39714
rect -27809 -39786 -27257 -39748
rect -27809 -39820 -27563 -39786
rect -27529 -39820 -27257 -39786
rect -27809 -39858 -27257 -39820
rect -27809 -39892 -27563 -39858
rect -27529 -39892 -27257 -39858
rect -27809 -39930 -27257 -39892
rect -27809 -39964 -27563 -39930
rect -27529 -39964 -27257 -39930
rect -27809 -40002 -27257 -39964
rect -27809 -40036 -27563 -40002
rect -27529 -40036 -27257 -40002
rect -27809 -40074 -27257 -40036
rect -27809 -40108 -27563 -40074
rect -27529 -40108 -27257 -40074
rect -27809 -40146 -27257 -40108
rect -27809 -40180 -27563 -40146
rect -27529 -40180 -27257 -40146
rect -27809 -40218 -27257 -40180
rect -27809 -40252 -27563 -40218
rect -27529 -40252 -27257 -40218
rect -27809 -40290 -27257 -40252
rect -27809 -40324 -27563 -40290
rect -27529 -40324 -27257 -40290
rect -27809 -40362 -27257 -40324
rect -27809 -40396 -27563 -40362
rect -27529 -40396 -27257 -40362
rect -27809 -40434 -27257 -40396
rect -27809 -40468 -27563 -40434
rect -27529 -40468 -27257 -40434
rect -27809 -40506 -27257 -40468
rect -27809 -40540 -27563 -40506
rect -27529 -40540 -27257 -40506
rect -27809 -40578 -27257 -40540
rect -27809 -40612 -27563 -40578
rect -27529 -40612 -27257 -40578
rect -27809 -40650 -27257 -40612
rect -27809 -40684 -27563 -40650
rect -27529 -40684 -27257 -40650
rect -27809 -40722 -27257 -40684
rect -27809 -40756 -27563 -40722
rect -27529 -40756 -27257 -40722
rect -27809 -40794 -27257 -40756
rect -27809 -40828 -27563 -40794
rect -27529 -40828 -27257 -40794
rect -27809 -40866 -27257 -40828
rect -27809 -40900 -27563 -40866
rect -27529 -40900 -27257 -40866
rect -27809 -40938 -27257 -40900
rect -27809 -40972 -27563 -40938
rect -27529 -40972 -27257 -40938
rect -27809 -41010 -27257 -40972
rect -27809 -41044 -27563 -41010
rect -27529 -41044 -27257 -41010
rect -27809 -41082 -27257 -41044
rect -27809 -41116 -27563 -41082
rect -27529 -41116 -27257 -41082
rect -27809 -42856 -27257 -41116
rect 90119 -34284 92731 -18574
rect 90119 -35110 90887 -34284
rect 91785 -35110 92731 -34284
rect -25977 -42849 -25639 -42789
rect -25977 -42856 -25880 -42849
rect -27809 -43027 -25880 -42856
rect -25702 -43027 -25639 -42849
rect -22415 -42924 -22111 -42864
rect -27809 -43047 -25639 -43027
rect -27809 -43351 -27257 -43047
rect -25977 -43127 -25639 -43047
rect -29580 -46337 -29421 -45439
rect -28307 -46337 -28157 -45439
rect -29580 -46472 -28157 -46337
rect 90119 -52499 92731 -35110
rect -29536 -54844 -29081 -52616
rect 90119 -53325 91497 -52499
rect 92395 -53325 92731 -52499
rect 90119 -54278 92731 -53325
rect -29536 -58982 -29370 -54844
rect -29264 -58982 -29081 -54844
rect -29536 -60594 -29081 -58982
rect -27322 -60583 -26810 -60453
rect -27322 -60594 -27227 -60583
rect -29536 -60977 -27227 -60594
rect -26905 -60977 -26810 -60583
rect -29536 -61049 -26810 -60977
rect -21712 -61035 -21354 -60975
rect -27322 -61078 -26810 -61049
rect -31679 -63836 -30520 -62597
rect -31679 -63855 -30522 -63836
rect -31679 -64753 -31520 -63855
rect -30694 -64753 -30522 -63855
rect -31679 -64865 -30522 -64753
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_0
timestamp 1726359333
transform 1 0 5174 0 1 -1085
box -887 -901 1886 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_1
timestamp 1726359333
transform 1 0 -2940 0 1 1429
box -887 -901 1886 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_2
timestamp 1726359333
transform 1 0 -4408 0 1 -943
box -887 -901 1886 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_3
timestamp 1726359333
transform 1 0 20610 0 1 -580
box -887 -901 1886 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_4
timestamp 1726359333
transform 1 0 5159 0 1 1605
box -887 -901 1886 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_5
timestamp 1726359333
transform 1 0 20438 0 1 2770
box -887 -901 1886 842
use ANALOG_MUX_MAG  ANALOG_MUX_MAG_6
timestamp 1726359333
transform 1 0 63037 0 1 -3446
box -887 -901 1886 842
use CP  CP_0
timestamp 1726361494
transform 0 -1 14952 1 0 9056
box -1443 -80648 80252 15146
use divider_top  divider_top_0
timestamp 1726359333
transform 1 0 9841 0 1 -30857
box -34598 -144 78159 15696
use divider_top  divider_top_1
timestamp 1726359333
transform 1 0 10539 0 1 -47448
box -34598 -144 78159 15696
use divider_top  divider_top_2
timestamp 1726359333
transform 0 1 -17326 1 0 43154
box -34598 -144 78159 15696
use divider_top  divider_top_3
timestamp 1726359333
transform 1 0 11242 0 1 -65559
box -34598 -144 78159 15696
use mirror_mag  mirror_mag_0
timestamp 1726359333
transform -1 0 14294 0 1 4889
box 1529 -557 6212 3030
use PFD  PFD_0
timestamp 1726359333
transform 1 0 540 0 1 474
box -539 -474 2730 2342
use Tapered_Buffer_mag  Tapered_Buffer_mag_0
timestamp 1726359333
transform -1 0 -5857 0 1 1513
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_1
timestamp 1726359333
transform 1 0 7529 0 1 -961
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_2
timestamp 1726359333
transform -1 0 -7497 0 -1 -16074
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_3
timestamp 1726359333
transform 1 0 50645 0 1 -3386
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_4
timestamp 1726359333
transform 1 0 50848 0 1 2572
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_5
timestamp 1726359333
transform 1 0 50645 0 1 -339
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_6
timestamp 1726359333
transform 1 0 7570 0 1 1795
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_7
timestamp 1726359333
transform 0 1 -27894 1 0 -59716
box -156 -982 7721 769
use Tapered_Buffer_mag  Tapered_Buffer_mag_8
timestamp 1726359333
transform 0 1 -26074 1 0 -41571
box -156 -982 7721 769
use VCO  VCO_0
timestamp 1726359333
transform 1 0 33690 0 1 -975
box -8117 -475 13984 4754
<< labels >>
flabel locali s -21980 -628 -21980 -628 0 FreeSans 2000 0 0 0 S6
flabel locali s -26239 -2019 -26239 -2019 0 FreeSans 2000 0 0 0 UP_INPUT
flabel locali s -26267 -2271 -26267 -2271 0 FreeSans 2000 0 0 0 DN_INPUT
flabel locali s -26048 -2492 -26048 -2492 0 FreeSans 2000 0 0 0 S2
flabel locali s -26089 -2778 -26089 -2778 0 FreeSans 2000 0 0 0 S3
flabel locali s -25937 -3111 -25937 -3111 0 FreeSans 2000 0 0 0 UP_OUT
flabel locali s -26013 -3482 -26013 -3482 0 FreeSans 2000 0 0 0 DN_OUT
flabel locali s -26050 -4594 -26050 -4594 0 FreeSans 2000 0 0 0 ITAIL
flabel locali s -26022 -5307 -26022 -5307 0 FreeSans 2000 0 0 0 S4
flabel locali s -26146 -6015 -26146 -6015 0 FreeSans 2000 0 0 0 VCTRL_IN
flabel locali s -26433 -6567 -26433 -6567 0 FreeSans 2000 0 0 0 LF_OFFCHIP
flabel locali s -26457 -7358 -26457 -7358 0 FreeSans 2000 0 0 0 S5
flabel locali s -32043 -33050 -32043 -33050 0 FreeSans 2000 0 0 0 OUT_CORE
flabel locali s -32436 -50788 -32436 -50788 0 FreeSans 2000 0 0 0 OUT_USB
flabel locali s -32358 -44578 -32358 -44578 0 FreeSans 2000 0 0 0 D12
flabel locali s -32366 -44780 -32366 -44780 0 FreeSans 2000 0 0 0 D13
flabel locali s -32390 -45015 -32390 -45015 0 FreeSans 2000 0 0 0 D14
flabel locali s -32390 -45265 -32390 -45265 0 FreeSans 2000 0 0 0 D15
flabel locali s -22154 405 -22154 405 0 FreeSans 2000 0 0 0 F_IN
flabel locali s -32479 -27992 -32479 -27992 0 FreeSans 2000 0 0 0 D0
flabel locali s -32448 -28196 -32448 -28196 0 FreeSans 2000 0 0 0 D1
flabel locali s -32417 -28414 -32417 -28414 0 FreeSans 2000 0 0 0 D2
flabel locali s -32504 -28656 -32504 -28656 0 FreeSans 2000 0 0 0 D3
flabel locali s -32907 -28960 -32907 -28960 0 FreeSans 2000 0 0 0 D4
flabel locali s -32684 -29264 -32684 -29264 0 FreeSans 2000 0 0 0 D5
flabel locali s -32808 -29624 -32808 -29624 0 FreeSans 2000 0 0 0 D6
flabel locali s -20443 4401 -20443 4401 0 FreeSans 2000 0 0 0 D7
flabel locali s -19883 5428 -19883 5428 0 FreeSans 2000 0 0 0 D8
flabel locali s -19736 7109 -19736 7109 0 FreeSans 2000 0 0 0 D9
flabel locali s -18882 7776 -18882 7776 0 FreeSans 2000 0 0 0 D10
flabel locali s -32966 -62696 -32966 -62696 0 FreeSans 2000 0 0 0 D16
flabel locali s -33364 -62901 -33364 -62901 0 FreeSans 2000 0 0 0 D17
flabel locali s -32912 -63121 -32912 -63121 0 FreeSans 2000 0 0 0 D18
flabel locali s -32843 -63367 -32843 -63367 0 FreeSans 2000 0 0 0 D19
flabel locali s -33957 -9382 -33957 -9382 0 FreeSans 2000 0 0 0 OUTB
flabel locali s -34119 -12958 -34119 -12958 0 FreeSans 2000 0 0 0 OUT
flabel locali s -22650 1410 -22650 1410 0 FreeSans 2000 0 0 0 PRE_SCALAR
flabel locali s -22938 181 -22938 181 0 FreeSans 2000 0 0 0 S1
flabel locali s -34376 -14319 -34376 -14319 0 FreeSans 2000 0 0 0 S7
flabel locali s -34232 -15974 -34232 -15974 0 FreeSans 2000 0 0 0 DIV_OUT
flabel locali s 97170 -15073 97170 -15073 0 FreeSans 20000 0 0 0 VDD
flabel locali s 79409 -6079 79409 -6079 0 FreeSans 20000 0 0 0 VSS
<< end >>
