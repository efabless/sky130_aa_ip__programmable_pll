magic
tech sky130A
magscale 1 2
timestamp 1726359333
<< metal3 >>
rect -9022 7952 -6650 8000
rect -9022 7888 -6734 7952
rect -6670 7888 -6650 7952
rect -9022 7872 -6650 7888
rect -9022 7808 -6734 7872
rect -6670 7808 -6650 7872
rect -9022 7792 -6650 7808
rect -9022 7728 -6734 7792
rect -6670 7728 -6650 7792
rect -9022 7712 -6650 7728
rect -9022 7648 -6734 7712
rect -6670 7648 -6650 7712
rect -9022 7632 -6650 7648
rect -9022 7568 -6734 7632
rect -6670 7568 -6650 7632
rect -9022 7552 -6650 7568
rect -9022 7488 -6734 7552
rect -6670 7488 -6650 7552
rect -9022 7472 -6650 7488
rect -9022 7408 -6734 7472
rect -6670 7408 -6650 7472
rect -9022 7392 -6650 7408
rect -9022 7328 -6734 7392
rect -6670 7328 -6650 7392
rect -9022 7312 -6650 7328
rect -9022 7248 -6734 7312
rect -6670 7248 -6650 7312
rect -9022 7232 -6650 7248
rect -9022 7168 -6734 7232
rect -6670 7168 -6650 7232
rect -9022 7152 -6650 7168
rect -9022 7088 -6734 7152
rect -6670 7088 -6650 7152
rect -9022 7072 -6650 7088
rect -9022 7008 -6734 7072
rect -6670 7008 -6650 7072
rect -9022 6992 -6650 7008
rect -9022 6928 -6734 6992
rect -6670 6928 -6650 6992
rect -9022 6912 -6650 6928
rect -9022 6848 -6734 6912
rect -6670 6848 -6650 6912
rect -9022 6832 -6650 6848
rect -9022 6768 -6734 6832
rect -6670 6768 -6650 6832
rect -9022 6752 -6650 6768
rect -9022 6688 -6734 6752
rect -6670 6688 -6650 6752
rect -9022 6672 -6650 6688
rect -9022 6608 -6734 6672
rect -6670 6608 -6650 6672
rect -9022 6592 -6650 6608
rect -9022 6528 -6734 6592
rect -6670 6528 -6650 6592
rect -9022 6512 -6650 6528
rect -9022 6448 -6734 6512
rect -6670 6448 -6650 6512
rect -9022 6432 -6650 6448
rect -9022 6368 -6734 6432
rect -6670 6368 -6650 6432
rect -9022 6352 -6650 6368
rect -9022 6288 -6734 6352
rect -6670 6288 -6650 6352
rect -9022 6272 -6650 6288
rect -9022 6208 -6734 6272
rect -6670 6208 -6650 6272
rect -9022 6192 -6650 6208
rect -9022 6128 -6734 6192
rect -6670 6128 -6650 6192
rect -9022 6112 -6650 6128
rect -9022 6048 -6734 6112
rect -6670 6048 -6650 6112
rect -9022 6032 -6650 6048
rect -9022 5968 -6734 6032
rect -6670 5968 -6650 6032
rect -9022 5920 -6650 5968
rect -6410 7952 -4038 8000
rect -6410 7888 -4122 7952
rect -4058 7888 -4038 7952
rect -6410 7872 -4038 7888
rect -6410 7808 -4122 7872
rect -4058 7808 -4038 7872
rect -6410 7792 -4038 7808
rect -6410 7728 -4122 7792
rect -4058 7728 -4038 7792
rect -6410 7712 -4038 7728
rect -6410 7648 -4122 7712
rect -4058 7648 -4038 7712
rect -6410 7632 -4038 7648
rect -6410 7568 -4122 7632
rect -4058 7568 -4038 7632
rect -6410 7552 -4038 7568
rect -6410 7488 -4122 7552
rect -4058 7488 -4038 7552
rect -6410 7472 -4038 7488
rect -6410 7408 -4122 7472
rect -4058 7408 -4038 7472
rect -6410 7392 -4038 7408
rect -6410 7328 -4122 7392
rect -4058 7328 -4038 7392
rect -6410 7312 -4038 7328
rect -6410 7248 -4122 7312
rect -4058 7248 -4038 7312
rect -6410 7232 -4038 7248
rect -6410 7168 -4122 7232
rect -4058 7168 -4038 7232
rect -6410 7152 -4038 7168
rect -6410 7088 -4122 7152
rect -4058 7088 -4038 7152
rect -6410 7072 -4038 7088
rect -6410 7008 -4122 7072
rect -4058 7008 -4038 7072
rect -6410 6992 -4038 7008
rect -6410 6928 -4122 6992
rect -4058 6928 -4038 6992
rect -6410 6912 -4038 6928
rect -6410 6848 -4122 6912
rect -4058 6848 -4038 6912
rect -6410 6832 -4038 6848
rect -6410 6768 -4122 6832
rect -4058 6768 -4038 6832
rect -6410 6752 -4038 6768
rect -6410 6688 -4122 6752
rect -4058 6688 -4038 6752
rect -6410 6672 -4038 6688
rect -6410 6608 -4122 6672
rect -4058 6608 -4038 6672
rect -6410 6592 -4038 6608
rect -6410 6528 -4122 6592
rect -4058 6528 -4038 6592
rect -6410 6512 -4038 6528
rect -6410 6448 -4122 6512
rect -4058 6448 -4038 6512
rect -6410 6432 -4038 6448
rect -6410 6368 -4122 6432
rect -4058 6368 -4038 6432
rect -6410 6352 -4038 6368
rect -6410 6288 -4122 6352
rect -4058 6288 -4038 6352
rect -6410 6272 -4038 6288
rect -6410 6208 -4122 6272
rect -4058 6208 -4038 6272
rect -6410 6192 -4038 6208
rect -6410 6128 -4122 6192
rect -4058 6128 -4038 6192
rect -6410 6112 -4038 6128
rect -6410 6048 -4122 6112
rect -4058 6048 -4038 6112
rect -6410 6032 -4038 6048
rect -6410 5968 -4122 6032
rect -4058 5968 -4038 6032
rect -6410 5920 -4038 5968
rect -3798 7952 -1426 8000
rect -3798 7888 -1510 7952
rect -1446 7888 -1426 7952
rect -3798 7872 -1426 7888
rect -3798 7808 -1510 7872
rect -1446 7808 -1426 7872
rect -3798 7792 -1426 7808
rect -3798 7728 -1510 7792
rect -1446 7728 -1426 7792
rect -3798 7712 -1426 7728
rect -3798 7648 -1510 7712
rect -1446 7648 -1426 7712
rect -3798 7632 -1426 7648
rect -3798 7568 -1510 7632
rect -1446 7568 -1426 7632
rect -3798 7552 -1426 7568
rect -3798 7488 -1510 7552
rect -1446 7488 -1426 7552
rect -3798 7472 -1426 7488
rect -3798 7408 -1510 7472
rect -1446 7408 -1426 7472
rect -3798 7392 -1426 7408
rect -3798 7328 -1510 7392
rect -1446 7328 -1426 7392
rect -3798 7312 -1426 7328
rect -3798 7248 -1510 7312
rect -1446 7248 -1426 7312
rect -3798 7232 -1426 7248
rect -3798 7168 -1510 7232
rect -1446 7168 -1426 7232
rect -3798 7152 -1426 7168
rect -3798 7088 -1510 7152
rect -1446 7088 -1426 7152
rect -3798 7072 -1426 7088
rect -3798 7008 -1510 7072
rect -1446 7008 -1426 7072
rect -3798 6992 -1426 7008
rect -3798 6928 -1510 6992
rect -1446 6928 -1426 6992
rect -3798 6912 -1426 6928
rect -3798 6848 -1510 6912
rect -1446 6848 -1426 6912
rect -3798 6832 -1426 6848
rect -3798 6768 -1510 6832
rect -1446 6768 -1426 6832
rect -3798 6752 -1426 6768
rect -3798 6688 -1510 6752
rect -1446 6688 -1426 6752
rect -3798 6672 -1426 6688
rect -3798 6608 -1510 6672
rect -1446 6608 -1426 6672
rect -3798 6592 -1426 6608
rect -3798 6528 -1510 6592
rect -1446 6528 -1426 6592
rect -3798 6512 -1426 6528
rect -3798 6448 -1510 6512
rect -1446 6448 -1426 6512
rect -3798 6432 -1426 6448
rect -3798 6368 -1510 6432
rect -1446 6368 -1426 6432
rect -3798 6352 -1426 6368
rect -3798 6288 -1510 6352
rect -1446 6288 -1426 6352
rect -3798 6272 -1426 6288
rect -3798 6208 -1510 6272
rect -1446 6208 -1426 6272
rect -3798 6192 -1426 6208
rect -3798 6128 -1510 6192
rect -1446 6128 -1426 6192
rect -3798 6112 -1426 6128
rect -3798 6048 -1510 6112
rect -1446 6048 -1426 6112
rect -3798 6032 -1426 6048
rect -3798 5968 -1510 6032
rect -1446 5968 -1426 6032
rect -3798 5920 -1426 5968
rect -1186 7952 1186 8000
rect -1186 7888 1102 7952
rect 1166 7888 1186 7952
rect -1186 7872 1186 7888
rect -1186 7808 1102 7872
rect 1166 7808 1186 7872
rect -1186 7792 1186 7808
rect -1186 7728 1102 7792
rect 1166 7728 1186 7792
rect -1186 7712 1186 7728
rect -1186 7648 1102 7712
rect 1166 7648 1186 7712
rect -1186 7632 1186 7648
rect -1186 7568 1102 7632
rect 1166 7568 1186 7632
rect -1186 7552 1186 7568
rect -1186 7488 1102 7552
rect 1166 7488 1186 7552
rect -1186 7472 1186 7488
rect -1186 7408 1102 7472
rect 1166 7408 1186 7472
rect -1186 7392 1186 7408
rect -1186 7328 1102 7392
rect 1166 7328 1186 7392
rect -1186 7312 1186 7328
rect -1186 7248 1102 7312
rect 1166 7248 1186 7312
rect -1186 7232 1186 7248
rect -1186 7168 1102 7232
rect 1166 7168 1186 7232
rect -1186 7152 1186 7168
rect -1186 7088 1102 7152
rect 1166 7088 1186 7152
rect -1186 7072 1186 7088
rect -1186 7008 1102 7072
rect 1166 7008 1186 7072
rect -1186 6992 1186 7008
rect -1186 6928 1102 6992
rect 1166 6928 1186 6992
rect -1186 6912 1186 6928
rect -1186 6848 1102 6912
rect 1166 6848 1186 6912
rect -1186 6832 1186 6848
rect -1186 6768 1102 6832
rect 1166 6768 1186 6832
rect -1186 6752 1186 6768
rect -1186 6688 1102 6752
rect 1166 6688 1186 6752
rect -1186 6672 1186 6688
rect -1186 6608 1102 6672
rect 1166 6608 1186 6672
rect -1186 6592 1186 6608
rect -1186 6528 1102 6592
rect 1166 6528 1186 6592
rect -1186 6512 1186 6528
rect -1186 6448 1102 6512
rect 1166 6448 1186 6512
rect -1186 6432 1186 6448
rect -1186 6368 1102 6432
rect 1166 6368 1186 6432
rect -1186 6352 1186 6368
rect -1186 6288 1102 6352
rect 1166 6288 1186 6352
rect -1186 6272 1186 6288
rect -1186 6208 1102 6272
rect 1166 6208 1186 6272
rect -1186 6192 1186 6208
rect -1186 6128 1102 6192
rect 1166 6128 1186 6192
rect -1186 6112 1186 6128
rect -1186 6048 1102 6112
rect 1166 6048 1186 6112
rect -1186 6032 1186 6048
rect -1186 5968 1102 6032
rect 1166 5968 1186 6032
rect -1186 5920 1186 5968
rect 1426 7952 3798 8000
rect 1426 7888 3714 7952
rect 3778 7888 3798 7952
rect 1426 7872 3798 7888
rect 1426 7808 3714 7872
rect 3778 7808 3798 7872
rect 1426 7792 3798 7808
rect 1426 7728 3714 7792
rect 3778 7728 3798 7792
rect 1426 7712 3798 7728
rect 1426 7648 3714 7712
rect 3778 7648 3798 7712
rect 1426 7632 3798 7648
rect 1426 7568 3714 7632
rect 3778 7568 3798 7632
rect 1426 7552 3798 7568
rect 1426 7488 3714 7552
rect 3778 7488 3798 7552
rect 1426 7472 3798 7488
rect 1426 7408 3714 7472
rect 3778 7408 3798 7472
rect 1426 7392 3798 7408
rect 1426 7328 3714 7392
rect 3778 7328 3798 7392
rect 1426 7312 3798 7328
rect 1426 7248 3714 7312
rect 3778 7248 3798 7312
rect 1426 7232 3798 7248
rect 1426 7168 3714 7232
rect 3778 7168 3798 7232
rect 1426 7152 3798 7168
rect 1426 7088 3714 7152
rect 3778 7088 3798 7152
rect 1426 7072 3798 7088
rect 1426 7008 3714 7072
rect 3778 7008 3798 7072
rect 1426 6992 3798 7008
rect 1426 6928 3714 6992
rect 3778 6928 3798 6992
rect 1426 6912 3798 6928
rect 1426 6848 3714 6912
rect 3778 6848 3798 6912
rect 1426 6832 3798 6848
rect 1426 6768 3714 6832
rect 3778 6768 3798 6832
rect 1426 6752 3798 6768
rect 1426 6688 3714 6752
rect 3778 6688 3798 6752
rect 1426 6672 3798 6688
rect 1426 6608 3714 6672
rect 3778 6608 3798 6672
rect 1426 6592 3798 6608
rect 1426 6528 3714 6592
rect 3778 6528 3798 6592
rect 1426 6512 3798 6528
rect 1426 6448 3714 6512
rect 3778 6448 3798 6512
rect 1426 6432 3798 6448
rect 1426 6368 3714 6432
rect 3778 6368 3798 6432
rect 1426 6352 3798 6368
rect 1426 6288 3714 6352
rect 3778 6288 3798 6352
rect 1426 6272 3798 6288
rect 1426 6208 3714 6272
rect 3778 6208 3798 6272
rect 1426 6192 3798 6208
rect 1426 6128 3714 6192
rect 3778 6128 3798 6192
rect 1426 6112 3798 6128
rect 1426 6048 3714 6112
rect 3778 6048 3798 6112
rect 1426 6032 3798 6048
rect 1426 5968 3714 6032
rect 3778 5968 3798 6032
rect 1426 5920 3798 5968
rect 4038 7952 6410 8000
rect 4038 7888 6326 7952
rect 6390 7888 6410 7952
rect 4038 7872 6410 7888
rect 4038 7808 6326 7872
rect 6390 7808 6410 7872
rect 4038 7792 6410 7808
rect 4038 7728 6326 7792
rect 6390 7728 6410 7792
rect 4038 7712 6410 7728
rect 4038 7648 6326 7712
rect 6390 7648 6410 7712
rect 4038 7632 6410 7648
rect 4038 7568 6326 7632
rect 6390 7568 6410 7632
rect 4038 7552 6410 7568
rect 4038 7488 6326 7552
rect 6390 7488 6410 7552
rect 4038 7472 6410 7488
rect 4038 7408 6326 7472
rect 6390 7408 6410 7472
rect 4038 7392 6410 7408
rect 4038 7328 6326 7392
rect 6390 7328 6410 7392
rect 4038 7312 6410 7328
rect 4038 7248 6326 7312
rect 6390 7248 6410 7312
rect 4038 7232 6410 7248
rect 4038 7168 6326 7232
rect 6390 7168 6410 7232
rect 4038 7152 6410 7168
rect 4038 7088 6326 7152
rect 6390 7088 6410 7152
rect 4038 7072 6410 7088
rect 4038 7008 6326 7072
rect 6390 7008 6410 7072
rect 4038 6992 6410 7008
rect 4038 6928 6326 6992
rect 6390 6928 6410 6992
rect 4038 6912 6410 6928
rect 4038 6848 6326 6912
rect 6390 6848 6410 6912
rect 4038 6832 6410 6848
rect 4038 6768 6326 6832
rect 6390 6768 6410 6832
rect 4038 6752 6410 6768
rect 4038 6688 6326 6752
rect 6390 6688 6410 6752
rect 4038 6672 6410 6688
rect 4038 6608 6326 6672
rect 6390 6608 6410 6672
rect 4038 6592 6410 6608
rect 4038 6528 6326 6592
rect 6390 6528 6410 6592
rect 4038 6512 6410 6528
rect 4038 6448 6326 6512
rect 6390 6448 6410 6512
rect 4038 6432 6410 6448
rect 4038 6368 6326 6432
rect 6390 6368 6410 6432
rect 4038 6352 6410 6368
rect 4038 6288 6326 6352
rect 6390 6288 6410 6352
rect 4038 6272 6410 6288
rect 4038 6208 6326 6272
rect 6390 6208 6410 6272
rect 4038 6192 6410 6208
rect 4038 6128 6326 6192
rect 6390 6128 6410 6192
rect 4038 6112 6410 6128
rect 4038 6048 6326 6112
rect 6390 6048 6410 6112
rect 4038 6032 6410 6048
rect 4038 5968 6326 6032
rect 6390 5968 6410 6032
rect 4038 5920 6410 5968
rect 6650 7952 9022 8000
rect 6650 7888 8938 7952
rect 9002 7888 9022 7952
rect 6650 7872 9022 7888
rect 6650 7808 8938 7872
rect 9002 7808 9022 7872
rect 6650 7792 9022 7808
rect 6650 7728 8938 7792
rect 9002 7728 9022 7792
rect 6650 7712 9022 7728
rect 6650 7648 8938 7712
rect 9002 7648 9022 7712
rect 6650 7632 9022 7648
rect 6650 7568 8938 7632
rect 9002 7568 9022 7632
rect 6650 7552 9022 7568
rect 6650 7488 8938 7552
rect 9002 7488 9022 7552
rect 6650 7472 9022 7488
rect 6650 7408 8938 7472
rect 9002 7408 9022 7472
rect 6650 7392 9022 7408
rect 6650 7328 8938 7392
rect 9002 7328 9022 7392
rect 6650 7312 9022 7328
rect 6650 7248 8938 7312
rect 9002 7248 9022 7312
rect 6650 7232 9022 7248
rect 6650 7168 8938 7232
rect 9002 7168 9022 7232
rect 6650 7152 9022 7168
rect 6650 7088 8938 7152
rect 9002 7088 9022 7152
rect 6650 7072 9022 7088
rect 6650 7008 8938 7072
rect 9002 7008 9022 7072
rect 6650 6992 9022 7008
rect 6650 6928 8938 6992
rect 9002 6928 9022 6992
rect 6650 6912 9022 6928
rect 6650 6848 8938 6912
rect 9002 6848 9022 6912
rect 6650 6832 9022 6848
rect 6650 6768 8938 6832
rect 9002 6768 9022 6832
rect 6650 6752 9022 6768
rect 6650 6688 8938 6752
rect 9002 6688 9022 6752
rect 6650 6672 9022 6688
rect 6650 6608 8938 6672
rect 9002 6608 9022 6672
rect 6650 6592 9022 6608
rect 6650 6528 8938 6592
rect 9002 6528 9022 6592
rect 6650 6512 9022 6528
rect 6650 6448 8938 6512
rect 9002 6448 9022 6512
rect 6650 6432 9022 6448
rect 6650 6368 8938 6432
rect 9002 6368 9022 6432
rect 6650 6352 9022 6368
rect 6650 6288 8938 6352
rect 9002 6288 9022 6352
rect 6650 6272 9022 6288
rect 6650 6208 8938 6272
rect 9002 6208 9022 6272
rect 6650 6192 9022 6208
rect 6650 6128 8938 6192
rect 9002 6128 9022 6192
rect 6650 6112 9022 6128
rect 6650 6048 8938 6112
rect 9002 6048 9022 6112
rect 6650 6032 9022 6048
rect 6650 5968 8938 6032
rect 9002 5968 9022 6032
rect 6650 5920 9022 5968
rect -9022 5632 -6650 5680
rect -9022 5568 -6734 5632
rect -6670 5568 -6650 5632
rect -9022 5552 -6650 5568
rect -9022 5488 -6734 5552
rect -6670 5488 -6650 5552
rect -9022 5472 -6650 5488
rect -9022 5408 -6734 5472
rect -6670 5408 -6650 5472
rect -9022 5392 -6650 5408
rect -9022 5328 -6734 5392
rect -6670 5328 -6650 5392
rect -9022 5312 -6650 5328
rect -9022 5248 -6734 5312
rect -6670 5248 -6650 5312
rect -9022 5232 -6650 5248
rect -9022 5168 -6734 5232
rect -6670 5168 -6650 5232
rect -9022 5152 -6650 5168
rect -9022 5088 -6734 5152
rect -6670 5088 -6650 5152
rect -9022 5072 -6650 5088
rect -9022 5008 -6734 5072
rect -6670 5008 -6650 5072
rect -9022 4992 -6650 5008
rect -9022 4928 -6734 4992
rect -6670 4928 -6650 4992
rect -9022 4912 -6650 4928
rect -9022 4848 -6734 4912
rect -6670 4848 -6650 4912
rect -9022 4832 -6650 4848
rect -9022 4768 -6734 4832
rect -6670 4768 -6650 4832
rect -9022 4752 -6650 4768
rect -9022 4688 -6734 4752
rect -6670 4688 -6650 4752
rect -9022 4672 -6650 4688
rect -9022 4608 -6734 4672
rect -6670 4608 -6650 4672
rect -9022 4592 -6650 4608
rect -9022 4528 -6734 4592
rect -6670 4528 -6650 4592
rect -9022 4512 -6650 4528
rect -9022 4448 -6734 4512
rect -6670 4448 -6650 4512
rect -9022 4432 -6650 4448
rect -9022 4368 -6734 4432
rect -6670 4368 -6650 4432
rect -9022 4352 -6650 4368
rect -9022 4288 -6734 4352
rect -6670 4288 -6650 4352
rect -9022 4272 -6650 4288
rect -9022 4208 -6734 4272
rect -6670 4208 -6650 4272
rect -9022 4192 -6650 4208
rect -9022 4128 -6734 4192
rect -6670 4128 -6650 4192
rect -9022 4112 -6650 4128
rect -9022 4048 -6734 4112
rect -6670 4048 -6650 4112
rect -9022 4032 -6650 4048
rect -9022 3968 -6734 4032
rect -6670 3968 -6650 4032
rect -9022 3952 -6650 3968
rect -9022 3888 -6734 3952
rect -6670 3888 -6650 3952
rect -9022 3872 -6650 3888
rect -9022 3808 -6734 3872
rect -6670 3808 -6650 3872
rect -9022 3792 -6650 3808
rect -9022 3728 -6734 3792
rect -6670 3728 -6650 3792
rect -9022 3712 -6650 3728
rect -9022 3648 -6734 3712
rect -6670 3648 -6650 3712
rect -9022 3600 -6650 3648
rect -6410 5632 -4038 5680
rect -6410 5568 -4122 5632
rect -4058 5568 -4038 5632
rect -6410 5552 -4038 5568
rect -6410 5488 -4122 5552
rect -4058 5488 -4038 5552
rect -6410 5472 -4038 5488
rect -6410 5408 -4122 5472
rect -4058 5408 -4038 5472
rect -6410 5392 -4038 5408
rect -6410 5328 -4122 5392
rect -4058 5328 -4038 5392
rect -6410 5312 -4038 5328
rect -6410 5248 -4122 5312
rect -4058 5248 -4038 5312
rect -6410 5232 -4038 5248
rect -6410 5168 -4122 5232
rect -4058 5168 -4038 5232
rect -6410 5152 -4038 5168
rect -6410 5088 -4122 5152
rect -4058 5088 -4038 5152
rect -6410 5072 -4038 5088
rect -6410 5008 -4122 5072
rect -4058 5008 -4038 5072
rect -6410 4992 -4038 5008
rect -6410 4928 -4122 4992
rect -4058 4928 -4038 4992
rect -6410 4912 -4038 4928
rect -6410 4848 -4122 4912
rect -4058 4848 -4038 4912
rect -6410 4832 -4038 4848
rect -6410 4768 -4122 4832
rect -4058 4768 -4038 4832
rect -6410 4752 -4038 4768
rect -6410 4688 -4122 4752
rect -4058 4688 -4038 4752
rect -6410 4672 -4038 4688
rect -6410 4608 -4122 4672
rect -4058 4608 -4038 4672
rect -6410 4592 -4038 4608
rect -6410 4528 -4122 4592
rect -4058 4528 -4038 4592
rect -6410 4512 -4038 4528
rect -6410 4448 -4122 4512
rect -4058 4448 -4038 4512
rect -6410 4432 -4038 4448
rect -6410 4368 -4122 4432
rect -4058 4368 -4038 4432
rect -6410 4352 -4038 4368
rect -6410 4288 -4122 4352
rect -4058 4288 -4038 4352
rect -6410 4272 -4038 4288
rect -6410 4208 -4122 4272
rect -4058 4208 -4038 4272
rect -6410 4192 -4038 4208
rect -6410 4128 -4122 4192
rect -4058 4128 -4038 4192
rect -6410 4112 -4038 4128
rect -6410 4048 -4122 4112
rect -4058 4048 -4038 4112
rect -6410 4032 -4038 4048
rect -6410 3968 -4122 4032
rect -4058 3968 -4038 4032
rect -6410 3952 -4038 3968
rect -6410 3888 -4122 3952
rect -4058 3888 -4038 3952
rect -6410 3872 -4038 3888
rect -6410 3808 -4122 3872
rect -4058 3808 -4038 3872
rect -6410 3792 -4038 3808
rect -6410 3728 -4122 3792
rect -4058 3728 -4038 3792
rect -6410 3712 -4038 3728
rect -6410 3648 -4122 3712
rect -4058 3648 -4038 3712
rect -6410 3600 -4038 3648
rect -3798 5632 -1426 5680
rect -3798 5568 -1510 5632
rect -1446 5568 -1426 5632
rect -3798 5552 -1426 5568
rect -3798 5488 -1510 5552
rect -1446 5488 -1426 5552
rect -3798 5472 -1426 5488
rect -3798 5408 -1510 5472
rect -1446 5408 -1426 5472
rect -3798 5392 -1426 5408
rect -3798 5328 -1510 5392
rect -1446 5328 -1426 5392
rect -3798 5312 -1426 5328
rect -3798 5248 -1510 5312
rect -1446 5248 -1426 5312
rect -3798 5232 -1426 5248
rect -3798 5168 -1510 5232
rect -1446 5168 -1426 5232
rect -3798 5152 -1426 5168
rect -3798 5088 -1510 5152
rect -1446 5088 -1426 5152
rect -3798 5072 -1426 5088
rect -3798 5008 -1510 5072
rect -1446 5008 -1426 5072
rect -3798 4992 -1426 5008
rect -3798 4928 -1510 4992
rect -1446 4928 -1426 4992
rect -3798 4912 -1426 4928
rect -3798 4848 -1510 4912
rect -1446 4848 -1426 4912
rect -3798 4832 -1426 4848
rect -3798 4768 -1510 4832
rect -1446 4768 -1426 4832
rect -3798 4752 -1426 4768
rect -3798 4688 -1510 4752
rect -1446 4688 -1426 4752
rect -3798 4672 -1426 4688
rect -3798 4608 -1510 4672
rect -1446 4608 -1426 4672
rect -3798 4592 -1426 4608
rect -3798 4528 -1510 4592
rect -1446 4528 -1426 4592
rect -3798 4512 -1426 4528
rect -3798 4448 -1510 4512
rect -1446 4448 -1426 4512
rect -3798 4432 -1426 4448
rect -3798 4368 -1510 4432
rect -1446 4368 -1426 4432
rect -3798 4352 -1426 4368
rect -3798 4288 -1510 4352
rect -1446 4288 -1426 4352
rect -3798 4272 -1426 4288
rect -3798 4208 -1510 4272
rect -1446 4208 -1426 4272
rect -3798 4192 -1426 4208
rect -3798 4128 -1510 4192
rect -1446 4128 -1426 4192
rect -3798 4112 -1426 4128
rect -3798 4048 -1510 4112
rect -1446 4048 -1426 4112
rect -3798 4032 -1426 4048
rect -3798 3968 -1510 4032
rect -1446 3968 -1426 4032
rect -3798 3952 -1426 3968
rect -3798 3888 -1510 3952
rect -1446 3888 -1426 3952
rect -3798 3872 -1426 3888
rect -3798 3808 -1510 3872
rect -1446 3808 -1426 3872
rect -3798 3792 -1426 3808
rect -3798 3728 -1510 3792
rect -1446 3728 -1426 3792
rect -3798 3712 -1426 3728
rect -3798 3648 -1510 3712
rect -1446 3648 -1426 3712
rect -3798 3600 -1426 3648
rect -1186 5632 1186 5680
rect -1186 5568 1102 5632
rect 1166 5568 1186 5632
rect -1186 5552 1186 5568
rect -1186 5488 1102 5552
rect 1166 5488 1186 5552
rect -1186 5472 1186 5488
rect -1186 5408 1102 5472
rect 1166 5408 1186 5472
rect -1186 5392 1186 5408
rect -1186 5328 1102 5392
rect 1166 5328 1186 5392
rect -1186 5312 1186 5328
rect -1186 5248 1102 5312
rect 1166 5248 1186 5312
rect -1186 5232 1186 5248
rect -1186 5168 1102 5232
rect 1166 5168 1186 5232
rect -1186 5152 1186 5168
rect -1186 5088 1102 5152
rect 1166 5088 1186 5152
rect -1186 5072 1186 5088
rect -1186 5008 1102 5072
rect 1166 5008 1186 5072
rect -1186 4992 1186 5008
rect -1186 4928 1102 4992
rect 1166 4928 1186 4992
rect -1186 4912 1186 4928
rect -1186 4848 1102 4912
rect 1166 4848 1186 4912
rect -1186 4832 1186 4848
rect -1186 4768 1102 4832
rect 1166 4768 1186 4832
rect -1186 4752 1186 4768
rect -1186 4688 1102 4752
rect 1166 4688 1186 4752
rect -1186 4672 1186 4688
rect -1186 4608 1102 4672
rect 1166 4608 1186 4672
rect -1186 4592 1186 4608
rect -1186 4528 1102 4592
rect 1166 4528 1186 4592
rect -1186 4512 1186 4528
rect -1186 4448 1102 4512
rect 1166 4448 1186 4512
rect -1186 4432 1186 4448
rect -1186 4368 1102 4432
rect 1166 4368 1186 4432
rect -1186 4352 1186 4368
rect -1186 4288 1102 4352
rect 1166 4288 1186 4352
rect -1186 4272 1186 4288
rect -1186 4208 1102 4272
rect 1166 4208 1186 4272
rect -1186 4192 1186 4208
rect -1186 4128 1102 4192
rect 1166 4128 1186 4192
rect -1186 4112 1186 4128
rect -1186 4048 1102 4112
rect 1166 4048 1186 4112
rect -1186 4032 1186 4048
rect -1186 3968 1102 4032
rect 1166 3968 1186 4032
rect -1186 3952 1186 3968
rect -1186 3888 1102 3952
rect 1166 3888 1186 3952
rect -1186 3872 1186 3888
rect -1186 3808 1102 3872
rect 1166 3808 1186 3872
rect -1186 3792 1186 3808
rect -1186 3728 1102 3792
rect 1166 3728 1186 3792
rect -1186 3712 1186 3728
rect -1186 3648 1102 3712
rect 1166 3648 1186 3712
rect -1186 3600 1186 3648
rect 1426 5632 3798 5680
rect 1426 5568 3714 5632
rect 3778 5568 3798 5632
rect 1426 5552 3798 5568
rect 1426 5488 3714 5552
rect 3778 5488 3798 5552
rect 1426 5472 3798 5488
rect 1426 5408 3714 5472
rect 3778 5408 3798 5472
rect 1426 5392 3798 5408
rect 1426 5328 3714 5392
rect 3778 5328 3798 5392
rect 1426 5312 3798 5328
rect 1426 5248 3714 5312
rect 3778 5248 3798 5312
rect 1426 5232 3798 5248
rect 1426 5168 3714 5232
rect 3778 5168 3798 5232
rect 1426 5152 3798 5168
rect 1426 5088 3714 5152
rect 3778 5088 3798 5152
rect 1426 5072 3798 5088
rect 1426 5008 3714 5072
rect 3778 5008 3798 5072
rect 1426 4992 3798 5008
rect 1426 4928 3714 4992
rect 3778 4928 3798 4992
rect 1426 4912 3798 4928
rect 1426 4848 3714 4912
rect 3778 4848 3798 4912
rect 1426 4832 3798 4848
rect 1426 4768 3714 4832
rect 3778 4768 3798 4832
rect 1426 4752 3798 4768
rect 1426 4688 3714 4752
rect 3778 4688 3798 4752
rect 1426 4672 3798 4688
rect 1426 4608 3714 4672
rect 3778 4608 3798 4672
rect 1426 4592 3798 4608
rect 1426 4528 3714 4592
rect 3778 4528 3798 4592
rect 1426 4512 3798 4528
rect 1426 4448 3714 4512
rect 3778 4448 3798 4512
rect 1426 4432 3798 4448
rect 1426 4368 3714 4432
rect 3778 4368 3798 4432
rect 1426 4352 3798 4368
rect 1426 4288 3714 4352
rect 3778 4288 3798 4352
rect 1426 4272 3798 4288
rect 1426 4208 3714 4272
rect 3778 4208 3798 4272
rect 1426 4192 3798 4208
rect 1426 4128 3714 4192
rect 3778 4128 3798 4192
rect 1426 4112 3798 4128
rect 1426 4048 3714 4112
rect 3778 4048 3798 4112
rect 1426 4032 3798 4048
rect 1426 3968 3714 4032
rect 3778 3968 3798 4032
rect 1426 3952 3798 3968
rect 1426 3888 3714 3952
rect 3778 3888 3798 3952
rect 1426 3872 3798 3888
rect 1426 3808 3714 3872
rect 3778 3808 3798 3872
rect 1426 3792 3798 3808
rect 1426 3728 3714 3792
rect 3778 3728 3798 3792
rect 1426 3712 3798 3728
rect 1426 3648 3714 3712
rect 3778 3648 3798 3712
rect 1426 3600 3798 3648
rect 4038 5632 6410 5680
rect 4038 5568 6326 5632
rect 6390 5568 6410 5632
rect 4038 5552 6410 5568
rect 4038 5488 6326 5552
rect 6390 5488 6410 5552
rect 4038 5472 6410 5488
rect 4038 5408 6326 5472
rect 6390 5408 6410 5472
rect 4038 5392 6410 5408
rect 4038 5328 6326 5392
rect 6390 5328 6410 5392
rect 4038 5312 6410 5328
rect 4038 5248 6326 5312
rect 6390 5248 6410 5312
rect 4038 5232 6410 5248
rect 4038 5168 6326 5232
rect 6390 5168 6410 5232
rect 4038 5152 6410 5168
rect 4038 5088 6326 5152
rect 6390 5088 6410 5152
rect 4038 5072 6410 5088
rect 4038 5008 6326 5072
rect 6390 5008 6410 5072
rect 4038 4992 6410 5008
rect 4038 4928 6326 4992
rect 6390 4928 6410 4992
rect 4038 4912 6410 4928
rect 4038 4848 6326 4912
rect 6390 4848 6410 4912
rect 4038 4832 6410 4848
rect 4038 4768 6326 4832
rect 6390 4768 6410 4832
rect 4038 4752 6410 4768
rect 4038 4688 6326 4752
rect 6390 4688 6410 4752
rect 4038 4672 6410 4688
rect 4038 4608 6326 4672
rect 6390 4608 6410 4672
rect 4038 4592 6410 4608
rect 4038 4528 6326 4592
rect 6390 4528 6410 4592
rect 4038 4512 6410 4528
rect 4038 4448 6326 4512
rect 6390 4448 6410 4512
rect 4038 4432 6410 4448
rect 4038 4368 6326 4432
rect 6390 4368 6410 4432
rect 4038 4352 6410 4368
rect 4038 4288 6326 4352
rect 6390 4288 6410 4352
rect 4038 4272 6410 4288
rect 4038 4208 6326 4272
rect 6390 4208 6410 4272
rect 4038 4192 6410 4208
rect 4038 4128 6326 4192
rect 6390 4128 6410 4192
rect 4038 4112 6410 4128
rect 4038 4048 6326 4112
rect 6390 4048 6410 4112
rect 4038 4032 6410 4048
rect 4038 3968 6326 4032
rect 6390 3968 6410 4032
rect 4038 3952 6410 3968
rect 4038 3888 6326 3952
rect 6390 3888 6410 3952
rect 4038 3872 6410 3888
rect 4038 3808 6326 3872
rect 6390 3808 6410 3872
rect 4038 3792 6410 3808
rect 4038 3728 6326 3792
rect 6390 3728 6410 3792
rect 4038 3712 6410 3728
rect 4038 3648 6326 3712
rect 6390 3648 6410 3712
rect 4038 3600 6410 3648
rect 6650 5632 9022 5680
rect 6650 5568 8938 5632
rect 9002 5568 9022 5632
rect 6650 5552 9022 5568
rect 6650 5488 8938 5552
rect 9002 5488 9022 5552
rect 6650 5472 9022 5488
rect 6650 5408 8938 5472
rect 9002 5408 9022 5472
rect 6650 5392 9022 5408
rect 6650 5328 8938 5392
rect 9002 5328 9022 5392
rect 6650 5312 9022 5328
rect 6650 5248 8938 5312
rect 9002 5248 9022 5312
rect 6650 5232 9022 5248
rect 6650 5168 8938 5232
rect 9002 5168 9022 5232
rect 6650 5152 9022 5168
rect 6650 5088 8938 5152
rect 9002 5088 9022 5152
rect 6650 5072 9022 5088
rect 6650 5008 8938 5072
rect 9002 5008 9022 5072
rect 6650 4992 9022 5008
rect 6650 4928 8938 4992
rect 9002 4928 9022 4992
rect 6650 4912 9022 4928
rect 6650 4848 8938 4912
rect 9002 4848 9022 4912
rect 6650 4832 9022 4848
rect 6650 4768 8938 4832
rect 9002 4768 9022 4832
rect 6650 4752 9022 4768
rect 6650 4688 8938 4752
rect 9002 4688 9022 4752
rect 6650 4672 9022 4688
rect 6650 4608 8938 4672
rect 9002 4608 9022 4672
rect 6650 4592 9022 4608
rect 6650 4528 8938 4592
rect 9002 4528 9022 4592
rect 6650 4512 9022 4528
rect 6650 4448 8938 4512
rect 9002 4448 9022 4512
rect 6650 4432 9022 4448
rect 6650 4368 8938 4432
rect 9002 4368 9022 4432
rect 6650 4352 9022 4368
rect 6650 4288 8938 4352
rect 9002 4288 9022 4352
rect 6650 4272 9022 4288
rect 6650 4208 8938 4272
rect 9002 4208 9022 4272
rect 6650 4192 9022 4208
rect 6650 4128 8938 4192
rect 9002 4128 9022 4192
rect 6650 4112 9022 4128
rect 6650 4048 8938 4112
rect 9002 4048 9022 4112
rect 6650 4032 9022 4048
rect 6650 3968 8938 4032
rect 9002 3968 9022 4032
rect 6650 3952 9022 3968
rect 6650 3888 8938 3952
rect 9002 3888 9022 3952
rect 6650 3872 9022 3888
rect 6650 3808 8938 3872
rect 9002 3808 9022 3872
rect 6650 3792 9022 3808
rect 6650 3728 8938 3792
rect 9002 3728 9022 3792
rect 6650 3712 9022 3728
rect 6650 3648 8938 3712
rect 9002 3648 9022 3712
rect 6650 3600 9022 3648
rect -9022 3312 -6650 3360
rect -9022 3248 -6734 3312
rect -6670 3248 -6650 3312
rect -9022 3232 -6650 3248
rect -9022 3168 -6734 3232
rect -6670 3168 -6650 3232
rect -9022 3152 -6650 3168
rect -9022 3088 -6734 3152
rect -6670 3088 -6650 3152
rect -9022 3072 -6650 3088
rect -9022 3008 -6734 3072
rect -6670 3008 -6650 3072
rect -9022 2992 -6650 3008
rect -9022 2928 -6734 2992
rect -6670 2928 -6650 2992
rect -9022 2912 -6650 2928
rect -9022 2848 -6734 2912
rect -6670 2848 -6650 2912
rect -9022 2832 -6650 2848
rect -9022 2768 -6734 2832
rect -6670 2768 -6650 2832
rect -9022 2752 -6650 2768
rect -9022 2688 -6734 2752
rect -6670 2688 -6650 2752
rect -9022 2672 -6650 2688
rect -9022 2608 -6734 2672
rect -6670 2608 -6650 2672
rect -9022 2592 -6650 2608
rect -9022 2528 -6734 2592
rect -6670 2528 -6650 2592
rect -9022 2512 -6650 2528
rect -9022 2448 -6734 2512
rect -6670 2448 -6650 2512
rect -9022 2432 -6650 2448
rect -9022 2368 -6734 2432
rect -6670 2368 -6650 2432
rect -9022 2352 -6650 2368
rect -9022 2288 -6734 2352
rect -6670 2288 -6650 2352
rect -9022 2272 -6650 2288
rect -9022 2208 -6734 2272
rect -6670 2208 -6650 2272
rect -9022 2192 -6650 2208
rect -9022 2128 -6734 2192
rect -6670 2128 -6650 2192
rect -9022 2112 -6650 2128
rect -9022 2048 -6734 2112
rect -6670 2048 -6650 2112
rect -9022 2032 -6650 2048
rect -9022 1968 -6734 2032
rect -6670 1968 -6650 2032
rect -9022 1952 -6650 1968
rect -9022 1888 -6734 1952
rect -6670 1888 -6650 1952
rect -9022 1872 -6650 1888
rect -9022 1808 -6734 1872
rect -6670 1808 -6650 1872
rect -9022 1792 -6650 1808
rect -9022 1728 -6734 1792
rect -6670 1728 -6650 1792
rect -9022 1712 -6650 1728
rect -9022 1648 -6734 1712
rect -6670 1648 -6650 1712
rect -9022 1632 -6650 1648
rect -9022 1568 -6734 1632
rect -6670 1568 -6650 1632
rect -9022 1552 -6650 1568
rect -9022 1488 -6734 1552
rect -6670 1488 -6650 1552
rect -9022 1472 -6650 1488
rect -9022 1408 -6734 1472
rect -6670 1408 -6650 1472
rect -9022 1392 -6650 1408
rect -9022 1328 -6734 1392
rect -6670 1328 -6650 1392
rect -9022 1280 -6650 1328
rect -6410 3312 -4038 3360
rect -6410 3248 -4122 3312
rect -4058 3248 -4038 3312
rect -6410 3232 -4038 3248
rect -6410 3168 -4122 3232
rect -4058 3168 -4038 3232
rect -6410 3152 -4038 3168
rect -6410 3088 -4122 3152
rect -4058 3088 -4038 3152
rect -6410 3072 -4038 3088
rect -6410 3008 -4122 3072
rect -4058 3008 -4038 3072
rect -6410 2992 -4038 3008
rect -6410 2928 -4122 2992
rect -4058 2928 -4038 2992
rect -6410 2912 -4038 2928
rect -6410 2848 -4122 2912
rect -4058 2848 -4038 2912
rect -6410 2832 -4038 2848
rect -6410 2768 -4122 2832
rect -4058 2768 -4038 2832
rect -6410 2752 -4038 2768
rect -6410 2688 -4122 2752
rect -4058 2688 -4038 2752
rect -6410 2672 -4038 2688
rect -6410 2608 -4122 2672
rect -4058 2608 -4038 2672
rect -6410 2592 -4038 2608
rect -6410 2528 -4122 2592
rect -4058 2528 -4038 2592
rect -6410 2512 -4038 2528
rect -6410 2448 -4122 2512
rect -4058 2448 -4038 2512
rect -6410 2432 -4038 2448
rect -6410 2368 -4122 2432
rect -4058 2368 -4038 2432
rect -6410 2352 -4038 2368
rect -6410 2288 -4122 2352
rect -4058 2288 -4038 2352
rect -6410 2272 -4038 2288
rect -6410 2208 -4122 2272
rect -4058 2208 -4038 2272
rect -6410 2192 -4038 2208
rect -6410 2128 -4122 2192
rect -4058 2128 -4038 2192
rect -6410 2112 -4038 2128
rect -6410 2048 -4122 2112
rect -4058 2048 -4038 2112
rect -6410 2032 -4038 2048
rect -6410 1968 -4122 2032
rect -4058 1968 -4038 2032
rect -6410 1952 -4038 1968
rect -6410 1888 -4122 1952
rect -4058 1888 -4038 1952
rect -6410 1872 -4038 1888
rect -6410 1808 -4122 1872
rect -4058 1808 -4038 1872
rect -6410 1792 -4038 1808
rect -6410 1728 -4122 1792
rect -4058 1728 -4038 1792
rect -6410 1712 -4038 1728
rect -6410 1648 -4122 1712
rect -4058 1648 -4038 1712
rect -6410 1632 -4038 1648
rect -6410 1568 -4122 1632
rect -4058 1568 -4038 1632
rect -6410 1552 -4038 1568
rect -6410 1488 -4122 1552
rect -4058 1488 -4038 1552
rect -6410 1472 -4038 1488
rect -6410 1408 -4122 1472
rect -4058 1408 -4038 1472
rect -6410 1392 -4038 1408
rect -6410 1328 -4122 1392
rect -4058 1328 -4038 1392
rect -6410 1280 -4038 1328
rect -3798 3312 -1426 3360
rect -3798 3248 -1510 3312
rect -1446 3248 -1426 3312
rect -3798 3232 -1426 3248
rect -3798 3168 -1510 3232
rect -1446 3168 -1426 3232
rect -3798 3152 -1426 3168
rect -3798 3088 -1510 3152
rect -1446 3088 -1426 3152
rect -3798 3072 -1426 3088
rect -3798 3008 -1510 3072
rect -1446 3008 -1426 3072
rect -3798 2992 -1426 3008
rect -3798 2928 -1510 2992
rect -1446 2928 -1426 2992
rect -3798 2912 -1426 2928
rect -3798 2848 -1510 2912
rect -1446 2848 -1426 2912
rect -3798 2832 -1426 2848
rect -3798 2768 -1510 2832
rect -1446 2768 -1426 2832
rect -3798 2752 -1426 2768
rect -3798 2688 -1510 2752
rect -1446 2688 -1426 2752
rect -3798 2672 -1426 2688
rect -3798 2608 -1510 2672
rect -1446 2608 -1426 2672
rect -3798 2592 -1426 2608
rect -3798 2528 -1510 2592
rect -1446 2528 -1426 2592
rect -3798 2512 -1426 2528
rect -3798 2448 -1510 2512
rect -1446 2448 -1426 2512
rect -3798 2432 -1426 2448
rect -3798 2368 -1510 2432
rect -1446 2368 -1426 2432
rect -3798 2352 -1426 2368
rect -3798 2288 -1510 2352
rect -1446 2288 -1426 2352
rect -3798 2272 -1426 2288
rect -3798 2208 -1510 2272
rect -1446 2208 -1426 2272
rect -3798 2192 -1426 2208
rect -3798 2128 -1510 2192
rect -1446 2128 -1426 2192
rect -3798 2112 -1426 2128
rect -3798 2048 -1510 2112
rect -1446 2048 -1426 2112
rect -3798 2032 -1426 2048
rect -3798 1968 -1510 2032
rect -1446 1968 -1426 2032
rect -3798 1952 -1426 1968
rect -3798 1888 -1510 1952
rect -1446 1888 -1426 1952
rect -3798 1872 -1426 1888
rect -3798 1808 -1510 1872
rect -1446 1808 -1426 1872
rect -3798 1792 -1426 1808
rect -3798 1728 -1510 1792
rect -1446 1728 -1426 1792
rect -3798 1712 -1426 1728
rect -3798 1648 -1510 1712
rect -1446 1648 -1426 1712
rect -3798 1632 -1426 1648
rect -3798 1568 -1510 1632
rect -1446 1568 -1426 1632
rect -3798 1552 -1426 1568
rect -3798 1488 -1510 1552
rect -1446 1488 -1426 1552
rect -3798 1472 -1426 1488
rect -3798 1408 -1510 1472
rect -1446 1408 -1426 1472
rect -3798 1392 -1426 1408
rect -3798 1328 -1510 1392
rect -1446 1328 -1426 1392
rect -3798 1280 -1426 1328
rect -1186 3312 1186 3360
rect -1186 3248 1102 3312
rect 1166 3248 1186 3312
rect -1186 3232 1186 3248
rect -1186 3168 1102 3232
rect 1166 3168 1186 3232
rect -1186 3152 1186 3168
rect -1186 3088 1102 3152
rect 1166 3088 1186 3152
rect -1186 3072 1186 3088
rect -1186 3008 1102 3072
rect 1166 3008 1186 3072
rect -1186 2992 1186 3008
rect -1186 2928 1102 2992
rect 1166 2928 1186 2992
rect -1186 2912 1186 2928
rect -1186 2848 1102 2912
rect 1166 2848 1186 2912
rect -1186 2832 1186 2848
rect -1186 2768 1102 2832
rect 1166 2768 1186 2832
rect -1186 2752 1186 2768
rect -1186 2688 1102 2752
rect 1166 2688 1186 2752
rect -1186 2672 1186 2688
rect -1186 2608 1102 2672
rect 1166 2608 1186 2672
rect -1186 2592 1186 2608
rect -1186 2528 1102 2592
rect 1166 2528 1186 2592
rect -1186 2512 1186 2528
rect -1186 2448 1102 2512
rect 1166 2448 1186 2512
rect -1186 2432 1186 2448
rect -1186 2368 1102 2432
rect 1166 2368 1186 2432
rect -1186 2352 1186 2368
rect -1186 2288 1102 2352
rect 1166 2288 1186 2352
rect -1186 2272 1186 2288
rect -1186 2208 1102 2272
rect 1166 2208 1186 2272
rect -1186 2192 1186 2208
rect -1186 2128 1102 2192
rect 1166 2128 1186 2192
rect -1186 2112 1186 2128
rect -1186 2048 1102 2112
rect 1166 2048 1186 2112
rect -1186 2032 1186 2048
rect -1186 1968 1102 2032
rect 1166 1968 1186 2032
rect -1186 1952 1186 1968
rect -1186 1888 1102 1952
rect 1166 1888 1186 1952
rect -1186 1872 1186 1888
rect -1186 1808 1102 1872
rect 1166 1808 1186 1872
rect -1186 1792 1186 1808
rect -1186 1728 1102 1792
rect 1166 1728 1186 1792
rect -1186 1712 1186 1728
rect -1186 1648 1102 1712
rect 1166 1648 1186 1712
rect -1186 1632 1186 1648
rect -1186 1568 1102 1632
rect 1166 1568 1186 1632
rect -1186 1552 1186 1568
rect -1186 1488 1102 1552
rect 1166 1488 1186 1552
rect -1186 1472 1186 1488
rect -1186 1408 1102 1472
rect 1166 1408 1186 1472
rect -1186 1392 1186 1408
rect -1186 1328 1102 1392
rect 1166 1328 1186 1392
rect -1186 1280 1186 1328
rect 1426 3312 3798 3360
rect 1426 3248 3714 3312
rect 3778 3248 3798 3312
rect 1426 3232 3798 3248
rect 1426 3168 3714 3232
rect 3778 3168 3798 3232
rect 1426 3152 3798 3168
rect 1426 3088 3714 3152
rect 3778 3088 3798 3152
rect 1426 3072 3798 3088
rect 1426 3008 3714 3072
rect 3778 3008 3798 3072
rect 1426 2992 3798 3008
rect 1426 2928 3714 2992
rect 3778 2928 3798 2992
rect 1426 2912 3798 2928
rect 1426 2848 3714 2912
rect 3778 2848 3798 2912
rect 1426 2832 3798 2848
rect 1426 2768 3714 2832
rect 3778 2768 3798 2832
rect 1426 2752 3798 2768
rect 1426 2688 3714 2752
rect 3778 2688 3798 2752
rect 1426 2672 3798 2688
rect 1426 2608 3714 2672
rect 3778 2608 3798 2672
rect 1426 2592 3798 2608
rect 1426 2528 3714 2592
rect 3778 2528 3798 2592
rect 1426 2512 3798 2528
rect 1426 2448 3714 2512
rect 3778 2448 3798 2512
rect 1426 2432 3798 2448
rect 1426 2368 3714 2432
rect 3778 2368 3798 2432
rect 1426 2352 3798 2368
rect 1426 2288 3714 2352
rect 3778 2288 3798 2352
rect 1426 2272 3798 2288
rect 1426 2208 3714 2272
rect 3778 2208 3798 2272
rect 1426 2192 3798 2208
rect 1426 2128 3714 2192
rect 3778 2128 3798 2192
rect 1426 2112 3798 2128
rect 1426 2048 3714 2112
rect 3778 2048 3798 2112
rect 1426 2032 3798 2048
rect 1426 1968 3714 2032
rect 3778 1968 3798 2032
rect 1426 1952 3798 1968
rect 1426 1888 3714 1952
rect 3778 1888 3798 1952
rect 1426 1872 3798 1888
rect 1426 1808 3714 1872
rect 3778 1808 3798 1872
rect 1426 1792 3798 1808
rect 1426 1728 3714 1792
rect 3778 1728 3798 1792
rect 1426 1712 3798 1728
rect 1426 1648 3714 1712
rect 3778 1648 3798 1712
rect 1426 1632 3798 1648
rect 1426 1568 3714 1632
rect 3778 1568 3798 1632
rect 1426 1552 3798 1568
rect 1426 1488 3714 1552
rect 3778 1488 3798 1552
rect 1426 1472 3798 1488
rect 1426 1408 3714 1472
rect 3778 1408 3798 1472
rect 1426 1392 3798 1408
rect 1426 1328 3714 1392
rect 3778 1328 3798 1392
rect 1426 1280 3798 1328
rect 4038 3312 6410 3360
rect 4038 3248 6326 3312
rect 6390 3248 6410 3312
rect 4038 3232 6410 3248
rect 4038 3168 6326 3232
rect 6390 3168 6410 3232
rect 4038 3152 6410 3168
rect 4038 3088 6326 3152
rect 6390 3088 6410 3152
rect 4038 3072 6410 3088
rect 4038 3008 6326 3072
rect 6390 3008 6410 3072
rect 4038 2992 6410 3008
rect 4038 2928 6326 2992
rect 6390 2928 6410 2992
rect 4038 2912 6410 2928
rect 4038 2848 6326 2912
rect 6390 2848 6410 2912
rect 4038 2832 6410 2848
rect 4038 2768 6326 2832
rect 6390 2768 6410 2832
rect 4038 2752 6410 2768
rect 4038 2688 6326 2752
rect 6390 2688 6410 2752
rect 4038 2672 6410 2688
rect 4038 2608 6326 2672
rect 6390 2608 6410 2672
rect 4038 2592 6410 2608
rect 4038 2528 6326 2592
rect 6390 2528 6410 2592
rect 4038 2512 6410 2528
rect 4038 2448 6326 2512
rect 6390 2448 6410 2512
rect 4038 2432 6410 2448
rect 4038 2368 6326 2432
rect 6390 2368 6410 2432
rect 4038 2352 6410 2368
rect 4038 2288 6326 2352
rect 6390 2288 6410 2352
rect 4038 2272 6410 2288
rect 4038 2208 6326 2272
rect 6390 2208 6410 2272
rect 4038 2192 6410 2208
rect 4038 2128 6326 2192
rect 6390 2128 6410 2192
rect 4038 2112 6410 2128
rect 4038 2048 6326 2112
rect 6390 2048 6410 2112
rect 4038 2032 6410 2048
rect 4038 1968 6326 2032
rect 6390 1968 6410 2032
rect 4038 1952 6410 1968
rect 4038 1888 6326 1952
rect 6390 1888 6410 1952
rect 4038 1872 6410 1888
rect 4038 1808 6326 1872
rect 6390 1808 6410 1872
rect 4038 1792 6410 1808
rect 4038 1728 6326 1792
rect 6390 1728 6410 1792
rect 4038 1712 6410 1728
rect 4038 1648 6326 1712
rect 6390 1648 6410 1712
rect 4038 1632 6410 1648
rect 4038 1568 6326 1632
rect 6390 1568 6410 1632
rect 4038 1552 6410 1568
rect 4038 1488 6326 1552
rect 6390 1488 6410 1552
rect 4038 1472 6410 1488
rect 4038 1408 6326 1472
rect 6390 1408 6410 1472
rect 4038 1392 6410 1408
rect 4038 1328 6326 1392
rect 6390 1328 6410 1392
rect 4038 1280 6410 1328
rect 6650 3312 9022 3360
rect 6650 3248 8938 3312
rect 9002 3248 9022 3312
rect 6650 3232 9022 3248
rect 6650 3168 8938 3232
rect 9002 3168 9022 3232
rect 6650 3152 9022 3168
rect 6650 3088 8938 3152
rect 9002 3088 9022 3152
rect 6650 3072 9022 3088
rect 6650 3008 8938 3072
rect 9002 3008 9022 3072
rect 6650 2992 9022 3008
rect 6650 2928 8938 2992
rect 9002 2928 9022 2992
rect 6650 2912 9022 2928
rect 6650 2848 8938 2912
rect 9002 2848 9022 2912
rect 6650 2832 9022 2848
rect 6650 2768 8938 2832
rect 9002 2768 9022 2832
rect 6650 2752 9022 2768
rect 6650 2688 8938 2752
rect 9002 2688 9022 2752
rect 6650 2672 9022 2688
rect 6650 2608 8938 2672
rect 9002 2608 9022 2672
rect 6650 2592 9022 2608
rect 6650 2528 8938 2592
rect 9002 2528 9022 2592
rect 6650 2512 9022 2528
rect 6650 2448 8938 2512
rect 9002 2448 9022 2512
rect 6650 2432 9022 2448
rect 6650 2368 8938 2432
rect 9002 2368 9022 2432
rect 6650 2352 9022 2368
rect 6650 2288 8938 2352
rect 9002 2288 9022 2352
rect 6650 2272 9022 2288
rect 6650 2208 8938 2272
rect 9002 2208 9022 2272
rect 6650 2192 9022 2208
rect 6650 2128 8938 2192
rect 9002 2128 9022 2192
rect 6650 2112 9022 2128
rect 6650 2048 8938 2112
rect 9002 2048 9022 2112
rect 6650 2032 9022 2048
rect 6650 1968 8938 2032
rect 9002 1968 9022 2032
rect 6650 1952 9022 1968
rect 6650 1888 8938 1952
rect 9002 1888 9022 1952
rect 6650 1872 9022 1888
rect 6650 1808 8938 1872
rect 9002 1808 9022 1872
rect 6650 1792 9022 1808
rect 6650 1728 8938 1792
rect 9002 1728 9022 1792
rect 6650 1712 9022 1728
rect 6650 1648 8938 1712
rect 9002 1648 9022 1712
rect 6650 1632 9022 1648
rect 6650 1568 8938 1632
rect 9002 1568 9022 1632
rect 6650 1552 9022 1568
rect 6650 1488 8938 1552
rect 9002 1488 9022 1552
rect 6650 1472 9022 1488
rect 6650 1408 8938 1472
rect 9002 1408 9022 1472
rect 6650 1392 9022 1408
rect 6650 1328 8938 1392
rect 9002 1328 9022 1392
rect 6650 1280 9022 1328
rect -9022 992 -6650 1040
rect -9022 928 -6734 992
rect -6670 928 -6650 992
rect -9022 912 -6650 928
rect -9022 848 -6734 912
rect -6670 848 -6650 912
rect -9022 832 -6650 848
rect -9022 768 -6734 832
rect -6670 768 -6650 832
rect -9022 752 -6650 768
rect -9022 688 -6734 752
rect -6670 688 -6650 752
rect -9022 672 -6650 688
rect -9022 608 -6734 672
rect -6670 608 -6650 672
rect -9022 592 -6650 608
rect -9022 528 -6734 592
rect -6670 528 -6650 592
rect -9022 512 -6650 528
rect -9022 448 -6734 512
rect -6670 448 -6650 512
rect -9022 432 -6650 448
rect -9022 368 -6734 432
rect -6670 368 -6650 432
rect -9022 352 -6650 368
rect -9022 288 -6734 352
rect -6670 288 -6650 352
rect -9022 272 -6650 288
rect -9022 208 -6734 272
rect -6670 208 -6650 272
rect -9022 192 -6650 208
rect -9022 128 -6734 192
rect -6670 128 -6650 192
rect -9022 112 -6650 128
rect -9022 48 -6734 112
rect -6670 48 -6650 112
rect -9022 32 -6650 48
rect -9022 -32 -6734 32
rect -6670 -32 -6650 32
rect -9022 -48 -6650 -32
rect -9022 -112 -6734 -48
rect -6670 -112 -6650 -48
rect -9022 -128 -6650 -112
rect -9022 -192 -6734 -128
rect -6670 -192 -6650 -128
rect -9022 -208 -6650 -192
rect -9022 -272 -6734 -208
rect -6670 -272 -6650 -208
rect -9022 -288 -6650 -272
rect -9022 -352 -6734 -288
rect -6670 -352 -6650 -288
rect -9022 -368 -6650 -352
rect -9022 -432 -6734 -368
rect -6670 -432 -6650 -368
rect -9022 -448 -6650 -432
rect -9022 -512 -6734 -448
rect -6670 -512 -6650 -448
rect -9022 -528 -6650 -512
rect -9022 -592 -6734 -528
rect -6670 -592 -6650 -528
rect -9022 -608 -6650 -592
rect -9022 -672 -6734 -608
rect -6670 -672 -6650 -608
rect -9022 -688 -6650 -672
rect -9022 -752 -6734 -688
rect -6670 -752 -6650 -688
rect -9022 -768 -6650 -752
rect -9022 -832 -6734 -768
rect -6670 -832 -6650 -768
rect -9022 -848 -6650 -832
rect -9022 -912 -6734 -848
rect -6670 -912 -6650 -848
rect -9022 -928 -6650 -912
rect -9022 -992 -6734 -928
rect -6670 -992 -6650 -928
rect -9022 -1040 -6650 -992
rect -6410 992 -4038 1040
rect -6410 928 -4122 992
rect -4058 928 -4038 992
rect -6410 912 -4038 928
rect -6410 848 -4122 912
rect -4058 848 -4038 912
rect -6410 832 -4038 848
rect -6410 768 -4122 832
rect -4058 768 -4038 832
rect -6410 752 -4038 768
rect -6410 688 -4122 752
rect -4058 688 -4038 752
rect -6410 672 -4038 688
rect -6410 608 -4122 672
rect -4058 608 -4038 672
rect -6410 592 -4038 608
rect -6410 528 -4122 592
rect -4058 528 -4038 592
rect -6410 512 -4038 528
rect -6410 448 -4122 512
rect -4058 448 -4038 512
rect -6410 432 -4038 448
rect -6410 368 -4122 432
rect -4058 368 -4038 432
rect -6410 352 -4038 368
rect -6410 288 -4122 352
rect -4058 288 -4038 352
rect -6410 272 -4038 288
rect -6410 208 -4122 272
rect -4058 208 -4038 272
rect -6410 192 -4038 208
rect -6410 128 -4122 192
rect -4058 128 -4038 192
rect -6410 112 -4038 128
rect -6410 48 -4122 112
rect -4058 48 -4038 112
rect -6410 32 -4038 48
rect -6410 -32 -4122 32
rect -4058 -32 -4038 32
rect -6410 -48 -4038 -32
rect -6410 -112 -4122 -48
rect -4058 -112 -4038 -48
rect -6410 -128 -4038 -112
rect -6410 -192 -4122 -128
rect -4058 -192 -4038 -128
rect -6410 -208 -4038 -192
rect -6410 -272 -4122 -208
rect -4058 -272 -4038 -208
rect -6410 -288 -4038 -272
rect -6410 -352 -4122 -288
rect -4058 -352 -4038 -288
rect -6410 -368 -4038 -352
rect -6410 -432 -4122 -368
rect -4058 -432 -4038 -368
rect -6410 -448 -4038 -432
rect -6410 -512 -4122 -448
rect -4058 -512 -4038 -448
rect -6410 -528 -4038 -512
rect -6410 -592 -4122 -528
rect -4058 -592 -4038 -528
rect -6410 -608 -4038 -592
rect -6410 -672 -4122 -608
rect -4058 -672 -4038 -608
rect -6410 -688 -4038 -672
rect -6410 -752 -4122 -688
rect -4058 -752 -4038 -688
rect -6410 -768 -4038 -752
rect -6410 -832 -4122 -768
rect -4058 -832 -4038 -768
rect -6410 -848 -4038 -832
rect -6410 -912 -4122 -848
rect -4058 -912 -4038 -848
rect -6410 -928 -4038 -912
rect -6410 -992 -4122 -928
rect -4058 -992 -4038 -928
rect -6410 -1040 -4038 -992
rect -3798 992 -1426 1040
rect -3798 928 -1510 992
rect -1446 928 -1426 992
rect -3798 912 -1426 928
rect -3798 848 -1510 912
rect -1446 848 -1426 912
rect -3798 832 -1426 848
rect -3798 768 -1510 832
rect -1446 768 -1426 832
rect -3798 752 -1426 768
rect -3798 688 -1510 752
rect -1446 688 -1426 752
rect -3798 672 -1426 688
rect -3798 608 -1510 672
rect -1446 608 -1426 672
rect -3798 592 -1426 608
rect -3798 528 -1510 592
rect -1446 528 -1426 592
rect -3798 512 -1426 528
rect -3798 448 -1510 512
rect -1446 448 -1426 512
rect -3798 432 -1426 448
rect -3798 368 -1510 432
rect -1446 368 -1426 432
rect -3798 352 -1426 368
rect -3798 288 -1510 352
rect -1446 288 -1426 352
rect -3798 272 -1426 288
rect -3798 208 -1510 272
rect -1446 208 -1426 272
rect -3798 192 -1426 208
rect -3798 128 -1510 192
rect -1446 128 -1426 192
rect -3798 112 -1426 128
rect -3798 48 -1510 112
rect -1446 48 -1426 112
rect -3798 32 -1426 48
rect -3798 -32 -1510 32
rect -1446 -32 -1426 32
rect -3798 -48 -1426 -32
rect -3798 -112 -1510 -48
rect -1446 -112 -1426 -48
rect -3798 -128 -1426 -112
rect -3798 -192 -1510 -128
rect -1446 -192 -1426 -128
rect -3798 -208 -1426 -192
rect -3798 -272 -1510 -208
rect -1446 -272 -1426 -208
rect -3798 -288 -1426 -272
rect -3798 -352 -1510 -288
rect -1446 -352 -1426 -288
rect -3798 -368 -1426 -352
rect -3798 -432 -1510 -368
rect -1446 -432 -1426 -368
rect -3798 -448 -1426 -432
rect -3798 -512 -1510 -448
rect -1446 -512 -1426 -448
rect -3798 -528 -1426 -512
rect -3798 -592 -1510 -528
rect -1446 -592 -1426 -528
rect -3798 -608 -1426 -592
rect -3798 -672 -1510 -608
rect -1446 -672 -1426 -608
rect -3798 -688 -1426 -672
rect -3798 -752 -1510 -688
rect -1446 -752 -1426 -688
rect -3798 -768 -1426 -752
rect -3798 -832 -1510 -768
rect -1446 -832 -1426 -768
rect -3798 -848 -1426 -832
rect -3798 -912 -1510 -848
rect -1446 -912 -1426 -848
rect -3798 -928 -1426 -912
rect -3798 -992 -1510 -928
rect -1446 -992 -1426 -928
rect -3798 -1040 -1426 -992
rect -1186 992 1186 1040
rect -1186 928 1102 992
rect 1166 928 1186 992
rect -1186 912 1186 928
rect -1186 848 1102 912
rect 1166 848 1186 912
rect -1186 832 1186 848
rect -1186 768 1102 832
rect 1166 768 1186 832
rect -1186 752 1186 768
rect -1186 688 1102 752
rect 1166 688 1186 752
rect -1186 672 1186 688
rect -1186 608 1102 672
rect 1166 608 1186 672
rect -1186 592 1186 608
rect -1186 528 1102 592
rect 1166 528 1186 592
rect -1186 512 1186 528
rect -1186 448 1102 512
rect 1166 448 1186 512
rect -1186 432 1186 448
rect -1186 368 1102 432
rect 1166 368 1186 432
rect -1186 352 1186 368
rect -1186 288 1102 352
rect 1166 288 1186 352
rect -1186 272 1186 288
rect -1186 208 1102 272
rect 1166 208 1186 272
rect -1186 192 1186 208
rect -1186 128 1102 192
rect 1166 128 1186 192
rect -1186 112 1186 128
rect -1186 48 1102 112
rect 1166 48 1186 112
rect -1186 32 1186 48
rect -1186 -32 1102 32
rect 1166 -32 1186 32
rect -1186 -48 1186 -32
rect -1186 -112 1102 -48
rect 1166 -112 1186 -48
rect -1186 -128 1186 -112
rect -1186 -192 1102 -128
rect 1166 -192 1186 -128
rect -1186 -208 1186 -192
rect -1186 -272 1102 -208
rect 1166 -272 1186 -208
rect -1186 -288 1186 -272
rect -1186 -352 1102 -288
rect 1166 -352 1186 -288
rect -1186 -368 1186 -352
rect -1186 -432 1102 -368
rect 1166 -432 1186 -368
rect -1186 -448 1186 -432
rect -1186 -512 1102 -448
rect 1166 -512 1186 -448
rect -1186 -528 1186 -512
rect -1186 -592 1102 -528
rect 1166 -592 1186 -528
rect -1186 -608 1186 -592
rect -1186 -672 1102 -608
rect 1166 -672 1186 -608
rect -1186 -688 1186 -672
rect -1186 -752 1102 -688
rect 1166 -752 1186 -688
rect -1186 -768 1186 -752
rect -1186 -832 1102 -768
rect 1166 -832 1186 -768
rect -1186 -848 1186 -832
rect -1186 -912 1102 -848
rect 1166 -912 1186 -848
rect -1186 -928 1186 -912
rect -1186 -992 1102 -928
rect 1166 -992 1186 -928
rect -1186 -1040 1186 -992
rect 1426 992 3798 1040
rect 1426 928 3714 992
rect 3778 928 3798 992
rect 1426 912 3798 928
rect 1426 848 3714 912
rect 3778 848 3798 912
rect 1426 832 3798 848
rect 1426 768 3714 832
rect 3778 768 3798 832
rect 1426 752 3798 768
rect 1426 688 3714 752
rect 3778 688 3798 752
rect 1426 672 3798 688
rect 1426 608 3714 672
rect 3778 608 3798 672
rect 1426 592 3798 608
rect 1426 528 3714 592
rect 3778 528 3798 592
rect 1426 512 3798 528
rect 1426 448 3714 512
rect 3778 448 3798 512
rect 1426 432 3798 448
rect 1426 368 3714 432
rect 3778 368 3798 432
rect 1426 352 3798 368
rect 1426 288 3714 352
rect 3778 288 3798 352
rect 1426 272 3798 288
rect 1426 208 3714 272
rect 3778 208 3798 272
rect 1426 192 3798 208
rect 1426 128 3714 192
rect 3778 128 3798 192
rect 1426 112 3798 128
rect 1426 48 3714 112
rect 3778 48 3798 112
rect 1426 32 3798 48
rect 1426 -32 3714 32
rect 3778 -32 3798 32
rect 1426 -48 3798 -32
rect 1426 -112 3714 -48
rect 3778 -112 3798 -48
rect 1426 -128 3798 -112
rect 1426 -192 3714 -128
rect 3778 -192 3798 -128
rect 1426 -208 3798 -192
rect 1426 -272 3714 -208
rect 3778 -272 3798 -208
rect 1426 -288 3798 -272
rect 1426 -352 3714 -288
rect 3778 -352 3798 -288
rect 1426 -368 3798 -352
rect 1426 -432 3714 -368
rect 3778 -432 3798 -368
rect 1426 -448 3798 -432
rect 1426 -512 3714 -448
rect 3778 -512 3798 -448
rect 1426 -528 3798 -512
rect 1426 -592 3714 -528
rect 3778 -592 3798 -528
rect 1426 -608 3798 -592
rect 1426 -672 3714 -608
rect 3778 -672 3798 -608
rect 1426 -688 3798 -672
rect 1426 -752 3714 -688
rect 3778 -752 3798 -688
rect 1426 -768 3798 -752
rect 1426 -832 3714 -768
rect 3778 -832 3798 -768
rect 1426 -848 3798 -832
rect 1426 -912 3714 -848
rect 3778 -912 3798 -848
rect 1426 -928 3798 -912
rect 1426 -992 3714 -928
rect 3778 -992 3798 -928
rect 1426 -1040 3798 -992
rect 4038 992 6410 1040
rect 4038 928 6326 992
rect 6390 928 6410 992
rect 4038 912 6410 928
rect 4038 848 6326 912
rect 6390 848 6410 912
rect 4038 832 6410 848
rect 4038 768 6326 832
rect 6390 768 6410 832
rect 4038 752 6410 768
rect 4038 688 6326 752
rect 6390 688 6410 752
rect 4038 672 6410 688
rect 4038 608 6326 672
rect 6390 608 6410 672
rect 4038 592 6410 608
rect 4038 528 6326 592
rect 6390 528 6410 592
rect 4038 512 6410 528
rect 4038 448 6326 512
rect 6390 448 6410 512
rect 4038 432 6410 448
rect 4038 368 6326 432
rect 6390 368 6410 432
rect 4038 352 6410 368
rect 4038 288 6326 352
rect 6390 288 6410 352
rect 4038 272 6410 288
rect 4038 208 6326 272
rect 6390 208 6410 272
rect 4038 192 6410 208
rect 4038 128 6326 192
rect 6390 128 6410 192
rect 4038 112 6410 128
rect 4038 48 6326 112
rect 6390 48 6410 112
rect 4038 32 6410 48
rect 4038 -32 6326 32
rect 6390 -32 6410 32
rect 4038 -48 6410 -32
rect 4038 -112 6326 -48
rect 6390 -112 6410 -48
rect 4038 -128 6410 -112
rect 4038 -192 6326 -128
rect 6390 -192 6410 -128
rect 4038 -208 6410 -192
rect 4038 -272 6326 -208
rect 6390 -272 6410 -208
rect 4038 -288 6410 -272
rect 4038 -352 6326 -288
rect 6390 -352 6410 -288
rect 4038 -368 6410 -352
rect 4038 -432 6326 -368
rect 6390 -432 6410 -368
rect 4038 -448 6410 -432
rect 4038 -512 6326 -448
rect 6390 -512 6410 -448
rect 4038 -528 6410 -512
rect 4038 -592 6326 -528
rect 6390 -592 6410 -528
rect 4038 -608 6410 -592
rect 4038 -672 6326 -608
rect 6390 -672 6410 -608
rect 4038 -688 6410 -672
rect 4038 -752 6326 -688
rect 6390 -752 6410 -688
rect 4038 -768 6410 -752
rect 4038 -832 6326 -768
rect 6390 -832 6410 -768
rect 4038 -848 6410 -832
rect 4038 -912 6326 -848
rect 6390 -912 6410 -848
rect 4038 -928 6410 -912
rect 4038 -992 6326 -928
rect 6390 -992 6410 -928
rect 4038 -1040 6410 -992
rect 6650 992 9022 1040
rect 6650 928 8938 992
rect 9002 928 9022 992
rect 6650 912 9022 928
rect 6650 848 8938 912
rect 9002 848 9022 912
rect 6650 832 9022 848
rect 6650 768 8938 832
rect 9002 768 9022 832
rect 6650 752 9022 768
rect 6650 688 8938 752
rect 9002 688 9022 752
rect 6650 672 9022 688
rect 6650 608 8938 672
rect 9002 608 9022 672
rect 6650 592 9022 608
rect 6650 528 8938 592
rect 9002 528 9022 592
rect 6650 512 9022 528
rect 6650 448 8938 512
rect 9002 448 9022 512
rect 6650 432 9022 448
rect 6650 368 8938 432
rect 9002 368 9022 432
rect 6650 352 9022 368
rect 6650 288 8938 352
rect 9002 288 9022 352
rect 6650 272 9022 288
rect 6650 208 8938 272
rect 9002 208 9022 272
rect 6650 192 9022 208
rect 6650 128 8938 192
rect 9002 128 9022 192
rect 6650 112 9022 128
rect 6650 48 8938 112
rect 9002 48 9022 112
rect 6650 32 9022 48
rect 6650 -32 8938 32
rect 9002 -32 9022 32
rect 6650 -48 9022 -32
rect 6650 -112 8938 -48
rect 9002 -112 9022 -48
rect 6650 -128 9022 -112
rect 6650 -192 8938 -128
rect 9002 -192 9022 -128
rect 6650 -208 9022 -192
rect 6650 -272 8938 -208
rect 9002 -272 9022 -208
rect 6650 -288 9022 -272
rect 6650 -352 8938 -288
rect 9002 -352 9022 -288
rect 6650 -368 9022 -352
rect 6650 -432 8938 -368
rect 9002 -432 9022 -368
rect 6650 -448 9022 -432
rect 6650 -512 8938 -448
rect 9002 -512 9022 -448
rect 6650 -528 9022 -512
rect 6650 -592 8938 -528
rect 9002 -592 9022 -528
rect 6650 -608 9022 -592
rect 6650 -672 8938 -608
rect 9002 -672 9022 -608
rect 6650 -688 9022 -672
rect 6650 -752 8938 -688
rect 9002 -752 9022 -688
rect 6650 -768 9022 -752
rect 6650 -832 8938 -768
rect 9002 -832 9022 -768
rect 6650 -848 9022 -832
rect 6650 -912 8938 -848
rect 9002 -912 9022 -848
rect 6650 -928 9022 -912
rect 6650 -992 8938 -928
rect 9002 -992 9022 -928
rect 6650 -1040 9022 -992
rect -9022 -1328 -6650 -1280
rect -9022 -1392 -6734 -1328
rect -6670 -1392 -6650 -1328
rect -9022 -1408 -6650 -1392
rect -9022 -1472 -6734 -1408
rect -6670 -1472 -6650 -1408
rect -9022 -1488 -6650 -1472
rect -9022 -1552 -6734 -1488
rect -6670 -1552 -6650 -1488
rect -9022 -1568 -6650 -1552
rect -9022 -1632 -6734 -1568
rect -6670 -1632 -6650 -1568
rect -9022 -1648 -6650 -1632
rect -9022 -1712 -6734 -1648
rect -6670 -1712 -6650 -1648
rect -9022 -1728 -6650 -1712
rect -9022 -1792 -6734 -1728
rect -6670 -1792 -6650 -1728
rect -9022 -1808 -6650 -1792
rect -9022 -1872 -6734 -1808
rect -6670 -1872 -6650 -1808
rect -9022 -1888 -6650 -1872
rect -9022 -1952 -6734 -1888
rect -6670 -1952 -6650 -1888
rect -9022 -1968 -6650 -1952
rect -9022 -2032 -6734 -1968
rect -6670 -2032 -6650 -1968
rect -9022 -2048 -6650 -2032
rect -9022 -2112 -6734 -2048
rect -6670 -2112 -6650 -2048
rect -9022 -2128 -6650 -2112
rect -9022 -2192 -6734 -2128
rect -6670 -2192 -6650 -2128
rect -9022 -2208 -6650 -2192
rect -9022 -2272 -6734 -2208
rect -6670 -2272 -6650 -2208
rect -9022 -2288 -6650 -2272
rect -9022 -2352 -6734 -2288
rect -6670 -2352 -6650 -2288
rect -9022 -2368 -6650 -2352
rect -9022 -2432 -6734 -2368
rect -6670 -2432 -6650 -2368
rect -9022 -2448 -6650 -2432
rect -9022 -2512 -6734 -2448
rect -6670 -2512 -6650 -2448
rect -9022 -2528 -6650 -2512
rect -9022 -2592 -6734 -2528
rect -6670 -2592 -6650 -2528
rect -9022 -2608 -6650 -2592
rect -9022 -2672 -6734 -2608
rect -6670 -2672 -6650 -2608
rect -9022 -2688 -6650 -2672
rect -9022 -2752 -6734 -2688
rect -6670 -2752 -6650 -2688
rect -9022 -2768 -6650 -2752
rect -9022 -2832 -6734 -2768
rect -6670 -2832 -6650 -2768
rect -9022 -2848 -6650 -2832
rect -9022 -2912 -6734 -2848
rect -6670 -2912 -6650 -2848
rect -9022 -2928 -6650 -2912
rect -9022 -2992 -6734 -2928
rect -6670 -2992 -6650 -2928
rect -9022 -3008 -6650 -2992
rect -9022 -3072 -6734 -3008
rect -6670 -3072 -6650 -3008
rect -9022 -3088 -6650 -3072
rect -9022 -3152 -6734 -3088
rect -6670 -3152 -6650 -3088
rect -9022 -3168 -6650 -3152
rect -9022 -3232 -6734 -3168
rect -6670 -3232 -6650 -3168
rect -9022 -3248 -6650 -3232
rect -9022 -3312 -6734 -3248
rect -6670 -3312 -6650 -3248
rect -9022 -3360 -6650 -3312
rect -6410 -1328 -4038 -1280
rect -6410 -1392 -4122 -1328
rect -4058 -1392 -4038 -1328
rect -6410 -1408 -4038 -1392
rect -6410 -1472 -4122 -1408
rect -4058 -1472 -4038 -1408
rect -6410 -1488 -4038 -1472
rect -6410 -1552 -4122 -1488
rect -4058 -1552 -4038 -1488
rect -6410 -1568 -4038 -1552
rect -6410 -1632 -4122 -1568
rect -4058 -1632 -4038 -1568
rect -6410 -1648 -4038 -1632
rect -6410 -1712 -4122 -1648
rect -4058 -1712 -4038 -1648
rect -6410 -1728 -4038 -1712
rect -6410 -1792 -4122 -1728
rect -4058 -1792 -4038 -1728
rect -6410 -1808 -4038 -1792
rect -6410 -1872 -4122 -1808
rect -4058 -1872 -4038 -1808
rect -6410 -1888 -4038 -1872
rect -6410 -1952 -4122 -1888
rect -4058 -1952 -4038 -1888
rect -6410 -1968 -4038 -1952
rect -6410 -2032 -4122 -1968
rect -4058 -2032 -4038 -1968
rect -6410 -2048 -4038 -2032
rect -6410 -2112 -4122 -2048
rect -4058 -2112 -4038 -2048
rect -6410 -2128 -4038 -2112
rect -6410 -2192 -4122 -2128
rect -4058 -2192 -4038 -2128
rect -6410 -2208 -4038 -2192
rect -6410 -2272 -4122 -2208
rect -4058 -2272 -4038 -2208
rect -6410 -2288 -4038 -2272
rect -6410 -2352 -4122 -2288
rect -4058 -2352 -4038 -2288
rect -6410 -2368 -4038 -2352
rect -6410 -2432 -4122 -2368
rect -4058 -2432 -4038 -2368
rect -6410 -2448 -4038 -2432
rect -6410 -2512 -4122 -2448
rect -4058 -2512 -4038 -2448
rect -6410 -2528 -4038 -2512
rect -6410 -2592 -4122 -2528
rect -4058 -2592 -4038 -2528
rect -6410 -2608 -4038 -2592
rect -6410 -2672 -4122 -2608
rect -4058 -2672 -4038 -2608
rect -6410 -2688 -4038 -2672
rect -6410 -2752 -4122 -2688
rect -4058 -2752 -4038 -2688
rect -6410 -2768 -4038 -2752
rect -6410 -2832 -4122 -2768
rect -4058 -2832 -4038 -2768
rect -6410 -2848 -4038 -2832
rect -6410 -2912 -4122 -2848
rect -4058 -2912 -4038 -2848
rect -6410 -2928 -4038 -2912
rect -6410 -2992 -4122 -2928
rect -4058 -2992 -4038 -2928
rect -6410 -3008 -4038 -2992
rect -6410 -3072 -4122 -3008
rect -4058 -3072 -4038 -3008
rect -6410 -3088 -4038 -3072
rect -6410 -3152 -4122 -3088
rect -4058 -3152 -4038 -3088
rect -6410 -3168 -4038 -3152
rect -6410 -3232 -4122 -3168
rect -4058 -3232 -4038 -3168
rect -6410 -3248 -4038 -3232
rect -6410 -3312 -4122 -3248
rect -4058 -3312 -4038 -3248
rect -6410 -3360 -4038 -3312
rect -3798 -1328 -1426 -1280
rect -3798 -1392 -1510 -1328
rect -1446 -1392 -1426 -1328
rect -3798 -1408 -1426 -1392
rect -3798 -1472 -1510 -1408
rect -1446 -1472 -1426 -1408
rect -3798 -1488 -1426 -1472
rect -3798 -1552 -1510 -1488
rect -1446 -1552 -1426 -1488
rect -3798 -1568 -1426 -1552
rect -3798 -1632 -1510 -1568
rect -1446 -1632 -1426 -1568
rect -3798 -1648 -1426 -1632
rect -3798 -1712 -1510 -1648
rect -1446 -1712 -1426 -1648
rect -3798 -1728 -1426 -1712
rect -3798 -1792 -1510 -1728
rect -1446 -1792 -1426 -1728
rect -3798 -1808 -1426 -1792
rect -3798 -1872 -1510 -1808
rect -1446 -1872 -1426 -1808
rect -3798 -1888 -1426 -1872
rect -3798 -1952 -1510 -1888
rect -1446 -1952 -1426 -1888
rect -3798 -1968 -1426 -1952
rect -3798 -2032 -1510 -1968
rect -1446 -2032 -1426 -1968
rect -3798 -2048 -1426 -2032
rect -3798 -2112 -1510 -2048
rect -1446 -2112 -1426 -2048
rect -3798 -2128 -1426 -2112
rect -3798 -2192 -1510 -2128
rect -1446 -2192 -1426 -2128
rect -3798 -2208 -1426 -2192
rect -3798 -2272 -1510 -2208
rect -1446 -2272 -1426 -2208
rect -3798 -2288 -1426 -2272
rect -3798 -2352 -1510 -2288
rect -1446 -2352 -1426 -2288
rect -3798 -2368 -1426 -2352
rect -3798 -2432 -1510 -2368
rect -1446 -2432 -1426 -2368
rect -3798 -2448 -1426 -2432
rect -3798 -2512 -1510 -2448
rect -1446 -2512 -1426 -2448
rect -3798 -2528 -1426 -2512
rect -3798 -2592 -1510 -2528
rect -1446 -2592 -1426 -2528
rect -3798 -2608 -1426 -2592
rect -3798 -2672 -1510 -2608
rect -1446 -2672 -1426 -2608
rect -3798 -2688 -1426 -2672
rect -3798 -2752 -1510 -2688
rect -1446 -2752 -1426 -2688
rect -3798 -2768 -1426 -2752
rect -3798 -2832 -1510 -2768
rect -1446 -2832 -1426 -2768
rect -3798 -2848 -1426 -2832
rect -3798 -2912 -1510 -2848
rect -1446 -2912 -1426 -2848
rect -3798 -2928 -1426 -2912
rect -3798 -2992 -1510 -2928
rect -1446 -2992 -1426 -2928
rect -3798 -3008 -1426 -2992
rect -3798 -3072 -1510 -3008
rect -1446 -3072 -1426 -3008
rect -3798 -3088 -1426 -3072
rect -3798 -3152 -1510 -3088
rect -1446 -3152 -1426 -3088
rect -3798 -3168 -1426 -3152
rect -3798 -3232 -1510 -3168
rect -1446 -3232 -1426 -3168
rect -3798 -3248 -1426 -3232
rect -3798 -3312 -1510 -3248
rect -1446 -3312 -1426 -3248
rect -3798 -3360 -1426 -3312
rect -1186 -1328 1186 -1280
rect -1186 -1392 1102 -1328
rect 1166 -1392 1186 -1328
rect -1186 -1408 1186 -1392
rect -1186 -1472 1102 -1408
rect 1166 -1472 1186 -1408
rect -1186 -1488 1186 -1472
rect -1186 -1552 1102 -1488
rect 1166 -1552 1186 -1488
rect -1186 -1568 1186 -1552
rect -1186 -1632 1102 -1568
rect 1166 -1632 1186 -1568
rect -1186 -1648 1186 -1632
rect -1186 -1712 1102 -1648
rect 1166 -1712 1186 -1648
rect -1186 -1728 1186 -1712
rect -1186 -1792 1102 -1728
rect 1166 -1792 1186 -1728
rect -1186 -1808 1186 -1792
rect -1186 -1872 1102 -1808
rect 1166 -1872 1186 -1808
rect -1186 -1888 1186 -1872
rect -1186 -1952 1102 -1888
rect 1166 -1952 1186 -1888
rect -1186 -1968 1186 -1952
rect -1186 -2032 1102 -1968
rect 1166 -2032 1186 -1968
rect -1186 -2048 1186 -2032
rect -1186 -2112 1102 -2048
rect 1166 -2112 1186 -2048
rect -1186 -2128 1186 -2112
rect -1186 -2192 1102 -2128
rect 1166 -2192 1186 -2128
rect -1186 -2208 1186 -2192
rect -1186 -2272 1102 -2208
rect 1166 -2272 1186 -2208
rect -1186 -2288 1186 -2272
rect -1186 -2352 1102 -2288
rect 1166 -2352 1186 -2288
rect -1186 -2368 1186 -2352
rect -1186 -2432 1102 -2368
rect 1166 -2432 1186 -2368
rect -1186 -2448 1186 -2432
rect -1186 -2512 1102 -2448
rect 1166 -2512 1186 -2448
rect -1186 -2528 1186 -2512
rect -1186 -2592 1102 -2528
rect 1166 -2592 1186 -2528
rect -1186 -2608 1186 -2592
rect -1186 -2672 1102 -2608
rect 1166 -2672 1186 -2608
rect -1186 -2688 1186 -2672
rect -1186 -2752 1102 -2688
rect 1166 -2752 1186 -2688
rect -1186 -2768 1186 -2752
rect -1186 -2832 1102 -2768
rect 1166 -2832 1186 -2768
rect -1186 -2848 1186 -2832
rect -1186 -2912 1102 -2848
rect 1166 -2912 1186 -2848
rect -1186 -2928 1186 -2912
rect -1186 -2992 1102 -2928
rect 1166 -2992 1186 -2928
rect -1186 -3008 1186 -2992
rect -1186 -3072 1102 -3008
rect 1166 -3072 1186 -3008
rect -1186 -3088 1186 -3072
rect -1186 -3152 1102 -3088
rect 1166 -3152 1186 -3088
rect -1186 -3168 1186 -3152
rect -1186 -3232 1102 -3168
rect 1166 -3232 1186 -3168
rect -1186 -3248 1186 -3232
rect -1186 -3312 1102 -3248
rect 1166 -3312 1186 -3248
rect -1186 -3360 1186 -3312
rect 1426 -1328 3798 -1280
rect 1426 -1392 3714 -1328
rect 3778 -1392 3798 -1328
rect 1426 -1408 3798 -1392
rect 1426 -1472 3714 -1408
rect 3778 -1472 3798 -1408
rect 1426 -1488 3798 -1472
rect 1426 -1552 3714 -1488
rect 3778 -1552 3798 -1488
rect 1426 -1568 3798 -1552
rect 1426 -1632 3714 -1568
rect 3778 -1632 3798 -1568
rect 1426 -1648 3798 -1632
rect 1426 -1712 3714 -1648
rect 3778 -1712 3798 -1648
rect 1426 -1728 3798 -1712
rect 1426 -1792 3714 -1728
rect 3778 -1792 3798 -1728
rect 1426 -1808 3798 -1792
rect 1426 -1872 3714 -1808
rect 3778 -1872 3798 -1808
rect 1426 -1888 3798 -1872
rect 1426 -1952 3714 -1888
rect 3778 -1952 3798 -1888
rect 1426 -1968 3798 -1952
rect 1426 -2032 3714 -1968
rect 3778 -2032 3798 -1968
rect 1426 -2048 3798 -2032
rect 1426 -2112 3714 -2048
rect 3778 -2112 3798 -2048
rect 1426 -2128 3798 -2112
rect 1426 -2192 3714 -2128
rect 3778 -2192 3798 -2128
rect 1426 -2208 3798 -2192
rect 1426 -2272 3714 -2208
rect 3778 -2272 3798 -2208
rect 1426 -2288 3798 -2272
rect 1426 -2352 3714 -2288
rect 3778 -2352 3798 -2288
rect 1426 -2368 3798 -2352
rect 1426 -2432 3714 -2368
rect 3778 -2432 3798 -2368
rect 1426 -2448 3798 -2432
rect 1426 -2512 3714 -2448
rect 3778 -2512 3798 -2448
rect 1426 -2528 3798 -2512
rect 1426 -2592 3714 -2528
rect 3778 -2592 3798 -2528
rect 1426 -2608 3798 -2592
rect 1426 -2672 3714 -2608
rect 3778 -2672 3798 -2608
rect 1426 -2688 3798 -2672
rect 1426 -2752 3714 -2688
rect 3778 -2752 3798 -2688
rect 1426 -2768 3798 -2752
rect 1426 -2832 3714 -2768
rect 3778 -2832 3798 -2768
rect 1426 -2848 3798 -2832
rect 1426 -2912 3714 -2848
rect 3778 -2912 3798 -2848
rect 1426 -2928 3798 -2912
rect 1426 -2992 3714 -2928
rect 3778 -2992 3798 -2928
rect 1426 -3008 3798 -2992
rect 1426 -3072 3714 -3008
rect 3778 -3072 3798 -3008
rect 1426 -3088 3798 -3072
rect 1426 -3152 3714 -3088
rect 3778 -3152 3798 -3088
rect 1426 -3168 3798 -3152
rect 1426 -3232 3714 -3168
rect 3778 -3232 3798 -3168
rect 1426 -3248 3798 -3232
rect 1426 -3312 3714 -3248
rect 3778 -3312 3798 -3248
rect 1426 -3360 3798 -3312
rect 4038 -1328 6410 -1280
rect 4038 -1392 6326 -1328
rect 6390 -1392 6410 -1328
rect 4038 -1408 6410 -1392
rect 4038 -1472 6326 -1408
rect 6390 -1472 6410 -1408
rect 4038 -1488 6410 -1472
rect 4038 -1552 6326 -1488
rect 6390 -1552 6410 -1488
rect 4038 -1568 6410 -1552
rect 4038 -1632 6326 -1568
rect 6390 -1632 6410 -1568
rect 4038 -1648 6410 -1632
rect 4038 -1712 6326 -1648
rect 6390 -1712 6410 -1648
rect 4038 -1728 6410 -1712
rect 4038 -1792 6326 -1728
rect 6390 -1792 6410 -1728
rect 4038 -1808 6410 -1792
rect 4038 -1872 6326 -1808
rect 6390 -1872 6410 -1808
rect 4038 -1888 6410 -1872
rect 4038 -1952 6326 -1888
rect 6390 -1952 6410 -1888
rect 4038 -1968 6410 -1952
rect 4038 -2032 6326 -1968
rect 6390 -2032 6410 -1968
rect 4038 -2048 6410 -2032
rect 4038 -2112 6326 -2048
rect 6390 -2112 6410 -2048
rect 4038 -2128 6410 -2112
rect 4038 -2192 6326 -2128
rect 6390 -2192 6410 -2128
rect 4038 -2208 6410 -2192
rect 4038 -2272 6326 -2208
rect 6390 -2272 6410 -2208
rect 4038 -2288 6410 -2272
rect 4038 -2352 6326 -2288
rect 6390 -2352 6410 -2288
rect 4038 -2368 6410 -2352
rect 4038 -2432 6326 -2368
rect 6390 -2432 6410 -2368
rect 4038 -2448 6410 -2432
rect 4038 -2512 6326 -2448
rect 6390 -2512 6410 -2448
rect 4038 -2528 6410 -2512
rect 4038 -2592 6326 -2528
rect 6390 -2592 6410 -2528
rect 4038 -2608 6410 -2592
rect 4038 -2672 6326 -2608
rect 6390 -2672 6410 -2608
rect 4038 -2688 6410 -2672
rect 4038 -2752 6326 -2688
rect 6390 -2752 6410 -2688
rect 4038 -2768 6410 -2752
rect 4038 -2832 6326 -2768
rect 6390 -2832 6410 -2768
rect 4038 -2848 6410 -2832
rect 4038 -2912 6326 -2848
rect 6390 -2912 6410 -2848
rect 4038 -2928 6410 -2912
rect 4038 -2992 6326 -2928
rect 6390 -2992 6410 -2928
rect 4038 -3008 6410 -2992
rect 4038 -3072 6326 -3008
rect 6390 -3072 6410 -3008
rect 4038 -3088 6410 -3072
rect 4038 -3152 6326 -3088
rect 6390 -3152 6410 -3088
rect 4038 -3168 6410 -3152
rect 4038 -3232 6326 -3168
rect 6390 -3232 6410 -3168
rect 4038 -3248 6410 -3232
rect 4038 -3312 6326 -3248
rect 6390 -3312 6410 -3248
rect 4038 -3360 6410 -3312
rect 6650 -1328 9022 -1280
rect 6650 -1392 8938 -1328
rect 9002 -1392 9022 -1328
rect 6650 -1408 9022 -1392
rect 6650 -1472 8938 -1408
rect 9002 -1472 9022 -1408
rect 6650 -1488 9022 -1472
rect 6650 -1552 8938 -1488
rect 9002 -1552 9022 -1488
rect 6650 -1568 9022 -1552
rect 6650 -1632 8938 -1568
rect 9002 -1632 9022 -1568
rect 6650 -1648 9022 -1632
rect 6650 -1712 8938 -1648
rect 9002 -1712 9022 -1648
rect 6650 -1728 9022 -1712
rect 6650 -1792 8938 -1728
rect 9002 -1792 9022 -1728
rect 6650 -1808 9022 -1792
rect 6650 -1872 8938 -1808
rect 9002 -1872 9022 -1808
rect 6650 -1888 9022 -1872
rect 6650 -1952 8938 -1888
rect 9002 -1952 9022 -1888
rect 6650 -1968 9022 -1952
rect 6650 -2032 8938 -1968
rect 9002 -2032 9022 -1968
rect 6650 -2048 9022 -2032
rect 6650 -2112 8938 -2048
rect 9002 -2112 9022 -2048
rect 6650 -2128 9022 -2112
rect 6650 -2192 8938 -2128
rect 9002 -2192 9022 -2128
rect 6650 -2208 9022 -2192
rect 6650 -2272 8938 -2208
rect 9002 -2272 9022 -2208
rect 6650 -2288 9022 -2272
rect 6650 -2352 8938 -2288
rect 9002 -2352 9022 -2288
rect 6650 -2368 9022 -2352
rect 6650 -2432 8938 -2368
rect 9002 -2432 9022 -2368
rect 6650 -2448 9022 -2432
rect 6650 -2512 8938 -2448
rect 9002 -2512 9022 -2448
rect 6650 -2528 9022 -2512
rect 6650 -2592 8938 -2528
rect 9002 -2592 9022 -2528
rect 6650 -2608 9022 -2592
rect 6650 -2672 8938 -2608
rect 9002 -2672 9022 -2608
rect 6650 -2688 9022 -2672
rect 6650 -2752 8938 -2688
rect 9002 -2752 9022 -2688
rect 6650 -2768 9022 -2752
rect 6650 -2832 8938 -2768
rect 9002 -2832 9022 -2768
rect 6650 -2848 9022 -2832
rect 6650 -2912 8938 -2848
rect 9002 -2912 9022 -2848
rect 6650 -2928 9022 -2912
rect 6650 -2992 8938 -2928
rect 9002 -2992 9022 -2928
rect 6650 -3008 9022 -2992
rect 6650 -3072 8938 -3008
rect 9002 -3072 9022 -3008
rect 6650 -3088 9022 -3072
rect 6650 -3152 8938 -3088
rect 9002 -3152 9022 -3088
rect 6650 -3168 9022 -3152
rect 6650 -3232 8938 -3168
rect 9002 -3232 9022 -3168
rect 6650 -3248 9022 -3232
rect 6650 -3312 8938 -3248
rect 9002 -3312 9022 -3248
rect 6650 -3360 9022 -3312
rect -9022 -3648 -6650 -3600
rect -9022 -3712 -6734 -3648
rect -6670 -3712 -6650 -3648
rect -9022 -3728 -6650 -3712
rect -9022 -3792 -6734 -3728
rect -6670 -3792 -6650 -3728
rect -9022 -3808 -6650 -3792
rect -9022 -3872 -6734 -3808
rect -6670 -3872 -6650 -3808
rect -9022 -3888 -6650 -3872
rect -9022 -3952 -6734 -3888
rect -6670 -3952 -6650 -3888
rect -9022 -3968 -6650 -3952
rect -9022 -4032 -6734 -3968
rect -6670 -4032 -6650 -3968
rect -9022 -4048 -6650 -4032
rect -9022 -4112 -6734 -4048
rect -6670 -4112 -6650 -4048
rect -9022 -4128 -6650 -4112
rect -9022 -4192 -6734 -4128
rect -6670 -4192 -6650 -4128
rect -9022 -4208 -6650 -4192
rect -9022 -4272 -6734 -4208
rect -6670 -4272 -6650 -4208
rect -9022 -4288 -6650 -4272
rect -9022 -4352 -6734 -4288
rect -6670 -4352 -6650 -4288
rect -9022 -4368 -6650 -4352
rect -9022 -4432 -6734 -4368
rect -6670 -4432 -6650 -4368
rect -9022 -4448 -6650 -4432
rect -9022 -4512 -6734 -4448
rect -6670 -4512 -6650 -4448
rect -9022 -4528 -6650 -4512
rect -9022 -4592 -6734 -4528
rect -6670 -4592 -6650 -4528
rect -9022 -4608 -6650 -4592
rect -9022 -4672 -6734 -4608
rect -6670 -4672 -6650 -4608
rect -9022 -4688 -6650 -4672
rect -9022 -4752 -6734 -4688
rect -6670 -4752 -6650 -4688
rect -9022 -4768 -6650 -4752
rect -9022 -4832 -6734 -4768
rect -6670 -4832 -6650 -4768
rect -9022 -4848 -6650 -4832
rect -9022 -4912 -6734 -4848
rect -6670 -4912 -6650 -4848
rect -9022 -4928 -6650 -4912
rect -9022 -4992 -6734 -4928
rect -6670 -4992 -6650 -4928
rect -9022 -5008 -6650 -4992
rect -9022 -5072 -6734 -5008
rect -6670 -5072 -6650 -5008
rect -9022 -5088 -6650 -5072
rect -9022 -5152 -6734 -5088
rect -6670 -5152 -6650 -5088
rect -9022 -5168 -6650 -5152
rect -9022 -5232 -6734 -5168
rect -6670 -5232 -6650 -5168
rect -9022 -5248 -6650 -5232
rect -9022 -5312 -6734 -5248
rect -6670 -5312 -6650 -5248
rect -9022 -5328 -6650 -5312
rect -9022 -5392 -6734 -5328
rect -6670 -5392 -6650 -5328
rect -9022 -5408 -6650 -5392
rect -9022 -5472 -6734 -5408
rect -6670 -5472 -6650 -5408
rect -9022 -5488 -6650 -5472
rect -9022 -5552 -6734 -5488
rect -6670 -5552 -6650 -5488
rect -9022 -5568 -6650 -5552
rect -9022 -5632 -6734 -5568
rect -6670 -5632 -6650 -5568
rect -9022 -5680 -6650 -5632
rect -6410 -3648 -4038 -3600
rect -6410 -3712 -4122 -3648
rect -4058 -3712 -4038 -3648
rect -6410 -3728 -4038 -3712
rect -6410 -3792 -4122 -3728
rect -4058 -3792 -4038 -3728
rect -6410 -3808 -4038 -3792
rect -6410 -3872 -4122 -3808
rect -4058 -3872 -4038 -3808
rect -6410 -3888 -4038 -3872
rect -6410 -3952 -4122 -3888
rect -4058 -3952 -4038 -3888
rect -6410 -3968 -4038 -3952
rect -6410 -4032 -4122 -3968
rect -4058 -4032 -4038 -3968
rect -6410 -4048 -4038 -4032
rect -6410 -4112 -4122 -4048
rect -4058 -4112 -4038 -4048
rect -6410 -4128 -4038 -4112
rect -6410 -4192 -4122 -4128
rect -4058 -4192 -4038 -4128
rect -6410 -4208 -4038 -4192
rect -6410 -4272 -4122 -4208
rect -4058 -4272 -4038 -4208
rect -6410 -4288 -4038 -4272
rect -6410 -4352 -4122 -4288
rect -4058 -4352 -4038 -4288
rect -6410 -4368 -4038 -4352
rect -6410 -4432 -4122 -4368
rect -4058 -4432 -4038 -4368
rect -6410 -4448 -4038 -4432
rect -6410 -4512 -4122 -4448
rect -4058 -4512 -4038 -4448
rect -6410 -4528 -4038 -4512
rect -6410 -4592 -4122 -4528
rect -4058 -4592 -4038 -4528
rect -6410 -4608 -4038 -4592
rect -6410 -4672 -4122 -4608
rect -4058 -4672 -4038 -4608
rect -6410 -4688 -4038 -4672
rect -6410 -4752 -4122 -4688
rect -4058 -4752 -4038 -4688
rect -6410 -4768 -4038 -4752
rect -6410 -4832 -4122 -4768
rect -4058 -4832 -4038 -4768
rect -6410 -4848 -4038 -4832
rect -6410 -4912 -4122 -4848
rect -4058 -4912 -4038 -4848
rect -6410 -4928 -4038 -4912
rect -6410 -4992 -4122 -4928
rect -4058 -4992 -4038 -4928
rect -6410 -5008 -4038 -4992
rect -6410 -5072 -4122 -5008
rect -4058 -5072 -4038 -5008
rect -6410 -5088 -4038 -5072
rect -6410 -5152 -4122 -5088
rect -4058 -5152 -4038 -5088
rect -6410 -5168 -4038 -5152
rect -6410 -5232 -4122 -5168
rect -4058 -5232 -4038 -5168
rect -6410 -5248 -4038 -5232
rect -6410 -5312 -4122 -5248
rect -4058 -5312 -4038 -5248
rect -6410 -5328 -4038 -5312
rect -6410 -5392 -4122 -5328
rect -4058 -5392 -4038 -5328
rect -6410 -5408 -4038 -5392
rect -6410 -5472 -4122 -5408
rect -4058 -5472 -4038 -5408
rect -6410 -5488 -4038 -5472
rect -6410 -5552 -4122 -5488
rect -4058 -5552 -4038 -5488
rect -6410 -5568 -4038 -5552
rect -6410 -5632 -4122 -5568
rect -4058 -5632 -4038 -5568
rect -6410 -5680 -4038 -5632
rect -3798 -3648 -1426 -3600
rect -3798 -3712 -1510 -3648
rect -1446 -3712 -1426 -3648
rect -3798 -3728 -1426 -3712
rect -3798 -3792 -1510 -3728
rect -1446 -3792 -1426 -3728
rect -3798 -3808 -1426 -3792
rect -3798 -3872 -1510 -3808
rect -1446 -3872 -1426 -3808
rect -3798 -3888 -1426 -3872
rect -3798 -3952 -1510 -3888
rect -1446 -3952 -1426 -3888
rect -3798 -3968 -1426 -3952
rect -3798 -4032 -1510 -3968
rect -1446 -4032 -1426 -3968
rect -3798 -4048 -1426 -4032
rect -3798 -4112 -1510 -4048
rect -1446 -4112 -1426 -4048
rect -3798 -4128 -1426 -4112
rect -3798 -4192 -1510 -4128
rect -1446 -4192 -1426 -4128
rect -3798 -4208 -1426 -4192
rect -3798 -4272 -1510 -4208
rect -1446 -4272 -1426 -4208
rect -3798 -4288 -1426 -4272
rect -3798 -4352 -1510 -4288
rect -1446 -4352 -1426 -4288
rect -3798 -4368 -1426 -4352
rect -3798 -4432 -1510 -4368
rect -1446 -4432 -1426 -4368
rect -3798 -4448 -1426 -4432
rect -3798 -4512 -1510 -4448
rect -1446 -4512 -1426 -4448
rect -3798 -4528 -1426 -4512
rect -3798 -4592 -1510 -4528
rect -1446 -4592 -1426 -4528
rect -3798 -4608 -1426 -4592
rect -3798 -4672 -1510 -4608
rect -1446 -4672 -1426 -4608
rect -3798 -4688 -1426 -4672
rect -3798 -4752 -1510 -4688
rect -1446 -4752 -1426 -4688
rect -3798 -4768 -1426 -4752
rect -3798 -4832 -1510 -4768
rect -1446 -4832 -1426 -4768
rect -3798 -4848 -1426 -4832
rect -3798 -4912 -1510 -4848
rect -1446 -4912 -1426 -4848
rect -3798 -4928 -1426 -4912
rect -3798 -4992 -1510 -4928
rect -1446 -4992 -1426 -4928
rect -3798 -5008 -1426 -4992
rect -3798 -5072 -1510 -5008
rect -1446 -5072 -1426 -5008
rect -3798 -5088 -1426 -5072
rect -3798 -5152 -1510 -5088
rect -1446 -5152 -1426 -5088
rect -3798 -5168 -1426 -5152
rect -3798 -5232 -1510 -5168
rect -1446 -5232 -1426 -5168
rect -3798 -5248 -1426 -5232
rect -3798 -5312 -1510 -5248
rect -1446 -5312 -1426 -5248
rect -3798 -5328 -1426 -5312
rect -3798 -5392 -1510 -5328
rect -1446 -5392 -1426 -5328
rect -3798 -5408 -1426 -5392
rect -3798 -5472 -1510 -5408
rect -1446 -5472 -1426 -5408
rect -3798 -5488 -1426 -5472
rect -3798 -5552 -1510 -5488
rect -1446 -5552 -1426 -5488
rect -3798 -5568 -1426 -5552
rect -3798 -5632 -1510 -5568
rect -1446 -5632 -1426 -5568
rect -3798 -5680 -1426 -5632
rect -1186 -3648 1186 -3600
rect -1186 -3712 1102 -3648
rect 1166 -3712 1186 -3648
rect -1186 -3728 1186 -3712
rect -1186 -3792 1102 -3728
rect 1166 -3792 1186 -3728
rect -1186 -3808 1186 -3792
rect -1186 -3872 1102 -3808
rect 1166 -3872 1186 -3808
rect -1186 -3888 1186 -3872
rect -1186 -3952 1102 -3888
rect 1166 -3952 1186 -3888
rect -1186 -3968 1186 -3952
rect -1186 -4032 1102 -3968
rect 1166 -4032 1186 -3968
rect -1186 -4048 1186 -4032
rect -1186 -4112 1102 -4048
rect 1166 -4112 1186 -4048
rect -1186 -4128 1186 -4112
rect -1186 -4192 1102 -4128
rect 1166 -4192 1186 -4128
rect -1186 -4208 1186 -4192
rect -1186 -4272 1102 -4208
rect 1166 -4272 1186 -4208
rect -1186 -4288 1186 -4272
rect -1186 -4352 1102 -4288
rect 1166 -4352 1186 -4288
rect -1186 -4368 1186 -4352
rect -1186 -4432 1102 -4368
rect 1166 -4432 1186 -4368
rect -1186 -4448 1186 -4432
rect -1186 -4512 1102 -4448
rect 1166 -4512 1186 -4448
rect -1186 -4528 1186 -4512
rect -1186 -4592 1102 -4528
rect 1166 -4592 1186 -4528
rect -1186 -4608 1186 -4592
rect -1186 -4672 1102 -4608
rect 1166 -4672 1186 -4608
rect -1186 -4688 1186 -4672
rect -1186 -4752 1102 -4688
rect 1166 -4752 1186 -4688
rect -1186 -4768 1186 -4752
rect -1186 -4832 1102 -4768
rect 1166 -4832 1186 -4768
rect -1186 -4848 1186 -4832
rect -1186 -4912 1102 -4848
rect 1166 -4912 1186 -4848
rect -1186 -4928 1186 -4912
rect -1186 -4992 1102 -4928
rect 1166 -4992 1186 -4928
rect -1186 -5008 1186 -4992
rect -1186 -5072 1102 -5008
rect 1166 -5072 1186 -5008
rect -1186 -5088 1186 -5072
rect -1186 -5152 1102 -5088
rect 1166 -5152 1186 -5088
rect -1186 -5168 1186 -5152
rect -1186 -5232 1102 -5168
rect 1166 -5232 1186 -5168
rect -1186 -5248 1186 -5232
rect -1186 -5312 1102 -5248
rect 1166 -5312 1186 -5248
rect -1186 -5328 1186 -5312
rect -1186 -5392 1102 -5328
rect 1166 -5392 1186 -5328
rect -1186 -5408 1186 -5392
rect -1186 -5472 1102 -5408
rect 1166 -5472 1186 -5408
rect -1186 -5488 1186 -5472
rect -1186 -5552 1102 -5488
rect 1166 -5552 1186 -5488
rect -1186 -5568 1186 -5552
rect -1186 -5632 1102 -5568
rect 1166 -5632 1186 -5568
rect -1186 -5680 1186 -5632
rect 1426 -3648 3798 -3600
rect 1426 -3712 3714 -3648
rect 3778 -3712 3798 -3648
rect 1426 -3728 3798 -3712
rect 1426 -3792 3714 -3728
rect 3778 -3792 3798 -3728
rect 1426 -3808 3798 -3792
rect 1426 -3872 3714 -3808
rect 3778 -3872 3798 -3808
rect 1426 -3888 3798 -3872
rect 1426 -3952 3714 -3888
rect 3778 -3952 3798 -3888
rect 1426 -3968 3798 -3952
rect 1426 -4032 3714 -3968
rect 3778 -4032 3798 -3968
rect 1426 -4048 3798 -4032
rect 1426 -4112 3714 -4048
rect 3778 -4112 3798 -4048
rect 1426 -4128 3798 -4112
rect 1426 -4192 3714 -4128
rect 3778 -4192 3798 -4128
rect 1426 -4208 3798 -4192
rect 1426 -4272 3714 -4208
rect 3778 -4272 3798 -4208
rect 1426 -4288 3798 -4272
rect 1426 -4352 3714 -4288
rect 3778 -4352 3798 -4288
rect 1426 -4368 3798 -4352
rect 1426 -4432 3714 -4368
rect 3778 -4432 3798 -4368
rect 1426 -4448 3798 -4432
rect 1426 -4512 3714 -4448
rect 3778 -4512 3798 -4448
rect 1426 -4528 3798 -4512
rect 1426 -4592 3714 -4528
rect 3778 -4592 3798 -4528
rect 1426 -4608 3798 -4592
rect 1426 -4672 3714 -4608
rect 3778 -4672 3798 -4608
rect 1426 -4688 3798 -4672
rect 1426 -4752 3714 -4688
rect 3778 -4752 3798 -4688
rect 1426 -4768 3798 -4752
rect 1426 -4832 3714 -4768
rect 3778 -4832 3798 -4768
rect 1426 -4848 3798 -4832
rect 1426 -4912 3714 -4848
rect 3778 -4912 3798 -4848
rect 1426 -4928 3798 -4912
rect 1426 -4992 3714 -4928
rect 3778 -4992 3798 -4928
rect 1426 -5008 3798 -4992
rect 1426 -5072 3714 -5008
rect 3778 -5072 3798 -5008
rect 1426 -5088 3798 -5072
rect 1426 -5152 3714 -5088
rect 3778 -5152 3798 -5088
rect 1426 -5168 3798 -5152
rect 1426 -5232 3714 -5168
rect 3778 -5232 3798 -5168
rect 1426 -5248 3798 -5232
rect 1426 -5312 3714 -5248
rect 3778 -5312 3798 -5248
rect 1426 -5328 3798 -5312
rect 1426 -5392 3714 -5328
rect 3778 -5392 3798 -5328
rect 1426 -5408 3798 -5392
rect 1426 -5472 3714 -5408
rect 3778 -5472 3798 -5408
rect 1426 -5488 3798 -5472
rect 1426 -5552 3714 -5488
rect 3778 -5552 3798 -5488
rect 1426 -5568 3798 -5552
rect 1426 -5632 3714 -5568
rect 3778 -5632 3798 -5568
rect 1426 -5680 3798 -5632
rect 4038 -3648 6410 -3600
rect 4038 -3712 6326 -3648
rect 6390 -3712 6410 -3648
rect 4038 -3728 6410 -3712
rect 4038 -3792 6326 -3728
rect 6390 -3792 6410 -3728
rect 4038 -3808 6410 -3792
rect 4038 -3872 6326 -3808
rect 6390 -3872 6410 -3808
rect 4038 -3888 6410 -3872
rect 4038 -3952 6326 -3888
rect 6390 -3952 6410 -3888
rect 4038 -3968 6410 -3952
rect 4038 -4032 6326 -3968
rect 6390 -4032 6410 -3968
rect 4038 -4048 6410 -4032
rect 4038 -4112 6326 -4048
rect 6390 -4112 6410 -4048
rect 4038 -4128 6410 -4112
rect 4038 -4192 6326 -4128
rect 6390 -4192 6410 -4128
rect 4038 -4208 6410 -4192
rect 4038 -4272 6326 -4208
rect 6390 -4272 6410 -4208
rect 4038 -4288 6410 -4272
rect 4038 -4352 6326 -4288
rect 6390 -4352 6410 -4288
rect 4038 -4368 6410 -4352
rect 4038 -4432 6326 -4368
rect 6390 -4432 6410 -4368
rect 4038 -4448 6410 -4432
rect 4038 -4512 6326 -4448
rect 6390 -4512 6410 -4448
rect 4038 -4528 6410 -4512
rect 4038 -4592 6326 -4528
rect 6390 -4592 6410 -4528
rect 4038 -4608 6410 -4592
rect 4038 -4672 6326 -4608
rect 6390 -4672 6410 -4608
rect 4038 -4688 6410 -4672
rect 4038 -4752 6326 -4688
rect 6390 -4752 6410 -4688
rect 4038 -4768 6410 -4752
rect 4038 -4832 6326 -4768
rect 6390 -4832 6410 -4768
rect 4038 -4848 6410 -4832
rect 4038 -4912 6326 -4848
rect 6390 -4912 6410 -4848
rect 4038 -4928 6410 -4912
rect 4038 -4992 6326 -4928
rect 6390 -4992 6410 -4928
rect 4038 -5008 6410 -4992
rect 4038 -5072 6326 -5008
rect 6390 -5072 6410 -5008
rect 4038 -5088 6410 -5072
rect 4038 -5152 6326 -5088
rect 6390 -5152 6410 -5088
rect 4038 -5168 6410 -5152
rect 4038 -5232 6326 -5168
rect 6390 -5232 6410 -5168
rect 4038 -5248 6410 -5232
rect 4038 -5312 6326 -5248
rect 6390 -5312 6410 -5248
rect 4038 -5328 6410 -5312
rect 4038 -5392 6326 -5328
rect 6390 -5392 6410 -5328
rect 4038 -5408 6410 -5392
rect 4038 -5472 6326 -5408
rect 6390 -5472 6410 -5408
rect 4038 -5488 6410 -5472
rect 4038 -5552 6326 -5488
rect 6390 -5552 6410 -5488
rect 4038 -5568 6410 -5552
rect 4038 -5632 6326 -5568
rect 6390 -5632 6410 -5568
rect 4038 -5680 6410 -5632
rect 6650 -3648 9022 -3600
rect 6650 -3712 8938 -3648
rect 9002 -3712 9022 -3648
rect 6650 -3728 9022 -3712
rect 6650 -3792 8938 -3728
rect 9002 -3792 9022 -3728
rect 6650 -3808 9022 -3792
rect 6650 -3872 8938 -3808
rect 9002 -3872 9022 -3808
rect 6650 -3888 9022 -3872
rect 6650 -3952 8938 -3888
rect 9002 -3952 9022 -3888
rect 6650 -3968 9022 -3952
rect 6650 -4032 8938 -3968
rect 9002 -4032 9022 -3968
rect 6650 -4048 9022 -4032
rect 6650 -4112 8938 -4048
rect 9002 -4112 9022 -4048
rect 6650 -4128 9022 -4112
rect 6650 -4192 8938 -4128
rect 9002 -4192 9022 -4128
rect 6650 -4208 9022 -4192
rect 6650 -4272 8938 -4208
rect 9002 -4272 9022 -4208
rect 6650 -4288 9022 -4272
rect 6650 -4352 8938 -4288
rect 9002 -4352 9022 -4288
rect 6650 -4368 9022 -4352
rect 6650 -4432 8938 -4368
rect 9002 -4432 9022 -4368
rect 6650 -4448 9022 -4432
rect 6650 -4512 8938 -4448
rect 9002 -4512 9022 -4448
rect 6650 -4528 9022 -4512
rect 6650 -4592 8938 -4528
rect 9002 -4592 9022 -4528
rect 6650 -4608 9022 -4592
rect 6650 -4672 8938 -4608
rect 9002 -4672 9022 -4608
rect 6650 -4688 9022 -4672
rect 6650 -4752 8938 -4688
rect 9002 -4752 9022 -4688
rect 6650 -4768 9022 -4752
rect 6650 -4832 8938 -4768
rect 9002 -4832 9022 -4768
rect 6650 -4848 9022 -4832
rect 6650 -4912 8938 -4848
rect 9002 -4912 9022 -4848
rect 6650 -4928 9022 -4912
rect 6650 -4992 8938 -4928
rect 9002 -4992 9022 -4928
rect 6650 -5008 9022 -4992
rect 6650 -5072 8938 -5008
rect 9002 -5072 9022 -5008
rect 6650 -5088 9022 -5072
rect 6650 -5152 8938 -5088
rect 9002 -5152 9022 -5088
rect 6650 -5168 9022 -5152
rect 6650 -5232 8938 -5168
rect 9002 -5232 9022 -5168
rect 6650 -5248 9022 -5232
rect 6650 -5312 8938 -5248
rect 9002 -5312 9022 -5248
rect 6650 -5328 9022 -5312
rect 6650 -5392 8938 -5328
rect 9002 -5392 9022 -5328
rect 6650 -5408 9022 -5392
rect 6650 -5472 8938 -5408
rect 9002 -5472 9022 -5408
rect 6650 -5488 9022 -5472
rect 6650 -5552 8938 -5488
rect 9002 -5552 9022 -5488
rect 6650 -5568 9022 -5552
rect 6650 -5632 8938 -5568
rect 9002 -5632 9022 -5568
rect 6650 -5680 9022 -5632
rect -9022 -5968 -6650 -5920
rect -9022 -6032 -6734 -5968
rect -6670 -6032 -6650 -5968
rect -9022 -6048 -6650 -6032
rect -9022 -6112 -6734 -6048
rect -6670 -6112 -6650 -6048
rect -9022 -6128 -6650 -6112
rect -9022 -6192 -6734 -6128
rect -6670 -6192 -6650 -6128
rect -9022 -6208 -6650 -6192
rect -9022 -6272 -6734 -6208
rect -6670 -6272 -6650 -6208
rect -9022 -6288 -6650 -6272
rect -9022 -6352 -6734 -6288
rect -6670 -6352 -6650 -6288
rect -9022 -6368 -6650 -6352
rect -9022 -6432 -6734 -6368
rect -6670 -6432 -6650 -6368
rect -9022 -6448 -6650 -6432
rect -9022 -6512 -6734 -6448
rect -6670 -6512 -6650 -6448
rect -9022 -6528 -6650 -6512
rect -9022 -6592 -6734 -6528
rect -6670 -6592 -6650 -6528
rect -9022 -6608 -6650 -6592
rect -9022 -6672 -6734 -6608
rect -6670 -6672 -6650 -6608
rect -9022 -6688 -6650 -6672
rect -9022 -6752 -6734 -6688
rect -6670 -6752 -6650 -6688
rect -9022 -6768 -6650 -6752
rect -9022 -6832 -6734 -6768
rect -6670 -6832 -6650 -6768
rect -9022 -6848 -6650 -6832
rect -9022 -6912 -6734 -6848
rect -6670 -6912 -6650 -6848
rect -9022 -6928 -6650 -6912
rect -9022 -6992 -6734 -6928
rect -6670 -6992 -6650 -6928
rect -9022 -7008 -6650 -6992
rect -9022 -7072 -6734 -7008
rect -6670 -7072 -6650 -7008
rect -9022 -7088 -6650 -7072
rect -9022 -7152 -6734 -7088
rect -6670 -7152 -6650 -7088
rect -9022 -7168 -6650 -7152
rect -9022 -7232 -6734 -7168
rect -6670 -7232 -6650 -7168
rect -9022 -7248 -6650 -7232
rect -9022 -7312 -6734 -7248
rect -6670 -7312 -6650 -7248
rect -9022 -7328 -6650 -7312
rect -9022 -7392 -6734 -7328
rect -6670 -7392 -6650 -7328
rect -9022 -7408 -6650 -7392
rect -9022 -7472 -6734 -7408
rect -6670 -7472 -6650 -7408
rect -9022 -7488 -6650 -7472
rect -9022 -7552 -6734 -7488
rect -6670 -7552 -6650 -7488
rect -9022 -7568 -6650 -7552
rect -9022 -7632 -6734 -7568
rect -6670 -7632 -6650 -7568
rect -9022 -7648 -6650 -7632
rect -9022 -7712 -6734 -7648
rect -6670 -7712 -6650 -7648
rect -9022 -7728 -6650 -7712
rect -9022 -7792 -6734 -7728
rect -6670 -7792 -6650 -7728
rect -9022 -7808 -6650 -7792
rect -9022 -7872 -6734 -7808
rect -6670 -7872 -6650 -7808
rect -9022 -7888 -6650 -7872
rect -9022 -7952 -6734 -7888
rect -6670 -7952 -6650 -7888
rect -9022 -8000 -6650 -7952
rect -6410 -5968 -4038 -5920
rect -6410 -6032 -4122 -5968
rect -4058 -6032 -4038 -5968
rect -6410 -6048 -4038 -6032
rect -6410 -6112 -4122 -6048
rect -4058 -6112 -4038 -6048
rect -6410 -6128 -4038 -6112
rect -6410 -6192 -4122 -6128
rect -4058 -6192 -4038 -6128
rect -6410 -6208 -4038 -6192
rect -6410 -6272 -4122 -6208
rect -4058 -6272 -4038 -6208
rect -6410 -6288 -4038 -6272
rect -6410 -6352 -4122 -6288
rect -4058 -6352 -4038 -6288
rect -6410 -6368 -4038 -6352
rect -6410 -6432 -4122 -6368
rect -4058 -6432 -4038 -6368
rect -6410 -6448 -4038 -6432
rect -6410 -6512 -4122 -6448
rect -4058 -6512 -4038 -6448
rect -6410 -6528 -4038 -6512
rect -6410 -6592 -4122 -6528
rect -4058 -6592 -4038 -6528
rect -6410 -6608 -4038 -6592
rect -6410 -6672 -4122 -6608
rect -4058 -6672 -4038 -6608
rect -6410 -6688 -4038 -6672
rect -6410 -6752 -4122 -6688
rect -4058 -6752 -4038 -6688
rect -6410 -6768 -4038 -6752
rect -6410 -6832 -4122 -6768
rect -4058 -6832 -4038 -6768
rect -6410 -6848 -4038 -6832
rect -6410 -6912 -4122 -6848
rect -4058 -6912 -4038 -6848
rect -6410 -6928 -4038 -6912
rect -6410 -6992 -4122 -6928
rect -4058 -6992 -4038 -6928
rect -6410 -7008 -4038 -6992
rect -6410 -7072 -4122 -7008
rect -4058 -7072 -4038 -7008
rect -6410 -7088 -4038 -7072
rect -6410 -7152 -4122 -7088
rect -4058 -7152 -4038 -7088
rect -6410 -7168 -4038 -7152
rect -6410 -7232 -4122 -7168
rect -4058 -7232 -4038 -7168
rect -6410 -7248 -4038 -7232
rect -6410 -7312 -4122 -7248
rect -4058 -7312 -4038 -7248
rect -6410 -7328 -4038 -7312
rect -6410 -7392 -4122 -7328
rect -4058 -7392 -4038 -7328
rect -6410 -7408 -4038 -7392
rect -6410 -7472 -4122 -7408
rect -4058 -7472 -4038 -7408
rect -6410 -7488 -4038 -7472
rect -6410 -7552 -4122 -7488
rect -4058 -7552 -4038 -7488
rect -6410 -7568 -4038 -7552
rect -6410 -7632 -4122 -7568
rect -4058 -7632 -4038 -7568
rect -6410 -7648 -4038 -7632
rect -6410 -7712 -4122 -7648
rect -4058 -7712 -4038 -7648
rect -6410 -7728 -4038 -7712
rect -6410 -7792 -4122 -7728
rect -4058 -7792 -4038 -7728
rect -6410 -7808 -4038 -7792
rect -6410 -7872 -4122 -7808
rect -4058 -7872 -4038 -7808
rect -6410 -7888 -4038 -7872
rect -6410 -7952 -4122 -7888
rect -4058 -7952 -4038 -7888
rect -6410 -8000 -4038 -7952
rect -3798 -5968 -1426 -5920
rect -3798 -6032 -1510 -5968
rect -1446 -6032 -1426 -5968
rect -3798 -6048 -1426 -6032
rect -3798 -6112 -1510 -6048
rect -1446 -6112 -1426 -6048
rect -3798 -6128 -1426 -6112
rect -3798 -6192 -1510 -6128
rect -1446 -6192 -1426 -6128
rect -3798 -6208 -1426 -6192
rect -3798 -6272 -1510 -6208
rect -1446 -6272 -1426 -6208
rect -3798 -6288 -1426 -6272
rect -3798 -6352 -1510 -6288
rect -1446 -6352 -1426 -6288
rect -3798 -6368 -1426 -6352
rect -3798 -6432 -1510 -6368
rect -1446 -6432 -1426 -6368
rect -3798 -6448 -1426 -6432
rect -3798 -6512 -1510 -6448
rect -1446 -6512 -1426 -6448
rect -3798 -6528 -1426 -6512
rect -3798 -6592 -1510 -6528
rect -1446 -6592 -1426 -6528
rect -3798 -6608 -1426 -6592
rect -3798 -6672 -1510 -6608
rect -1446 -6672 -1426 -6608
rect -3798 -6688 -1426 -6672
rect -3798 -6752 -1510 -6688
rect -1446 -6752 -1426 -6688
rect -3798 -6768 -1426 -6752
rect -3798 -6832 -1510 -6768
rect -1446 -6832 -1426 -6768
rect -3798 -6848 -1426 -6832
rect -3798 -6912 -1510 -6848
rect -1446 -6912 -1426 -6848
rect -3798 -6928 -1426 -6912
rect -3798 -6992 -1510 -6928
rect -1446 -6992 -1426 -6928
rect -3798 -7008 -1426 -6992
rect -3798 -7072 -1510 -7008
rect -1446 -7072 -1426 -7008
rect -3798 -7088 -1426 -7072
rect -3798 -7152 -1510 -7088
rect -1446 -7152 -1426 -7088
rect -3798 -7168 -1426 -7152
rect -3798 -7232 -1510 -7168
rect -1446 -7232 -1426 -7168
rect -3798 -7248 -1426 -7232
rect -3798 -7312 -1510 -7248
rect -1446 -7312 -1426 -7248
rect -3798 -7328 -1426 -7312
rect -3798 -7392 -1510 -7328
rect -1446 -7392 -1426 -7328
rect -3798 -7408 -1426 -7392
rect -3798 -7472 -1510 -7408
rect -1446 -7472 -1426 -7408
rect -3798 -7488 -1426 -7472
rect -3798 -7552 -1510 -7488
rect -1446 -7552 -1426 -7488
rect -3798 -7568 -1426 -7552
rect -3798 -7632 -1510 -7568
rect -1446 -7632 -1426 -7568
rect -3798 -7648 -1426 -7632
rect -3798 -7712 -1510 -7648
rect -1446 -7712 -1426 -7648
rect -3798 -7728 -1426 -7712
rect -3798 -7792 -1510 -7728
rect -1446 -7792 -1426 -7728
rect -3798 -7808 -1426 -7792
rect -3798 -7872 -1510 -7808
rect -1446 -7872 -1426 -7808
rect -3798 -7888 -1426 -7872
rect -3798 -7952 -1510 -7888
rect -1446 -7952 -1426 -7888
rect -3798 -8000 -1426 -7952
rect -1186 -5968 1186 -5920
rect -1186 -6032 1102 -5968
rect 1166 -6032 1186 -5968
rect -1186 -6048 1186 -6032
rect -1186 -6112 1102 -6048
rect 1166 -6112 1186 -6048
rect -1186 -6128 1186 -6112
rect -1186 -6192 1102 -6128
rect 1166 -6192 1186 -6128
rect -1186 -6208 1186 -6192
rect -1186 -6272 1102 -6208
rect 1166 -6272 1186 -6208
rect -1186 -6288 1186 -6272
rect -1186 -6352 1102 -6288
rect 1166 -6352 1186 -6288
rect -1186 -6368 1186 -6352
rect -1186 -6432 1102 -6368
rect 1166 -6432 1186 -6368
rect -1186 -6448 1186 -6432
rect -1186 -6512 1102 -6448
rect 1166 -6512 1186 -6448
rect -1186 -6528 1186 -6512
rect -1186 -6592 1102 -6528
rect 1166 -6592 1186 -6528
rect -1186 -6608 1186 -6592
rect -1186 -6672 1102 -6608
rect 1166 -6672 1186 -6608
rect -1186 -6688 1186 -6672
rect -1186 -6752 1102 -6688
rect 1166 -6752 1186 -6688
rect -1186 -6768 1186 -6752
rect -1186 -6832 1102 -6768
rect 1166 -6832 1186 -6768
rect -1186 -6848 1186 -6832
rect -1186 -6912 1102 -6848
rect 1166 -6912 1186 -6848
rect -1186 -6928 1186 -6912
rect -1186 -6992 1102 -6928
rect 1166 -6992 1186 -6928
rect -1186 -7008 1186 -6992
rect -1186 -7072 1102 -7008
rect 1166 -7072 1186 -7008
rect -1186 -7088 1186 -7072
rect -1186 -7152 1102 -7088
rect 1166 -7152 1186 -7088
rect -1186 -7168 1186 -7152
rect -1186 -7232 1102 -7168
rect 1166 -7232 1186 -7168
rect -1186 -7248 1186 -7232
rect -1186 -7312 1102 -7248
rect 1166 -7312 1186 -7248
rect -1186 -7328 1186 -7312
rect -1186 -7392 1102 -7328
rect 1166 -7392 1186 -7328
rect -1186 -7408 1186 -7392
rect -1186 -7472 1102 -7408
rect 1166 -7472 1186 -7408
rect -1186 -7488 1186 -7472
rect -1186 -7552 1102 -7488
rect 1166 -7552 1186 -7488
rect -1186 -7568 1186 -7552
rect -1186 -7632 1102 -7568
rect 1166 -7632 1186 -7568
rect -1186 -7648 1186 -7632
rect -1186 -7712 1102 -7648
rect 1166 -7712 1186 -7648
rect -1186 -7728 1186 -7712
rect -1186 -7792 1102 -7728
rect 1166 -7792 1186 -7728
rect -1186 -7808 1186 -7792
rect -1186 -7872 1102 -7808
rect 1166 -7872 1186 -7808
rect -1186 -7888 1186 -7872
rect -1186 -7952 1102 -7888
rect 1166 -7952 1186 -7888
rect -1186 -8000 1186 -7952
rect 1426 -5968 3798 -5920
rect 1426 -6032 3714 -5968
rect 3778 -6032 3798 -5968
rect 1426 -6048 3798 -6032
rect 1426 -6112 3714 -6048
rect 3778 -6112 3798 -6048
rect 1426 -6128 3798 -6112
rect 1426 -6192 3714 -6128
rect 3778 -6192 3798 -6128
rect 1426 -6208 3798 -6192
rect 1426 -6272 3714 -6208
rect 3778 -6272 3798 -6208
rect 1426 -6288 3798 -6272
rect 1426 -6352 3714 -6288
rect 3778 -6352 3798 -6288
rect 1426 -6368 3798 -6352
rect 1426 -6432 3714 -6368
rect 3778 -6432 3798 -6368
rect 1426 -6448 3798 -6432
rect 1426 -6512 3714 -6448
rect 3778 -6512 3798 -6448
rect 1426 -6528 3798 -6512
rect 1426 -6592 3714 -6528
rect 3778 -6592 3798 -6528
rect 1426 -6608 3798 -6592
rect 1426 -6672 3714 -6608
rect 3778 -6672 3798 -6608
rect 1426 -6688 3798 -6672
rect 1426 -6752 3714 -6688
rect 3778 -6752 3798 -6688
rect 1426 -6768 3798 -6752
rect 1426 -6832 3714 -6768
rect 3778 -6832 3798 -6768
rect 1426 -6848 3798 -6832
rect 1426 -6912 3714 -6848
rect 3778 -6912 3798 -6848
rect 1426 -6928 3798 -6912
rect 1426 -6992 3714 -6928
rect 3778 -6992 3798 -6928
rect 1426 -7008 3798 -6992
rect 1426 -7072 3714 -7008
rect 3778 -7072 3798 -7008
rect 1426 -7088 3798 -7072
rect 1426 -7152 3714 -7088
rect 3778 -7152 3798 -7088
rect 1426 -7168 3798 -7152
rect 1426 -7232 3714 -7168
rect 3778 -7232 3798 -7168
rect 1426 -7248 3798 -7232
rect 1426 -7312 3714 -7248
rect 3778 -7312 3798 -7248
rect 1426 -7328 3798 -7312
rect 1426 -7392 3714 -7328
rect 3778 -7392 3798 -7328
rect 1426 -7408 3798 -7392
rect 1426 -7472 3714 -7408
rect 3778 -7472 3798 -7408
rect 1426 -7488 3798 -7472
rect 1426 -7552 3714 -7488
rect 3778 -7552 3798 -7488
rect 1426 -7568 3798 -7552
rect 1426 -7632 3714 -7568
rect 3778 -7632 3798 -7568
rect 1426 -7648 3798 -7632
rect 1426 -7712 3714 -7648
rect 3778 -7712 3798 -7648
rect 1426 -7728 3798 -7712
rect 1426 -7792 3714 -7728
rect 3778 -7792 3798 -7728
rect 1426 -7808 3798 -7792
rect 1426 -7872 3714 -7808
rect 3778 -7872 3798 -7808
rect 1426 -7888 3798 -7872
rect 1426 -7952 3714 -7888
rect 3778 -7952 3798 -7888
rect 1426 -8000 3798 -7952
rect 4038 -5968 6410 -5920
rect 4038 -6032 6326 -5968
rect 6390 -6032 6410 -5968
rect 4038 -6048 6410 -6032
rect 4038 -6112 6326 -6048
rect 6390 -6112 6410 -6048
rect 4038 -6128 6410 -6112
rect 4038 -6192 6326 -6128
rect 6390 -6192 6410 -6128
rect 4038 -6208 6410 -6192
rect 4038 -6272 6326 -6208
rect 6390 -6272 6410 -6208
rect 4038 -6288 6410 -6272
rect 4038 -6352 6326 -6288
rect 6390 -6352 6410 -6288
rect 4038 -6368 6410 -6352
rect 4038 -6432 6326 -6368
rect 6390 -6432 6410 -6368
rect 4038 -6448 6410 -6432
rect 4038 -6512 6326 -6448
rect 6390 -6512 6410 -6448
rect 4038 -6528 6410 -6512
rect 4038 -6592 6326 -6528
rect 6390 -6592 6410 -6528
rect 4038 -6608 6410 -6592
rect 4038 -6672 6326 -6608
rect 6390 -6672 6410 -6608
rect 4038 -6688 6410 -6672
rect 4038 -6752 6326 -6688
rect 6390 -6752 6410 -6688
rect 4038 -6768 6410 -6752
rect 4038 -6832 6326 -6768
rect 6390 -6832 6410 -6768
rect 4038 -6848 6410 -6832
rect 4038 -6912 6326 -6848
rect 6390 -6912 6410 -6848
rect 4038 -6928 6410 -6912
rect 4038 -6992 6326 -6928
rect 6390 -6992 6410 -6928
rect 4038 -7008 6410 -6992
rect 4038 -7072 6326 -7008
rect 6390 -7072 6410 -7008
rect 4038 -7088 6410 -7072
rect 4038 -7152 6326 -7088
rect 6390 -7152 6410 -7088
rect 4038 -7168 6410 -7152
rect 4038 -7232 6326 -7168
rect 6390 -7232 6410 -7168
rect 4038 -7248 6410 -7232
rect 4038 -7312 6326 -7248
rect 6390 -7312 6410 -7248
rect 4038 -7328 6410 -7312
rect 4038 -7392 6326 -7328
rect 6390 -7392 6410 -7328
rect 4038 -7408 6410 -7392
rect 4038 -7472 6326 -7408
rect 6390 -7472 6410 -7408
rect 4038 -7488 6410 -7472
rect 4038 -7552 6326 -7488
rect 6390 -7552 6410 -7488
rect 4038 -7568 6410 -7552
rect 4038 -7632 6326 -7568
rect 6390 -7632 6410 -7568
rect 4038 -7648 6410 -7632
rect 4038 -7712 6326 -7648
rect 6390 -7712 6410 -7648
rect 4038 -7728 6410 -7712
rect 4038 -7792 6326 -7728
rect 6390 -7792 6410 -7728
rect 4038 -7808 6410 -7792
rect 4038 -7872 6326 -7808
rect 6390 -7872 6410 -7808
rect 4038 -7888 6410 -7872
rect 4038 -7952 6326 -7888
rect 6390 -7952 6410 -7888
rect 4038 -8000 6410 -7952
rect 6650 -5968 9022 -5920
rect 6650 -6032 8938 -5968
rect 9002 -6032 9022 -5968
rect 6650 -6048 9022 -6032
rect 6650 -6112 8938 -6048
rect 9002 -6112 9022 -6048
rect 6650 -6128 9022 -6112
rect 6650 -6192 8938 -6128
rect 9002 -6192 9022 -6128
rect 6650 -6208 9022 -6192
rect 6650 -6272 8938 -6208
rect 9002 -6272 9022 -6208
rect 6650 -6288 9022 -6272
rect 6650 -6352 8938 -6288
rect 9002 -6352 9022 -6288
rect 6650 -6368 9022 -6352
rect 6650 -6432 8938 -6368
rect 9002 -6432 9022 -6368
rect 6650 -6448 9022 -6432
rect 6650 -6512 8938 -6448
rect 9002 -6512 9022 -6448
rect 6650 -6528 9022 -6512
rect 6650 -6592 8938 -6528
rect 9002 -6592 9022 -6528
rect 6650 -6608 9022 -6592
rect 6650 -6672 8938 -6608
rect 9002 -6672 9022 -6608
rect 6650 -6688 9022 -6672
rect 6650 -6752 8938 -6688
rect 9002 -6752 9022 -6688
rect 6650 -6768 9022 -6752
rect 6650 -6832 8938 -6768
rect 9002 -6832 9022 -6768
rect 6650 -6848 9022 -6832
rect 6650 -6912 8938 -6848
rect 9002 -6912 9022 -6848
rect 6650 -6928 9022 -6912
rect 6650 -6992 8938 -6928
rect 9002 -6992 9022 -6928
rect 6650 -7008 9022 -6992
rect 6650 -7072 8938 -7008
rect 9002 -7072 9022 -7008
rect 6650 -7088 9022 -7072
rect 6650 -7152 8938 -7088
rect 9002 -7152 9022 -7088
rect 6650 -7168 9022 -7152
rect 6650 -7232 8938 -7168
rect 9002 -7232 9022 -7168
rect 6650 -7248 9022 -7232
rect 6650 -7312 8938 -7248
rect 9002 -7312 9022 -7248
rect 6650 -7328 9022 -7312
rect 6650 -7392 8938 -7328
rect 9002 -7392 9022 -7328
rect 6650 -7408 9022 -7392
rect 6650 -7472 8938 -7408
rect 9002 -7472 9022 -7408
rect 6650 -7488 9022 -7472
rect 6650 -7552 8938 -7488
rect 9002 -7552 9022 -7488
rect 6650 -7568 9022 -7552
rect 6650 -7632 8938 -7568
rect 9002 -7632 9022 -7568
rect 6650 -7648 9022 -7632
rect 6650 -7712 8938 -7648
rect 9002 -7712 9022 -7648
rect 6650 -7728 9022 -7712
rect 6650 -7792 8938 -7728
rect 9002 -7792 9022 -7728
rect 6650 -7808 9022 -7792
rect 6650 -7872 8938 -7808
rect 9002 -7872 9022 -7808
rect 6650 -7888 9022 -7872
rect 6650 -7952 8938 -7888
rect 9002 -7952 9022 -7888
rect 6650 -8000 9022 -7952
<< via3 >>
rect -6734 7888 -6670 7952
rect -6734 7808 -6670 7872
rect -6734 7728 -6670 7792
rect -6734 7648 -6670 7712
rect -6734 7568 -6670 7632
rect -6734 7488 -6670 7552
rect -6734 7408 -6670 7472
rect -6734 7328 -6670 7392
rect -6734 7248 -6670 7312
rect -6734 7168 -6670 7232
rect -6734 7088 -6670 7152
rect -6734 7008 -6670 7072
rect -6734 6928 -6670 6992
rect -6734 6848 -6670 6912
rect -6734 6768 -6670 6832
rect -6734 6688 -6670 6752
rect -6734 6608 -6670 6672
rect -6734 6528 -6670 6592
rect -6734 6448 -6670 6512
rect -6734 6368 -6670 6432
rect -6734 6288 -6670 6352
rect -6734 6208 -6670 6272
rect -6734 6128 -6670 6192
rect -6734 6048 -6670 6112
rect -6734 5968 -6670 6032
rect -4122 7888 -4058 7952
rect -4122 7808 -4058 7872
rect -4122 7728 -4058 7792
rect -4122 7648 -4058 7712
rect -4122 7568 -4058 7632
rect -4122 7488 -4058 7552
rect -4122 7408 -4058 7472
rect -4122 7328 -4058 7392
rect -4122 7248 -4058 7312
rect -4122 7168 -4058 7232
rect -4122 7088 -4058 7152
rect -4122 7008 -4058 7072
rect -4122 6928 -4058 6992
rect -4122 6848 -4058 6912
rect -4122 6768 -4058 6832
rect -4122 6688 -4058 6752
rect -4122 6608 -4058 6672
rect -4122 6528 -4058 6592
rect -4122 6448 -4058 6512
rect -4122 6368 -4058 6432
rect -4122 6288 -4058 6352
rect -4122 6208 -4058 6272
rect -4122 6128 -4058 6192
rect -4122 6048 -4058 6112
rect -4122 5968 -4058 6032
rect -1510 7888 -1446 7952
rect -1510 7808 -1446 7872
rect -1510 7728 -1446 7792
rect -1510 7648 -1446 7712
rect -1510 7568 -1446 7632
rect -1510 7488 -1446 7552
rect -1510 7408 -1446 7472
rect -1510 7328 -1446 7392
rect -1510 7248 -1446 7312
rect -1510 7168 -1446 7232
rect -1510 7088 -1446 7152
rect -1510 7008 -1446 7072
rect -1510 6928 -1446 6992
rect -1510 6848 -1446 6912
rect -1510 6768 -1446 6832
rect -1510 6688 -1446 6752
rect -1510 6608 -1446 6672
rect -1510 6528 -1446 6592
rect -1510 6448 -1446 6512
rect -1510 6368 -1446 6432
rect -1510 6288 -1446 6352
rect -1510 6208 -1446 6272
rect -1510 6128 -1446 6192
rect -1510 6048 -1446 6112
rect -1510 5968 -1446 6032
rect 1102 7888 1166 7952
rect 1102 7808 1166 7872
rect 1102 7728 1166 7792
rect 1102 7648 1166 7712
rect 1102 7568 1166 7632
rect 1102 7488 1166 7552
rect 1102 7408 1166 7472
rect 1102 7328 1166 7392
rect 1102 7248 1166 7312
rect 1102 7168 1166 7232
rect 1102 7088 1166 7152
rect 1102 7008 1166 7072
rect 1102 6928 1166 6992
rect 1102 6848 1166 6912
rect 1102 6768 1166 6832
rect 1102 6688 1166 6752
rect 1102 6608 1166 6672
rect 1102 6528 1166 6592
rect 1102 6448 1166 6512
rect 1102 6368 1166 6432
rect 1102 6288 1166 6352
rect 1102 6208 1166 6272
rect 1102 6128 1166 6192
rect 1102 6048 1166 6112
rect 1102 5968 1166 6032
rect 3714 7888 3778 7952
rect 3714 7808 3778 7872
rect 3714 7728 3778 7792
rect 3714 7648 3778 7712
rect 3714 7568 3778 7632
rect 3714 7488 3778 7552
rect 3714 7408 3778 7472
rect 3714 7328 3778 7392
rect 3714 7248 3778 7312
rect 3714 7168 3778 7232
rect 3714 7088 3778 7152
rect 3714 7008 3778 7072
rect 3714 6928 3778 6992
rect 3714 6848 3778 6912
rect 3714 6768 3778 6832
rect 3714 6688 3778 6752
rect 3714 6608 3778 6672
rect 3714 6528 3778 6592
rect 3714 6448 3778 6512
rect 3714 6368 3778 6432
rect 3714 6288 3778 6352
rect 3714 6208 3778 6272
rect 3714 6128 3778 6192
rect 3714 6048 3778 6112
rect 3714 5968 3778 6032
rect 6326 7888 6390 7952
rect 6326 7808 6390 7872
rect 6326 7728 6390 7792
rect 6326 7648 6390 7712
rect 6326 7568 6390 7632
rect 6326 7488 6390 7552
rect 6326 7408 6390 7472
rect 6326 7328 6390 7392
rect 6326 7248 6390 7312
rect 6326 7168 6390 7232
rect 6326 7088 6390 7152
rect 6326 7008 6390 7072
rect 6326 6928 6390 6992
rect 6326 6848 6390 6912
rect 6326 6768 6390 6832
rect 6326 6688 6390 6752
rect 6326 6608 6390 6672
rect 6326 6528 6390 6592
rect 6326 6448 6390 6512
rect 6326 6368 6390 6432
rect 6326 6288 6390 6352
rect 6326 6208 6390 6272
rect 6326 6128 6390 6192
rect 6326 6048 6390 6112
rect 6326 5968 6390 6032
rect 8938 7888 9002 7952
rect 8938 7808 9002 7872
rect 8938 7728 9002 7792
rect 8938 7648 9002 7712
rect 8938 7568 9002 7632
rect 8938 7488 9002 7552
rect 8938 7408 9002 7472
rect 8938 7328 9002 7392
rect 8938 7248 9002 7312
rect 8938 7168 9002 7232
rect 8938 7088 9002 7152
rect 8938 7008 9002 7072
rect 8938 6928 9002 6992
rect 8938 6848 9002 6912
rect 8938 6768 9002 6832
rect 8938 6688 9002 6752
rect 8938 6608 9002 6672
rect 8938 6528 9002 6592
rect 8938 6448 9002 6512
rect 8938 6368 9002 6432
rect 8938 6288 9002 6352
rect 8938 6208 9002 6272
rect 8938 6128 9002 6192
rect 8938 6048 9002 6112
rect 8938 5968 9002 6032
rect -6734 5568 -6670 5632
rect -6734 5488 -6670 5552
rect -6734 5408 -6670 5472
rect -6734 5328 -6670 5392
rect -6734 5248 -6670 5312
rect -6734 5168 -6670 5232
rect -6734 5088 -6670 5152
rect -6734 5008 -6670 5072
rect -6734 4928 -6670 4992
rect -6734 4848 -6670 4912
rect -6734 4768 -6670 4832
rect -6734 4688 -6670 4752
rect -6734 4608 -6670 4672
rect -6734 4528 -6670 4592
rect -6734 4448 -6670 4512
rect -6734 4368 -6670 4432
rect -6734 4288 -6670 4352
rect -6734 4208 -6670 4272
rect -6734 4128 -6670 4192
rect -6734 4048 -6670 4112
rect -6734 3968 -6670 4032
rect -6734 3888 -6670 3952
rect -6734 3808 -6670 3872
rect -6734 3728 -6670 3792
rect -6734 3648 -6670 3712
rect -4122 5568 -4058 5632
rect -4122 5488 -4058 5552
rect -4122 5408 -4058 5472
rect -4122 5328 -4058 5392
rect -4122 5248 -4058 5312
rect -4122 5168 -4058 5232
rect -4122 5088 -4058 5152
rect -4122 5008 -4058 5072
rect -4122 4928 -4058 4992
rect -4122 4848 -4058 4912
rect -4122 4768 -4058 4832
rect -4122 4688 -4058 4752
rect -4122 4608 -4058 4672
rect -4122 4528 -4058 4592
rect -4122 4448 -4058 4512
rect -4122 4368 -4058 4432
rect -4122 4288 -4058 4352
rect -4122 4208 -4058 4272
rect -4122 4128 -4058 4192
rect -4122 4048 -4058 4112
rect -4122 3968 -4058 4032
rect -4122 3888 -4058 3952
rect -4122 3808 -4058 3872
rect -4122 3728 -4058 3792
rect -4122 3648 -4058 3712
rect -1510 5568 -1446 5632
rect -1510 5488 -1446 5552
rect -1510 5408 -1446 5472
rect -1510 5328 -1446 5392
rect -1510 5248 -1446 5312
rect -1510 5168 -1446 5232
rect -1510 5088 -1446 5152
rect -1510 5008 -1446 5072
rect -1510 4928 -1446 4992
rect -1510 4848 -1446 4912
rect -1510 4768 -1446 4832
rect -1510 4688 -1446 4752
rect -1510 4608 -1446 4672
rect -1510 4528 -1446 4592
rect -1510 4448 -1446 4512
rect -1510 4368 -1446 4432
rect -1510 4288 -1446 4352
rect -1510 4208 -1446 4272
rect -1510 4128 -1446 4192
rect -1510 4048 -1446 4112
rect -1510 3968 -1446 4032
rect -1510 3888 -1446 3952
rect -1510 3808 -1446 3872
rect -1510 3728 -1446 3792
rect -1510 3648 -1446 3712
rect 1102 5568 1166 5632
rect 1102 5488 1166 5552
rect 1102 5408 1166 5472
rect 1102 5328 1166 5392
rect 1102 5248 1166 5312
rect 1102 5168 1166 5232
rect 1102 5088 1166 5152
rect 1102 5008 1166 5072
rect 1102 4928 1166 4992
rect 1102 4848 1166 4912
rect 1102 4768 1166 4832
rect 1102 4688 1166 4752
rect 1102 4608 1166 4672
rect 1102 4528 1166 4592
rect 1102 4448 1166 4512
rect 1102 4368 1166 4432
rect 1102 4288 1166 4352
rect 1102 4208 1166 4272
rect 1102 4128 1166 4192
rect 1102 4048 1166 4112
rect 1102 3968 1166 4032
rect 1102 3888 1166 3952
rect 1102 3808 1166 3872
rect 1102 3728 1166 3792
rect 1102 3648 1166 3712
rect 3714 5568 3778 5632
rect 3714 5488 3778 5552
rect 3714 5408 3778 5472
rect 3714 5328 3778 5392
rect 3714 5248 3778 5312
rect 3714 5168 3778 5232
rect 3714 5088 3778 5152
rect 3714 5008 3778 5072
rect 3714 4928 3778 4992
rect 3714 4848 3778 4912
rect 3714 4768 3778 4832
rect 3714 4688 3778 4752
rect 3714 4608 3778 4672
rect 3714 4528 3778 4592
rect 3714 4448 3778 4512
rect 3714 4368 3778 4432
rect 3714 4288 3778 4352
rect 3714 4208 3778 4272
rect 3714 4128 3778 4192
rect 3714 4048 3778 4112
rect 3714 3968 3778 4032
rect 3714 3888 3778 3952
rect 3714 3808 3778 3872
rect 3714 3728 3778 3792
rect 3714 3648 3778 3712
rect 6326 5568 6390 5632
rect 6326 5488 6390 5552
rect 6326 5408 6390 5472
rect 6326 5328 6390 5392
rect 6326 5248 6390 5312
rect 6326 5168 6390 5232
rect 6326 5088 6390 5152
rect 6326 5008 6390 5072
rect 6326 4928 6390 4992
rect 6326 4848 6390 4912
rect 6326 4768 6390 4832
rect 6326 4688 6390 4752
rect 6326 4608 6390 4672
rect 6326 4528 6390 4592
rect 6326 4448 6390 4512
rect 6326 4368 6390 4432
rect 6326 4288 6390 4352
rect 6326 4208 6390 4272
rect 6326 4128 6390 4192
rect 6326 4048 6390 4112
rect 6326 3968 6390 4032
rect 6326 3888 6390 3952
rect 6326 3808 6390 3872
rect 6326 3728 6390 3792
rect 6326 3648 6390 3712
rect 8938 5568 9002 5632
rect 8938 5488 9002 5552
rect 8938 5408 9002 5472
rect 8938 5328 9002 5392
rect 8938 5248 9002 5312
rect 8938 5168 9002 5232
rect 8938 5088 9002 5152
rect 8938 5008 9002 5072
rect 8938 4928 9002 4992
rect 8938 4848 9002 4912
rect 8938 4768 9002 4832
rect 8938 4688 9002 4752
rect 8938 4608 9002 4672
rect 8938 4528 9002 4592
rect 8938 4448 9002 4512
rect 8938 4368 9002 4432
rect 8938 4288 9002 4352
rect 8938 4208 9002 4272
rect 8938 4128 9002 4192
rect 8938 4048 9002 4112
rect 8938 3968 9002 4032
rect 8938 3888 9002 3952
rect 8938 3808 9002 3872
rect 8938 3728 9002 3792
rect 8938 3648 9002 3712
rect -6734 3248 -6670 3312
rect -6734 3168 -6670 3232
rect -6734 3088 -6670 3152
rect -6734 3008 -6670 3072
rect -6734 2928 -6670 2992
rect -6734 2848 -6670 2912
rect -6734 2768 -6670 2832
rect -6734 2688 -6670 2752
rect -6734 2608 -6670 2672
rect -6734 2528 -6670 2592
rect -6734 2448 -6670 2512
rect -6734 2368 -6670 2432
rect -6734 2288 -6670 2352
rect -6734 2208 -6670 2272
rect -6734 2128 -6670 2192
rect -6734 2048 -6670 2112
rect -6734 1968 -6670 2032
rect -6734 1888 -6670 1952
rect -6734 1808 -6670 1872
rect -6734 1728 -6670 1792
rect -6734 1648 -6670 1712
rect -6734 1568 -6670 1632
rect -6734 1488 -6670 1552
rect -6734 1408 -6670 1472
rect -6734 1328 -6670 1392
rect -4122 3248 -4058 3312
rect -4122 3168 -4058 3232
rect -4122 3088 -4058 3152
rect -4122 3008 -4058 3072
rect -4122 2928 -4058 2992
rect -4122 2848 -4058 2912
rect -4122 2768 -4058 2832
rect -4122 2688 -4058 2752
rect -4122 2608 -4058 2672
rect -4122 2528 -4058 2592
rect -4122 2448 -4058 2512
rect -4122 2368 -4058 2432
rect -4122 2288 -4058 2352
rect -4122 2208 -4058 2272
rect -4122 2128 -4058 2192
rect -4122 2048 -4058 2112
rect -4122 1968 -4058 2032
rect -4122 1888 -4058 1952
rect -4122 1808 -4058 1872
rect -4122 1728 -4058 1792
rect -4122 1648 -4058 1712
rect -4122 1568 -4058 1632
rect -4122 1488 -4058 1552
rect -4122 1408 -4058 1472
rect -4122 1328 -4058 1392
rect -1510 3248 -1446 3312
rect -1510 3168 -1446 3232
rect -1510 3088 -1446 3152
rect -1510 3008 -1446 3072
rect -1510 2928 -1446 2992
rect -1510 2848 -1446 2912
rect -1510 2768 -1446 2832
rect -1510 2688 -1446 2752
rect -1510 2608 -1446 2672
rect -1510 2528 -1446 2592
rect -1510 2448 -1446 2512
rect -1510 2368 -1446 2432
rect -1510 2288 -1446 2352
rect -1510 2208 -1446 2272
rect -1510 2128 -1446 2192
rect -1510 2048 -1446 2112
rect -1510 1968 -1446 2032
rect -1510 1888 -1446 1952
rect -1510 1808 -1446 1872
rect -1510 1728 -1446 1792
rect -1510 1648 -1446 1712
rect -1510 1568 -1446 1632
rect -1510 1488 -1446 1552
rect -1510 1408 -1446 1472
rect -1510 1328 -1446 1392
rect 1102 3248 1166 3312
rect 1102 3168 1166 3232
rect 1102 3088 1166 3152
rect 1102 3008 1166 3072
rect 1102 2928 1166 2992
rect 1102 2848 1166 2912
rect 1102 2768 1166 2832
rect 1102 2688 1166 2752
rect 1102 2608 1166 2672
rect 1102 2528 1166 2592
rect 1102 2448 1166 2512
rect 1102 2368 1166 2432
rect 1102 2288 1166 2352
rect 1102 2208 1166 2272
rect 1102 2128 1166 2192
rect 1102 2048 1166 2112
rect 1102 1968 1166 2032
rect 1102 1888 1166 1952
rect 1102 1808 1166 1872
rect 1102 1728 1166 1792
rect 1102 1648 1166 1712
rect 1102 1568 1166 1632
rect 1102 1488 1166 1552
rect 1102 1408 1166 1472
rect 1102 1328 1166 1392
rect 3714 3248 3778 3312
rect 3714 3168 3778 3232
rect 3714 3088 3778 3152
rect 3714 3008 3778 3072
rect 3714 2928 3778 2992
rect 3714 2848 3778 2912
rect 3714 2768 3778 2832
rect 3714 2688 3778 2752
rect 3714 2608 3778 2672
rect 3714 2528 3778 2592
rect 3714 2448 3778 2512
rect 3714 2368 3778 2432
rect 3714 2288 3778 2352
rect 3714 2208 3778 2272
rect 3714 2128 3778 2192
rect 3714 2048 3778 2112
rect 3714 1968 3778 2032
rect 3714 1888 3778 1952
rect 3714 1808 3778 1872
rect 3714 1728 3778 1792
rect 3714 1648 3778 1712
rect 3714 1568 3778 1632
rect 3714 1488 3778 1552
rect 3714 1408 3778 1472
rect 3714 1328 3778 1392
rect 6326 3248 6390 3312
rect 6326 3168 6390 3232
rect 6326 3088 6390 3152
rect 6326 3008 6390 3072
rect 6326 2928 6390 2992
rect 6326 2848 6390 2912
rect 6326 2768 6390 2832
rect 6326 2688 6390 2752
rect 6326 2608 6390 2672
rect 6326 2528 6390 2592
rect 6326 2448 6390 2512
rect 6326 2368 6390 2432
rect 6326 2288 6390 2352
rect 6326 2208 6390 2272
rect 6326 2128 6390 2192
rect 6326 2048 6390 2112
rect 6326 1968 6390 2032
rect 6326 1888 6390 1952
rect 6326 1808 6390 1872
rect 6326 1728 6390 1792
rect 6326 1648 6390 1712
rect 6326 1568 6390 1632
rect 6326 1488 6390 1552
rect 6326 1408 6390 1472
rect 6326 1328 6390 1392
rect 8938 3248 9002 3312
rect 8938 3168 9002 3232
rect 8938 3088 9002 3152
rect 8938 3008 9002 3072
rect 8938 2928 9002 2992
rect 8938 2848 9002 2912
rect 8938 2768 9002 2832
rect 8938 2688 9002 2752
rect 8938 2608 9002 2672
rect 8938 2528 9002 2592
rect 8938 2448 9002 2512
rect 8938 2368 9002 2432
rect 8938 2288 9002 2352
rect 8938 2208 9002 2272
rect 8938 2128 9002 2192
rect 8938 2048 9002 2112
rect 8938 1968 9002 2032
rect 8938 1888 9002 1952
rect 8938 1808 9002 1872
rect 8938 1728 9002 1792
rect 8938 1648 9002 1712
rect 8938 1568 9002 1632
rect 8938 1488 9002 1552
rect 8938 1408 9002 1472
rect 8938 1328 9002 1392
rect -6734 928 -6670 992
rect -6734 848 -6670 912
rect -6734 768 -6670 832
rect -6734 688 -6670 752
rect -6734 608 -6670 672
rect -6734 528 -6670 592
rect -6734 448 -6670 512
rect -6734 368 -6670 432
rect -6734 288 -6670 352
rect -6734 208 -6670 272
rect -6734 128 -6670 192
rect -6734 48 -6670 112
rect -6734 -32 -6670 32
rect -6734 -112 -6670 -48
rect -6734 -192 -6670 -128
rect -6734 -272 -6670 -208
rect -6734 -352 -6670 -288
rect -6734 -432 -6670 -368
rect -6734 -512 -6670 -448
rect -6734 -592 -6670 -528
rect -6734 -672 -6670 -608
rect -6734 -752 -6670 -688
rect -6734 -832 -6670 -768
rect -6734 -912 -6670 -848
rect -6734 -992 -6670 -928
rect -4122 928 -4058 992
rect -4122 848 -4058 912
rect -4122 768 -4058 832
rect -4122 688 -4058 752
rect -4122 608 -4058 672
rect -4122 528 -4058 592
rect -4122 448 -4058 512
rect -4122 368 -4058 432
rect -4122 288 -4058 352
rect -4122 208 -4058 272
rect -4122 128 -4058 192
rect -4122 48 -4058 112
rect -4122 -32 -4058 32
rect -4122 -112 -4058 -48
rect -4122 -192 -4058 -128
rect -4122 -272 -4058 -208
rect -4122 -352 -4058 -288
rect -4122 -432 -4058 -368
rect -4122 -512 -4058 -448
rect -4122 -592 -4058 -528
rect -4122 -672 -4058 -608
rect -4122 -752 -4058 -688
rect -4122 -832 -4058 -768
rect -4122 -912 -4058 -848
rect -4122 -992 -4058 -928
rect -1510 928 -1446 992
rect -1510 848 -1446 912
rect -1510 768 -1446 832
rect -1510 688 -1446 752
rect -1510 608 -1446 672
rect -1510 528 -1446 592
rect -1510 448 -1446 512
rect -1510 368 -1446 432
rect -1510 288 -1446 352
rect -1510 208 -1446 272
rect -1510 128 -1446 192
rect -1510 48 -1446 112
rect -1510 -32 -1446 32
rect -1510 -112 -1446 -48
rect -1510 -192 -1446 -128
rect -1510 -272 -1446 -208
rect -1510 -352 -1446 -288
rect -1510 -432 -1446 -368
rect -1510 -512 -1446 -448
rect -1510 -592 -1446 -528
rect -1510 -672 -1446 -608
rect -1510 -752 -1446 -688
rect -1510 -832 -1446 -768
rect -1510 -912 -1446 -848
rect -1510 -992 -1446 -928
rect 1102 928 1166 992
rect 1102 848 1166 912
rect 1102 768 1166 832
rect 1102 688 1166 752
rect 1102 608 1166 672
rect 1102 528 1166 592
rect 1102 448 1166 512
rect 1102 368 1166 432
rect 1102 288 1166 352
rect 1102 208 1166 272
rect 1102 128 1166 192
rect 1102 48 1166 112
rect 1102 -32 1166 32
rect 1102 -112 1166 -48
rect 1102 -192 1166 -128
rect 1102 -272 1166 -208
rect 1102 -352 1166 -288
rect 1102 -432 1166 -368
rect 1102 -512 1166 -448
rect 1102 -592 1166 -528
rect 1102 -672 1166 -608
rect 1102 -752 1166 -688
rect 1102 -832 1166 -768
rect 1102 -912 1166 -848
rect 1102 -992 1166 -928
rect 3714 928 3778 992
rect 3714 848 3778 912
rect 3714 768 3778 832
rect 3714 688 3778 752
rect 3714 608 3778 672
rect 3714 528 3778 592
rect 3714 448 3778 512
rect 3714 368 3778 432
rect 3714 288 3778 352
rect 3714 208 3778 272
rect 3714 128 3778 192
rect 3714 48 3778 112
rect 3714 -32 3778 32
rect 3714 -112 3778 -48
rect 3714 -192 3778 -128
rect 3714 -272 3778 -208
rect 3714 -352 3778 -288
rect 3714 -432 3778 -368
rect 3714 -512 3778 -448
rect 3714 -592 3778 -528
rect 3714 -672 3778 -608
rect 3714 -752 3778 -688
rect 3714 -832 3778 -768
rect 3714 -912 3778 -848
rect 3714 -992 3778 -928
rect 6326 928 6390 992
rect 6326 848 6390 912
rect 6326 768 6390 832
rect 6326 688 6390 752
rect 6326 608 6390 672
rect 6326 528 6390 592
rect 6326 448 6390 512
rect 6326 368 6390 432
rect 6326 288 6390 352
rect 6326 208 6390 272
rect 6326 128 6390 192
rect 6326 48 6390 112
rect 6326 -32 6390 32
rect 6326 -112 6390 -48
rect 6326 -192 6390 -128
rect 6326 -272 6390 -208
rect 6326 -352 6390 -288
rect 6326 -432 6390 -368
rect 6326 -512 6390 -448
rect 6326 -592 6390 -528
rect 6326 -672 6390 -608
rect 6326 -752 6390 -688
rect 6326 -832 6390 -768
rect 6326 -912 6390 -848
rect 6326 -992 6390 -928
rect 8938 928 9002 992
rect 8938 848 9002 912
rect 8938 768 9002 832
rect 8938 688 9002 752
rect 8938 608 9002 672
rect 8938 528 9002 592
rect 8938 448 9002 512
rect 8938 368 9002 432
rect 8938 288 9002 352
rect 8938 208 9002 272
rect 8938 128 9002 192
rect 8938 48 9002 112
rect 8938 -32 9002 32
rect 8938 -112 9002 -48
rect 8938 -192 9002 -128
rect 8938 -272 9002 -208
rect 8938 -352 9002 -288
rect 8938 -432 9002 -368
rect 8938 -512 9002 -448
rect 8938 -592 9002 -528
rect 8938 -672 9002 -608
rect 8938 -752 9002 -688
rect 8938 -832 9002 -768
rect 8938 -912 9002 -848
rect 8938 -992 9002 -928
rect -6734 -1392 -6670 -1328
rect -6734 -1472 -6670 -1408
rect -6734 -1552 -6670 -1488
rect -6734 -1632 -6670 -1568
rect -6734 -1712 -6670 -1648
rect -6734 -1792 -6670 -1728
rect -6734 -1872 -6670 -1808
rect -6734 -1952 -6670 -1888
rect -6734 -2032 -6670 -1968
rect -6734 -2112 -6670 -2048
rect -6734 -2192 -6670 -2128
rect -6734 -2272 -6670 -2208
rect -6734 -2352 -6670 -2288
rect -6734 -2432 -6670 -2368
rect -6734 -2512 -6670 -2448
rect -6734 -2592 -6670 -2528
rect -6734 -2672 -6670 -2608
rect -6734 -2752 -6670 -2688
rect -6734 -2832 -6670 -2768
rect -6734 -2912 -6670 -2848
rect -6734 -2992 -6670 -2928
rect -6734 -3072 -6670 -3008
rect -6734 -3152 -6670 -3088
rect -6734 -3232 -6670 -3168
rect -6734 -3312 -6670 -3248
rect -4122 -1392 -4058 -1328
rect -4122 -1472 -4058 -1408
rect -4122 -1552 -4058 -1488
rect -4122 -1632 -4058 -1568
rect -4122 -1712 -4058 -1648
rect -4122 -1792 -4058 -1728
rect -4122 -1872 -4058 -1808
rect -4122 -1952 -4058 -1888
rect -4122 -2032 -4058 -1968
rect -4122 -2112 -4058 -2048
rect -4122 -2192 -4058 -2128
rect -4122 -2272 -4058 -2208
rect -4122 -2352 -4058 -2288
rect -4122 -2432 -4058 -2368
rect -4122 -2512 -4058 -2448
rect -4122 -2592 -4058 -2528
rect -4122 -2672 -4058 -2608
rect -4122 -2752 -4058 -2688
rect -4122 -2832 -4058 -2768
rect -4122 -2912 -4058 -2848
rect -4122 -2992 -4058 -2928
rect -4122 -3072 -4058 -3008
rect -4122 -3152 -4058 -3088
rect -4122 -3232 -4058 -3168
rect -4122 -3312 -4058 -3248
rect -1510 -1392 -1446 -1328
rect -1510 -1472 -1446 -1408
rect -1510 -1552 -1446 -1488
rect -1510 -1632 -1446 -1568
rect -1510 -1712 -1446 -1648
rect -1510 -1792 -1446 -1728
rect -1510 -1872 -1446 -1808
rect -1510 -1952 -1446 -1888
rect -1510 -2032 -1446 -1968
rect -1510 -2112 -1446 -2048
rect -1510 -2192 -1446 -2128
rect -1510 -2272 -1446 -2208
rect -1510 -2352 -1446 -2288
rect -1510 -2432 -1446 -2368
rect -1510 -2512 -1446 -2448
rect -1510 -2592 -1446 -2528
rect -1510 -2672 -1446 -2608
rect -1510 -2752 -1446 -2688
rect -1510 -2832 -1446 -2768
rect -1510 -2912 -1446 -2848
rect -1510 -2992 -1446 -2928
rect -1510 -3072 -1446 -3008
rect -1510 -3152 -1446 -3088
rect -1510 -3232 -1446 -3168
rect -1510 -3312 -1446 -3248
rect 1102 -1392 1166 -1328
rect 1102 -1472 1166 -1408
rect 1102 -1552 1166 -1488
rect 1102 -1632 1166 -1568
rect 1102 -1712 1166 -1648
rect 1102 -1792 1166 -1728
rect 1102 -1872 1166 -1808
rect 1102 -1952 1166 -1888
rect 1102 -2032 1166 -1968
rect 1102 -2112 1166 -2048
rect 1102 -2192 1166 -2128
rect 1102 -2272 1166 -2208
rect 1102 -2352 1166 -2288
rect 1102 -2432 1166 -2368
rect 1102 -2512 1166 -2448
rect 1102 -2592 1166 -2528
rect 1102 -2672 1166 -2608
rect 1102 -2752 1166 -2688
rect 1102 -2832 1166 -2768
rect 1102 -2912 1166 -2848
rect 1102 -2992 1166 -2928
rect 1102 -3072 1166 -3008
rect 1102 -3152 1166 -3088
rect 1102 -3232 1166 -3168
rect 1102 -3312 1166 -3248
rect 3714 -1392 3778 -1328
rect 3714 -1472 3778 -1408
rect 3714 -1552 3778 -1488
rect 3714 -1632 3778 -1568
rect 3714 -1712 3778 -1648
rect 3714 -1792 3778 -1728
rect 3714 -1872 3778 -1808
rect 3714 -1952 3778 -1888
rect 3714 -2032 3778 -1968
rect 3714 -2112 3778 -2048
rect 3714 -2192 3778 -2128
rect 3714 -2272 3778 -2208
rect 3714 -2352 3778 -2288
rect 3714 -2432 3778 -2368
rect 3714 -2512 3778 -2448
rect 3714 -2592 3778 -2528
rect 3714 -2672 3778 -2608
rect 3714 -2752 3778 -2688
rect 3714 -2832 3778 -2768
rect 3714 -2912 3778 -2848
rect 3714 -2992 3778 -2928
rect 3714 -3072 3778 -3008
rect 3714 -3152 3778 -3088
rect 3714 -3232 3778 -3168
rect 3714 -3312 3778 -3248
rect 6326 -1392 6390 -1328
rect 6326 -1472 6390 -1408
rect 6326 -1552 6390 -1488
rect 6326 -1632 6390 -1568
rect 6326 -1712 6390 -1648
rect 6326 -1792 6390 -1728
rect 6326 -1872 6390 -1808
rect 6326 -1952 6390 -1888
rect 6326 -2032 6390 -1968
rect 6326 -2112 6390 -2048
rect 6326 -2192 6390 -2128
rect 6326 -2272 6390 -2208
rect 6326 -2352 6390 -2288
rect 6326 -2432 6390 -2368
rect 6326 -2512 6390 -2448
rect 6326 -2592 6390 -2528
rect 6326 -2672 6390 -2608
rect 6326 -2752 6390 -2688
rect 6326 -2832 6390 -2768
rect 6326 -2912 6390 -2848
rect 6326 -2992 6390 -2928
rect 6326 -3072 6390 -3008
rect 6326 -3152 6390 -3088
rect 6326 -3232 6390 -3168
rect 6326 -3312 6390 -3248
rect 8938 -1392 9002 -1328
rect 8938 -1472 9002 -1408
rect 8938 -1552 9002 -1488
rect 8938 -1632 9002 -1568
rect 8938 -1712 9002 -1648
rect 8938 -1792 9002 -1728
rect 8938 -1872 9002 -1808
rect 8938 -1952 9002 -1888
rect 8938 -2032 9002 -1968
rect 8938 -2112 9002 -2048
rect 8938 -2192 9002 -2128
rect 8938 -2272 9002 -2208
rect 8938 -2352 9002 -2288
rect 8938 -2432 9002 -2368
rect 8938 -2512 9002 -2448
rect 8938 -2592 9002 -2528
rect 8938 -2672 9002 -2608
rect 8938 -2752 9002 -2688
rect 8938 -2832 9002 -2768
rect 8938 -2912 9002 -2848
rect 8938 -2992 9002 -2928
rect 8938 -3072 9002 -3008
rect 8938 -3152 9002 -3088
rect 8938 -3232 9002 -3168
rect 8938 -3312 9002 -3248
rect -6734 -3712 -6670 -3648
rect -6734 -3792 -6670 -3728
rect -6734 -3872 -6670 -3808
rect -6734 -3952 -6670 -3888
rect -6734 -4032 -6670 -3968
rect -6734 -4112 -6670 -4048
rect -6734 -4192 -6670 -4128
rect -6734 -4272 -6670 -4208
rect -6734 -4352 -6670 -4288
rect -6734 -4432 -6670 -4368
rect -6734 -4512 -6670 -4448
rect -6734 -4592 -6670 -4528
rect -6734 -4672 -6670 -4608
rect -6734 -4752 -6670 -4688
rect -6734 -4832 -6670 -4768
rect -6734 -4912 -6670 -4848
rect -6734 -4992 -6670 -4928
rect -6734 -5072 -6670 -5008
rect -6734 -5152 -6670 -5088
rect -6734 -5232 -6670 -5168
rect -6734 -5312 -6670 -5248
rect -6734 -5392 -6670 -5328
rect -6734 -5472 -6670 -5408
rect -6734 -5552 -6670 -5488
rect -6734 -5632 -6670 -5568
rect -4122 -3712 -4058 -3648
rect -4122 -3792 -4058 -3728
rect -4122 -3872 -4058 -3808
rect -4122 -3952 -4058 -3888
rect -4122 -4032 -4058 -3968
rect -4122 -4112 -4058 -4048
rect -4122 -4192 -4058 -4128
rect -4122 -4272 -4058 -4208
rect -4122 -4352 -4058 -4288
rect -4122 -4432 -4058 -4368
rect -4122 -4512 -4058 -4448
rect -4122 -4592 -4058 -4528
rect -4122 -4672 -4058 -4608
rect -4122 -4752 -4058 -4688
rect -4122 -4832 -4058 -4768
rect -4122 -4912 -4058 -4848
rect -4122 -4992 -4058 -4928
rect -4122 -5072 -4058 -5008
rect -4122 -5152 -4058 -5088
rect -4122 -5232 -4058 -5168
rect -4122 -5312 -4058 -5248
rect -4122 -5392 -4058 -5328
rect -4122 -5472 -4058 -5408
rect -4122 -5552 -4058 -5488
rect -4122 -5632 -4058 -5568
rect -1510 -3712 -1446 -3648
rect -1510 -3792 -1446 -3728
rect -1510 -3872 -1446 -3808
rect -1510 -3952 -1446 -3888
rect -1510 -4032 -1446 -3968
rect -1510 -4112 -1446 -4048
rect -1510 -4192 -1446 -4128
rect -1510 -4272 -1446 -4208
rect -1510 -4352 -1446 -4288
rect -1510 -4432 -1446 -4368
rect -1510 -4512 -1446 -4448
rect -1510 -4592 -1446 -4528
rect -1510 -4672 -1446 -4608
rect -1510 -4752 -1446 -4688
rect -1510 -4832 -1446 -4768
rect -1510 -4912 -1446 -4848
rect -1510 -4992 -1446 -4928
rect -1510 -5072 -1446 -5008
rect -1510 -5152 -1446 -5088
rect -1510 -5232 -1446 -5168
rect -1510 -5312 -1446 -5248
rect -1510 -5392 -1446 -5328
rect -1510 -5472 -1446 -5408
rect -1510 -5552 -1446 -5488
rect -1510 -5632 -1446 -5568
rect 1102 -3712 1166 -3648
rect 1102 -3792 1166 -3728
rect 1102 -3872 1166 -3808
rect 1102 -3952 1166 -3888
rect 1102 -4032 1166 -3968
rect 1102 -4112 1166 -4048
rect 1102 -4192 1166 -4128
rect 1102 -4272 1166 -4208
rect 1102 -4352 1166 -4288
rect 1102 -4432 1166 -4368
rect 1102 -4512 1166 -4448
rect 1102 -4592 1166 -4528
rect 1102 -4672 1166 -4608
rect 1102 -4752 1166 -4688
rect 1102 -4832 1166 -4768
rect 1102 -4912 1166 -4848
rect 1102 -4992 1166 -4928
rect 1102 -5072 1166 -5008
rect 1102 -5152 1166 -5088
rect 1102 -5232 1166 -5168
rect 1102 -5312 1166 -5248
rect 1102 -5392 1166 -5328
rect 1102 -5472 1166 -5408
rect 1102 -5552 1166 -5488
rect 1102 -5632 1166 -5568
rect 3714 -3712 3778 -3648
rect 3714 -3792 3778 -3728
rect 3714 -3872 3778 -3808
rect 3714 -3952 3778 -3888
rect 3714 -4032 3778 -3968
rect 3714 -4112 3778 -4048
rect 3714 -4192 3778 -4128
rect 3714 -4272 3778 -4208
rect 3714 -4352 3778 -4288
rect 3714 -4432 3778 -4368
rect 3714 -4512 3778 -4448
rect 3714 -4592 3778 -4528
rect 3714 -4672 3778 -4608
rect 3714 -4752 3778 -4688
rect 3714 -4832 3778 -4768
rect 3714 -4912 3778 -4848
rect 3714 -4992 3778 -4928
rect 3714 -5072 3778 -5008
rect 3714 -5152 3778 -5088
rect 3714 -5232 3778 -5168
rect 3714 -5312 3778 -5248
rect 3714 -5392 3778 -5328
rect 3714 -5472 3778 -5408
rect 3714 -5552 3778 -5488
rect 3714 -5632 3778 -5568
rect 6326 -3712 6390 -3648
rect 6326 -3792 6390 -3728
rect 6326 -3872 6390 -3808
rect 6326 -3952 6390 -3888
rect 6326 -4032 6390 -3968
rect 6326 -4112 6390 -4048
rect 6326 -4192 6390 -4128
rect 6326 -4272 6390 -4208
rect 6326 -4352 6390 -4288
rect 6326 -4432 6390 -4368
rect 6326 -4512 6390 -4448
rect 6326 -4592 6390 -4528
rect 6326 -4672 6390 -4608
rect 6326 -4752 6390 -4688
rect 6326 -4832 6390 -4768
rect 6326 -4912 6390 -4848
rect 6326 -4992 6390 -4928
rect 6326 -5072 6390 -5008
rect 6326 -5152 6390 -5088
rect 6326 -5232 6390 -5168
rect 6326 -5312 6390 -5248
rect 6326 -5392 6390 -5328
rect 6326 -5472 6390 -5408
rect 6326 -5552 6390 -5488
rect 6326 -5632 6390 -5568
rect 8938 -3712 9002 -3648
rect 8938 -3792 9002 -3728
rect 8938 -3872 9002 -3808
rect 8938 -3952 9002 -3888
rect 8938 -4032 9002 -3968
rect 8938 -4112 9002 -4048
rect 8938 -4192 9002 -4128
rect 8938 -4272 9002 -4208
rect 8938 -4352 9002 -4288
rect 8938 -4432 9002 -4368
rect 8938 -4512 9002 -4448
rect 8938 -4592 9002 -4528
rect 8938 -4672 9002 -4608
rect 8938 -4752 9002 -4688
rect 8938 -4832 9002 -4768
rect 8938 -4912 9002 -4848
rect 8938 -4992 9002 -4928
rect 8938 -5072 9002 -5008
rect 8938 -5152 9002 -5088
rect 8938 -5232 9002 -5168
rect 8938 -5312 9002 -5248
rect 8938 -5392 9002 -5328
rect 8938 -5472 9002 -5408
rect 8938 -5552 9002 -5488
rect 8938 -5632 9002 -5568
rect -6734 -6032 -6670 -5968
rect -6734 -6112 -6670 -6048
rect -6734 -6192 -6670 -6128
rect -6734 -6272 -6670 -6208
rect -6734 -6352 -6670 -6288
rect -6734 -6432 -6670 -6368
rect -6734 -6512 -6670 -6448
rect -6734 -6592 -6670 -6528
rect -6734 -6672 -6670 -6608
rect -6734 -6752 -6670 -6688
rect -6734 -6832 -6670 -6768
rect -6734 -6912 -6670 -6848
rect -6734 -6992 -6670 -6928
rect -6734 -7072 -6670 -7008
rect -6734 -7152 -6670 -7088
rect -6734 -7232 -6670 -7168
rect -6734 -7312 -6670 -7248
rect -6734 -7392 -6670 -7328
rect -6734 -7472 -6670 -7408
rect -6734 -7552 -6670 -7488
rect -6734 -7632 -6670 -7568
rect -6734 -7712 -6670 -7648
rect -6734 -7792 -6670 -7728
rect -6734 -7872 -6670 -7808
rect -6734 -7952 -6670 -7888
rect -4122 -6032 -4058 -5968
rect -4122 -6112 -4058 -6048
rect -4122 -6192 -4058 -6128
rect -4122 -6272 -4058 -6208
rect -4122 -6352 -4058 -6288
rect -4122 -6432 -4058 -6368
rect -4122 -6512 -4058 -6448
rect -4122 -6592 -4058 -6528
rect -4122 -6672 -4058 -6608
rect -4122 -6752 -4058 -6688
rect -4122 -6832 -4058 -6768
rect -4122 -6912 -4058 -6848
rect -4122 -6992 -4058 -6928
rect -4122 -7072 -4058 -7008
rect -4122 -7152 -4058 -7088
rect -4122 -7232 -4058 -7168
rect -4122 -7312 -4058 -7248
rect -4122 -7392 -4058 -7328
rect -4122 -7472 -4058 -7408
rect -4122 -7552 -4058 -7488
rect -4122 -7632 -4058 -7568
rect -4122 -7712 -4058 -7648
rect -4122 -7792 -4058 -7728
rect -4122 -7872 -4058 -7808
rect -4122 -7952 -4058 -7888
rect -1510 -6032 -1446 -5968
rect -1510 -6112 -1446 -6048
rect -1510 -6192 -1446 -6128
rect -1510 -6272 -1446 -6208
rect -1510 -6352 -1446 -6288
rect -1510 -6432 -1446 -6368
rect -1510 -6512 -1446 -6448
rect -1510 -6592 -1446 -6528
rect -1510 -6672 -1446 -6608
rect -1510 -6752 -1446 -6688
rect -1510 -6832 -1446 -6768
rect -1510 -6912 -1446 -6848
rect -1510 -6992 -1446 -6928
rect -1510 -7072 -1446 -7008
rect -1510 -7152 -1446 -7088
rect -1510 -7232 -1446 -7168
rect -1510 -7312 -1446 -7248
rect -1510 -7392 -1446 -7328
rect -1510 -7472 -1446 -7408
rect -1510 -7552 -1446 -7488
rect -1510 -7632 -1446 -7568
rect -1510 -7712 -1446 -7648
rect -1510 -7792 -1446 -7728
rect -1510 -7872 -1446 -7808
rect -1510 -7952 -1446 -7888
rect 1102 -6032 1166 -5968
rect 1102 -6112 1166 -6048
rect 1102 -6192 1166 -6128
rect 1102 -6272 1166 -6208
rect 1102 -6352 1166 -6288
rect 1102 -6432 1166 -6368
rect 1102 -6512 1166 -6448
rect 1102 -6592 1166 -6528
rect 1102 -6672 1166 -6608
rect 1102 -6752 1166 -6688
rect 1102 -6832 1166 -6768
rect 1102 -6912 1166 -6848
rect 1102 -6992 1166 -6928
rect 1102 -7072 1166 -7008
rect 1102 -7152 1166 -7088
rect 1102 -7232 1166 -7168
rect 1102 -7312 1166 -7248
rect 1102 -7392 1166 -7328
rect 1102 -7472 1166 -7408
rect 1102 -7552 1166 -7488
rect 1102 -7632 1166 -7568
rect 1102 -7712 1166 -7648
rect 1102 -7792 1166 -7728
rect 1102 -7872 1166 -7808
rect 1102 -7952 1166 -7888
rect 3714 -6032 3778 -5968
rect 3714 -6112 3778 -6048
rect 3714 -6192 3778 -6128
rect 3714 -6272 3778 -6208
rect 3714 -6352 3778 -6288
rect 3714 -6432 3778 -6368
rect 3714 -6512 3778 -6448
rect 3714 -6592 3778 -6528
rect 3714 -6672 3778 -6608
rect 3714 -6752 3778 -6688
rect 3714 -6832 3778 -6768
rect 3714 -6912 3778 -6848
rect 3714 -6992 3778 -6928
rect 3714 -7072 3778 -7008
rect 3714 -7152 3778 -7088
rect 3714 -7232 3778 -7168
rect 3714 -7312 3778 -7248
rect 3714 -7392 3778 -7328
rect 3714 -7472 3778 -7408
rect 3714 -7552 3778 -7488
rect 3714 -7632 3778 -7568
rect 3714 -7712 3778 -7648
rect 3714 -7792 3778 -7728
rect 3714 -7872 3778 -7808
rect 3714 -7952 3778 -7888
rect 6326 -6032 6390 -5968
rect 6326 -6112 6390 -6048
rect 6326 -6192 6390 -6128
rect 6326 -6272 6390 -6208
rect 6326 -6352 6390 -6288
rect 6326 -6432 6390 -6368
rect 6326 -6512 6390 -6448
rect 6326 -6592 6390 -6528
rect 6326 -6672 6390 -6608
rect 6326 -6752 6390 -6688
rect 6326 -6832 6390 -6768
rect 6326 -6912 6390 -6848
rect 6326 -6992 6390 -6928
rect 6326 -7072 6390 -7008
rect 6326 -7152 6390 -7088
rect 6326 -7232 6390 -7168
rect 6326 -7312 6390 -7248
rect 6326 -7392 6390 -7328
rect 6326 -7472 6390 -7408
rect 6326 -7552 6390 -7488
rect 6326 -7632 6390 -7568
rect 6326 -7712 6390 -7648
rect 6326 -7792 6390 -7728
rect 6326 -7872 6390 -7808
rect 6326 -7952 6390 -7888
rect 8938 -6032 9002 -5968
rect 8938 -6112 9002 -6048
rect 8938 -6192 9002 -6128
rect 8938 -6272 9002 -6208
rect 8938 -6352 9002 -6288
rect 8938 -6432 9002 -6368
rect 8938 -6512 9002 -6448
rect 8938 -6592 9002 -6528
rect 8938 -6672 9002 -6608
rect 8938 -6752 9002 -6688
rect 8938 -6832 9002 -6768
rect 8938 -6912 9002 -6848
rect 8938 -6992 9002 -6928
rect 8938 -7072 9002 -7008
rect 8938 -7152 9002 -7088
rect 8938 -7232 9002 -7168
rect 8938 -7312 9002 -7248
rect 8938 -7392 9002 -7328
rect 8938 -7472 9002 -7408
rect 8938 -7552 9002 -7488
rect 8938 -7632 9002 -7568
rect 8938 -7712 9002 -7648
rect 8938 -7792 9002 -7728
rect 8938 -7872 9002 -7808
rect 8938 -7952 9002 -7888
<< mimcap >>
rect -8982 7912 -6982 7960
rect -8982 6008 -8934 7912
rect -7030 6008 -6982 7912
rect -8982 5960 -6982 6008
rect -6370 7912 -4370 7960
rect -6370 6008 -6322 7912
rect -4418 6008 -4370 7912
rect -6370 5960 -4370 6008
rect -3758 7912 -1758 7960
rect -3758 6008 -3710 7912
rect -1806 6008 -1758 7912
rect -3758 5960 -1758 6008
rect -1146 7912 854 7960
rect -1146 6008 -1098 7912
rect 806 6008 854 7912
rect -1146 5960 854 6008
rect 1466 7912 3466 7960
rect 1466 6008 1514 7912
rect 3418 6008 3466 7912
rect 1466 5960 3466 6008
rect 4078 7912 6078 7960
rect 4078 6008 4126 7912
rect 6030 6008 6078 7912
rect 4078 5960 6078 6008
rect 6690 7912 8690 7960
rect 6690 6008 6738 7912
rect 8642 6008 8690 7912
rect 6690 5960 8690 6008
rect -8982 5592 -6982 5640
rect -8982 3688 -8934 5592
rect -7030 3688 -6982 5592
rect -8982 3640 -6982 3688
rect -6370 5592 -4370 5640
rect -6370 3688 -6322 5592
rect -4418 3688 -4370 5592
rect -6370 3640 -4370 3688
rect -3758 5592 -1758 5640
rect -3758 3688 -3710 5592
rect -1806 3688 -1758 5592
rect -3758 3640 -1758 3688
rect -1146 5592 854 5640
rect -1146 3688 -1098 5592
rect 806 3688 854 5592
rect -1146 3640 854 3688
rect 1466 5592 3466 5640
rect 1466 3688 1514 5592
rect 3418 3688 3466 5592
rect 1466 3640 3466 3688
rect 4078 5592 6078 5640
rect 4078 3688 4126 5592
rect 6030 3688 6078 5592
rect 4078 3640 6078 3688
rect 6690 5592 8690 5640
rect 6690 3688 6738 5592
rect 8642 3688 8690 5592
rect 6690 3640 8690 3688
rect -8982 3272 -6982 3320
rect -8982 1368 -8934 3272
rect -7030 1368 -6982 3272
rect -8982 1320 -6982 1368
rect -6370 3272 -4370 3320
rect -6370 1368 -6322 3272
rect -4418 1368 -4370 3272
rect -6370 1320 -4370 1368
rect -3758 3272 -1758 3320
rect -3758 1368 -3710 3272
rect -1806 1368 -1758 3272
rect -3758 1320 -1758 1368
rect -1146 3272 854 3320
rect -1146 1368 -1098 3272
rect 806 1368 854 3272
rect -1146 1320 854 1368
rect 1466 3272 3466 3320
rect 1466 1368 1514 3272
rect 3418 1368 3466 3272
rect 1466 1320 3466 1368
rect 4078 3272 6078 3320
rect 4078 1368 4126 3272
rect 6030 1368 6078 3272
rect 4078 1320 6078 1368
rect 6690 3272 8690 3320
rect 6690 1368 6738 3272
rect 8642 1368 8690 3272
rect 6690 1320 8690 1368
rect -8982 952 -6982 1000
rect -8982 -952 -8934 952
rect -7030 -952 -6982 952
rect -8982 -1000 -6982 -952
rect -6370 952 -4370 1000
rect -6370 -952 -6322 952
rect -4418 -952 -4370 952
rect -6370 -1000 -4370 -952
rect -3758 952 -1758 1000
rect -3758 -952 -3710 952
rect -1806 -952 -1758 952
rect -3758 -1000 -1758 -952
rect -1146 952 854 1000
rect -1146 -952 -1098 952
rect 806 -952 854 952
rect -1146 -1000 854 -952
rect 1466 952 3466 1000
rect 1466 -952 1514 952
rect 3418 -952 3466 952
rect 1466 -1000 3466 -952
rect 4078 952 6078 1000
rect 4078 -952 4126 952
rect 6030 -952 6078 952
rect 4078 -1000 6078 -952
rect 6690 952 8690 1000
rect 6690 -952 6738 952
rect 8642 -952 8690 952
rect 6690 -1000 8690 -952
rect -8982 -1368 -6982 -1320
rect -8982 -3272 -8934 -1368
rect -7030 -3272 -6982 -1368
rect -8982 -3320 -6982 -3272
rect -6370 -1368 -4370 -1320
rect -6370 -3272 -6322 -1368
rect -4418 -3272 -4370 -1368
rect -6370 -3320 -4370 -3272
rect -3758 -1368 -1758 -1320
rect -3758 -3272 -3710 -1368
rect -1806 -3272 -1758 -1368
rect -3758 -3320 -1758 -3272
rect -1146 -1368 854 -1320
rect -1146 -3272 -1098 -1368
rect 806 -3272 854 -1368
rect -1146 -3320 854 -3272
rect 1466 -1368 3466 -1320
rect 1466 -3272 1514 -1368
rect 3418 -3272 3466 -1368
rect 1466 -3320 3466 -3272
rect 4078 -1368 6078 -1320
rect 4078 -3272 4126 -1368
rect 6030 -3272 6078 -1368
rect 4078 -3320 6078 -3272
rect 6690 -1368 8690 -1320
rect 6690 -3272 6738 -1368
rect 8642 -3272 8690 -1368
rect 6690 -3320 8690 -3272
rect -8982 -3688 -6982 -3640
rect -8982 -5592 -8934 -3688
rect -7030 -5592 -6982 -3688
rect -8982 -5640 -6982 -5592
rect -6370 -3688 -4370 -3640
rect -6370 -5592 -6322 -3688
rect -4418 -5592 -4370 -3688
rect -6370 -5640 -4370 -5592
rect -3758 -3688 -1758 -3640
rect -3758 -5592 -3710 -3688
rect -1806 -5592 -1758 -3688
rect -3758 -5640 -1758 -5592
rect -1146 -3688 854 -3640
rect -1146 -5592 -1098 -3688
rect 806 -5592 854 -3688
rect -1146 -5640 854 -5592
rect 1466 -3688 3466 -3640
rect 1466 -5592 1514 -3688
rect 3418 -5592 3466 -3688
rect 1466 -5640 3466 -5592
rect 4078 -3688 6078 -3640
rect 4078 -5592 4126 -3688
rect 6030 -5592 6078 -3688
rect 4078 -5640 6078 -5592
rect 6690 -3688 8690 -3640
rect 6690 -5592 6738 -3688
rect 8642 -5592 8690 -3688
rect 6690 -5640 8690 -5592
rect -8982 -6008 -6982 -5960
rect -8982 -7912 -8934 -6008
rect -7030 -7912 -6982 -6008
rect -8982 -7960 -6982 -7912
rect -6370 -6008 -4370 -5960
rect -6370 -7912 -6322 -6008
rect -4418 -7912 -4370 -6008
rect -6370 -7960 -4370 -7912
rect -3758 -6008 -1758 -5960
rect -3758 -7912 -3710 -6008
rect -1806 -7912 -1758 -6008
rect -3758 -7960 -1758 -7912
rect -1146 -6008 854 -5960
rect -1146 -7912 -1098 -6008
rect 806 -7912 854 -6008
rect -1146 -7960 854 -7912
rect 1466 -6008 3466 -5960
rect 1466 -7912 1514 -6008
rect 3418 -7912 3466 -6008
rect 1466 -7960 3466 -7912
rect 4078 -6008 6078 -5960
rect 4078 -7912 4126 -6008
rect 6030 -7912 6078 -6008
rect 4078 -7960 6078 -7912
rect 6690 -6008 8690 -5960
rect 6690 -7912 6738 -6008
rect 8642 -7912 8690 -6008
rect 6690 -7960 8690 -7912
<< mimcapcontact >>
rect -8934 6008 -7030 7912
rect -6322 6008 -4418 7912
rect -3710 6008 -1806 7912
rect -1098 6008 806 7912
rect 1514 6008 3418 7912
rect 4126 6008 6030 7912
rect 6738 6008 8642 7912
rect -8934 3688 -7030 5592
rect -6322 3688 -4418 5592
rect -3710 3688 -1806 5592
rect -1098 3688 806 5592
rect 1514 3688 3418 5592
rect 4126 3688 6030 5592
rect 6738 3688 8642 5592
rect -8934 1368 -7030 3272
rect -6322 1368 -4418 3272
rect -3710 1368 -1806 3272
rect -1098 1368 806 3272
rect 1514 1368 3418 3272
rect 4126 1368 6030 3272
rect 6738 1368 8642 3272
rect -8934 -952 -7030 952
rect -6322 -952 -4418 952
rect -3710 -952 -1806 952
rect -1098 -952 806 952
rect 1514 -952 3418 952
rect 4126 -952 6030 952
rect 6738 -952 8642 952
rect -8934 -3272 -7030 -1368
rect -6322 -3272 -4418 -1368
rect -3710 -3272 -1806 -1368
rect -1098 -3272 806 -1368
rect 1514 -3272 3418 -1368
rect 4126 -3272 6030 -1368
rect 6738 -3272 8642 -1368
rect -8934 -5592 -7030 -3688
rect -6322 -5592 -4418 -3688
rect -3710 -5592 -1806 -3688
rect -1098 -5592 806 -3688
rect 1514 -5592 3418 -3688
rect 4126 -5592 6030 -3688
rect 6738 -5592 8642 -3688
rect -8934 -7912 -7030 -6008
rect -6322 -7912 -4418 -6008
rect -3710 -7912 -1806 -6008
rect -1098 -7912 806 -6008
rect 1514 -7912 3418 -6008
rect 4126 -7912 6030 -6008
rect 6738 -7912 8642 -6008
<< metal4 >>
rect -8034 7921 -7930 8120
rect -6754 7952 -6650 8120
rect -8943 7912 -7021 7921
rect -8943 6008 -8934 7912
rect -7030 6008 -7021 7912
rect -8943 5999 -7021 6008
rect -6754 7888 -6734 7952
rect -6670 7888 -6650 7952
rect -5422 7921 -5318 8120
rect -4142 7952 -4038 8120
rect -6754 7872 -6650 7888
rect -6754 7808 -6734 7872
rect -6670 7808 -6650 7872
rect -6754 7792 -6650 7808
rect -6754 7728 -6734 7792
rect -6670 7728 -6650 7792
rect -6754 7712 -6650 7728
rect -6754 7648 -6734 7712
rect -6670 7648 -6650 7712
rect -6754 7632 -6650 7648
rect -6754 7568 -6734 7632
rect -6670 7568 -6650 7632
rect -6754 7552 -6650 7568
rect -6754 7488 -6734 7552
rect -6670 7488 -6650 7552
rect -6754 7472 -6650 7488
rect -6754 7408 -6734 7472
rect -6670 7408 -6650 7472
rect -6754 7392 -6650 7408
rect -6754 7328 -6734 7392
rect -6670 7328 -6650 7392
rect -6754 7312 -6650 7328
rect -6754 7248 -6734 7312
rect -6670 7248 -6650 7312
rect -6754 7232 -6650 7248
rect -6754 7168 -6734 7232
rect -6670 7168 -6650 7232
rect -6754 7152 -6650 7168
rect -6754 7088 -6734 7152
rect -6670 7088 -6650 7152
rect -6754 7072 -6650 7088
rect -6754 7008 -6734 7072
rect -6670 7008 -6650 7072
rect -6754 6992 -6650 7008
rect -6754 6928 -6734 6992
rect -6670 6928 -6650 6992
rect -6754 6912 -6650 6928
rect -6754 6848 -6734 6912
rect -6670 6848 -6650 6912
rect -6754 6832 -6650 6848
rect -6754 6768 -6734 6832
rect -6670 6768 -6650 6832
rect -6754 6752 -6650 6768
rect -6754 6688 -6734 6752
rect -6670 6688 -6650 6752
rect -6754 6672 -6650 6688
rect -6754 6608 -6734 6672
rect -6670 6608 -6650 6672
rect -6754 6592 -6650 6608
rect -6754 6528 -6734 6592
rect -6670 6528 -6650 6592
rect -6754 6512 -6650 6528
rect -6754 6448 -6734 6512
rect -6670 6448 -6650 6512
rect -6754 6432 -6650 6448
rect -6754 6368 -6734 6432
rect -6670 6368 -6650 6432
rect -6754 6352 -6650 6368
rect -6754 6288 -6734 6352
rect -6670 6288 -6650 6352
rect -6754 6272 -6650 6288
rect -6754 6208 -6734 6272
rect -6670 6208 -6650 6272
rect -6754 6192 -6650 6208
rect -6754 6128 -6734 6192
rect -6670 6128 -6650 6192
rect -6754 6112 -6650 6128
rect -6754 6048 -6734 6112
rect -6670 6048 -6650 6112
rect -6754 6032 -6650 6048
rect -8034 5601 -7930 5999
rect -6754 5968 -6734 6032
rect -6670 5968 -6650 6032
rect -6331 7912 -4409 7921
rect -6331 6008 -6322 7912
rect -4418 6008 -4409 7912
rect -6331 5999 -4409 6008
rect -4142 7888 -4122 7952
rect -4058 7888 -4038 7952
rect -2810 7921 -2706 8120
rect -1530 7952 -1426 8120
rect -4142 7872 -4038 7888
rect -4142 7808 -4122 7872
rect -4058 7808 -4038 7872
rect -4142 7792 -4038 7808
rect -4142 7728 -4122 7792
rect -4058 7728 -4038 7792
rect -4142 7712 -4038 7728
rect -4142 7648 -4122 7712
rect -4058 7648 -4038 7712
rect -4142 7632 -4038 7648
rect -4142 7568 -4122 7632
rect -4058 7568 -4038 7632
rect -4142 7552 -4038 7568
rect -4142 7488 -4122 7552
rect -4058 7488 -4038 7552
rect -4142 7472 -4038 7488
rect -4142 7408 -4122 7472
rect -4058 7408 -4038 7472
rect -4142 7392 -4038 7408
rect -4142 7328 -4122 7392
rect -4058 7328 -4038 7392
rect -4142 7312 -4038 7328
rect -4142 7248 -4122 7312
rect -4058 7248 -4038 7312
rect -4142 7232 -4038 7248
rect -4142 7168 -4122 7232
rect -4058 7168 -4038 7232
rect -4142 7152 -4038 7168
rect -4142 7088 -4122 7152
rect -4058 7088 -4038 7152
rect -4142 7072 -4038 7088
rect -4142 7008 -4122 7072
rect -4058 7008 -4038 7072
rect -4142 6992 -4038 7008
rect -4142 6928 -4122 6992
rect -4058 6928 -4038 6992
rect -4142 6912 -4038 6928
rect -4142 6848 -4122 6912
rect -4058 6848 -4038 6912
rect -4142 6832 -4038 6848
rect -4142 6768 -4122 6832
rect -4058 6768 -4038 6832
rect -4142 6752 -4038 6768
rect -4142 6688 -4122 6752
rect -4058 6688 -4038 6752
rect -4142 6672 -4038 6688
rect -4142 6608 -4122 6672
rect -4058 6608 -4038 6672
rect -4142 6592 -4038 6608
rect -4142 6528 -4122 6592
rect -4058 6528 -4038 6592
rect -4142 6512 -4038 6528
rect -4142 6448 -4122 6512
rect -4058 6448 -4038 6512
rect -4142 6432 -4038 6448
rect -4142 6368 -4122 6432
rect -4058 6368 -4038 6432
rect -4142 6352 -4038 6368
rect -4142 6288 -4122 6352
rect -4058 6288 -4038 6352
rect -4142 6272 -4038 6288
rect -4142 6208 -4122 6272
rect -4058 6208 -4038 6272
rect -4142 6192 -4038 6208
rect -4142 6128 -4122 6192
rect -4058 6128 -4038 6192
rect -4142 6112 -4038 6128
rect -4142 6048 -4122 6112
rect -4058 6048 -4038 6112
rect -4142 6032 -4038 6048
rect -6754 5632 -6650 5968
rect -8943 5592 -7021 5601
rect -8943 3688 -8934 5592
rect -7030 3688 -7021 5592
rect -8943 3679 -7021 3688
rect -6754 5568 -6734 5632
rect -6670 5568 -6650 5632
rect -5422 5601 -5318 5999
rect -4142 5968 -4122 6032
rect -4058 5968 -4038 6032
rect -3719 7912 -1797 7921
rect -3719 6008 -3710 7912
rect -1806 6008 -1797 7912
rect -3719 5999 -1797 6008
rect -1530 7888 -1510 7952
rect -1446 7888 -1426 7952
rect -198 7921 -94 8120
rect 1082 7952 1186 8120
rect -1530 7872 -1426 7888
rect -1530 7808 -1510 7872
rect -1446 7808 -1426 7872
rect -1530 7792 -1426 7808
rect -1530 7728 -1510 7792
rect -1446 7728 -1426 7792
rect -1530 7712 -1426 7728
rect -1530 7648 -1510 7712
rect -1446 7648 -1426 7712
rect -1530 7632 -1426 7648
rect -1530 7568 -1510 7632
rect -1446 7568 -1426 7632
rect -1530 7552 -1426 7568
rect -1530 7488 -1510 7552
rect -1446 7488 -1426 7552
rect -1530 7472 -1426 7488
rect -1530 7408 -1510 7472
rect -1446 7408 -1426 7472
rect -1530 7392 -1426 7408
rect -1530 7328 -1510 7392
rect -1446 7328 -1426 7392
rect -1530 7312 -1426 7328
rect -1530 7248 -1510 7312
rect -1446 7248 -1426 7312
rect -1530 7232 -1426 7248
rect -1530 7168 -1510 7232
rect -1446 7168 -1426 7232
rect -1530 7152 -1426 7168
rect -1530 7088 -1510 7152
rect -1446 7088 -1426 7152
rect -1530 7072 -1426 7088
rect -1530 7008 -1510 7072
rect -1446 7008 -1426 7072
rect -1530 6992 -1426 7008
rect -1530 6928 -1510 6992
rect -1446 6928 -1426 6992
rect -1530 6912 -1426 6928
rect -1530 6848 -1510 6912
rect -1446 6848 -1426 6912
rect -1530 6832 -1426 6848
rect -1530 6768 -1510 6832
rect -1446 6768 -1426 6832
rect -1530 6752 -1426 6768
rect -1530 6688 -1510 6752
rect -1446 6688 -1426 6752
rect -1530 6672 -1426 6688
rect -1530 6608 -1510 6672
rect -1446 6608 -1426 6672
rect -1530 6592 -1426 6608
rect -1530 6528 -1510 6592
rect -1446 6528 -1426 6592
rect -1530 6512 -1426 6528
rect -1530 6448 -1510 6512
rect -1446 6448 -1426 6512
rect -1530 6432 -1426 6448
rect -1530 6368 -1510 6432
rect -1446 6368 -1426 6432
rect -1530 6352 -1426 6368
rect -1530 6288 -1510 6352
rect -1446 6288 -1426 6352
rect -1530 6272 -1426 6288
rect -1530 6208 -1510 6272
rect -1446 6208 -1426 6272
rect -1530 6192 -1426 6208
rect -1530 6128 -1510 6192
rect -1446 6128 -1426 6192
rect -1530 6112 -1426 6128
rect -1530 6048 -1510 6112
rect -1446 6048 -1426 6112
rect -1530 6032 -1426 6048
rect -4142 5632 -4038 5968
rect -6754 5552 -6650 5568
rect -6754 5488 -6734 5552
rect -6670 5488 -6650 5552
rect -6754 5472 -6650 5488
rect -6754 5408 -6734 5472
rect -6670 5408 -6650 5472
rect -6754 5392 -6650 5408
rect -6754 5328 -6734 5392
rect -6670 5328 -6650 5392
rect -6754 5312 -6650 5328
rect -6754 5248 -6734 5312
rect -6670 5248 -6650 5312
rect -6754 5232 -6650 5248
rect -6754 5168 -6734 5232
rect -6670 5168 -6650 5232
rect -6754 5152 -6650 5168
rect -6754 5088 -6734 5152
rect -6670 5088 -6650 5152
rect -6754 5072 -6650 5088
rect -6754 5008 -6734 5072
rect -6670 5008 -6650 5072
rect -6754 4992 -6650 5008
rect -6754 4928 -6734 4992
rect -6670 4928 -6650 4992
rect -6754 4912 -6650 4928
rect -6754 4848 -6734 4912
rect -6670 4848 -6650 4912
rect -6754 4832 -6650 4848
rect -6754 4768 -6734 4832
rect -6670 4768 -6650 4832
rect -6754 4752 -6650 4768
rect -6754 4688 -6734 4752
rect -6670 4688 -6650 4752
rect -6754 4672 -6650 4688
rect -6754 4608 -6734 4672
rect -6670 4608 -6650 4672
rect -6754 4592 -6650 4608
rect -6754 4528 -6734 4592
rect -6670 4528 -6650 4592
rect -6754 4512 -6650 4528
rect -6754 4448 -6734 4512
rect -6670 4448 -6650 4512
rect -6754 4432 -6650 4448
rect -6754 4368 -6734 4432
rect -6670 4368 -6650 4432
rect -6754 4352 -6650 4368
rect -6754 4288 -6734 4352
rect -6670 4288 -6650 4352
rect -6754 4272 -6650 4288
rect -6754 4208 -6734 4272
rect -6670 4208 -6650 4272
rect -6754 4192 -6650 4208
rect -6754 4128 -6734 4192
rect -6670 4128 -6650 4192
rect -6754 4112 -6650 4128
rect -6754 4048 -6734 4112
rect -6670 4048 -6650 4112
rect -6754 4032 -6650 4048
rect -6754 3968 -6734 4032
rect -6670 3968 -6650 4032
rect -6754 3952 -6650 3968
rect -6754 3888 -6734 3952
rect -6670 3888 -6650 3952
rect -6754 3872 -6650 3888
rect -6754 3808 -6734 3872
rect -6670 3808 -6650 3872
rect -6754 3792 -6650 3808
rect -6754 3728 -6734 3792
rect -6670 3728 -6650 3792
rect -6754 3712 -6650 3728
rect -8034 3281 -7930 3679
rect -6754 3648 -6734 3712
rect -6670 3648 -6650 3712
rect -6331 5592 -4409 5601
rect -6331 3688 -6322 5592
rect -4418 3688 -4409 5592
rect -6331 3679 -4409 3688
rect -4142 5568 -4122 5632
rect -4058 5568 -4038 5632
rect -2810 5601 -2706 5999
rect -1530 5968 -1510 6032
rect -1446 5968 -1426 6032
rect -1107 7912 815 7921
rect -1107 6008 -1098 7912
rect 806 6008 815 7912
rect -1107 5999 815 6008
rect 1082 7888 1102 7952
rect 1166 7888 1186 7952
rect 2414 7921 2518 8120
rect 3694 7952 3798 8120
rect 1082 7872 1186 7888
rect 1082 7808 1102 7872
rect 1166 7808 1186 7872
rect 1082 7792 1186 7808
rect 1082 7728 1102 7792
rect 1166 7728 1186 7792
rect 1082 7712 1186 7728
rect 1082 7648 1102 7712
rect 1166 7648 1186 7712
rect 1082 7632 1186 7648
rect 1082 7568 1102 7632
rect 1166 7568 1186 7632
rect 1082 7552 1186 7568
rect 1082 7488 1102 7552
rect 1166 7488 1186 7552
rect 1082 7472 1186 7488
rect 1082 7408 1102 7472
rect 1166 7408 1186 7472
rect 1082 7392 1186 7408
rect 1082 7328 1102 7392
rect 1166 7328 1186 7392
rect 1082 7312 1186 7328
rect 1082 7248 1102 7312
rect 1166 7248 1186 7312
rect 1082 7232 1186 7248
rect 1082 7168 1102 7232
rect 1166 7168 1186 7232
rect 1082 7152 1186 7168
rect 1082 7088 1102 7152
rect 1166 7088 1186 7152
rect 1082 7072 1186 7088
rect 1082 7008 1102 7072
rect 1166 7008 1186 7072
rect 1082 6992 1186 7008
rect 1082 6928 1102 6992
rect 1166 6928 1186 6992
rect 1082 6912 1186 6928
rect 1082 6848 1102 6912
rect 1166 6848 1186 6912
rect 1082 6832 1186 6848
rect 1082 6768 1102 6832
rect 1166 6768 1186 6832
rect 1082 6752 1186 6768
rect 1082 6688 1102 6752
rect 1166 6688 1186 6752
rect 1082 6672 1186 6688
rect 1082 6608 1102 6672
rect 1166 6608 1186 6672
rect 1082 6592 1186 6608
rect 1082 6528 1102 6592
rect 1166 6528 1186 6592
rect 1082 6512 1186 6528
rect 1082 6448 1102 6512
rect 1166 6448 1186 6512
rect 1082 6432 1186 6448
rect 1082 6368 1102 6432
rect 1166 6368 1186 6432
rect 1082 6352 1186 6368
rect 1082 6288 1102 6352
rect 1166 6288 1186 6352
rect 1082 6272 1186 6288
rect 1082 6208 1102 6272
rect 1166 6208 1186 6272
rect 1082 6192 1186 6208
rect 1082 6128 1102 6192
rect 1166 6128 1186 6192
rect 1082 6112 1186 6128
rect 1082 6048 1102 6112
rect 1166 6048 1186 6112
rect 1082 6032 1186 6048
rect -1530 5632 -1426 5968
rect -4142 5552 -4038 5568
rect -4142 5488 -4122 5552
rect -4058 5488 -4038 5552
rect -4142 5472 -4038 5488
rect -4142 5408 -4122 5472
rect -4058 5408 -4038 5472
rect -4142 5392 -4038 5408
rect -4142 5328 -4122 5392
rect -4058 5328 -4038 5392
rect -4142 5312 -4038 5328
rect -4142 5248 -4122 5312
rect -4058 5248 -4038 5312
rect -4142 5232 -4038 5248
rect -4142 5168 -4122 5232
rect -4058 5168 -4038 5232
rect -4142 5152 -4038 5168
rect -4142 5088 -4122 5152
rect -4058 5088 -4038 5152
rect -4142 5072 -4038 5088
rect -4142 5008 -4122 5072
rect -4058 5008 -4038 5072
rect -4142 4992 -4038 5008
rect -4142 4928 -4122 4992
rect -4058 4928 -4038 4992
rect -4142 4912 -4038 4928
rect -4142 4848 -4122 4912
rect -4058 4848 -4038 4912
rect -4142 4832 -4038 4848
rect -4142 4768 -4122 4832
rect -4058 4768 -4038 4832
rect -4142 4752 -4038 4768
rect -4142 4688 -4122 4752
rect -4058 4688 -4038 4752
rect -4142 4672 -4038 4688
rect -4142 4608 -4122 4672
rect -4058 4608 -4038 4672
rect -4142 4592 -4038 4608
rect -4142 4528 -4122 4592
rect -4058 4528 -4038 4592
rect -4142 4512 -4038 4528
rect -4142 4448 -4122 4512
rect -4058 4448 -4038 4512
rect -4142 4432 -4038 4448
rect -4142 4368 -4122 4432
rect -4058 4368 -4038 4432
rect -4142 4352 -4038 4368
rect -4142 4288 -4122 4352
rect -4058 4288 -4038 4352
rect -4142 4272 -4038 4288
rect -4142 4208 -4122 4272
rect -4058 4208 -4038 4272
rect -4142 4192 -4038 4208
rect -4142 4128 -4122 4192
rect -4058 4128 -4038 4192
rect -4142 4112 -4038 4128
rect -4142 4048 -4122 4112
rect -4058 4048 -4038 4112
rect -4142 4032 -4038 4048
rect -4142 3968 -4122 4032
rect -4058 3968 -4038 4032
rect -4142 3952 -4038 3968
rect -4142 3888 -4122 3952
rect -4058 3888 -4038 3952
rect -4142 3872 -4038 3888
rect -4142 3808 -4122 3872
rect -4058 3808 -4038 3872
rect -4142 3792 -4038 3808
rect -4142 3728 -4122 3792
rect -4058 3728 -4038 3792
rect -4142 3712 -4038 3728
rect -6754 3312 -6650 3648
rect -8943 3272 -7021 3281
rect -8943 1368 -8934 3272
rect -7030 1368 -7021 3272
rect -8943 1359 -7021 1368
rect -6754 3248 -6734 3312
rect -6670 3248 -6650 3312
rect -5422 3281 -5318 3679
rect -4142 3648 -4122 3712
rect -4058 3648 -4038 3712
rect -3719 5592 -1797 5601
rect -3719 3688 -3710 5592
rect -1806 3688 -1797 5592
rect -3719 3679 -1797 3688
rect -1530 5568 -1510 5632
rect -1446 5568 -1426 5632
rect -198 5601 -94 5999
rect 1082 5968 1102 6032
rect 1166 5968 1186 6032
rect 1505 7912 3427 7921
rect 1505 6008 1514 7912
rect 3418 6008 3427 7912
rect 1505 5999 3427 6008
rect 3694 7888 3714 7952
rect 3778 7888 3798 7952
rect 5026 7921 5130 8120
rect 6306 7952 6410 8120
rect 3694 7872 3798 7888
rect 3694 7808 3714 7872
rect 3778 7808 3798 7872
rect 3694 7792 3798 7808
rect 3694 7728 3714 7792
rect 3778 7728 3798 7792
rect 3694 7712 3798 7728
rect 3694 7648 3714 7712
rect 3778 7648 3798 7712
rect 3694 7632 3798 7648
rect 3694 7568 3714 7632
rect 3778 7568 3798 7632
rect 3694 7552 3798 7568
rect 3694 7488 3714 7552
rect 3778 7488 3798 7552
rect 3694 7472 3798 7488
rect 3694 7408 3714 7472
rect 3778 7408 3798 7472
rect 3694 7392 3798 7408
rect 3694 7328 3714 7392
rect 3778 7328 3798 7392
rect 3694 7312 3798 7328
rect 3694 7248 3714 7312
rect 3778 7248 3798 7312
rect 3694 7232 3798 7248
rect 3694 7168 3714 7232
rect 3778 7168 3798 7232
rect 3694 7152 3798 7168
rect 3694 7088 3714 7152
rect 3778 7088 3798 7152
rect 3694 7072 3798 7088
rect 3694 7008 3714 7072
rect 3778 7008 3798 7072
rect 3694 6992 3798 7008
rect 3694 6928 3714 6992
rect 3778 6928 3798 6992
rect 3694 6912 3798 6928
rect 3694 6848 3714 6912
rect 3778 6848 3798 6912
rect 3694 6832 3798 6848
rect 3694 6768 3714 6832
rect 3778 6768 3798 6832
rect 3694 6752 3798 6768
rect 3694 6688 3714 6752
rect 3778 6688 3798 6752
rect 3694 6672 3798 6688
rect 3694 6608 3714 6672
rect 3778 6608 3798 6672
rect 3694 6592 3798 6608
rect 3694 6528 3714 6592
rect 3778 6528 3798 6592
rect 3694 6512 3798 6528
rect 3694 6448 3714 6512
rect 3778 6448 3798 6512
rect 3694 6432 3798 6448
rect 3694 6368 3714 6432
rect 3778 6368 3798 6432
rect 3694 6352 3798 6368
rect 3694 6288 3714 6352
rect 3778 6288 3798 6352
rect 3694 6272 3798 6288
rect 3694 6208 3714 6272
rect 3778 6208 3798 6272
rect 3694 6192 3798 6208
rect 3694 6128 3714 6192
rect 3778 6128 3798 6192
rect 3694 6112 3798 6128
rect 3694 6048 3714 6112
rect 3778 6048 3798 6112
rect 3694 6032 3798 6048
rect 1082 5632 1186 5968
rect -1530 5552 -1426 5568
rect -1530 5488 -1510 5552
rect -1446 5488 -1426 5552
rect -1530 5472 -1426 5488
rect -1530 5408 -1510 5472
rect -1446 5408 -1426 5472
rect -1530 5392 -1426 5408
rect -1530 5328 -1510 5392
rect -1446 5328 -1426 5392
rect -1530 5312 -1426 5328
rect -1530 5248 -1510 5312
rect -1446 5248 -1426 5312
rect -1530 5232 -1426 5248
rect -1530 5168 -1510 5232
rect -1446 5168 -1426 5232
rect -1530 5152 -1426 5168
rect -1530 5088 -1510 5152
rect -1446 5088 -1426 5152
rect -1530 5072 -1426 5088
rect -1530 5008 -1510 5072
rect -1446 5008 -1426 5072
rect -1530 4992 -1426 5008
rect -1530 4928 -1510 4992
rect -1446 4928 -1426 4992
rect -1530 4912 -1426 4928
rect -1530 4848 -1510 4912
rect -1446 4848 -1426 4912
rect -1530 4832 -1426 4848
rect -1530 4768 -1510 4832
rect -1446 4768 -1426 4832
rect -1530 4752 -1426 4768
rect -1530 4688 -1510 4752
rect -1446 4688 -1426 4752
rect -1530 4672 -1426 4688
rect -1530 4608 -1510 4672
rect -1446 4608 -1426 4672
rect -1530 4592 -1426 4608
rect -1530 4528 -1510 4592
rect -1446 4528 -1426 4592
rect -1530 4512 -1426 4528
rect -1530 4448 -1510 4512
rect -1446 4448 -1426 4512
rect -1530 4432 -1426 4448
rect -1530 4368 -1510 4432
rect -1446 4368 -1426 4432
rect -1530 4352 -1426 4368
rect -1530 4288 -1510 4352
rect -1446 4288 -1426 4352
rect -1530 4272 -1426 4288
rect -1530 4208 -1510 4272
rect -1446 4208 -1426 4272
rect -1530 4192 -1426 4208
rect -1530 4128 -1510 4192
rect -1446 4128 -1426 4192
rect -1530 4112 -1426 4128
rect -1530 4048 -1510 4112
rect -1446 4048 -1426 4112
rect -1530 4032 -1426 4048
rect -1530 3968 -1510 4032
rect -1446 3968 -1426 4032
rect -1530 3952 -1426 3968
rect -1530 3888 -1510 3952
rect -1446 3888 -1426 3952
rect -1530 3872 -1426 3888
rect -1530 3808 -1510 3872
rect -1446 3808 -1426 3872
rect -1530 3792 -1426 3808
rect -1530 3728 -1510 3792
rect -1446 3728 -1426 3792
rect -1530 3712 -1426 3728
rect -4142 3312 -4038 3648
rect -6754 3232 -6650 3248
rect -6754 3168 -6734 3232
rect -6670 3168 -6650 3232
rect -6754 3152 -6650 3168
rect -6754 3088 -6734 3152
rect -6670 3088 -6650 3152
rect -6754 3072 -6650 3088
rect -6754 3008 -6734 3072
rect -6670 3008 -6650 3072
rect -6754 2992 -6650 3008
rect -6754 2928 -6734 2992
rect -6670 2928 -6650 2992
rect -6754 2912 -6650 2928
rect -6754 2848 -6734 2912
rect -6670 2848 -6650 2912
rect -6754 2832 -6650 2848
rect -6754 2768 -6734 2832
rect -6670 2768 -6650 2832
rect -6754 2752 -6650 2768
rect -6754 2688 -6734 2752
rect -6670 2688 -6650 2752
rect -6754 2672 -6650 2688
rect -6754 2608 -6734 2672
rect -6670 2608 -6650 2672
rect -6754 2592 -6650 2608
rect -6754 2528 -6734 2592
rect -6670 2528 -6650 2592
rect -6754 2512 -6650 2528
rect -6754 2448 -6734 2512
rect -6670 2448 -6650 2512
rect -6754 2432 -6650 2448
rect -6754 2368 -6734 2432
rect -6670 2368 -6650 2432
rect -6754 2352 -6650 2368
rect -6754 2288 -6734 2352
rect -6670 2288 -6650 2352
rect -6754 2272 -6650 2288
rect -6754 2208 -6734 2272
rect -6670 2208 -6650 2272
rect -6754 2192 -6650 2208
rect -6754 2128 -6734 2192
rect -6670 2128 -6650 2192
rect -6754 2112 -6650 2128
rect -6754 2048 -6734 2112
rect -6670 2048 -6650 2112
rect -6754 2032 -6650 2048
rect -6754 1968 -6734 2032
rect -6670 1968 -6650 2032
rect -6754 1952 -6650 1968
rect -6754 1888 -6734 1952
rect -6670 1888 -6650 1952
rect -6754 1872 -6650 1888
rect -6754 1808 -6734 1872
rect -6670 1808 -6650 1872
rect -6754 1792 -6650 1808
rect -6754 1728 -6734 1792
rect -6670 1728 -6650 1792
rect -6754 1712 -6650 1728
rect -6754 1648 -6734 1712
rect -6670 1648 -6650 1712
rect -6754 1632 -6650 1648
rect -6754 1568 -6734 1632
rect -6670 1568 -6650 1632
rect -6754 1552 -6650 1568
rect -6754 1488 -6734 1552
rect -6670 1488 -6650 1552
rect -6754 1472 -6650 1488
rect -6754 1408 -6734 1472
rect -6670 1408 -6650 1472
rect -6754 1392 -6650 1408
rect -8034 961 -7930 1359
rect -6754 1328 -6734 1392
rect -6670 1328 -6650 1392
rect -6331 3272 -4409 3281
rect -6331 1368 -6322 3272
rect -4418 1368 -4409 3272
rect -6331 1359 -4409 1368
rect -4142 3248 -4122 3312
rect -4058 3248 -4038 3312
rect -2810 3281 -2706 3679
rect -1530 3648 -1510 3712
rect -1446 3648 -1426 3712
rect -1107 5592 815 5601
rect -1107 3688 -1098 5592
rect 806 3688 815 5592
rect -1107 3679 815 3688
rect 1082 5568 1102 5632
rect 1166 5568 1186 5632
rect 2414 5601 2518 5999
rect 3694 5968 3714 6032
rect 3778 5968 3798 6032
rect 4117 7912 6039 7921
rect 4117 6008 4126 7912
rect 6030 6008 6039 7912
rect 4117 5999 6039 6008
rect 6306 7888 6326 7952
rect 6390 7888 6410 7952
rect 7638 7921 7742 8120
rect 8918 7952 9022 8120
rect 6306 7872 6410 7888
rect 6306 7808 6326 7872
rect 6390 7808 6410 7872
rect 6306 7792 6410 7808
rect 6306 7728 6326 7792
rect 6390 7728 6410 7792
rect 6306 7712 6410 7728
rect 6306 7648 6326 7712
rect 6390 7648 6410 7712
rect 6306 7632 6410 7648
rect 6306 7568 6326 7632
rect 6390 7568 6410 7632
rect 6306 7552 6410 7568
rect 6306 7488 6326 7552
rect 6390 7488 6410 7552
rect 6306 7472 6410 7488
rect 6306 7408 6326 7472
rect 6390 7408 6410 7472
rect 6306 7392 6410 7408
rect 6306 7328 6326 7392
rect 6390 7328 6410 7392
rect 6306 7312 6410 7328
rect 6306 7248 6326 7312
rect 6390 7248 6410 7312
rect 6306 7232 6410 7248
rect 6306 7168 6326 7232
rect 6390 7168 6410 7232
rect 6306 7152 6410 7168
rect 6306 7088 6326 7152
rect 6390 7088 6410 7152
rect 6306 7072 6410 7088
rect 6306 7008 6326 7072
rect 6390 7008 6410 7072
rect 6306 6992 6410 7008
rect 6306 6928 6326 6992
rect 6390 6928 6410 6992
rect 6306 6912 6410 6928
rect 6306 6848 6326 6912
rect 6390 6848 6410 6912
rect 6306 6832 6410 6848
rect 6306 6768 6326 6832
rect 6390 6768 6410 6832
rect 6306 6752 6410 6768
rect 6306 6688 6326 6752
rect 6390 6688 6410 6752
rect 6306 6672 6410 6688
rect 6306 6608 6326 6672
rect 6390 6608 6410 6672
rect 6306 6592 6410 6608
rect 6306 6528 6326 6592
rect 6390 6528 6410 6592
rect 6306 6512 6410 6528
rect 6306 6448 6326 6512
rect 6390 6448 6410 6512
rect 6306 6432 6410 6448
rect 6306 6368 6326 6432
rect 6390 6368 6410 6432
rect 6306 6352 6410 6368
rect 6306 6288 6326 6352
rect 6390 6288 6410 6352
rect 6306 6272 6410 6288
rect 6306 6208 6326 6272
rect 6390 6208 6410 6272
rect 6306 6192 6410 6208
rect 6306 6128 6326 6192
rect 6390 6128 6410 6192
rect 6306 6112 6410 6128
rect 6306 6048 6326 6112
rect 6390 6048 6410 6112
rect 6306 6032 6410 6048
rect 3694 5632 3798 5968
rect 1082 5552 1186 5568
rect 1082 5488 1102 5552
rect 1166 5488 1186 5552
rect 1082 5472 1186 5488
rect 1082 5408 1102 5472
rect 1166 5408 1186 5472
rect 1082 5392 1186 5408
rect 1082 5328 1102 5392
rect 1166 5328 1186 5392
rect 1082 5312 1186 5328
rect 1082 5248 1102 5312
rect 1166 5248 1186 5312
rect 1082 5232 1186 5248
rect 1082 5168 1102 5232
rect 1166 5168 1186 5232
rect 1082 5152 1186 5168
rect 1082 5088 1102 5152
rect 1166 5088 1186 5152
rect 1082 5072 1186 5088
rect 1082 5008 1102 5072
rect 1166 5008 1186 5072
rect 1082 4992 1186 5008
rect 1082 4928 1102 4992
rect 1166 4928 1186 4992
rect 1082 4912 1186 4928
rect 1082 4848 1102 4912
rect 1166 4848 1186 4912
rect 1082 4832 1186 4848
rect 1082 4768 1102 4832
rect 1166 4768 1186 4832
rect 1082 4752 1186 4768
rect 1082 4688 1102 4752
rect 1166 4688 1186 4752
rect 1082 4672 1186 4688
rect 1082 4608 1102 4672
rect 1166 4608 1186 4672
rect 1082 4592 1186 4608
rect 1082 4528 1102 4592
rect 1166 4528 1186 4592
rect 1082 4512 1186 4528
rect 1082 4448 1102 4512
rect 1166 4448 1186 4512
rect 1082 4432 1186 4448
rect 1082 4368 1102 4432
rect 1166 4368 1186 4432
rect 1082 4352 1186 4368
rect 1082 4288 1102 4352
rect 1166 4288 1186 4352
rect 1082 4272 1186 4288
rect 1082 4208 1102 4272
rect 1166 4208 1186 4272
rect 1082 4192 1186 4208
rect 1082 4128 1102 4192
rect 1166 4128 1186 4192
rect 1082 4112 1186 4128
rect 1082 4048 1102 4112
rect 1166 4048 1186 4112
rect 1082 4032 1186 4048
rect 1082 3968 1102 4032
rect 1166 3968 1186 4032
rect 1082 3952 1186 3968
rect 1082 3888 1102 3952
rect 1166 3888 1186 3952
rect 1082 3872 1186 3888
rect 1082 3808 1102 3872
rect 1166 3808 1186 3872
rect 1082 3792 1186 3808
rect 1082 3728 1102 3792
rect 1166 3728 1186 3792
rect 1082 3712 1186 3728
rect -1530 3312 -1426 3648
rect -4142 3232 -4038 3248
rect -4142 3168 -4122 3232
rect -4058 3168 -4038 3232
rect -4142 3152 -4038 3168
rect -4142 3088 -4122 3152
rect -4058 3088 -4038 3152
rect -4142 3072 -4038 3088
rect -4142 3008 -4122 3072
rect -4058 3008 -4038 3072
rect -4142 2992 -4038 3008
rect -4142 2928 -4122 2992
rect -4058 2928 -4038 2992
rect -4142 2912 -4038 2928
rect -4142 2848 -4122 2912
rect -4058 2848 -4038 2912
rect -4142 2832 -4038 2848
rect -4142 2768 -4122 2832
rect -4058 2768 -4038 2832
rect -4142 2752 -4038 2768
rect -4142 2688 -4122 2752
rect -4058 2688 -4038 2752
rect -4142 2672 -4038 2688
rect -4142 2608 -4122 2672
rect -4058 2608 -4038 2672
rect -4142 2592 -4038 2608
rect -4142 2528 -4122 2592
rect -4058 2528 -4038 2592
rect -4142 2512 -4038 2528
rect -4142 2448 -4122 2512
rect -4058 2448 -4038 2512
rect -4142 2432 -4038 2448
rect -4142 2368 -4122 2432
rect -4058 2368 -4038 2432
rect -4142 2352 -4038 2368
rect -4142 2288 -4122 2352
rect -4058 2288 -4038 2352
rect -4142 2272 -4038 2288
rect -4142 2208 -4122 2272
rect -4058 2208 -4038 2272
rect -4142 2192 -4038 2208
rect -4142 2128 -4122 2192
rect -4058 2128 -4038 2192
rect -4142 2112 -4038 2128
rect -4142 2048 -4122 2112
rect -4058 2048 -4038 2112
rect -4142 2032 -4038 2048
rect -4142 1968 -4122 2032
rect -4058 1968 -4038 2032
rect -4142 1952 -4038 1968
rect -4142 1888 -4122 1952
rect -4058 1888 -4038 1952
rect -4142 1872 -4038 1888
rect -4142 1808 -4122 1872
rect -4058 1808 -4038 1872
rect -4142 1792 -4038 1808
rect -4142 1728 -4122 1792
rect -4058 1728 -4038 1792
rect -4142 1712 -4038 1728
rect -4142 1648 -4122 1712
rect -4058 1648 -4038 1712
rect -4142 1632 -4038 1648
rect -4142 1568 -4122 1632
rect -4058 1568 -4038 1632
rect -4142 1552 -4038 1568
rect -4142 1488 -4122 1552
rect -4058 1488 -4038 1552
rect -4142 1472 -4038 1488
rect -4142 1408 -4122 1472
rect -4058 1408 -4038 1472
rect -4142 1392 -4038 1408
rect -6754 992 -6650 1328
rect -8943 952 -7021 961
rect -8943 -952 -8934 952
rect -7030 -952 -7021 952
rect -8943 -961 -7021 -952
rect -6754 928 -6734 992
rect -6670 928 -6650 992
rect -5422 961 -5318 1359
rect -4142 1328 -4122 1392
rect -4058 1328 -4038 1392
rect -3719 3272 -1797 3281
rect -3719 1368 -3710 3272
rect -1806 1368 -1797 3272
rect -3719 1359 -1797 1368
rect -1530 3248 -1510 3312
rect -1446 3248 -1426 3312
rect -198 3281 -94 3679
rect 1082 3648 1102 3712
rect 1166 3648 1186 3712
rect 1505 5592 3427 5601
rect 1505 3688 1514 5592
rect 3418 3688 3427 5592
rect 1505 3679 3427 3688
rect 3694 5568 3714 5632
rect 3778 5568 3798 5632
rect 5026 5601 5130 5999
rect 6306 5968 6326 6032
rect 6390 5968 6410 6032
rect 6729 7912 8651 7921
rect 6729 6008 6738 7912
rect 8642 6008 8651 7912
rect 6729 5999 8651 6008
rect 8918 7888 8938 7952
rect 9002 7888 9022 7952
rect 8918 7872 9022 7888
rect 8918 7808 8938 7872
rect 9002 7808 9022 7872
rect 8918 7792 9022 7808
rect 8918 7728 8938 7792
rect 9002 7728 9022 7792
rect 8918 7712 9022 7728
rect 8918 7648 8938 7712
rect 9002 7648 9022 7712
rect 8918 7632 9022 7648
rect 8918 7568 8938 7632
rect 9002 7568 9022 7632
rect 8918 7552 9022 7568
rect 8918 7488 8938 7552
rect 9002 7488 9022 7552
rect 8918 7472 9022 7488
rect 8918 7408 8938 7472
rect 9002 7408 9022 7472
rect 8918 7392 9022 7408
rect 8918 7328 8938 7392
rect 9002 7328 9022 7392
rect 8918 7312 9022 7328
rect 8918 7248 8938 7312
rect 9002 7248 9022 7312
rect 8918 7232 9022 7248
rect 8918 7168 8938 7232
rect 9002 7168 9022 7232
rect 8918 7152 9022 7168
rect 8918 7088 8938 7152
rect 9002 7088 9022 7152
rect 8918 7072 9022 7088
rect 8918 7008 8938 7072
rect 9002 7008 9022 7072
rect 8918 6992 9022 7008
rect 8918 6928 8938 6992
rect 9002 6928 9022 6992
rect 8918 6912 9022 6928
rect 8918 6848 8938 6912
rect 9002 6848 9022 6912
rect 8918 6832 9022 6848
rect 8918 6768 8938 6832
rect 9002 6768 9022 6832
rect 8918 6752 9022 6768
rect 8918 6688 8938 6752
rect 9002 6688 9022 6752
rect 8918 6672 9022 6688
rect 8918 6608 8938 6672
rect 9002 6608 9022 6672
rect 8918 6592 9022 6608
rect 8918 6528 8938 6592
rect 9002 6528 9022 6592
rect 8918 6512 9022 6528
rect 8918 6448 8938 6512
rect 9002 6448 9022 6512
rect 8918 6432 9022 6448
rect 8918 6368 8938 6432
rect 9002 6368 9022 6432
rect 8918 6352 9022 6368
rect 8918 6288 8938 6352
rect 9002 6288 9022 6352
rect 8918 6272 9022 6288
rect 8918 6208 8938 6272
rect 9002 6208 9022 6272
rect 8918 6192 9022 6208
rect 8918 6128 8938 6192
rect 9002 6128 9022 6192
rect 8918 6112 9022 6128
rect 8918 6048 8938 6112
rect 9002 6048 9022 6112
rect 8918 6032 9022 6048
rect 6306 5632 6410 5968
rect 3694 5552 3798 5568
rect 3694 5488 3714 5552
rect 3778 5488 3798 5552
rect 3694 5472 3798 5488
rect 3694 5408 3714 5472
rect 3778 5408 3798 5472
rect 3694 5392 3798 5408
rect 3694 5328 3714 5392
rect 3778 5328 3798 5392
rect 3694 5312 3798 5328
rect 3694 5248 3714 5312
rect 3778 5248 3798 5312
rect 3694 5232 3798 5248
rect 3694 5168 3714 5232
rect 3778 5168 3798 5232
rect 3694 5152 3798 5168
rect 3694 5088 3714 5152
rect 3778 5088 3798 5152
rect 3694 5072 3798 5088
rect 3694 5008 3714 5072
rect 3778 5008 3798 5072
rect 3694 4992 3798 5008
rect 3694 4928 3714 4992
rect 3778 4928 3798 4992
rect 3694 4912 3798 4928
rect 3694 4848 3714 4912
rect 3778 4848 3798 4912
rect 3694 4832 3798 4848
rect 3694 4768 3714 4832
rect 3778 4768 3798 4832
rect 3694 4752 3798 4768
rect 3694 4688 3714 4752
rect 3778 4688 3798 4752
rect 3694 4672 3798 4688
rect 3694 4608 3714 4672
rect 3778 4608 3798 4672
rect 3694 4592 3798 4608
rect 3694 4528 3714 4592
rect 3778 4528 3798 4592
rect 3694 4512 3798 4528
rect 3694 4448 3714 4512
rect 3778 4448 3798 4512
rect 3694 4432 3798 4448
rect 3694 4368 3714 4432
rect 3778 4368 3798 4432
rect 3694 4352 3798 4368
rect 3694 4288 3714 4352
rect 3778 4288 3798 4352
rect 3694 4272 3798 4288
rect 3694 4208 3714 4272
rect 3778 4208 3798 4272
rect 3694 4192 3798 4208
rect 3694 4128 3714 4192
rect 3778 4128 3798 4192
rect 3694 4112 3798 4128
rect 3694 4048 3714 4112
rect 3778 4048 3798 4112
rect 3694 4032 3798 4048
rect 3694 3968 3714 4032
rect 3778 3968 3798 4032
rect 3694 3952 3798 3968
rect 3694 3888 3714 3952
rect 3778 3888 3798 3952
rect 3694 3872 3798 3888
rect 3694 3808 3714 3872
rect 3778 3808 3798 3872
rect 3694 3792 3798 3808
rect 3694 3728 3714 3792
rect 3778 3728 3798 3792
rect 3694 3712 3798 3728
rect 1082 3312 1186 3648
rect -1530 3232 -1426 3248
rect -1530 3168 -1510 3232
rect -1446 3168 -1426 3232
rect -1530 3152 -1426 3168
rect -1530 3088 -1510 3152
rect -1446 3088 -1426 3152
rect -1530 3072 -1426 3088
rect -1530 3008 -1510 3072
rect -1446 3008 -1426 3072
rect -1530 2992 -1426 3008
rect -1530 2928 -1510 2992
rect -1446 2928 -1426 2992
rect -1530 2912 -1426 2928
rect -1530 2848 -1510 2912
rect -1446 2848 -1426 2912
rect -1530 2832 -1426 2848
rect -1530 2768 -1510 2832
rect -1446 2768 -1426 2832
rect -1530 2752 -1426 2768
rect -1530 2688 -1510 2752
rect -1446 2688 -1426 2752
rect -1530 2672 -1426 2688
rect -1530 2608 -1510 2672
rect -1446 2608 -1426 2672
rect -1530 2592 -1426 2608
rect -1530 2528 -1510 2592
rect -1446 2528 -1426 2592
rect -1530 2512 -1426 2528
rect -1530 2448 -1510 2512
rect -1446 2448 -1426 2512
rect -1530 2432 -1426 2448
rect -1530 2368 -1510 2432
rect -1446 2368 -1426 2432
rect -1530 2352 -1426 2368
rect -1530 2288 -1510 2352
rect -1446 2288 -1426 2352
rect -1530 2272 -1426 2288
rect -1530 2208 -1510 2272
rect -1446 2208 -1426 2272
rect -1530 2192 -1426 2208
rect -1530 2128 -1510 2192
rect -1446 2128 -1426 2192
rect -1530 2112 -1426 2128
rect -1530 2048 -1510 2112
rect -1446 2048 -1426 2112
rect -1530 2032 -1426 2048
rect -1530 1968 -1510 2032
rect -1446 1968 -1426 2032
rect -1530 1952 -1426 1968
rect -1530 1888 -1510 1952
rect -1446 1888 -1426 1952
rect -1530 1872 -1426 1888
rect -1530 1808 -1510 1872
rect -1446 1808 -1426 1872
rect -1530 1792 -1426 1808
rect -1530 1728 -1510 1792
rect -1446 1728 -1426 1792
rect -1530 1712 -1426 1728
rect -1530 1648 -1510 1712
rect -1446 1648 -1426 1712
rect -1530 1632 -1426 1648
rect -1530 1568 -1510 1632
rect -1446 1568 -1426 1632
rect -1530 1552 -1426 1568
rect -1530 1488 -1510 1552
rect -1446 1488 -1426 1552
rect -1530 1472 -1426 1488
rect -1530 1408 -1510 1472
rect -1446 1408 -1426 1472
rect -1530 1392 -1426 1408
rect -4142 992 -4038 1328
rect -6754 912 -6650 928
rect -6754 848 -6734 912
rect -6670 848 -6650 912
rect -6754 832 -6650 848
rect -6754 768 -6734 832
rect -6670 768 -6650 832
rect -6754 752 -6650 768
rect -6754 688 -6734 752
rect -6670 688 -6650 752
rect -6754 672 -6650 688
rect -6754 608 -6734 672
rect -6670 608 -6650 672
rect -6754 592 -6650 608
rect -6754 528 -6734 592
rect -6670 528 -6650 592
rect -6754 512 -6650 528
rect -6754 448 -6734 512
rect -6670 448 -6650 512
rect -6754 432 -6650 448
rect -6754 368 -6734 432
rect -6670 368 -6650 432
rect -6754 352 -6650 368
rect -6754 288 -6734 352
rect -6670 288 -6650 352
rect -6754 272 -6650 288
rect -6754 208 -6734 272
rect -6670 208 -6650 272
rect -6754 192 -6650 208
rect -6754 128 -6734 192
rect -6670 128 -6650 192
rect -6754 112 -6650 128
rect -6754 48 -6734 112
rect -6670 48 -6650 112
rect -6754 32 -6650 48
rect -6754 -32 -6734 32
rect -6670 -32 -6650 32
rect -6754 -48 -6650 -32
rect -6754 -112 -6734 -48
rect -6670 -112 -6650 -48
rect -6754 -128 -6650 -112
rect -6754 -192 -6734 -128
rect -6670 -192 -6650 -128
rect -6754 -208 -6650 -192
rect -6754 -272 -6734 -208
rect -6670 -272 -6650 -208
rect -6754 -288 -6650 -272
rect -6754 -352 -6734 -288
rect -6670 -352 -6650 -288
rect -6754 -368 -6650 -352
rect -6754 -432 -6734 -368
rect -6670 -432 -6650 -368
rect -6754 -448 -6650 -432
rect -6754 -512 -6734 -448
rect -6670 -512 -6650 -448
rect -6754 -528 -6650 -512
rect -6754 -592 -6734 -528
rect -6670 -592 -6650 -528
rect -6754 -608 -6650 -592
rect -6754 -672 -6734 -608
rect -6670 -672 -6650 -608
rect -6754 -688 -6650 -672
rect -6754 -752 -6734 -688
rect -6670 -752 -6650 -688
rect -6754 -768 -6650 -752
rect -6754 -832 -6734 -768
rect -6670 -832 -6650 -768
rect -6754 -848 -6650 -832
rect -6754 -912 -6734 -848
rect -6670 -912 -6650 -848
rect -6754 -928 -6650 -912
rect -8034 -1359 -7930 -961
rect -6754 -992 -6734 -928
rect -6670 -992 -6650 -928
rect -6331 952 -4409 961
rect -6331 -952 -6322 952
rect -4418 -952 -4409 952
rect -6331 -961 -4409 -952
rect -4142 928 -4122 992
rect -4058 928 -4038 992
rect -2810 961 -2706 1359
rect -1530 1328 -1510 1392
rect -1446 1328 -1426 1392
rect -1107 3272 815 3281
rect -1107 1368 -1098 3272
rect 806 1368 815 3272
rect -1107 1359 815 1368
rect 1082 3248 1102 3312
rect 1166 3248 1186 3312
rect 2414 3281 2518 3679
rect 3694 3648 3714 3712
rect 3778 3648 3798 3712
rect 4117 5592 6039 5601
rect 4117 3688 4126 5592
rect 6030 3688 6039 5592
rect 4117 3679 6039 3688
rect 6306 5568 6326 5632
rect 6390 5568 6410 5632
rect 7638 5601 7742 5999
rect 8918 5968 8938 6032
rect 9002 5968 9022 6032
rect 8918 5632 9022 5968
rect 6306 5552 6410 5568
rect 6306 5488 6326 5552
rect 6390 5488 6410 5552
rect 6306 5472 6410 5488
rect 6306 5408 6326 5472
rect 6390 5408 6410 5472
rect 6306 5392 6410 5408
rect 6306 5328 6326 5392
rect 6390 5328 6410 5392
rect 6306 5312 6410 5328
rect 6306 5248 6326 5312
rect 6390 5248 6410 5312
rect 6306 5232 6410 5248
rect 6306 5168 6326 5232
rect 6390 5168 6410 5232
rect 6306 5152 6410 5168
rect 6306 5088 6326 5152
rect 6390 5088 6410 5152
rect 6306 5072 6410 5088
rect 6306 5008 6326 5072
rect 6390 5008 6410 5072
rect 6306 4992 6410 5008
rect 6306 4928 6326 4992
rect 6390 4928 6410 4992
rect 6306 4912 6410 4928
rect 6306 4848 6326 4912
rect 6390 4848 6410 4912
rect 6306 4832 6410 4848
rect 6306 4768 6326 4832
rect 6390 4768 6410 4832
rect 6306 4752 6410 4768
rect 6306 4688 6326 4752
rect 6390 4688 6410 4752
rect 6306 4672 6410 4688
rect 6306 4608 6326 4672
rect 6390 4608 6410 4672
rect 6306 4592 6410 4608
rect 6306 4528 6326 4592
rect 6390 4528 6410 4592
rect 6306 4512 6410 4528
rect 6306 4448 6326 4512
rect 6390 4448 6410 4512
rect 6306 4432 6410 4448
rect 6306 4368 6326 4432
rect 6390 4368 6410 4432
rect 6306 4352 6410 4368
rect 6306 4288 6326 4352
rect 6390 4288 6410 4352
rect 6306 4272 6410 4288
rect 6306 4208 6326 4272
rect 6390 4208 6410 4272
rect 6306 4192 6410 4208
rect 6306 4128 6326 4192
rect 6390 4128 6410 4192
rect 6306 4112 6410 4128
rect 6306 4048 6326 4112
rect 6390 4048 6410 4112
rect 6306 4032 6410 4048
rect 6306 3968 6326 4032
rect 6390 3968 6410 4032
rect 6306 3952 6410 3968
rect 6306 3888 6326 3952
rect 6390 3888 6410 3952
rect 6306 3872 6410 3888
rect 6306 3808 6326 3872
rect 6390 3808 6410 3872
rect 6306 3792 6410 3808
rect 6306 3728 6326 3792
rect 6390 3728 6410 3792
rect 6306 3712 6410 3728
rect 3694 3312 3798 3648
rect 1082 3232 1186 3248
rect 1082 3168 1102 3232
rect 1166 3168 1186 3232
rect 1082 3152 1186 3168
rect 1082 3088 1102 3152
rect 1166 3088 1186 3152
rect 1082 3072 1186 3088
rect 1082 3008 1102 3072
rect 1166 3008 1186 3072
rect 1082 2992 1186 3008
rect 1082 2928 1102 2992
rect 1166 2928 1186 2992
rect 1082 2912 1186 2928
rect 1082 2848 1102 2912
rect 1166 2848 1186 2912
rect 1082 2832 1186 2848
rect 1082 2768 1102 2832
rect 1166 2768 1186 2832
rect 1082 2752 1186 2768
rect 1082 2688 1102 2752
rect 1166 2688 1186 2752
rect 1082 2672 1186 2688
rect 1082 2608 1102 2672
rect 1166 2608 1186 2672
rect 1082 2592 1186 2608
rect 1082 2528 1102 2592
rect 1166 2528 1186 2592
rect 1082 2512 1186 2528
rect 1082 2448 1102 2512
rect 1166 2448 1186 2512
rect 1082 2432 1186 2448
rect 1082 2368 1102 2432
rect 1166 2368 1186 2432
rect 1082 2352 1186 2368
rect 1082 2288 1102 2352
rect 1166 2288 1186 2352
rect 1082 2272 1186 2288
rect 1082 2208 1102 2272
rect 1166 2208 1186 2272
rect 1082 2192 1186 2208
rect 1082 2128 1102 2192
rect 1166 2128 1186 2192
rect 1082 2112 1186 2128
rect 1082 2048 1102 2112
rect 1166 2048 1186 2112
rect 1082 2032 1186 2048
rect 1082 1968 1102 2032
rect 1166 1968 1186 2032
rect 1082 1952 1186 1968
rect 1082 1888 1102 1952
rect 1166 1888 1186 1952
rect 1082 1872 1186 1888
rect 1082 1808 1102 1872
rect 1166 1808 1186 1872
rect 1082 1792 1186 1808
rect 1082 1728 1102 1792
rect 1166 1728 1186 1792
rect 1082 1712 1186 1728
rect 1082 1648 1102 1712
rect 1166 1648 1186 1712
rect 1082 1632 1186 1648
rect 1082 1568 1102 1632
rect 1166 1568 1186 1632
rect 1082 1552 1186 1568
rect 1082 1488 1102 1552
rect 1166 1488 1186 1552
rect 1082 1472 1186 1488
rect 1082 1408 1102 1472
rect 1166 1408 1186 1472
rect 1082 1392 1186 1408
rect -1530 992 -1426 1328
rect -4142 912 -4038 928
rect -4142 848 -4122 912
rect -4058 848 -4038 912
rect -4142 832 -4038 848
rect -4142 768 -4122 832
rect -4058 768 -4038 832
rect -4142 752 -4038 768
rect -4142 688 -4122 752
rect -4058 688 -4038 752
rect -4142 672 -4038 688
rect -4142 608 -4122 672
rect -4058 608 -4038 672
rect -4142 592 -4038 608
rect -4142 528 -4122 592
rect -4058 528 -4038 592
rect -4142 512 -4038 528
rect -4142 448 -4122 512
rect -4058 448 -4038 512
rect -4142 432 -4038 448
rect -4142 368 -4122 432
rect -4058 368 -4038 432
rect -4142 352 -4038 368
rect -4142 288 -4122 352
rect -4058 288 -4038 352
rect -4142 272 -4038 288
rect -4142 208 -4122 272
rect -4058 208 -4038 272
rect -4142 192 -4038 208
rect -4142 128 -4122 192
rect -4058 128 -4038 192
rect -4142 112 -4038 128
rect -4142 48 -4122 112
rect -4058 48 -4038 112
rect -4142 32 -4038 48
rect -4142 -32 -4122 32
rect -4058 -32 -4038 32
rect -4142 -48 -4038 -32
rect -4142 -112 -4122 -48
rect -4058 -112 -4038 -48
rect -4142 -128 -4038 -112
rect -4142 -192 -4122 -128
rect -4058 -192 -4038 -128
rect -4142 -208 -4038 -192
rect -4142 -272 -4122 -208
rect -4058 -272 -4038 -208
rect -4142 -288 -4038 -272
rect -4142 -352 -4122 -288
rect -4058 -352 -4038 -288
rect -4142 -368 -4038 -352
rect -4142 -432 -4122 -368
rect -4058 -432 -4038 -368
rect -4142 -448 -4038 -432
rect -4142 -512 -4122 -448
rect -4058 -512 -4038 -448
rect -4142 -528 -4038 -512
rect -4142 -592 -4122 -528
rect -4058 -592 -4038 -528
rect -4142 -608 -4038 -592
rect -4142 -672 -4122 -608
rect -4058 -672 -4038 -608
rect -4142 -688 -4038 -672
rect -4142 -752 -4122 -688
rect -4058 -752 -4038 -688
rect -4142 -768 -4038 -752
rect -4142 -832 -4122 -768
rect -4058 -832 -4038 -768
rect -4142 -848 -4038 -832
rect -4142 -912 -4122 -848
rect -4058 -912 -4038 -848
rect -4142 -928 -4038 -912
rect -6754 -1328 -6650 -992
rect -8943 -1368 -7021 -1359
rect -8943 -3272 -8934 -1368
rect -7030 -3272 -7021 -1368
rect -8943 -3281 -7021 -3272
rect -6754 -1392 -6734 -1328
rect -6670 -1392 -6650 -1328
rect -5422 -1359 -5318 -961
rect -4142 -992 -4122 -928
rect -4058 -992 -4038 -928
rect -3719 952 -1797 961
rect -3719 -952 -3710 952
rect -1806 -952 -1797 952
rect -3719 -961 -1797 -952
rect -1530 928 -1510 992
rect -1446 928 -1426 992
rect -198 961 -94 1359
rect 1082 1328 1102 1392
rect 1166 1328 1186 1392
rect 1505 3272 3427 3281
rect 1505 1368 1514 3272
rect 3418 1368 3427 3272
rect 1505 1359 3427 1368
rect 3694 3248 3714 3312
rect 3778 3248 3798 3312
rect 5026 3281 5130 3679
rect 6306 3648 6326 3712
rect 6390 3648 6410 3712
rect 6729 5592 8651 5601
rect 6729 3688 6738 5592
rect 8642 3688 8651 5592
rect 6729 3679 8651 3688
rect 8918 5568 8938 5632
rect 9002 5568 9022 5632
rect 8918 5552 9022 5568
rect 8918 5488 8938 5552
rect 9002 5488 9022 5552
rect 8918 5472 9022 5488
rect 8918 5408 8938 5472
rect 9002 5408 9022 5472
rect 8918 5392 9022 5408
rect 8918 5328 8938 5392
rect 9002 5328 9022 5392
rect 8918 5312 9022 5328
rect 8918 5248 8938 5312
rect 9002 5248 9022 5312
rect 8918 5232 9022 5248
rect 8918 5168 8938 5232
rect 9002 5168 9022 5232
rect 8918 5152 9022 5168
rect 8918 5088 8938 5152
rect 9002 5088 9022 5152
rect 8918 5072 9022 5088
rect 8918 5008 8938 5072
rect 9002 5008 9022 5072
rect 8918 4992 9022 5008
rect 8918 4928 8938 4992
rect 9002 4928 9022 4992
rect 8918 4912 9022 4928
rect 8918 4848 8938 4912
rect 9002 4848 9022 4912
rect 8918 4832 9022 4848
rect 8918 4768 8938 4832
rect 9002 4768 9022 4832
rect 8918 4752 9022 4768
rect 8918 4688 8938 4752
rect 9002 4688 9022 4752
rect 8918 4672 9022 4688
rect 8918 4608 8938 4672
rect 9002 4608 9022 4672
rect 8918 4592 9022 4608
rect 8918 4528 8938 4592
rect 9002 4528 9022 4592
rect 8918 4512 9022 4528
rect 8918 4448 8938 4512
rect 9002 4448 9022 4512
rect 8918 4432 9022 4448
rect 8918 4368 8938 4432
rect 9002 4368 9022 4432
rect 8918 4352 9022 4368
rect 8918 4288 8938 4352
rect 9002 4288 9022 4352
rect 8918 4272 9022 4288
rect 8918 4208 8938 4272
rect 9002 4208 9022 4272
rect 8918 4192 9022 4208
rect 8918 4128 8938 4192
rect 9002 4128 9022 4192
rect 8918 4112 9022 4128
rect 8918 4048 8938 4112
rect 9002 4048 9022 4112
rect 8918 4032 9022 4048
rect 8918 3968 8938 4032
rect 9002 3968 9022 4032
rect 8918 3952 9022 3968
rect 8918 3888 8938 3952
rect 9002 3888 9022 3952
rect 8918 3872 9022 3888
rect 8918 3808 8938 3872
rect 9002 3808 9022 3872
rect 8918 3792 9022 3808
rect 8918 3728 8938 3792
rect 9002 3728 9022 3792
rect 8918 3712 9022 3728
rect 6306 3312 6410 3648
rect 3694 3232 3798 3248
rect 3694 3168 3714 3232
rect 3778 3168 3798 3232
rect 3694 3152 3798 3168
rect 3694 3088 3714 3152
rect 3778 3088 3798 3152
rect 3694 3072 3798 3088
rect 3694 3008 3714 3072
rect 3778 3008 3798 3072
rect 3694 2992 3798 3008
rect 3694 2928 3714 2992
rect 3778 2928 3798 2992
rect 3694 2912 3798 2928
rect 3694 2848 3714 2912
rect 3778 2848 3798 2912
rect 3694 2832 3798 2848
rect 3694 2768 3714 2832
rect 3778 2768 3798 2832
rect 3694 2752 3798 2768
rect 3694 2688 3714 2752
rect 3778 2688 3798 2752
rect 3694 2672 3798 2688
rect 3694 2608 3714 2672
rect 3778 2608 3798 2672
rect 3694 2592 3798 2608
rect 3694 2528 3714 2592
rect 3778 2528 3798 2592
rect 3694 2512 3798 2528
rect 3694 2448 3714 2512
rect 3778 2448 3798 2512
rect 3694 2432 3798 2448
rect 3694 2368 3714 2432
rect 3778 2368 3798 2432
rect 3694 2352 3798 2368
rect 3694 2288 3714 2352
rect 3778 2288 3798 2352
rect 3694 2272 3798 2288
rect 3694 2208 3714 2272
rect 3778 2208 3798 2272
rect 3694 2192 3798 2208
rect 3694 2128 3714 2192
rect 3778 2128 3798 2192
rect 3694 2112 3798 2128
rect 3694 2048 3714 2112
rect 3778 2048 3798 2112
rect 3694 2032 3798 2048
rect 3694 1968 3714 2032
rect 3778 1968 3798 2032
rect 3694 1952 3798 1968
rect 3694 1888 3714 1952
rect 3778 1888 3798 1952
rect 3694 1872 3798 1888
rect 3694 1808 3714 1872
rect 3778 1808 3798 1872
rect 3694 1792 3798 1808
rect 3694 1728 3714 1792
rect 3778 1728 3798 1792
rect 3694 1712 3798 1728
rect 3694 1648 3714 1712
rect 3778 1648 3798 1712
rect 3694 1632 3798 1648
rect 3694 1568 3714 1632
rect 3778 1568 3798 1632
rect 3694 1552 3798 1568
rect 3694 1488 3714 1552
rect 3778 1488 3798 1552
rect 3694 1472 3798 1488
rect 3694 1408 3714 1472
rect 3778 1408 3798 1472
rect 3694 1392 3798 1408
rect 1082 992 1186 1328
rect -1530 912 -1426 928
rect -1530 848 -1510 912
rect -1446 848 -1426 912
rect -1530 832 -1426 848
rect -1530 768 -1510 832
rect -1446 768 -1426 832
rect -1530 752 -1426 768
rect -1530 688 -1510 752
rect -1446 688 -1426 752
rect -1530 672 -1426 688
rect -1530 608 -1510 672
rect -1446 608 -1426 672
rect -1530 592 -1426 608
rect -1530 528 -1510 592
rect -1446 528 -1426 592
rect -1530 512 -1426 528
rect -1530 448 -1510 512
rect -1446 448 -1426 512
rect -1530 432 -1426 448
rect -1530 368 -1510 432
rect -1446 368 -1426 432
rect -1530 352 -1426 368
rect -1530 288 -1510 352
rect -1446 288 -1426 352
rect -1530 272 -1426 288
rect -1530 208 -1510 272
rect -1446 208 -1426 272
rect -1530 192 -1426 208
rect -1530 128 -1510 192
rect -1446 128 -1426 192
rect -1530 112 -1426 128
rect -1530 48 -1510 112
rect -1446 48 -1426 112
rect -1530 32 -1426 48
rect -1530 -32 -1510 32
rect -1446 -32 -1426 32
rect -1530 -48 -1426 -32
rect -1530 -112 -1510 -48
rect -1446 -112 -1426 -48
rect -1530 -128 -1426 -112
rect -1530 -192 -1510 -128
rect -1446 -192 -1426 -128
rect -1530 -208 -1426 -192
rect -1530 -272 -1510 -208
rect -1446 -272 -1426 -208
rect -1530 -288 -1426 -272
rect -1530 -352 -1510 -288
rect -1446 -352 -1426 -288
rect -1530 -368 -1426 -352
rect -1530 -432 -1510 -368
rect -1446 -432 -1426 -368
rect -1530 -448 -1426 -432
rect -1530 -512 -1510 -448
rect -1446 -512 -1426 -448
rect -1530 -528 -1426 -512
rect -1530 -592 -1510 -528
rect -1446 -592 -1426 -528
rect -1530 -608 -1426 -592
rect -1530 -672 -1510 -608
rect -1446 -672 -1426 -608
rect -1530 -688 -1426 -672
rect -1530 -752 -1510 -688
rect -1446 -752 -1426 -688
rect -1530 -768 -1426 -752
rect -1530 -832 -1510 -768
rect -1446 -832 -1426 -768
rect -1530 -848 -1426 -832
rect -1530 -912 -1510 -848
rect -1446 -912 -1426 -848
rect -1530 -928 -1426 -912
rect -4142 -1328 -4038 -992
rect -6754 -1408 -6650 -1392
rect -6754 -1472 -6734 -1408
rect -6670 -1472 -6650 -1408
rect -6754 -1488 -6650 -1472
rect -6754 -1552 -6734 -1488
rect -6670 -1552 -6650 -1488
rect -6754 -1568 -6650 -1552
rect -6754 -1632 -6734 -1568
rect -6670 -1632 -6650 -1568
rect -6754 -1648 -6650 -1632
rect -6754 -1712 -6734 -1648
rect -6670 -1712 -6650 -1648
rect -6754 -1728 -6650 -1712
rect -6754 -1792 -6734 -1728
rect -6670 -1792 -6650 -1728
rect -6754 -1808 -6650 -1792
rect -6754 -1872 -6734 -1808
rect -6670 -1872 -6650 -1808
rect -6754 -1888 -6650 -1872
rect -6754 -1952 -6734 -1888
rect -6670 -1952 -6650 -1888
rect -6754 -1968 -6650 -1952
rect -6754 -2032 -6734 -1968
rect -6670 -2032 -6650 -1968
rect -6754 -2048 -6650 -2032
rect -6754 -2112 -6734 -2048
rect -6670 -2112 -6650 -2048
rect -6754 -2128 -6650 -2112
rect -6754 -2192 -6734 -2128
rect -6670 -2192 -6650 -2128
rect -6754 -2208 -6650 -2192
rect -6754 -2272 -6734 -2208
rect -6670 -2272 -6650 -2208
rect -6754 -2288 -6650 -2272
rect -6754 -2352 -6734 -2288
rect -6670 -2352 -6650 -2288
rect -6754 -2368 -6650 -2352
rect -6754 -2432 -6734 -2368
rect -6670 -2432 -6650 -2368
rect -6754 -2448 -6650 -2432
rect -6754 -2512 -6734 -2448
rect -6670 -2512 -6650 -2448
rect -6754 -2528 -6650 -2512
rect -6754 -2592 -6734 -2528
rect -6670 -2592 -6650 -2528
rect -6754 -2608 -6650 -2592
rect -6754 -2672 -6734 -2608
rect -6670 -2672 -6650 -2608
rect -6754 -2688 -6650 -2672
rect -6754 -2752 -6734 -2688
rect -6670 -2752 -6650 -2688
rect -6754 -2768 -6650 -2752
rect -6754 -2832 -6734 -2768
rect -6670 -2832 -6650 -2768
rect -6754 -2848 -6650 -2832
rect -6754 -2912 -6734 -2848
rect -6670 -2912 -6650 -2848
rect -6754 -2928 -6650 -2912
rect -6754 -2992 -6734 -2928
rect -6670 -2992 -6650 -2928
rect -6754 -3008 -6650 -2992
rect -6754 -3072 -6734 -3008
rect -6670 -3072 -6650 -3008
rect -6754 -3088 -6650 -3072
rect -6754 -3152 -6734 -3088
rect -6670 -3152 -6650 -3088
rect -6754 -3168 -6650 -3152
rect -6754 -3232 -6734 -3168
rect -6670 -3232 -6650 -3168
rect -6754 -3248 -6650 -3232
rect -8034 -3679 -7930 -3281
rect -6754 -3312 -6734 -3248
rect -6670 -3312 -6650 -3248
rect -6331 -1368 -4409 -1359
rect -6331 -3272 -6322 -1368
rect -4418 -3272 -4409 -1368
rect -6331 -3281 -4409 -3272
rect -4142 -1392 -4122 -1328
rect -4058 -1392 -4038 -1328
rect -2810 -1359 -2706 -961
rect -1530 -992 -1510 -928
rect -1446 -992 -1426 -928
rect -1107 952 815 961
rect -1107 -952 -1098 952
rect 806 -952 815 952
rect -1107 -961 815 -952
rect 1082 928 1102 992
rect 1166 928 1186 992
rect 2414 961 2518 1359
rect 3694 1328 3714 1392
rect 3778 1328 3798 1392
rect 4117 3272 6039 3281
rect 4117 1368 4126 3272
rect 6030 1368 6039 3272
rect 4117 1359 6039 1368
rect 6306 3248 6326 3312
rect 6390 3248 6410 3312
rect 7638 3281 7742 3679
rect 8918 3648 8938 3712
rect 9002 3648 9022 3712
rect 8918 3312 9022 3648
rect 6306 3232 6410 3248
rect 6306 3168 6326 3232
rect 6390 3168 6410 3232
rect 6306 3152 6410 3168
rect 6306 3088 6326 3152
rect 6390 3088 6410 3152
rect 6306 3072 6410 3088
rect 6306 3008 6326 3072
rect 6390 3008 6410 3072
rect 6306 2992 6410 3008
rect 6306 2928 6326 2992
rect 6390 2928 6410 2992
rect 6306 2912 6410 2928
rect 6306 2848 6326 2912
rect 6390 2848 6410 2912
rect 6306 2832 6410 2848
rect 6306 2768 6326 2832
rect 6390 2768 6410 2832
rect 6306 2752 6410 2768
rect 6306 2688 6326 2752
rect 6390 2688 6410 2752
rect 6306 2672 6410 2688
rect 6306 2608 6326 2672
rect 6390 2608 6410 2672
rect 6306 2592 6410 2608
rect 6306 2528 6326 2592
rect 6390 2528 6410 2592
rect 6306 2512 6410 2528
rect 6306 2448 6326 2512
rect 6390 2448 6410 2512
rect 6306 2432 6410 2448
rect 6306 2368 6326 2432
rect 6390 2368 6410 2432
rect 6306 2352 6410 2368
rect 6306 2288 6326 2352
rect 6390 2288 6410 2352
rect 6306 2272 6410 2288
rect 6306 2208 6326 2272
rect 6390 2208 6410 2272
rect 6306 2192 6410 2208
rect 6306 2128 6326 2192
rect 6390 2128 6410 2192
rect 6306 2112 6410 2128
rect 6306 2048 6326 2112
rect 6390 2048 6410 2112
rect 6306 2032 6410 2048
rect 6306 1968 6326 2032
rect 6390 1968 6410 2032
rect 6306 1952 6410 1968
rect 6306 1888 6326 1952
rect 6390 1888 6410 1952
rect 6306 1872 6410 1888
rect 6306 1808 6326 1872
rect 6390 1808 6410 1872
rect 6306 1792 6410 1808
rect 6306 1728 6326 1792
rect 6390 1728 6410 1792
rect 6306 1712 6410 1728
rect 6306 1648 6326 1712
rect 6390 1648 6410 1712
rect 6306 1632 6410 1648
rect 6306 1568 6326 1632
rect 6390 1568 6410 1632
rect 6306 1552 6410 1568
rect 6306 1488 6326 1552
rect 6390 1488 6410 1552
rect 6306 1472 6410 1488
rect 6306 1408 6326 1472
rect 6390 1408 6410 1472
rect 6306 1392 6410 1408
rect 3694 992 3798 1328
rect 1082 912 1186 928
rect 1082 848 1102 912
rect 1166 848 1186 912
rect 1082 832 1186 848
rect 1082 768 1102 832
rect 1166 768 1186 832
rect 1082 752 1186 768
rect 1082 688 1102 752
rect 1166 688 1186 752
rect 1082 672 1186 688
rect 1082 608 1102 672
rect 1166 608 1186 672
rect 1082 592 1186 608
rect 1082 528 1102 592
rect 1166 528 1186 592
rect 1082 512 1186 528
rect 1082 448 1102 512
rect 1166 448 1186 512
rect 1082 432 1186 448
rect 1082 368 1102 432
rect 1166 368 1186 432
rect 1082 352 1186 368
rect 1082 288 1102 352
rect 1166 288 1186 352
rect 1082 272 1186 288
rect 1082 208 1102 272
rect 1166 208 1186 272
rect 1082 192 1186 208
rect 1082 128 1102 192
rect 1166 128 1186 192
rect 1082 112 1186 128
rect 1082 48 1102 112
rect 1166 48 1186 112
rect 1082 32 1186 48
rect 1082 -32 1102 32
rect 1166 -32 1186 32
rect 1082 -48 1186 -32
rect 1082 -112 1102 -48
rect 1166 -112 1186 -48
rect 1082 -128 1186 -112
rect 1082 -192 1102 -128
rect 1166 -192 1186 -128
rect 1082 -208 1186 -192
rect 1082 -272 1102 -208
rect 1166 -272 1186 -208
rect 1082 -288 1186 -272
rect 1082 -352 1102 -288
rect 1166 -352 1186 -288
rect 1082 -368 1186 -352
rect 1082 -432 1102 -368
rect 1166 -432 1186 -368
rect 1082 -448 1186 -432
rect 1082 -512 1102 -448
rect 1166 -512 1186 -448
rect 1082 -528 1186 -512
rect 1082 -592 1102 -528
rect 1166 -592 1186 -528
rect 1082 -608 1186 -592
rect 1082 -672 1102 -608
rect 1166 -672 1186 -608
rect 1082 -688 1186 -672
rect 1082 -752 1102 -688
rect 1166 -752 1186 -688
rect 1082 -768 1186 -752
rect 1082 -832 1102 -768
rect 1166 -832 1186 -768
rect 1082 -848 1186 -832
rect 1082 -912 1102 -848
rect 1166 -912 1186 -848
rect 1082 -928 1186 -912
rect -1530 -1328 -1426 -992
rect -4142 -1408 -4038 -1392
rect -4142 -1472 -4122 -1408
rect -4058 -1472 -4038 -1408
rect -4142 -1488 -4038 -1472
rect -4142 -1552 -4122 -1488
rect -4058 -1552 -4038 -1488
rect -4142 -1568 -4038 -1552
rect -4142 -1632 -4122 -1568
rect -4058 -1632 -4038 -1568
rect -4142 -1648 -4038 -1632
rect -4142 -1712 -4122 -1648
rect -4058 -1712 -4038 -1648
rect -4142 -1728 -4038 -1712
rect -4142 -1792 -4122 -1728
rect -4058 -1792 -4038 -1728
rect -4142 -1808 -4038 -1792
rect -4142 -1872 -4122 -1808
rect -4058 -1872 -4038 -1808
rect -4142 -1888 -4038 -1872
rect -4142 -1952 -4122 -1888
rect -4058 -1952 -4038 -1888
rect -4142 -1968 -4038 -1952
rect -4142 -2032 -4122 -1968
rect -4058 -2032 -4038 -1968
rect -4142 -2048 -4038 -2032
rect -4142 -2112 -4122 -2048
rect -4058 -2112 -4038 -2048
rect -4142 -2128 -4038 -2112
rect -4142 -2192 -4122 -2128
rect -4058 -2192 -4038 -2128
rect -4142 -2208 -4038 -2192
rect -4142 -2272 -4122 -2208
rect -4058 -2272 -4038 -2208
rect -4142 -2288 -4038 -2272
rect -4142 -2352 -4122 -2288
rect -4058 -2352 -4038 -2288
rect -4142 -2368 -4038 -2352
rect -4142 -2432 -4122 -2368
rect -4058 -2432 -4038 -2368
rect -4142 -2448 -4038 -2432
rect -4142 -2512 -4122 -2448
rect -4058 -2512 -4038 -2448
rect -4142 -2528 -4038 -2512
rect -4142 -2592 -4122 -2528
rect -4058 -2592 -4038 -2528
rect -4142 -2608 -4038 -2592
rect -4142 -2672 -4122 -2608
rect -4058 -2672 -4038 -2608
rect -4142 -2688 -4038 -2672
rect -4142 -2752 -4122 -2688
rect -4058 -2752 -4038 -2688
rect -4142 -2768 -4038 -2752
rect -4142 -2832 -4122 -2768
rect -4058 -2832 -4038 -2768
rect -4142 -2848 -4038 -2832
rect -4142 -2912 -4122 -2848
rect -4058 -2912 -4038 -2848
rect -4142 -2928 -4038 -2912
rect -4142 -2992 -4122 -2928
rect -4058 -2992 -4038 -2928
rect -4142 -3008 -4038 -2992
rect -4142 -3072 -4122 -3008
rect -4058 -3072 -4038 -3008
rect -4142 -3088 -4038 -3072
rect -4142 -3152 -4122 -3088
rect -4058 -3152 -4038 -3088
rect -4142 -3168 -4038 -3152
rect -4142 -3232 -4122 -3168
rect -4058 -3232 -4038 -3168
rect -4142 -3248 -4038 -3232
rect -6754 -3648 -6650 -3312
rect -8943 -3688 -7021 -3679
rect -8943 -5592 -8934 -3688
rect -7030 -5592 -7021 -3688
rect -8943 -5601 -7021 -5592
rect -6754 -3712 -6734 -3648
rect -6670 -3712 -6650 -3648
rect -5422 -3679 -5318 -3281
rect -4142 -3312 -4122 -3248
rect -4058 -3312 -4038 -3248
rect -3719 -1368 -1797 -1359
rect -3719 -3272 -3710 -1368
rect -1806 -3272 -1797 -1368
rect -3719 -3281 -1797 -3272
rect -1530 -1392 -1510 -1328
rect -1446 -1392 -1426 -1328
rect -198 -1359 -94 -961
rect 1082 -992 1102 -928
rect 1166 -992 1186 -928
rect 1505 952 3427 961
rect 1505 -952 1514 952
rect 3418 -952 3427 952
rect 1505 -961 3427 -952
rect 3694 928 3714 992
rect 3778 928 3798 992
rect 5026 961 5130 1359
rect 6306 1328 6326 1392
rect 6390 1328 6410 1392
rect 6729 3272 8651 3281
rect 6729 1368 6738 3272
rect 8642 1368 8651 3272
rect 6729 1359 8651 1368
rect 8918 3248 8938 3312
rect 9002 3248 9022 3312
rect 8918 3232 9022 3248
rect 8918 3168 8938 3232
rect 9002 3168 9022 3232
rect 8918 3152 9022 3168
rect 8918 3088 8938 3152
rect 9002 3088 9022 3152
rect 8918 3072 9022 3088
rect 8918 3008 8938 3072
rect 9002 3008 9022 3072
rect 8918 2992 9022 3008
rect 8918 2928 8938 2992
rect 9002 2928 9022 2992
rect 8918 2912 9022 2928
rect 8918 2848 8938 2912
rect 9002 2848 9022 2912
rect 8918 2832 9022 2848
rect 8918 2768 8938 2832
rect 9002 2768 9022 2832
rect 8918 2752 9022 2768
rect 8918 2688 8938 2752
rect 9002 2688 9022 2752
rect 8918 2672 9022 2688
rect 8918 2608 8938 2672
rect 9002 2608 9022 2672
rect 8918 2592 9022 2608
rect 8918 2528 8938 2592
rect 9002 2528 9022 2592
rect 8918 2512 9022 2528
rect 8918 2448 8938 2512
rect 9002 2448 9022 2512
rect 8918 2432 9022 2448
rect 8918 2368 8938 2432
rect 9002 2368 9022 2432
rect 8918 2352 9022 2368
rect 8918 2288 8938 2352
rect 9002 2288 9022 2352
rect 8918 2272 9022 2288
rect 8918 2208 8938 2272
rect 9002 2208 9022 2272
rect 8918 2192 9022 2208
rect 8918 2128 8938 2192
rect 9002 2128 9022 2192
rect 8918 2112 9022 2128
rect 8918 2048 8938 2112
rect 9002 2048 9022 2112
rect 8918 2032 9022 2048
rect 8918 1968 8938 2032
rect 9002 1968 9022 2032
rect 8918 1952 9022 1968
rect 8918 1888 8938 1952
rect 9002 1888 9022 1952
rect 8918 1872 9022 1888
rect 8918 1808 8938 1872
rect 9002 1808 9022 1872
rect 8918 1792 9022 1808
rect 8918 1728 8938 1792
rect 9002 1728 9022 1792
rect 8918 1712 9022 1728
rect 8918 1648 8938 1712
rect 9002 1648 9022 1712
rect 8918 1632 9022 1648
rect 8918 1568 8938 1632
rect 9002 1568 9022 1632
rect 8918 1552 9022 1568
rect 8918 1488 8938 1552
rect 9002 1488 9022 1552
rect 8918 1472 9022 1488
rect 8918 1408 8938 1472
rect 9002 1408 9022 1472
rect 8918 1392 9022 1408
rect 6306 992 6410 1328
rect 3694 912 3798 928
rect 3694 848 3714 912
rect 3778 848 3798 912
rect 3694 832 3798 848
rect 3694 768 3714 832
rect 3778 768 3798 832
rect 3694 752 3798 768
rect 3694 688 3714 752
rect 3778 688 3798 752
rect 3694 672 3798 688
rect 3694 608 3714 672
rect 3778 608 3798 672
rect 3694 592 3798 608
rect 3694 528 3714 592
rect 3778 528 3798 592
rect 3694 512 3798 528
rect 3694 448 3714 512
rect 3778 448 3798 512
rect 3694 432 3798 448
rect 3694 368 3714 432
rect 3778 368 3798 432
rect 3694 352 3798 368
rect 3694 288 3714 352
rect 3778 288 3798 352
rect 3694 272 3798 288
rect 3694 208 3714 272
rect 3778 208 3798 272
rect 3694 192 3798 208
rect 3694 128 3714 192
rect 3778 128 3798 192
rect 3694 112 3798 128
rect 3694 48 3714 112
rect 3778 48 3798 112
rect 3694 32 3798 48
rect 3694 -32 3714 32
rect 3778 -32 3798 32
rect 3694 -48 3798 -32
rect 3694 -112 3714 -48
rect 3778 -112 3798 -48
rect 3694 -128 3798 -112
rect 3694 -192 3714 -128
rect 3778 -192 3798 -128
rect 3694 -208 3798 -192
rect 3694 -272 3714 -208
rect 3778 -272 3798 -208
rect 3694 -288 3798 -272
rect 3694 -352 3714 -288
rect 3778 -352 3798 -288
rect 3694 -368 3798 -352
rect 3694 -432 3714 -368
rect 3778 -432 3798 -368
rect 3694 -448 3798 -432
rect 3694 -512 3714 -448
rect 3778 -512 3798 -448
rect 3694 -528 3798 -512
rect 3694 -592 3714 -528
rect 3778 -592 3798 -528
rect 3694 -608 3798 -592
rect 3694 -672 3714 -608
rect 3778 -672 3798 -608
rect 3694 -688 3798 -672
rect 3694 -752 3714 -688
rect 3778 -752 3798 -688
rect 3694 -768 3798 -752
rect 3694 -832 3714 -768
rect 3778 -832 3798 -768
rect 3694 -848 3798 -832
rect 3694 -912 3714 -848
rect 3778 -912 3798 -848
rect 3694 -928 3798 -912
rect 1082 -1328 1186 -992
rect -1530 -1408 -1426 -1392
rect -1530 -1472 -1510 -1408
rect -1446 -1472 -1426 -1408
rect -1530 -1488 -1426 -1472
rect -1530 -1552 -1510 -1488
rect -1446 -1552 -1426 -1488
rect -1530 -1568 -1426 -1552
rect -1530 -1632 -1510 -1568
rect -1446 -1632 -1426 -1568
rect -1530 -1648 -1426 -1632
rect -1530 -1712 -1510 -1648
rect -1446 -1712 -1426 -1648
rect -1530 -1728 -1426 -1712
rect -1530 -1792 -1510 -1728
rect -1446 -1792 -1426 -1728
rect -1530 -1808 -1426 -1792
rect -1530 -1872 -1510 -1808
rect -1446 -1872 -1426 -1808
rect -1530 -1888 -1426 -1872
rect -1530 -1952 -1510 -1888
rect -1446 -1952 -1426 -1888
rect -1530 -1968 -1426 -1952
rect -1530 -2032 -1510 -1968
rect -1446 -2032 -1426 -1968
rect -1530 -2048 -1426 -2032
rect -1530 -2112 -1510 -2048
rect -1446 -2112 -1426 -2048
rect -1530 -2128 -1426 -2112
rect -1530 -2192 -1510 -2128
rect -1446 -2192 -1426 -2128
rect -1530 -2208 -1426 -2192
rect -1530 -2272 -1510 -2208
rect -1446 -2272 -1426 -2208
rect -1530 -2288 -1426 -2272
rect -1530 -2352 -1510 -2288
rect -1446 -2352 -1426 -2288
rect -1530 -2368 -1426 -2352
rect -1530 -2432 -1510 -2368
rect -1446 -2432 -1426 -2368
rect -1530 -2448 -1426 -2432
rect -1530 -2512 -1510 -2448
rect -1446 -2512 -1426 -2448
rect -1530 -2528 -1426 -2512
rect -1530 -2592 -1510 -2528
rect -1446 -2592 -1426 -2528
rect -1530 -2608 -1426 -2592
rect -1530 -2672 -1510 -2608
rect -1446 -2672 -1426 -2608
rect -1530 -2688 -1426 -2672
rect -1530 -2752 -1510 -2688
rect -1446 -2752 -1426 -2688
rect -1530 -2768 -1426 -2752
rect -1530 -2832 -1510 -2768
rect -1446 -2832 -1426 -2768
rect -1530 -2848 -1426 -2832
rect -1530 -2912 -1510 -2848
rect -1446 -2912 -1426 -2848
rect -1530 -2928 -1426 -2912
rect -1530 -2992 -1510 -2928
rect -1446 -2992 -1426 -2928
rect -1530 -3008 -1426 -2992
rect -1530 -3072 -1510 -3008
rect -1446 -3072 -1426 -3008
rect -1530 -3088 -1426 -3072
rect -1530 -3152 -1510 -3088
rect -1446 -3152 -1426 -3088
rect -1530 -3168 -1426 -3152
rect -1530 -3232 -1510 -3168
rect -1446 -3232 -1426 -3168
rect -1530 -3248 -1426 -3232
rect -4142 -3648 -4038 -3312
rect -6754 -3728 -6650 -3712
rect -6754 -3792 -6734 -3728
rect -6670 -3792 -6650 -3728
rect -6754 -3808 -6650 -3792
rect -6754 -3872 -6734 -3808
rect -6670 -3872 -6650 -3808
rect -6754 -3888 -6650 -3872
rect -6754 -3952 -6734 -3888
rect -6670 -3952 -6650 -3888
rect -6754 -3968 -6650 -3952
rect -6754 -4032 -6734 -3968
rect -6670 -4032 -6650 -3968
rect -6754 -4048 -6650 -4032
rect -6754 -4112 -6734 -4048
rect -6670 -4112 -6650 -4048
rect -6754 -4128 -6650 -4112
rect -6754 -4192 -6734 -4128
rect -6670 -4192 -6650 -4128
rect -6754 -4208 -6650 -4192
rect -6754 -4272 -6734 -4208
rect -6670 -4272 -6650 -4208
rect -6754 -4288 -6650 -4272
rect -6754 -4352 -6734 -4288
rect -6670 -4352 -6650 -4288
rect -6754 -4368 -6650 -4352
rect -6754 -4432 -6734 -4368
rect -6670 -4432 -6650 -4368
rect -6754 -4448 -6650 -4432
rect -6754 -4512 -6734 -4448
rect -6670 -4512 -6650 -4448
rect -6754 -4528 -6650 -4512
rect -6754 -4592 -6734 -4528
rect -6670 -4592 -6650 -4528
rect -6754 -4608 -6650 -4592
rect -6754 -4672 -6734 -4608
rect -6670 -4672 -6650 -4608
rect -6754 -4688 -6650 -4672
rect -6754 -4752 -6734 -4688
rect -6670 -4752 -6650 -4688
rect -6754 -4768 -6650 -4752
rect -6754 -4832 -6734 -4768
rect -6670 -4832 -6650 -4768
rect -6754 -4848 -6650 -4832
rect -6754 -4912 -6734 -4848
rect -6670 -4912 -6650 -4848
rect -6754 -4928 -6650 -4912
rect -6754 -4992 -6734 -4928
rect -6670 -4992 -6650 -4928
rect -6754 -5008 -6650 -4992
rect -6754 -5072 -6734 -5008
rect -6670 -5072 -6650 -5008
rect -6754 -5088 -6650 -5072
rect -6754 -5152 -6734 -5088
rect -6670 -5152 -6650 -5088
rect -6754 -5168 -6650 -5152
rect -6754 -5232 -6734 -5168
rect -6670 -5232 -6650 -5168
rect -6754 -5248 -6650 -5232
rect -6754 -5312 -6734 -5248
rect -6670 -5312 -6650 -5248
rect -6754 -5328 -6650 -5312
rect -6754 -5392 -6734 -5328
rect -6670 -5392 -6650 -5328
rect -6754 -5408 -6650 -5392
rect -6754 -5472 -6734 -5408
rect -6670 -5472 -6650 -5408
rect -6754 -5488 -6650 -5472
rect -6754 -5552 -6734 -5488
rect -6670 -5552 -6650 -5488
rect -6754 -5568 -6650 -5552
rect -8034 -5999 -7930 -5601
rect -6754 -5632 -6734 -5568
rect -6670 -5632 -6650 -5568
rect -6331 -3688 -4409 -3679
rect -6331 -5592 -6322 -3688
rect -4418 -5592 -4409 -3688
rect -6331 -5601 -4409 -5592
rect -4142 -3712 -4122 -3648
rect -4058 -3712 -4038 -3648
rect -2810 -3679 -2706 -3281
rect -1530 -3312 -1510 -3248
rect -1446 -3312 -1426 -3248
rect -1107 -1368 815 -1359
rect -1107 -3272 -1098 -1368
rect 806 -3272 815 -1368
rect -1107 -3281 815 -3272
rect 1082 -1392 1102 -1328
rect 1166 -1392 1186 -1328
rect 2414 -1359 2518 -961
rect 3694 -992 3714 -928
rect 3778 -992 3798 -928
rect 4117 952 6039 961
rect 4117 -952 4126 952
rect 6030 -952 6039 952
rect 4117 -961 6039 -952
rect 6306 928 6326 992
rect 6390 928 6410 992
rect 7638 961 7742 1359
rect 8918 1328 8938 1392
rect 9002 1328 9022 1392
rect 8918 992 9022 1328
rect 6306 912 6410 928
rect 6306 848 6326 912
rect 6390 848 6410 912
rect 6306 832 6410 848
rect 6306 768 6326 832
rect 6390 768 6410 832
rect 6306 752 6410 768
rect 6306 688 6326 752
rect 6390 688 6410 752
rect 6306 672 6410 688
rect 6306 608 6326 672
rect 6390 608 6410 672
rect 6306 592 6410 608
rect 6306 528 6326 592
rect 6390 528 6410 592
rect 6306 512 6410 528
rect 6306 448 6326 512
rect 6390 448 6410 512
rect 6306 432 6410 448
rect 6306 368 6326 432
rect 6390 368 6410 432
rect 6306 352 6410 368
rect 6306 288 6326 352
rect 6390 288 6410 352
rect 6306 272 6410 288
rect 6306 208 6326 272
rect 6390 208 6410 272
rect 6306 192 6410 208
rect 6306 128 6326 192
rect 6390 128 6410 192
rect 6306 112 6410 128
rect 6306 48 6326 112
rect 6390 48 6410 112
rect 6306 32 6410 48
rect 6306 -32 6326 32
rect 6390 -32 6410 32
rect 6306 -48 6410 -32
rect 6306 -112 6326 -48
rect 6390 -112 6410 -48
rect 6306 -128 6410 -112
rect 6306 -192 6326 -128
rect 6390 -192 6410 -128
rect 6306 -208 6410 -192
rect 6306 -272 6326 -208
rect 6390 -272 6410 -208
rect 6306 -288 6410 -272
rect 6306 -352 6326 -288
rect 6390 -352 6410 -288
rect 6306 -368 6410 -352
rect 6306 -432 6326 -368
rect 6390 -432 6410 -368
rect 6306 -448 6410 -432
rect 6306 -512 6326 -448
rect 6390 -512 6410 -448
rect 6306 -528 6410 -512
rect 6306 -592 6326 -528
rect 6390 -592 6410 -528
rect 6306 -608 6410 -592
rect 6306 -672 6326 -608
rect 6390 -672 6410 -608
rect 6306 -688 6410 -672
rect 6306 -752 6326 -688
rect 6390 -752 6410 -688
rect 6306 -768 6410 -752
rect 6306 -832 6326 -768
rect 6390 -832 6410 -768
rect 6306 -848 6410 -832
rect 6306 -912 6326 -848
rect 6390 -912 6410 -848
rect 6306 -928 6410 -912
rect 3694 -1328 3798 -992
rect 1082 -1408 1186 -1392
rect 1082 -1472 1102 -1408
rect 1166 -1472 1186 -1408
rect 1082 -1488 1186 -1472
rect 1082 -1552 1102 -1488
rect 1166 -1552 1186 -1488
rect 1082 -1568 1186 -1552
rect 1082 -1632 1102 -1568
rect 1166 -1632 1186 -1568
rect 1082 -1648 1186 -1632
rect 1082 -1712 1102 -1648
rect 1166 -1712 1186 -1648
rect 1082 -1728 1186 -1712
rect 1082 -1792 1102 -1728
rect 1166 -1792 1186 -1728
rect 1082 -1808 1186 -1792
rect 1082 -1872 1102 -1808
rect 1166 -1872 1186 -1808
rect 1082 -1888 1186 -1872
rect 1082 -1952 1102 -1888
rect 1166 -1952 1186 -1888
rect 1082 -1968 1186 -1952
rect 1082 -2032 1102 -1968
rect 1166 -2032 1186 -1968
rect 1082 -2048 1186 -2032
rect 1082 -2112 1102 -2048
rect 1166 -2112 1186 -2048
rect 1082 -2128 1186 -2112
rect 1082 -2192 1102 -2128
rect 1166 -2192 1186 -2128
rect 1082 -2208 1186 -2192
rect 1082 -2272 1102 -2208
rect 1166 -2272 1186 -2208
rect 1082 -2288 1186 -2272
rect 1082 -2352 1102 -2288
rect 1166 -2352 1186 -2288
rect 1082 -2368 1186 -2352
rect 1082 -2432 1102 -2368
rect 1166 -2432 1186 -2368
rect 1082 -2448 1186 -2432
rect 1082 -2512 1102 -2448
rect 1166 -2512 1186 -2448
rect 1082 -2528 1186 -2512
rect 1082 -2592 1102 -2528
rect 1166 -2592 1186 -2528
rect 1082 -2608 1186 -2592
rect 1082 -2672 1102 -2608
rect 1166 -2672 1186 -2608
rect 1082 -2688 1186 -2672
rect 1082 -2752 1102 -2688
rect 1166 -2752 1186 -2688
rect 1082 -2768 1186 -2752
rect 1082 -2832 1102 -2768
rect 1166 -2832 1186 -2768
rect 1082 -2848 1186 -2832
rect 1082 -2912 1102 -2848
rect 1166 -2912 1186 -2848
rect 1082 -2928 1186 -2912
rect 1082 -2992 1102 -2928
rect 1166 -2992 1186 -2928
rect 1082 -3008 1186 -2992
rect 1082 -3072 1102 -3008
rect 1166 -3072 1186 -3008
rect 1082 -3088 1186 -3072
rect 1082 -3152 1102 -3088
rect 1166 -3152 1186 -3088
rect 1082 -3168 1186 -3152
rect 1082 -3232 1102 -3168
rect 1166 -3232 1186 -3168
rect 1082 -3248 1186 -3232
rect -1530 -3648 -1426 -3312
rect -4142 -3728 -4038 -3712
rect -4142 -3792 -4122 -3728
rect -4058 -3792 -4038 -3728
rect -4142 -3808 -4038 -3792
rect -4142 -3872 -4122 -3808
rect -4058 -3872 -4038 -3808
rect -4142 -3888 -4038 -3872
rect -4142 -3952 -4122 -3888
rect -4058 -3952 -4038 -3888
rect -4142 -3968 -4038 -3952
rect -4142 -4032 -4122 -3968
rect -4058 -4032 -4038 -3968
rect -4142 -4048 -4038 -4032
rect -4142 -4112 -4122 -4048
rect -4058 -4112 -4038 -4048
rect -4142 -4128 -4038 -4112
rect -4142 -4192 -4122 -4128
rect -4058 -4192 -4038 -4128
rect -4142 -4208 -4038 -4192
rect -4142 -4272 -4122 -4208
rect -4058 -4272 -4038 -4208
rect -4142 -4288 -4038 -4272
rect -4142 -4352 -4122 -4288
rect -4058 -4352 -4038 -4288
rect -4142 -4368 -4038 -4352
rect -4142 -4432 -4122 -4368
rect -4058 -4432 -4038 -4368
rect -4142 -4448 -4038 -4432
rect -4142 -4512 -4122 -4448
rect -4058 -4512 -4038 -4448
rect -4142 -4528 -4038 -4512
rect -4142 -4592 -4122 -4528
rect -4058 -4592 -4038 -4528
rect -4142 -4608 -4038 -4592
rect -4142 -4672 -4122 -4608
rect -4058 -4672 -4038 -4608
rect -4142 -4688 -4038 -4672
rect -4142 -4752 -4122 -4688
rect -4058 -4752 -4038 -4688
rect -4142 -4768 -4038 -4752
rect -4142 -4832 -4122 -4768
rect -4058 -4832 -4038 -4768
rect -4142 -4848 -4038 -4832
rect -4142 -4912 -4122 -4848
rect -4058 -4912 -4038 -4848
rect -4142 -4928 -4038 -4912
rect -4142 -4992 -4122 -4928
rect -4058 -4992 -4038 -4928
rect -4142 -5008 -4038 -4992
rect -4142 -5072 -4122 -5008
rect -4058 -5072 -4038 -5008
rect -4142 -5088 -4038 -5072
rect -4142 -5152 -4122 -5088
rect -4058 -5152 -4038 -5088
rect -4142 -5168 -4038 -5152
rect -4142 -5232 -4122 -5168
rect -4058 -5232 -4038 -5168
rect -4142 -5248 -4038 -5232
rect -4142 -5312 -4122 -5248
rect -4058 -5312 -4038 -5248
rect -4142 -5328 -4038 -5312
rect -4142 -5392 -4122 -5328
rect -4058 -5392 -4038 -5328
rect -4142 -5408 -4038 -5392
rect -4142 -5472 -4122 -5408
rect -4058 -5472 -4038 -5408
rect -4142 -5488 -4038 -5472
rect -4142 -5552 -4122 -5488
rect -4058 -5552 -4038 -5488
rect -4142 -5568 -4038 -5552
rect -6754 -5968 -6650 -5632
rect -8943 -6008 -7021 -5999
rect -8943 -7912 -8934 -6008
rect -7030 -7912 -7021 -6008
rect -8943 -7921 -7021 -7912
rect -6754 -6032 -6734 -5968
rect -6670 -6032 -6650 -5968
rect -5422 -5999 -5318 -5601
rect -4142 -5632 -4122 -5568
rect -4058 -5632 -4038 -5568
rect -3719 -3688 -1797 -3679
rect -3719 -5592 -3710 -3688
rect -1806 -5592 -1797 -3688
rect -3719 -5601 -1797 -5592
rect -1530 -3712 -1510 -3648
rect -1446 -3712 -1426 -3648
rect -198 -3679 -94 -3281
rect 1082 -3312 1102 -3248
rect 1166 -3312 1186 -3248
rect 1505 -1368 3427 -1359
rect 1505 -3272 1514 -1368
rect 3418 -3272 3427 -1368
rect 1505 -3281 3427 -3272
rect 3694 -1392 3714 -1328
rect 3778 -1392 3798 -1328
rect 5026 -1359 5130 -961
rect 6306 -992 6326 -928
rect 6390 -992 6410 -928
rect 6729 952 8651 961
rect 6729 -952 6738 952
rect 8642 -952 8651 952
rect 6729 -961 8651 -952
rect 8918 928 8938 992
rect 9002 928 9022 992
rect 8918 912 9022 928
rect 8918 848 8938 912
rect 9002 848 9022 912
rect 8918 832 9022 848
rect 8918 768 8938 832
rect 9002 768 9022 832
rect 8918 752 9022 768
rect 8918 688 8938 752
rect 9002 688 9022 752
rect 8918 672 9022 688
rect 8918 608 8938 672
rect 9002 608 9022 672
rect 8918 592 9022 608
rect 8918 528 8938 592
rect 9002 528 9022 592
rect 8918 512 9022 528
rect 8918 448 8938 512
rect 9002 448 9022 512
rect 8918 432 9022 448
rect 8918 368 8938 432
rect 9002 368 9022 432
rect 8918 352 9022 368
rect 8918 288 8938 352
rect 9002 288 9022 352
rect 8918 272 9022 288
rect 8918 208 8938 272
rect 9002 208 9022 272
rect 8918 192 9022 208
rect 8918 128 8938 192
rect 9002 128 9022 192
rect 8918 112 9022 128
rect 8918 48 8938 112
rect 9002 48 9022 112
rect 8918 32 9022 48
rect 8918 -32 8938 32
rect 9002 -32 9022 32
rect 8918 -48 9022 -32
rect 8918 -112 8938 -48
rect 9002 -112 9022 -48
rect 8918 -128 9022 -112
rect 8918 -192 8938 -128
rect 9002 -192 9022 -128
rect 8918 -208 9022 -192
rect 8918 -272 8938 -208
rect 9002 -272 9022 -208
rect 8918 -288 9022 -272
rect 8918 -352 8938 -288
rect 9002 -352 9022 -288
rect 8918 -368 9022 -352
rect 8918 -432 8938 -368
rect 9002 -432 9022 -368
rect 8918 -448 9022 -432
rect 8918 -512 8938 -448
rect 9002 -512 9022 -448
rect 8918 -528 9022 -512
rect 8918 -592 8938 -528
rect 9002 -592 9022 -528
rect 8918 -608 9022 -592
rect 8918 -672 8938 -608
rect 9002 -672 9022 -608
rect 8918 -688 9022 -672
rect 8918 -752 8938 -688
rect 9002 -752 9022 -688
rect 8918 -768 9022 -752
rect 8918 -832 8938 -768
rect 9002 -832 9022 -768
rect 8918 -848 9022 -832
rect 8918 -912 8938 -848
rect 9002 -912 9022 -848
rect 8918 -928 9022 -912
rect 6306 -1328 6410 -992
rect 3694 -1408 3798 -1392
rect 3694 -1472 3714 -1408
rect 3778 -1472 3798 -1408
rect 3694 -1488 3798 -1472
rect 3694 -1552 3714 -1488
rect 3778 -1552 3798 -1488
rect 3694 -1568 3798 -1552
rect 3694 -1632 3714 -1568
rect 3778 -1632 3798 -1568
rect 3694 -1648 3798 -1632
rect 3694 -1712 3714 -1648
rect 3778 -1712 3798 -1648
rect 3694 -1728 3798 -1712
rect 3694 -1792 3714 -1728
rect 3778 -1792 3798 -1728
rect 3694 -1808 3798 -1792
rect 3694 -1872 3714 -1808
rect 3778 -1872 3798 -1808
rect 3694 -1888 3798 -1872
rect 3694 -1952 3714 -1888
rect 3778 -1952 3798 -1888
rect 3694 -1968 3798 -1952
rect 3694 -2032 3714 -1968
rect 3778 -2032 3798 -1968
rect 3694 -2048 3798 -2032
rect 3694 -2112 3714 -2048
rect 3778 -2112 3798 -2048
rect 3694 -2128 3798 -2112
rect 3694 -2192 3714 -2128
rect 3778 -2192 3798 -2128
rect 3694 -2208 3798 -2192
rect 3694 -2272 3714 -2208
rect 3778 -2272 3798 -2208
rect 3694 -2288 3798 -2272
rect 3694 -2352 3714 -2288
rect 3778 -2352 3798 -2288
rect 3694 -2368 3798 -2352
rect 3694 -2432 3714 -2368
rect 3778 -2432 3798 -2368
rect 3694 -2448 3798 -2432
rect 3694 -2512 3714 -2448
rect 3778 -2512 3798 -2448
rect 3694 -2528 3798 -2512
rect 3694 -2592 3714 -2528
rect 3778 -2592 3798 -2528
rect 3694 -2608 3798 -2592
rect 3694 -2672 3714 -2608
rect 3778 -2672 3798 -2608
rect 3694 -2688 3798 -2672
rect 3694 -2752 3714 -2688
rect 3778 -2752 3798 -2688
rect 3694 -2768 3798 -2752
rect 3694 -2832 3714 -2768
rect 3778 -2832 3798 -2768
rect 3694 -2848 3798 -2832
rect 3694 -2912 3714 -2848
rect 3778 -2912 3798 -2848
rect 3694 -2928 3798 -2912
rect 3694 -2992 3714 -2928
rect 3778 -2992 3798 -2928
rect 3694 -3008 3798 -2992
rect 3694 -3072 3714 -3008
rect 3778 -3072 3798 -3008
rect 3694 -3088 3798 -3072
rect 3694 -3152 3714 -3088
rect 3778 -3152 3798 -3088
rect 3694 -3168 3798 -3152
rect 3694 -3232 3714 -3168
rect 3778 -3232 3798 -3168
rect 3694 -3248 3798 -3232
rect 1082 -3648 1186 -3312
rect -1530 -3728 -1426 -3712
rect -1530 -3792 -1510 -3728
rect -1446 -3792 -1426 -3728
rect -1530 -3808 -1426 -3792
rect -1530 -3872 -1510 -3808
rect -1446 -3872 -1426 -3808
rect -1530 -3888 -1426 -3872
rect -1530 -3952 -1510 -3888
rect -1446 -3952 -1426 -3888
rect -1530 -3968 -1426 -3952
rect -1530 -4032 -1510 -3968
rect -1446 -4032 -1426 -3968
rect -1530 -4048 -1426 -4032
rect -1530 -4112 -1510 -4048
rect -1446 -4112 -1426 -4048
rect -1530 -4128 -1426 -4112
rect -1530 -4192 -1510 -4128
rect -1446 -4192 -1426 -4128
rect -1530 -4208 -1426 -4192
rect -1530 -4272 -1510 -4208
rect -1446 -4272 -1426 -4208
rect -1530 -4288 -1426 -4272
rect -1530 -4352 -1510 -4288
rect -1446 -4352 -1426 -4288
rect -1530 -4368 -1426 -4352
rect -1530 -4432 -1510 -4368
rect -1446 -4432 -1426 -4368
rect -1530 -4448 -1426 -4432
rect -1530 -4512 -1510 -4448
rect -1446 -4512 -1426 -4448
rect -1530 -4528 -1426 -4512
rect -1530 -4592 -1510 -4528
rect -1446 -4592 -1426 -4528
rect -1530 -4608 -1426 -4592
rect -1530 -4672 -1510 -4608
rect -1446 -4672 -1426 -4608
rect -1530 -4688 -1426 -4672
rect -1530 -4752 -1510 -4688
rect -1446 -4752 -1426 -4688
rect -1530 -4768 -1426 -4752
rect -1530 -4832 -1510 -4768
rect -1446 -4832 -1426 -4768
rect -1530 -4848 -1426 -4832
rect -1530 -4912 -1510 -4848
rect -1446 -4912 -1426 -4848
rect -1530 -4928 -1426 -4912
rect -1530 -4992 -1510 -4928
rect -1446 -4992 -1426 -4928
rect -1530 -5008 -1426 -4992
rect -1530 -5072 -1510 -5008
rect -1446 -5072 -1426 -5008
rect -1530 -5088 -1426 -5072
rect -1530 -5152 -1510 -5088
rect -1446 -5152 -1426 -5088
rect -1530 -5168 -1426 -5152
rect -1530 -5232 -1510 -5168
rect -1446 -5232 -1426 -5168
rect -1530 -5248 -1426 -5232
rect -1530 -5312 -1510 -5248
rect -1446 -5312 -1426 -5248
rect -1530 -5328 -1426 -5312
rect -1530 -5392 -1510 -5328
rect -1446 -5392 -1426 -5328
rect -1530 -5408 -1426 -5392
rect -1530 -5472 -1510 -5408
rect -1446 -5472 -1426 -5408
rect -1530 -5488 -1426 -5472
rect -1530 -5552 -1510 -5488
rect -1446 -5552 -1426 -5488
rect -1530 -5568 -1426 -5552
rect -4142 -5968 -4038 -5632
rect -6754 -6048 -6650 -6032
rect -6754 -6112 -6734 -6048
rect -6670 -6112 -6650 -6048
rect -6754 -6128 -6650 -6112
rect -6754 -6192 -6734 -6128
rect -6670 -6192 -6650 -6128
rect -6754 -6208 -6650 -6192
rect -6754 -6272 -6734 -6208
rect -6670 -6272 -6650 -6208
rect -6754 -6288 -6650 -6272
rect -6754 -6352 -6734 -6288
rect -6670 -6352 -6650 -6288
rect -6754 -6368 -6650 -6352
rect -6754 -6432 -6734 -6368
rect -6670 -6432 -6650 -6368
rect -6754 -6448 -6650 -6432
rect -6754 -6512 -6734 -6448
rect -6670 -6512 -6650 -6448
rect -6754 -6528 -6650 -6512
rect -6754 -6592 -6734 -6528
rect -6670 -6592 -6650 -6528
rect -6754 -6608 -6650 -6592
rect -6754 -6672 -6734 -6608
rect -6670 -6672 -6650 -6608
rect -6754 -6688 -6650 -6672
rect -6754 -6752 -6734 -6688
rect -6670 -6752 -6650 -6688
rect -6754 -6768 -6650 -6752
rect -6754 -6832 -6734 -6768
rect -6670 -6832 -6650 -6768
rect -6754 -6848 -6650 -6832
rect -6754 -6912 -6734 -6848
rect -6670 -6912 -6650 -6848
rect -6754 -6928 -6650 -6912
rect -6754 -6992 -6734 -6928
rect -6670 -6992 -6650 -6928
rect -6754 -7008 -6650 -6992
rect -6754 -7072 -6734 -7008
rect -6670 -7072 -6650 -7008
rect -6754 -7088 -6650 -7072
rect -6754 -7152 -6734 -7088
rect -6670 -7152 -6650 -7088
rect -6754 -7168 -6650 -7152
rect -6754 -7232 -6734 -7168
rect -6670 -7232 -6650 -7168
rect -6754 -7248 -6650 -7232
rect -6754 -7312 -6734 -7248
rect -6670 -7312 -6650 -7248
rect -6754 -7328 -6650 -7312
rect -6754 -7392 -6734 -7328
rect -6670 -7392 -6650 -7328
rect -6754 -7408 -6650 -7392
rect -6754 -7472 -6734 -7408
rect -6670 -7472 -6650 -7408
rect -6754 -7488 -6650 -7472
rect -6754 -7552 -6734 -7488
rect -6670 -7552 -6650 -7488
rect -6754 -7568 -6650 -7552
rect -6754 -7632 -6734 -7568
rect -6670 -7632 -6650 -7568
rect -6754 -7648 -6650 -7632
rect -6754 -7712 -6734 -7648
rect -6670 -7712 -6650 -7648
rect -6754 -7728 -6650 -7712
rect -6754 -7792 -6734 -7728
rect -6670 -7792 -6650 -7728
rect -6754 -7808 -6650 -7792
rect -6754 -7872 -6734 -7808
rect -6670 -7872 -6650 -7808
rect -6754 -7888 -6650 -7872
rect -8034 -8120 -7930 -7921
rect -6754 -7952 -6734 -7888
rect -6670 -7952 -6650 -7888
rect -6331 -6008 -4409 -5999
rect -6331 -7912 -6322 -6008
rect -4418 -7912 -4409 -6008
rect -6331 -7921 -4409 -7912
rect -4142 -6032 -4122 -5968
rect -4058 -6032 -4038 -5968
rect -2810 -5999 -2706 -5601
rect -1530 -5632 -1510 -5568
rect -1446 -5632 -1426 -5568
rect -1107 -3688 815 -3679
rect -1107 -5592 -1098 -3688
rect 806 -5592 815 -3688
rect -1107 -5601 815 -5592
rect 1082 -3712 1102 -3648
rect 1166 -3712 1186 -3648
rect 2414 -3679 2518 -3281
rect 3694 -3312 3714 -3248
rect 3778 -3312 3798 -3248
rect 4117 -1368 6039 -1359
rect 4117 -3272 4126 -1368
rect 6030 -3272 6039 -1368
rect 4117 -3281 6039 -3272
rect 6306 -1392 6326 -1328
rect 6390 -1392 6410 -1328
rect 7638 -1359 7742 -961
rect 8918 -992 8938 -928
rect 9002 -992 9022 -928
rect 8918 -1328 9022 -992
rect 6306 -1408 6410 -1392
rect 6306 -1472 6326 -1408
rect 6390 -1472 6410 -1408
rect 6306 -1488 6410 -1472
rect 6306 -1552 6326 -1488
rect 6390 -1552 6410 -1488
rect 6306 -1568 6410 -1552
rect 6306 -1632 6326 -1568
rect 6390 -1632 6410 -1568
rect 6306 -1648 6410 -1632
rect 6306 -1712 6326 -1648
rect 6390 -1712 6410 -1648
rect 6306 -1728 6410 -1712
rect 6306 -1792 6326 -1728
rect 6390 -1792 6410 -1728
rect 6306 -1808 6410 -1792
rect 6306 -1872 6326 -1808
rect 6390 -1872 6410 -1808
rect 6306 -1888 6410 -1872
rect 6306 -1952 6326 -1888
rect 6390 -1952 6410 -1888
rect 6306 -1968 6410 -1952
rect 6306 -2032 6326 -1968
rect 6390 -2032 6410 -1968
rect 6306 -2048 6410 -2032
rect 6306 -2112 6326 -2048
rect 6390 -2112 6410 -2048
rect 6306 -2128 6410 -2112
rect 6306 -2192 6326 -2128
rect 6390 -2192 6410 -2128
rect 6306 -2208 6410 -2192
rect 6306 -2272 6326 -2208
rect 6390 -2272 6410 -2208
rect 6306 -2288 6410 -2272
rect 6306 -2352 6326 -2288
rect 6390 -2352 6410 -2288
rect 6306 -2368 6410 -2352
rect 6306 -2432 6326 -2368
rect 6390 -2432 6410 -2368
rect 6306 -2448 6410 -2432
rect 6306 -2512 6326 -2448
rect 6390 -2512 6410 -2448
rect 6306 -2528 6410 -2512
rect 6306 -2592 6326 -2528
rect 6390 -2592 6410 -2528
rect 6306 -2608 6410 -2592
rect 6306 -2672 6326 -2608
rect 6390 -2672 6410 -2608
rect 6306 -2688 6410 -2672
rect 6306 -2752 6326 -2688
rect 6390 -2752 6410 -2688
rect 6306 -2768 6410 -2752
rect 6306 -2832 6326 -2768
rect 6390 -2832 6410 -2768
rect 6306 -2848 6410 -2832
rect 6306 -2912 6326 -2848
rect 6390 -2912 6410 -2848
rect 6306 -2928 6410 -2912
rect 6306 -2992 6326 -2928
rect 6390 -2992 6410 -2928
rect 6306 -3008 6410 -2992
rect 6306 -3072 6326 -3008
rect 6390 -3072 6410 -3008
rect 6306 -3088 6410 -3072
rect 6306 -3152 6326 -3088
rect 6390 -3152 6410 -3088
rect 6306 -3168 6410 -3152
rect 6306 -3232 6326 -3168
rect 6390 -3232 6410 -3168
rect 6306 -3248 6410 -3232
rect 3694 -3648 3798 -3312
rect 1082 -3728 1186 -3712
rect 1082 -3792 1102 -3728
rect 1166 -3792 1186 -3728
rect 1082 -3808 1186 -3792
rect 1082 -3872 1102 -3808
rect 1166 -3872 1186 -3808
rect 1082 -3888 1186 -3872
rect 1082 -3952 1102 -3888
rect 1166 -3952 1186 -3888
rect 1082 -3968 1186 -3952
rect 1082 -4032 1102 -3968
rect 1166 -4032 1186 -3968
rect 1082 -4048 1186 -4032
rect 1082 -4112 1102 -4048
rect 1166 -4112 1186 -4048
rect 1082 -4128 1186 -4112
rect 1082 -4192 1102 -4128
rect 1166 -4192 1186 -4128
rect 1082 -4208 1186 -4192
rect 1082 -4272 1102 -4208
rect 1166 -4272 1186 -4208
rect 1082 -4288 1186 -4272
rect 1082 -4352 1102 -4288
rect 1166 -4352 1186 -4288
rect 1082 -4368 1186 -4352
rect 1082 -4432 1102 -4368
rect 1166 -4432 1186 -4368
rect 1082 -4448 1186 -4432
rect 1082 -4512 1102 -4448
rect 1166 -4512 1186 -4448
rect 1082 -4528 1186 -4512
rect 1082 -4592 1102 -4528
rect 1166 -4592 1186 -4528
rect 1082 -4608 1186 -4592
rect 1082 -4672 1102 -4608
rect 1166 -4672 1186 -4608
rect 1082 -4688 1186 -4672
rect 1082 -4752 1102 -4688
rect 1166 -4752 1186 -4688
rect 1082 -4768 1186 -4752
rect 1082 -4832 1102 -4768
rect 1166 -4832 1186 -4768
rect 1082 -4848 1186 -4832
rect 1082 -4912 1102 -4848
rect 1166 -4912 1186 -4848
rect 1082 -4928 1186 -4912
rect 1082 -4992 1102 -4928
rect 1166 -4992 1186 -4928
rect 1082 -5008 1186 -4992
rect 1082 -5072 1102 -5008
rect 1166 -5072 1186 -5008
rect 1082 -5088 1186 -5072
rect 1082 -5152 1102 -5088
rect 1166 -5152 1186 -5088
rect 1082 -5168 1186 -5152
rect 1082 -5232 1102 -5168
rect 1166 -5232 1186 -5168
rect 1082 -5248 1186 -5232
rect 1082 -5312 1102 -5248
rect 1166 -5312 1186 -5248
rect 1082 -5328 1186 -5312
rect 1082 -5392 1102 -5328
rect 1166 -5392 1186 -5328
rect 1082 -5408 1186 -5392
rect 1082 -5472 1102 -5408
rect 1166 -5472 1186 -5408
rect 1082 -5488 1186 -5472
rect 1082 -5552 1102 -5488
rect 1166 -5552 1186 -5488
rect 1082 -5568 1186 -5552
rect -1530 -5968 -1426 -5632
rect -4142 -6048 -4038 -6032
rect -4142 -6112 -4122 -6048
rect -4058 -6112 -4038 -6048
rect -4142 -6128 -4038 -6112
rect -4142 -6192 -4122 -6128
rect -4058 -6192 -4038 -6128
rect -4142 -6208 -4038 -6192
rect -4142 -6272 -4122 -6208
rect -4058 -6272 -4038 -6208
rect -4142 -6288 -4038 -6272
rect -4142 -6352 -4122 -6288
rect -4058 -6352 -4038 -6288
rect -4142 -6368 -4038 -6352
rect -4142 -6432 -4122 -6368
rect -4058 -6432 -4038 -6368
rect -4142 -6448 -4038 -6432
rect -4142 -6512 -4122 -6448
rect -4058 -6512 -4038 -6448
rect -4142 -6528 -4038 -6512
rect -4142 -6592 -4122 -6528
rect -4058 -6592 -4038 -6528
rect -4142 -6608 -4038 -6592
rect -4142 -6672 -4122 -6608
rect -4058 -6672 -4038 -6608
rect -4142 -6688 -4038 -6672
rect -4142 -6752 -4122 -6688
rect -4058 -6752 -4038 -6688
rect -4142 -6768 -4038 -6752
rect -4142 -6832 -4122 -6768
rect -4058 -6832 -4038 -6768
rect -4142 -6848 -4038 -6832
rect -4142 -6912 -4122 -6848
rect -4058 -6912 -4038 -6848
rect -4142 -6928 -4038 -6912
rect -4142 -6992 -4122 -6928
rect -4058 -6992 -4038 -6928
rect -4142 -7008 -4038 -6992
rect -4142 -7072 -4122 -7008
rect -4058 -7072 -4038 -7008
rect -4142 -7088 -4038 -7072
rect -4142 -7152 -4122 -7088
rect -4058 -7152 -4038 -7088
rect -4142 -7168 -4038 -7152
rect -4142 -7232 -4122 -7168
rect -4058 -7232 -4038 -7168
rect -4142 -7248 -4038 -7232
rect -4142 -7312 -4122 -7248
rect -4058 -7312 -4038 -7248
rect -4142 -7328 -4038 -7312
rect -4142 -7392 -4122 -7328
rect -4058 -7392 -4038 -7328
rect -4142 -7408 -4038 -7392
rect -4142 -7472 -4122 -7408
rect -4058 -7472 -4038 -7408
rect -4142 -7488 -4038 -7472
rect -4142 -7552 -4122 -7488
rect -4058 -7552 -4038 -7488
rect -4142 -7568 -4038 -7552
rect -4142 -7632 -4122 -7568
rect -4058 -7632 -4038 -7568
rect -4142 -7648 -4038 -7632
rect -4142 -7712 -4122 -7648
rect -4058 -7712 -4038 -7648
rect -4142 -7728 -4038 -7712
rect -4142 -7792 -4122 -7728
rect -4058 -7792 -4038 -7728
rect -4142 -7808 -4038 -7792
rect -4142 -7872 -4122 -7808
rect -4058 -7872 -4038 -7808
rect -4142 -7888 -4038 -7872
rect -6754 -8120 -6650 -7952
rect -5422 -8120 -5318 -7921
rect -4142 -7952 -4122 -7888
rect -4058 -7952 -4038 -7888
rect -3719 -6008 -1797 -5999
rect -3719 -7912 -3710 -6008
rect -1806 -7912 -1797 -6008
rect -3719 -7921 -1797 -7912
rect -1530 -6032 -1510 -5968
rect -1446 -6032 -1426 -5968
rect -198 -5999 -94 -5601
rect 1082 -5632 1102 -5568
rect 1166 -5632 1186 -5568
rect 1505 -3688 3427 -3679
rect 1505 -5592 1514 -3688
rect 3418 -5592 3427 -3688
rect 1505 -5601 3427 -5592
rect 3694 -3712 3714 -3648
rect 3778 -3712 3798 -3648
rect 5026 -3679 5130 -3281
rect 6306 -3312 6326 -3248
rect 6390 -3312 6410 -3248
rect 6729 -1368 8651 -1359
rect 6729 -3272 6738 -1368
rect 8642 -3272 8651 -1368
rect 6729 -3281 8651 -3272
rect 8918 -1392 8938 -1328
rect 9002 -1392 9022 -1328
rect 8918 -1408 9022 -1392
rect 8918 -1472 8938 -1408
rect 9002 -1472 9022 -1408
rect 8918 -1488 9022 -1472
rect 8918 -1552 8938 -1488
rect 9002 -1552 9022 -1488
rect 8918 -1568 9022 -1552
rect 8918 -1632 8938 -1568
rect 9002 -1632 9022 -1568
rect 8918 -1648 9022 -1632
rect 8918 -1712 8938 -1648
rect 9002 -1712 9022 -1648
rect 8918 -1728 9022 -1712
rect 8918 -1792 8938 -1728
rect 9002 -1792 9022 -1728
rect 8918 -1808 9022 -1792
rect 8918 -1872 8938 -1808
rect 9002 -1872 9022 -1808
rect 8918 -1888 9022 -1872
rect 8918 -1952 8938 -1888
rect 9002 -1952 9022 -1888
rect 8918 -1968 9022 -1952
rect 8918 -2032 8938 -1968
rect 9002 -2032 9022 -1968
rect 8918 -2048 9022 -2032
rect 8918 -2112 8938 -2048
rect 9002 -2112 9022 -2048
rect 8918 -2128 9022 -2112
rect 8918 -2192 8938 -2128
rect 9002 -2192 9022 -2128
rect 8918 -2208 9022 -2192
rect 8918 -2272 8938 -2208
rect 9002 -2272 9022 -2208
rect 8918 -2288 9022 -2272
rect 8918 -2352 8938 -2288
rect 9002 -2352 9022 -2288
rect 8918 -2368 9022 -2352
rect 8918 -2432 8938 -2368
rect 9002 -2432 9022 -2368
rect 8918 -2448 9022 -2432
rect 8918 -2512 8938 -2448
rect 9002 -2512 9022 -2448
rect 8918 -2528 9022 -2512
rect 8918 -2592 8938 -2528
rect 9002 -2592 9022 -2528
rect 8918 -2608 9022 -2592
rect 8918 -2672 8938 -2608
rect 9002 -2672 9022 -2608
rect 8918 -2688 9022 -2672
rect 8918 -2752 8938 -2688
rect 9002 -2752 9022 -2688
rect 8918 -2768 9022 -2752
rect 8918 -2832 8938 -2768
rect 9002 -2832 9022 -2768
rect 8918 -2848 9022 -2832
rect 8918 -2912 8938 -2848
rect 9002 -2912 9022 -2848
rect 8918 -2928 9022 -2912
rect 8918 -2992 8938 -2928
rect 9002 -2992 9022 -2928
rect 8918 -3008 9022 -2992
rect 8918 -3072 8938 -3008
rect 9002 -3072 9022 -3008
rect 8918 -3088 9022 -3072
rect 8918 -3152 8938 -3088
rect 9002 -3152 9022 -3088
rect 8918 -3168 9022 -3152
rect 8918 -3232 8938 -3168
rect 9002 -3232 9022 -3168
rect 8918 -3248 9022 -3232
rect 6306 -3648 6410 -3312
rect 3694 -3728 3798 -3712
rect 3694 -3792 3714 -3728
rect 3778 -3792 3798 -3728
rect 3694 -3808 3798 -3792
rect 3694 -3872 3714 -3808
rect 3778 -3872 3798 -3808
rect 3694 -3888 3798 -3872
rect 3694 -3952 3714 -3888
rect 3778 -3952 3798 -3888
rect 3694 -3968 3798 -3952
rect 3694 -4032 3714 -3968
rect 3778 -4032 3798 -3968
rect 3694 -4048 3798 -4032
rect 3694 -4112 3714 -4048
rect 3778 -4112 3798 -4048
rect 3694 -4128 3798 -4112
rect 3694 -4192 3714 -4128
rect 3778 -4192 3798 -4128
rect 3694 -4208 3798 -4192
rect 3694 -4272 3714 -4208
rect 3778 -4272 3798 -4208
rect 3694 -4288 3798 -4272
rect 3694 -4352 3714 -4288
rect 3778 -4352 3798 -4288
rect 3694 -4368 3798 -4352
rect 3694 -4432 3714 -4368
rect 3778 -4432 3798 -4368
rect 3694 -4448 3798 -4432
rect 3694 -4512 3714 -4448
rect 3778 -4512 3798 -4448
rect 3694 -4528 3798 -4512
rect 3694 -4592 3714 -4528
rect 3778 -4592 3798 -4528
rect 3694 -4608 3798 -4592
rect 3694 -4672 3714 -4608
rect 3778 -4672 3798 -4608
rect 3694 -4688 3798 -4672
rect 3694 -4752 3714 -4688
rect 3778 -4752 3798 -4688
rect 3694 -4768 3798 -4752
rect 3694 -4832 3714 -4768
rect 3778 -4832 3798 -4768
rect 3694 -4848 3798 -4832
rect 3694 -4912 3714 -4848
rect 3778 -4912 3798 -4848
rect 3694 -4928 3798 -4912
rect 3694 -4992 3714 -4928
rect 3778 -4992 3798 -4928
rect 3694 -5008 3798 -4992
rect 3694 -5072 3714 -5008
rect 3778 -5072 3798 -5008
rect 3694 -5088 3798 -5072
rect 3694 -5152 3714 -5088
rect 3778 -5152 3798 -5088
rect 3694 -5168 3798 -5152
rect 3694 -5232 3714 -5168
rect 3778 -5232 3798 -5168
rect 3694 -5248 3798 -5232
rect 3694 -5312 3714 -5248
rect 3778 -5312 3798 -5248
rect 3694 -5328 3798 -5312
rect 3694 -5392 3714 -5328
rect 3778 -5392 3798 -5328
rect 3694 -5408 3798 -5392
rect 3694 -5472 3714 -5408
rect 3778 -5472 3798 -5408
rect 3694 -5488 3798 -5472
rect 3694 -5552 3714 -5488
rect 3778 -5552 3798 -5488
rect 3694 -5568 3798 -5552
rect 1082 -5968 1186 -5632
rect -1530 -6048 -1426 -6032
rect -1530 -6112 -1510 -6048
rect -1446 -6112 -1426 -6048
rect -1530 -6128 -1426 -6112
rect -1530 -6192 -1510 -6128
rect -1446 -6192 -1426 -6128
rect -1530 -6208 -1426 -6192
rect -1530 -6272 -1510 -6208
rect -1446 -6272 -1426 -6208
rect -1530 -6288 -1426 -6272
rect -1530 -6352 -1510 -6288
rect -1446 -6352 -1426 -6288
rect -1530 -6368 -1426 -6352
rect -1530 -6432 -1510 -6368
rect -1446 -6432 -1426 -6368
rect -1530 -6448 -1426 -6432
rect -1530 -6512 -1510 -6448
rect -1446 -6512 -1426 -6448
rect -1530 -6528 -1426 -6512
rect -1530 -6592 -1510 -6528
rect -1446 -6592 -1426 -6528
rect -1530 -6608 -1426 -6592
rect -1530 -6672 -1510 -6608
rect -1446 -6672 -1426 -6608
rect -1530 -6688 -1426 -6672
rect -1530 -6752 -1510 -6688
rect -1446 -6752 -1426 -6688
rect -1530 -6768 -1426 -6752
rect -1530 -6832 -1510 -6768
rect -1446 -6832 -1426 -6768
rect -1530 -6848 -1426 -6832
rect -1530 -6912 -1510 -6848
rect -1446 -6912 -1426 -6848
rect -1530 -6928 -1426 -6912
rect -1530 -6992 -1510 -6928
rect -1446 -6992 -1426 -6928
rect -1530 -7008 -1426 -6992
rect -1530 -7072 -1510 -7008
rect -1446 -7072 -1426 -7008
rect -1530 -7088 -1426 -7072
rect -1530 -7152 -1510 -7088
rect -1446 -7152 -1426 -7088
rect -1530 -7168 -1426 -7152
rect -1530 -7232 -1510 -7168
rect -1446 -7232 -1426 -7168
rect -1530 -7248 -1426 -7232
rect -1530 -7312 -1510 -7248
rect -1446 -7312 -1426 -7248
rect -1530 -7328 -1426 -7312
rect -1530 -7392 -1510 -7328
rect -1446 -7392 -1426 -7328
rect -1530 -7408 -1426 -7392
rect -1530 -7472 -1510 -7408
rect -1446 -7472 -1426 -7408
rect -1530 -7488 -1426 -7472
rect -1530 -7552 -1510 -7488
rect -1446 -7552 -1426 -7488
rect -1530 -7568 -1426 -7552
rect -1530 -7632 -1510 -7568
rect -1446 -7632 -1426 -7568
rect -1530 -7648 -1426 -7632
rect -1530 -7712 -1510 -7648
rect -1446 -7712 -1426 -7648
rect -1530 -7728 -1426 -7712
rect -1530 -7792 -1510 -7728
rect -1446 -7792 -1426 -7728
rect -1530 -7808 -1426 -7792
rect -1530 -7872 -1510 -7808
rect -1446 -7872 -1426 -7808
rect -1530 -7888 -1426 -7872
rect -4142 -8120 -4038 -7952
rect -2810 -8120 -2706 -7921
rect -1530 -7952 -1510 -7888
rect -1446 -7952 -1426 -7888
rect -1107 -6008 815 -5999
rect -1107 -7912 -1098 -6008
rect 806 -7912 815 -6008
rect -1107 -7921 815 -7912
rect 1082 -6032 1102 -5968
rect 1166 -6032 1186 -5968
rect 2414 -5999 2518 -5601
rect 3694 -5632 3714 -5568
rect 3778 -5632 3798 -5568
rect 4117 -3688 6039 -3679
rect 4117 -5592 4126 -3688
rect 6030 -5592 6039 -3688
rect 4117 -5601 6039 -5592
rect 6306 -3712 6326 -3648
rect 6390 -3712 6410 -3648
rect 7638 -3679 7742 -3281
rect 8918 -3312 8938 -3248
rect 9002 -3312 9022 -3248
rect 8918 -3648 9022 -3312
rect 6306 -3728 6410 -3712
rect 6306 -3792 6326 -3728
rect 6390 -3792 6410 -3728
rect 6306 -3808 6410 -3792
rect 6306 -3872 6326 -3808
rect 6390 -3872 6410 -3808
rect 6306 -3888 6410 -3872
rect 6306 -3952 6326 -3888
rect 6390 -3952 6410 -3888
rect 6306 -3968 6410 -3952
rect 6306 -4032 6326 -3968
rect 6390 -4032 6410 -3968
rect 6306 -4048 6410 -4032
rect 6306 -4112 6326 -4048
rect 6390 -4112 6410 -4048
rect 6306 -4128 6410 -4112
rect 6306 -4192 6326 -4128
rect 6390 -4192 6410 -4128
rect 6306 -4208 6410 -4192
rect 6306 -4272 6326 -4208
rect 6390 -4272 6410 -4208
rect 6306 -4288 6410 -4272
rect 6306 -4352 6326 -4288
rect 6390 -4352 6410 -4288
rect 6306 -4368 6410 -4352
rect 6306 -4432 6326 -4368
rect 6390 -4432 6410 -4368
rect 6306 -4448 6410 -4432
rect 6306 -4512 6326 -4448
rect 6390 -4512 6410 -4448
rect 6306 -4528 6410 -4512
rect 6306 -4592 6326 -4528
rect 6390 -4592 6410 -4528
rect 6306 -4608 6410 -4592
rect 6306 -4672 6326 -4608
rect 6390 -4672 6410 -4608
rect 6306 -4688 6410 -4672
rect 6306 -4752 6326 -4688
rect 6390 -4752 6410 -4688
rect 6306 -4768 6410 -4752
rect 6306 -4832 6326 -4768
rect 6390 -4832 6410 -4768
rect 6306 -4848 6410 -4832
rect 6306 -4912 6326 -4848
rect 6390 -4912 6410 -4848
rect 6306 -4928 6410 -4912
rect 6306 -4992 6326 -4928
rect 6390 -4992 6410 -4928
rect 6306 -5008 6410 -4992
rect 6306 -5072 6326 -5008
rect 6390 -5072 6410 -5008
rect 6306 -5088 6410 -5072
rect 6306 -5152 6326 -5088
rect 6390 -5152 6410 -5088
rect 6306 -5168 6410 -5152
rect 6306 -5232 6326 -5168
rect 6390 -5232 6410 -5168
rect 6306 -5248 6410 -5232
rect 6306 -5312 6326 -5248
rect 6390 -5312 6410 -5248
rect 6306 -5328 6410 -5312
rect 6306 -5392 6326 -5328
rect 6390 -5392 6410 -5328
rect 6306 -5408 6410 -5392
rect 6306 -5472 6326 -5408
rect 6390 -5472 6410 -5408
rect 6306 -5488 6410 -5472
rect 6306 -5552 6326 -5488
rect 6390 -5552 6410 -5488
rect 6306 -5568 6410 -5552
rect 3694 -5968 3798 -5632
rect 1082 -6048 1186 -6032
rect 1082 -6112 1102 -6048
rect 1166 -6112 1186 -6048
rect 1082 -6128 1186 -6112
rect 1082 -6192 1102 -6128
rect 1166 -6192 1186 -6128
rect 1082 -6208 1186 -6192
rect 1082 -6272 1102 -6208
rect 1166 -6272 1186 -6208
rect 1082 -6288 1186 -6272
rect 1082 -6352 1102 -6288
rect 1166 -6352 1186 -6288
rect 1082 -6368 1186 -6352
rect 1082 -6432 1102 -6368
rect 1166 -6432 1186 -6368
rect 1082 -6448 1186 -6432
rect 1082 -6512 1102 -6448
rect 1166 -6512 1186 -6448
rect 1082 -6528 1186 -6512
rect 1082 -6592 1102 -6528
rect 1166 -6592 1186 -6528
rect 1082 -6608 1186 -6592
rect 1082 -6672 1102 -6608
rect 1166 -6672 1186 -6608
rect 1082 -6688 1186 -6672
rect 1082 -6752 1102 -6688
rect 1166 -6752 1186 -6688
rect 1082 -6768 1186 -6752
rect 1082 -6832 1102 -6768
rect 1166 -6832 1186 -6768
rect 1082 -6848 1186 -6832
rect 1082 -6912 1102 -6848
rect 1166 -6912 1186 -6848
rect 1082 -6928 1186 -6912
rect 1082 -6992 1102 -6928
rect 1166 -6992 1186 -6928
rect 1082 -7008 1186 -6992
rect 1082 -7072 1102 -7008
rect 1166 -7072 1186 -7008
rect 1082 -7088 1186 -7072
rect 1082 -7152 1102 -7088
rect 1166 -7152 1186 -7088
rect 1082 -7168 1186 -7152
rect 1082 -7232 1102 -7168
rect 1166 -7232 1186 -7168
rect 1082 -7248 1186 -7232
rect 1082 -7312 1102 -7248
rect 1166 -7312 1186 -7248
rect 1082 -7328 1186 -7312
rect 1082 -7392 1102 -7328
rect 1166 -7392 1186 -7328
rect 1082 -7408 1186 -7392
rect 1082 -7472 1102 -7408
rect 1166 -7472 1186 -7408
rect 1082 -7488 1186 -7472
rect 1082 -7552 1102 -7488
rect 1166 -7552 1186 -7488
rect 1082 -7568 1186 -7552
rect 1082 -7632 1102 -7568
rect 1166 -7632 1186 -7568
rect 1082 -7648 1186 -7632
rect 1082 -7712 1102 -7648
rect 1166 -7712 1186 -7648
rect 1082 -7728 1186 -7712
rect 1082 -7792 1102 -7728
rect 1166 -7792 1186 -7728
rect 1082 -7808 1186 -7792
rect 1082 -7872 1102 -7808
rect 1166 -7872 1186 -7808
rect 1082 -7888 1186 -7872
rect -1530 -8120 -1426 -7952
rect -198 -8120 -94 -7921
rect 1082 -7952 1102 -7888
rect 1166 -7952 1186 -7888
rect 1505 -6008 3427 -5999
rect 1505 -7912 1514 -6008
rect 3418 -7912 3427 -6008
rect 1505 -7921 3427 -7912
rect 3694 -6032 3714 -5968
rect 3778 -6032 3798 -5968
rect 5026 -5999 5130 -5601
rect 6306 -5632 6326 -5568
rect 6390 -5632 6410 -5568
rect 6729 -3688 8651 -3679
rect 6729 -5592 6738 -3688
rect 8642 -5592 8651 -3688
rect 6729 -5601 8651 -5592
rect 8918 -3712 8938 -3648
rect 9002 -3712 9022 -3648
rect 8918 -3728 9022 -3712
rect 8918 -3792 8938 -3728
rect 9002 -3792 9022 -3728
rect 8918 -3808 9022 -3792
rect 8918 -3872 8938 -3808
rect 9002 -3872 9022 -3808
rect 8918 -3888 9022 -3872
rect 8918 -3952 8938 -3888
rect 9002 -3952 9022 -3888
rect 8918 -3968 9022 -3952
rect 8918 -4032 8938 -3968
rect 9002 -4032 9022 -3968
rect 8918 -4048 9022 -4032
rect 8918 -4112 8938 -4048
rect 9002 -4112 9022 -4048
rect 8918 -4128 9022 -4112
rect 8918 -4192 8938 -4128
rect 9002 -4192 9022 -4128
rect 8918 -4208 9022 -4192
rect 8918 -4272 8938 -4208
rect 9002 -4272 9022 -4208
rect 8918 -4288 9022 -4272
rect 8918 -4352 8938 -4288
rect 9002 -4352 9022 -4288
rect 8918 -4368 9022 -4352
rect 8918 -4432 8938 -4368
rect 9002 -4432 9022 -4368
rect 8918 -4448 9022 -4432
rect 8918 -4512 8938 -4448
rect 9002 -4512 9022 -4448
rect 8918 -4528 9022 -4512
rect 8918 -4592 8938 -4528
rect 9002 -4592 9022 -4528
rect 8918 -4608 9022 -4592
rect 8918 -4672 8938 -4608
rect 9002 -4672 9022 -4608
rect 8918 -4688 9022 -4672
rect 8918 -4752 8938 -4688
rect 9002 -4752 9022 -4688
rect 8918 -4768 9022 -4752
rect 8918 -4832 8938 -4768
rect 9002 -4832 9022 -4768
rect 8918 -4848 9022 -4832
rect 8918 -4912 8938 -4848
rect 9002 -4912 9022 -4848
rect 8918 -4928 9022 -4912
rect 8918 -4992 8938 -4928
rect 9002 -4992 9022 -4928
rect 8918 -5008 9022 -4992
rect 8918 -5072 8938 -5008
rect 9002 -5072 9022 -5008
rect 8918 -5088 9022 -5072
rect 8918 -5152 8938 -5088
rect 9002 -5152 9022 -5088
rect 8918 -5168 9022 -5152
rect 8918 -5232 8938 -5168
rect 9002 -5232 9022 -5168
rect 8918 -5248 9022 -5232
rect 8918 -5312 8938 -5248
rect 9002 -5312 9022 -5248
rect 8918 -5328 9022 -5312
rect 8918 -5392 8938 -5328
rect 9002 -5392 9022 -5328
rect 8918 -5408 9022 -5392
rect 8918 -5472 8938 -5408
rect 9002 -5472 9022 -5408
rect 8918 -5488 9022 -5472
rect 8918 -5552 8938 -5488
rect 9002 -5552 9022 -5488
rect 8918 -5568 9022 -5552
rect 6306 -5968 6410 -5632
rect 3694 -6048 3798 -6032
rect 3694 -6112 3714 -6048
rect 3778 -6112 3798 -6048
rect 3694 -6128 3798 -6112
rect 3694 -6192 3714 -6128
rect 3778 -6192 3798 -6128
rect 3694 -6208 3798 -6192
rect 3694 -6272 3714 -6208
rect 3778 -6272 3798 -6208
rect 3694 -6288 3798 -6272
rect 3694 -6352 3714 -6288
rect 3778 -6352 3798 -6288
rect 3694 -6368 3798 -6352
rect 3694 -6432 3714 -6368
rect 3778 -6432 3798 -6368
rect 3694 -6448 3798 -6432
rect 3694 -6512 3714 -6448
rect 3778 -6512 3798 -6448
rect 3694 -6528 3798 -6512
rect 3694 -6592 3714 -6528
rect 3778 -6592 3798 -6528
rect 3694 -6608 3798 -6592
rect 3694 -6672 3714 -6608
rect 3778 -6672 3798 -6608
rect 3694 -6688 3798 -6672
rect 3694 -6752 3714 -6688
rect 3778 -6752 3798 -6688
rect 3694 -6768 3798 -6752
rect 3694 -6832 3714 -6768
rect 3778 -6832 3798 -6768
rect 3694 -6848 3798 -6832
rect 3694 -6912 3714 -6848
rect 3778 -6912 3798 -6848
rect 3694 -6928 3798 -6912
rect 3694 -6992 3714 -6928
rect 3778 -6992 3798 -6928
rect 3694 -7008 3798 -6992
rect 3694 -7072 3714 -7008
rect 3778 -7072 3798 -7008
rect 3694 -7088 3798 -7072
rect 3694 -7152 3714 -7088
rect 3778 -7152 3798 -7088
rect 3694 -7168 3798 -7152
rect 3694 -7232 3714 -7168
rect 3778 -7232 3798 -7168
rect 3694 -7248 3798 -7232
rect 3694 -7312 3714 -7248
rect 3778 -7312 3798 -7248
rect 3694 -7328 3798 -7312
rect 3694 -7392 3714 -7328
rect 3778 -7392 3798 -7328
rect 3694 -7408 3798 -7392
rect 3694 -7472 3714 -7408
rect 3778 -7472 3798 -7408
rect 3694 -7488 3798 -7472
rect 3694 -7552 3714 -7488
rect 3778 -7552 3798 -7488
rect 3694 -7568 3798 -7552
rect 3694 -7632 3714 -7568
rect 3778 -7632 3798 -7568
rect 3694 -7648 3798 -7632
rect 3694 -7712 3714 -7648
rect 3778 -7712 3798 -7648
rect 3694 -7728 3798 -7712
rect 3694 -7792 3714 -7728
rect 3778 -7792 3798 -7728
rect 3694 -7808 3798 -7792
rect 3694 -7872 3714 -7808
rect 3778 -7872 3798 -7808
rect 3694 -7888 3798 -7872
rect 1082 -8120 1186 -7952
rect 2414 -8120 2518 -7921
rect 3694 -7952 3714 -7888
rect 3778 -7952 3798 -7888
rect 4117 -6008 6039 -5999
rect 4117 -7912 4126 -6008
rect 6030 -7912 6039 -6008
rect 4117 -7921 6039 -7912
rect 6306 -6032 6326 -5968
rect 6390 -6032 6410 -5968
rect 7638 -5999 7742 -5601
rect 8918 -5632 8938 -5568
rect 9002 -5632 9022 -5568
rect 8918 -5968 9022 -5632
rect 6306 -6048 6410 -6032
rect 6306 -6112 6326 -6048
rect 6390 -6112 6410 -6048
rect 6306 -6128 6410 -6112
rect 6306 -6192 6326 -6128
rect 6390 -6192 6410 -6128
rect 6306 -6208 6410 -6192
rect 6306 -6272 6326 -6208
rect 6390 -6272 6410 -6208
rect 6306 -6288 6410 -6272
rect 6306 -6352 6326 -6288
rect 6390 -6352 6410 -6288
rect 6306 -6368 6410 -6352
rect 6306 -6432 6326 -6368
rect 6390 -6432 6410 -6368
rect 6306 -6448 6410 -6432
rect 6306 -6512 6326 -6448
rect 6390 -6512 6410 -6448
rect 6306 -6528 6410 -6512
rect 6306 -6592 6326 -6528
rect 6390 -6592 6410 -6528
rect 6306 -6608 6410 -6592
rect 6306 -6672 6326 -6608
rect 6390 -6672 6410 -6608
rect 6306 -6688 6410 -6672
rect 6306 -6752 6326 -6688
rect 6390 -6752 6410 -6688
rect 6306 -6768 6410 -6752
rect 6306 -6832 6326 -6768
rect 6390 -6832 6410 -6768
rect 6306 -6848 6410 -6832
rect 6306 -6912 6326 -6848
rect 6390 -6912 6410 -6848
rect 6306 -6928 6410 -6912
rect 6306 -6992 6326 -6928
rect 6390 -6992 6410 -6928
rect 6306 -7008 6410 -6992
rect 6306 -7072 6326 -7008
rect 6390 -7072 6410 -7008
rect 6306 -7088 6410 -7072
rect 6306 -7152 6326 -7088
rect 6390 -7152 6410 -7088
rect 6306 -7168 6410 -7152
rect 6306 -7232 6326 -7168
rect 6390 -7232 6410 -7168
rect 6306 -7248 6410 -7232
rect 6306 -7312 6326 -7248
rect 6390 -7312 6410 -7248
rect 6306 -7328 6410 -7312
rect 6306 -7392 6326 -7328
rect 6390 -7392 6410 -7328
rect 6306 -7408 6410 -7392
rect 6306 -7472 6326 -7408
rect 6390 -7472 6410 -7408
rect 6306 -7488 6410 -7472
rect 6306 -7552 6326 -7488
rect 6390 -7552 6410 -7488
rect 6306 -7568 6410 -7552
rect 6306 -7632 6326 -7568
rect 6390 -7632 6410 -7568
rect 6306 -7648 6410 -7632
rect 6306 -7712 6326 -7648
rect 6390 -7712 6410 -7648
rect 6306 -7728 6410 -7712
rect 6306 -7792 6326 -7728
rect 6390 -7792 6410 -7728
rect 6306 -7808 6410 -7792
rect 6306 -7872 6326 -7808
rect 6390 -7872 6410 -7808
rect 6306 -7888 6410 -7872
rect 3694 -8120 3798 -7952
rect 5026 -8120 5130 -7921
rect 6306 -7952 6326 -7888
rect 6390 -7952 6410 -7888
rect 6729 -6008 8651 -5999
rect 6729 -7912 6738 -6008
rect 8642 -7912 8651 -6008
rect 6729 -7921 8651 -7912
rect 8918 -6032 8938 -5968
rect 9002 -6032 9022 -5968
rect 8918 -6048 9022 -6032
rect 8918 -6112 8938 -6048
rect 9002 -6112 9022 -6048
rect 8918 -6128 9022 -6112
rect 8918 -6192 8938 -6128
rect 9002 -6192 9022 -6128
rect 8918 -6208 9022 -6192
rect 8918 -6272 8938 -6208
rect 9002 -6272 9022 -6208
rect 8918 -6288 9022 -6272
rect 8918 -6352 8938 -6288
rect 9002 -6352 9022 -6288
rect 8918 -6368 9022 -6352
rect 8918 -6432 8938 -6368
rect 9002 -6432 9022 -6368
rect 8918 -6448 9022 -6432
rect 8918 -6512 8938 -6448
rect 9002 -6512 9022 -6448
rect 8918 -6528 9022 -6512
rect 8918 -6592 8938 -6528
rect 9002 -6592 9022 -6528
rect 8918 -6608 9022 -6592
rect 8918 -6672 8938 -6608
rect 9002 -6672 9022 -6608
rect 8918 -6688 9022 -6672
rect 8918 -6752 8938 -6688
rect 9002 -6752 9022 -6688
rect 8918 -6768 9022 -6752
rect 8918 -6832 8938 -6768
rect 9002 -6832 9022 -6768
rect 8918 -6848 9022 -6832
rect 8918 -6912 8938 -6848
rect 9002 -6912 9022 -6848
rect 8918 -6928 9022 -6912
rect 8918 -6992 8938 -6928
rect 9002 -6992 9022 -6928
rect 8918 -7008 9022 -6992
rect 8918 -7072 8938 -7008
rect 9002 -7072 9022 -7008
rect 8918 -7088 9022 -7072
rect 8918 -7152 8938 -7088
rect 9002 -7152 9022 -7088
rect 8918 -7168 9022 -7152
rect 8918 -7232 8938 -7168
rect 9002 -7232 9022 -7168
rect 8918 -7248 9022 -7232
rect 8918 -7312 8938 -7248
rect 9002 -7312 9022 -7248
rect 8918 -7328 9022 -7312
rect 8918 -7392 8938 -7328
rect 9002 -7392 9022 -7328
rect 8918 -7408 9022 -7392
rect 8918 -7472 8938 -7408
rect 9002 -7472 9022 -7408
rect 8918 -7488 9022 -7472
rect 8918 -7552 8938 -7488
rect 9002 -7552 9022 -7488
rect 8918 -7568 9022 -7552
rect 8918 -7632 8938 -7568
rect 9002 -7632 9022 -7568
rect 8918 -7648 9022 -7632
rect 8918 -7712 8938 -7648
rect 9002 -7712 9022 -7648
rect 8918 -7728 9022 -7712
rect 8918 -7792 8938 -7728
rect 9002 -7792 9022 -7728
rect 8918 -7808 9022 -7792
rect 8918 -7872 8938 -7808
rect 9002 -7872 9022 -7808
rect 8918 -7888 9022 -7872
rect 6306 -8120 6410 -7952
rect 7638 -8120 7742 -7921
rect 8918 -7952 8938 -7888
rect 9002 -7952 9022 -7888
rect 8918 -8120 9022 -7952
<< properties >>
string FIXED_BBOX 6650 5920 8730 8000
<< end >>
